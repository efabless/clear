magic
tech sky130A
magscale 1 2
timestamp 1682506994
<< viali >>
rect 16865 24361 16899 24395
rect 24869 24361 24903 24395
rect 29009 24361 29043 24395
rect 39589 24361 39623 24395
rect 47041 24361 47075 24395
rect 47961 24361 47995 24395
rect 19441 24293 19475 24327
rect 26433 24293 26467 24327
rect 30481 24293 30515 24327
rect 39313 24293 39347 24327
rect 46765 24293 46799 24327
rect 3249 24225 3283 24259
rect 5825 24225 5859 24259
rect 6561 24225 6595 24259
rect 8217 24225 8251 24259
rect 13553 24225 13587 24259
rect 16129 24225 16163 24259
rect 18705 24225 18739 24259
rect 20913 24225 20947 24259
rect 34069 24225 34103 24259
rect 34253 24225 34287 24259
rect 35357 24225 35391 24259
rect 35541 24225 35575 24259
rect 36553 24225 36587 24259
rect 36737 24225 36771 24259
rect 37933 24225 37967 24259
rect 38117 24225 38151 24259
rect 41153 24225 41187 24259
rect 41429 24225 41463 24259
rect 45477 24225 45511 24259
rect 48513 24225 48547 24259
rect 48789 24225 48823 24259
rect 2237 24157 2271 24191
rect 4169 24157 4203 24191
rect 4813 24157 4847 24191
rect 7389 24157 7423 24191
rect 9321 24157 9355 24191
rect 9965 24157 9999 24191
rect 11897 24157 11931 24191
rect 12357 24157 12391 24191
rect 15117 24157 15151 24191
rect 17049 24157 17083 24191
rect 17693 24157 17727 24191
rect 19625 24157 19659 24191
rect 20085 24157 20119 24191
rect 22201 24157 22235 24191
rect 22937 24157 22971 24191
rect 24041 24157 24075 24191
rect 24777 24157 24811 24191
rect 25421 24157 25455 24191
rect 27261 24157 27295 24191
rect 28365 24157 28399 24191
rect 30849 24157 30883 24191
rect 32505 24157 32539 24191
rect 35265 24157 35299 24191
rect 37841 24157 37875 24191
rect 38669 24157 38703 24191
rect 40049 24157 40083 24191
rect 45201 24157 45235 24191
rect 47225 24157 47259 24191
rect 47869 24157 47903 24191
rect 10977 24089 11011 24123
rect 29837 24089 29871 24123
rect 30389 24089 30423 24123
rect 31769 24089 31803 24123
rect 33149 24089 33183 24123
rect 33977 24089 34011 24123
rect 40693 24089 40727 24123
rect 42625 24089 42659 24123
rect 46581 24089 46615 24123
rect 3985 24021 4019 24055
rect 9137 24021 9171 24055
rect 11713 24021 11747 24055
rect 14289 24021 14323 24055
rect 23857 24021 23891 24055
rect 26065 24021 26099 24055
rect 26525 24021 26559 24055
rect 26709 24021 26743 24055
rect 27905 24021 27939 24055
rect 29285 24021 29319 24055
rect 29929 24021 29963 24055
rect 31493 24021 31527 24055
rect 32137 24021 32171 24055
rect 33609 24021 33643 24055
rect 34897 24021 34931 24055
rect 36093 24021 36127 24055
rect 36461 24021 36495 24055
rect 37473 24021 37507 24055
rect 44097 24021 44131 24055
rect 44741 24021 44775 24055
rect 20545 23817 20579 23851
rect 20913 23817 20947 23851
rect 22385 23817 22419 23851
rect 22477 23817 22511 23851
rect 23489 23817 23523 23851
rect 29377 23817 29411 23851
rect 32321 23817 32355 23851
rect 35265 23817 35299 23851
rect 35633 23817 35667 23851
rect 36277 23817 36311 23851
rect 38853 23817 38887 23851
rect 47961 23817 47995 23851
rect 1777 23749 1811 23783
rect 2145 23749 2179 23783
rect 9137 23749 9171 23783
rect 10701 23749 10735 23783
rect 14289 23749 14323 23783
rect 16129 23749 16163 23783
rect 18153 23749 18187 23783
rect 21281 23749 21315 23783
rect 24409 23749 24443 23783
rect 25145 23749 25179 23783
rect 33793 23749 33827 23783
rect 37933 23749 37967 23783
rect 40693 23749 40727 23783
rect 47869 23749 47903 23783
rect 2973 23681 3007 23715
rect 4813 23681 4847 23715
rect 6837 23681 6871 23715
rect 7941 23681 7975 23715
rect 9965 23681 9999 23715
rect 11805 23681 11839 23715
rect 12081 23681 12115 23715
rect 13277 23681 13311 23715
rect 14933 23681 14967 23715
rect 17141 23681 17175 23715
rect 18797 23681 18831 23715
rect 23799 23681 23833 23715
rect 27169 23681 27203 23715
rect 28273 23681 28307 23715
rect 29561 23681 29595 23715
rect 32689 23681 32723 23715
rect 37841 23681 37875 23715
rect 39221 23681 39255 23715
rect 39313 23681 39347 23715
rect 40049 23681 40083 23715
rect 41429 23681 41463 23715
rect 42625 23681 42659 23715
rect 44189 23681 44223 23715
rect 45477 23681 45511 23715
rect 46489 23681 46523 23715
rect 48513 23681 48547 23715
rect 3985 23613 4019 23647
rect 5457 23613 5491 23647
rect 19073 23613 19107 23647
rect 22569 23613 22603 23647
rect 23121 23613 23155 23647
rect 24869 23613 24903 23647
rect 30021 23613 30055 23647
rect 30297 23613 30331 23647
rect 32781 23613 32815 23647
rect 32965 23613 32999 23647
rect 33517 23613 33551 23647
rect 36369 23613 36403 23647
rect 36461 23613 36495 23647
rect 38025 23613 38059 23647
rect 39405 23613 39439 23647
rect 41153 23613 41187 23647
rect 42901 23613 42935 23647
rect 43913 23613 43947 23647
rect 45201 23613 45235 23647
rect 47225 23613 47259 23647
rect 49249 23613 49283 23647
rect 2329 23545 2363 23579
rect 6561 23545 6595 23579
rect 21465 23545 21499 23579
rect 22017 23545 22051 23579
rect 28917 23545 28951 23579
rect 37473 23545 37507 23579
rect 49433 23545 49467 23579
rect 7481 23477 7515 23511
rect 23305 23477 23339 23511
rect 26617 23477 26651 23511
rect 27813 23477 27847 23511
rect 31769 23477 31803 23511
rect 35909 23477 35943 23511
rect 36921 23477 36955 23511
rect 38485 23477 38519 23511
rect 46673 23477 46707 23511
rect 47133 23477 47167 23511
rect 48697 23477 48731 23511
rect 49065 23477 49099 23511
rect 3617 23273 3651 23307
rect 19717 23273 19751 23307
rect 27905 23273 27939 23307
rect 29745 23273 29779 23307
rect 38945 23273 38979 23307
rect 40049 23273 40083 23307
rect 41061 23273 41095 23307
rect 43913 23273 43947 23307
rect 44833 23273 44867 23307
rect 47593 23273 47627 23307
rect 47961 23273 47995 23307
rect 48513 23273 48547 23307
rect 49249 23273 49283 23307
rect 24041 23205 24075 23239
rect 30941 23205 30975 23239
rect 39497 23205 39531 23239
rect 39681 23205 39715 23239
rect 47869 23205 47903 23239
rect 4261 23137 4295 23171
rect 6101 23137 6135 23171
rect 7849 23137 7883 23171
rect 9413 23137 9447 23171
rect 11253 23137 11287 23171
rect 13369 23137 13403 23171
rect 14289 23137 14323 23171
rect 16405 23137 16439 23171
rect 17417 23137 17451 23171
rect 20361 23137 20395 23171
rect 23029 23137 23063 23171
rect 23121 23137 23155 23171
rect 25697 23137 25731 23171
rect 25973 23137 26007 23171
rect 28365 23137 28399 23171
rect 28457 23137 28491 23171
rect 30205 23137 30239 23171
rect 30297 23137 30331 23171
rect 31677 23137 31711 23171
rect 34345 23137 34379 23171
rect 34989 23137 35023 23171
rect 37197 23137 37231 23171
rect 40693 23137 40727 23171
rect 41521 23137 41555 23171
rect 45201 23137 45235 23171
rect 1777 23069 1811 23103
rect 3433 23069 3467 23103
rect 3985 23069 4019 23103
rect 5365 23069 5399 23103
rect 7205 23069 7239 23103
rect 9137 23069 9171 23103
rect 10701 23069 10735 23103
rect 12449 23069 12483 23103
rect 15485 23069 15519 23103
rect 17141 23069 17175 23103
rect 19901 23069 19935 23103
rect 23857 23069 23891 23103
rect 24593 23069 24627 23103
rect 31401 23069 31435 23103
rect 33701 23069 33735 23103
rect 40417 23069 40451 23103
rect 44281 23069 44315 23103
rect 45477 23069 45511 23103
rect 46489 23069 46523 23103
rect 46765 23069 46799 23103
rect 48329 23069 48363 23103
rect 49065 23069 49099 23103
rect 2789 23001 2823 23035
rect 14657 23001 14691 23035
rect 14841 23001 14875 23035
rect 19441 23001 19475 23035
rect 20637 23001 20671 23035
rect 35265 23001 35299 23035
rect 37473 23001 37507 23035
rect 40509 23001 40543 23035
rect 41797 23001 41831 23035
rect 43545 23001 43579 23035
rect 44465 23001 44499 23035
rect 18889 22933 18923 22967
rect 22109 22933 22143 22967
rect 22569 22933 22603 22967
rect 22937 22933 22971 22967
rect 25237 22933 25271 22967
rect 27445 22933 27479 22967
rect 28273 22933 28307 22967
rect 29009 22933 29043 22967
rect 29193 22933 29227 22967
rect 29377 22933 29411 22967
rect 30113 22933 30147 22967
rect 30757 22933 30791 22967
rect 33149 22933 33183 22967
rect 36737 22933 36771 22967
rect 39313 22933 39347 22967
rect 18613 22729 18647 22763
rect 19073 22729 19107 22763
rect 27353 22729 27387 22763
rect 31585 22729 31619 22763
rect 32321 22729 32355 22763
rect 33425 22729 33459 22763
rect 36093 22729 36127 22763
rect 41521 22729 41555 22763
rect 46949 22729 46983 22763
rect 47777 22729 47811 22763
rect 48513 22729 48547 22763
rect 49249 22729 49283 22763
rect 15853 22661 15887 22695
rect 17141 22661 17175 22695
rect 22293 22661 22327 22695
rect 27813 22661 27847 22695
rect 30665 22661 30699 22695
rect 33977 22661 34011 22695
rect 37749 22661 37783 22695
rect 41889 22661 41923 22695
rect 42073 22661 42107 22695
rect 42257 22661 42291 22695
rect 47593 22661 47627 22695
rect 1777 22593 1811 22627
rect 3617 22593 3651 22627
rect 3985 22593 4019 22627
rect 4629 22593 4663 22627
rect 6837 22593 6871 22627
rect 7481 22593 7515 22627
rect 9781 22593 9815 22627
rect 13093 22593 13127 22627
rect 15117 22593 15151 22627
rect 16865 22593 16899 22627
rect 22017 22593 22051 22627
rect 24869 22593 24903 22627
rect 27261 22593 27295 22627
rect 30757 22593 30791 22627
rect 32689 22593 32723 22627
rect 33701 22593 33735 22627
rect 36461 22593 36495 22627
rect 37473 22593 37507 22627
rect 40049 22593 40083 22627
rect 40877 22593 40911 22627
rect 42809 22593 42843 22627
rect 43545 22593 43579 22627
rect 44833 22593 44867 22627
rect 45845 22593 45879 22627
rect 47133 22593 47167 22627
rect 48329 22593 48363 22627
rect 49065 22593 49099 22627
rect 2789 22525 2823 22559
rect 4169 22525 4203 22559
rect 5089 22525 5123 22559
rect 7941 22525 7975 22559
rect 10241 22525 10275 22559
rect 11713 22525 11747 22559
rect 11989 22525 12023 22559
rect 13829 22525 13863 22559
rect 19533 22525 19567 22559
rect 19809 22525 19843 22559
rect 21281 22525 21315 22559
rect 23765 22525 23799 22559
rect 24225 22525 24259 22559
rect 25145 22525 25179 22559
rect 28089 22525 28123 22559
rect 28365 22525 28399 22559
rect 30849 22525 30883 22559
rect 32781 22525 32815 22559
rect 32873 22525 32907 22559
rect 36553 22525 36587 22559
rect 36737 22525 36771 22559
rect 39221 22525 39255 22559
rect 40141 22525 40175 22559
rect 40233 22525 40267 22559
rect 43269 22525 43303 22559
rect 44557 22525 44591 22559
rect 46121 22525 46155 22559
rect 47317 22525 47351 22559
rect 6469 22457 6503 22491
rect 35449 22457 35483 22491
rect 42625 22457 42659 22491
rect 48053 22457 48087 22491
rect 6929 22389 6963 22423
rect 9321 22389 9355 22423
rect 9505 22389 9539 22423
rect 19257 22389 19291 22423
rect 24317 22389 24351 22423
rect 24593 22389 24627 22423
rect 26617 22389 26651 22423
rect 29837 22389 29871 22423
rect 30297 22389 30331 22423
rect 35817 22389 35851 22423
rect 39681 22389 39715 22423
rect 15466 22185 15500 22219
rect 21452 22185 21486 22219
rect 24593 22185 24627 22219
rect 30389 22185 30423 22219
rect 37552 22185 37586 22219
rect 41245 22185 41279 22219
rect 44557 22185 44591 22219
rect 44833 22185 44867 22219
rect 47869 22185 47903 22219
rect 28365 22117 28399 22151
rect 32597 22117 32631 22151
rect 42901 22117 42935 22151
rect 45201 22117 45235 22151
rect 47593 22117 47627 22151
rect 2053 22049 2087 22083
rect 4445 22049 4479 22083
rect 6745 22049 6779 22083
rect 8585 22049 8619 22083
rect 9873 22049 9907 22083
rect 11253 22049 11287 22083
rect 11713 22049 11747 22083
rect 12449 22049 12483 22083
rect 13921 22049 13955 22083
rect 14749 22049 14783 22083
rect 20545 22049 20579 22083
rect 25145 22049 25179 22083
rect 26525 22049 26559 22083
rect 27721 22049 27755 22083
rect 28963 22049 28997 22083
rect 30849 22049 30883 22083
rect 33517 22049 33551 22083
rect 33609 22049 33643 22083
rect 34069 22049 34103 22083
rect 35357 22049 35391 22083
rect 35541 22049 35575 22083
rect 36737 22049 36771 22083
rect 39037 22049 39071 22083
rect 40601 22049 40635 22083
rect 41797 22049 41831 22083
rect 42441 22049 42475 22083
rect 43545 22049 43579 22083
rect 45845 22049 45879 22083
rect 48053 22049 48087 22083
rect 1777 21981 1811 22015
rect 4077 21981 4111 22015
rect 6009 21981 6043 22015
rect 7941 21981 7975 22015
rect 9137 21981 9171 22015
rect 11989 21981 12023 22015
rect 15209 21981 15243 22015
rect 17509 21981 17543 22015
rect 19533 21981 19567 22015
rect 19717 21981 19751 22015
rect 21189 21981 21223 22015
rect 23397 21981 23431 22015
rect 24041 21981 24075 22015
rect 25053 21981 25087 22015
rect 28733 21981 28767 22015
rect 29745 21981 29779 22015
rect 37289 21981 37323 22015
rect 39497 21981 39531 22015
rect 43269 21981 43303 22015
rect 45385 21981 45419 22015
rect 46121 21981 46155 22015
rect 47317 21981 47351 22015
rect 48329 21981 48363 22015
rect 7573 21913 7607 21947
rect 11069 21913 11103 21947
rect 13737 21913 13771 21947
rect 14565 21913 14599 21947
rect 18429 21913 18463 21947
rect 20361 21913 20395 21947
rect 26433 21913 26467 21947
rect 31125 21913 31159 21947
rect 33425 21913 33459 21947
rect 34345 21913 34379 21947
rect 39589 21913 39623 21947
rect 40417 21913 40451 21947
rect 44465 21913 44499 21947
rect 49157 21913 49191 21947
rect 49341 21913 49375 21947
rect 14197 21845 14231 21879
rect 16957 21845 16991 21879
rect 19349 21845 19383 21879
rect 19993 21845 20027 21879
rect 20453 21845 20487 21879
rect 22937 21845 22971 21879
rect 24961 21845 24995 21879
rect 25605 21845 25639 21879
rect 25973 21845 26007 21879
rect 26341 21845 26375 21879
rect 27169 21845 27203 21879
rect 27537 21845 27571 21879
rect 27629 21845 27663 21879
rect 28825 21845 28859 21879
rect 33057 21845 33091 21879
rect 34529 21845 34563 21879
rect 34897 21845 34931 21879
rect 35265 21845 35299 21879
rect 36093 21845 36127 21879
rect 36461 21845 36495 21879
rect 36553 21845 36587 21879
rect 40049 21845 40083 21879
rect 40509 21845 40543 21879
rect 41613 21845 41647 21879
rect 41705 21845 41739 21879
rect 47133 21845 47167 21879
rect 48513 21845 48547 21879
rect 5273 21641 5307 21675
rect 11805 21641 11839 21675
rect 13185 21641 13219 21675
rect 14749 21641 14783 21675
rect 15117 21641 15151 21675
rect 16221 21641 16255 21675
rect 17325 21641 17359 21675
rect 21097 21641 21131 21675
rect 25145 21641 25179 21675
rect 27169 21641 27203 21675
rect 28365 21641 28399 21675
rect 28733 21641 28767 21675
rect 29929 21641 29963 21675
rect 31861 21641 31895 21675
rect 36093 21641 36127 21675
rect 40233 21641 40267 21675
rect 46305 21641 46339 21675
rect 47961 21641 47995 21675
rect 4353 21573 4387 21607
rect 27629 21573 27663 21607
rect 30021 21573 30055 21607
rect 31125 21573 31159 21607
rect 34897 21573 34931 21607
rect 36921 21573 36955 21607
rect 37657 21573 37691 21607
rect 47593 21573 47627 21607
rect 48421 21573 48455 21607
rect 1685 21505 1719 21539
rect 3617 21505 3651 21539
rect 5825 21505 5859 21539
rect 6561 21505 6595 21539
rect 8401 21505 8435 21539
rect 10517 21505 10551 21539
rect 11989 21505 12023 21539
rect 12541 21505 12575 21539
rect 13645 21505 13679 21539
rect 15209 21505 15243 21539
rect 16129 21505 16163 21539
rect 17233 21505 17267 21539
rect 21189 21505 21223 21539
rect 21925 21505 21959 21539
rect 22477 21505 22511 21539
rect 25973 21505 26007 21539
rect 26617 21505 26651 21539
rect 27537 21505 27571 21539
rect 31217 21505 31251 21539
rect 33609 21505 33643 21539
rect 34805 21505 34839 21539
rect 40601 21505 40635 21539
rect 41429 21505 41463 21539
rect 42625 21505 42659 21539
rect 43913 21505 43947 21539
rect 44557 21505 44591 21539
rect 45201 21505 45235 21539
rect 45845 21505 45879 21539
rect 46489 21505 46523 21539
rect 47133 21505 47167 21539
rect 47777 21505 47811 21539
rect 49065 21505 49099 21539
rect 2053 21437 2087 21471
rect 6009 21437 6043 21471
rect 7021 21437 7055 21471
rect 8861 21437 8895 21471
rect 11161 21437 11195 21471
rect 15301 21437 15335 21471
rect 17417 21437 17451 21471
rect 18061 21437 18095 21471
rect 18337 21437 18371 21471
rect 21373 21437 21407 21471
rect 22753 21437 22787 21471
rect 25237 21437 25271 21471
rect 25329 21437 25363 21471
rect 27721 21437 27755 21471
rect 28825 21437 28859 21471
rect 28917 21437 28951 21471
rect 30113 21437 30147 21471
rect 31309 21437 31343 21471
rect 32321 21437 32355 21471
rect 33701 21437 33735 21471
rect 33885 21437 33919 21471
rect 35081 21437 35115 21471
rect 36185 21437 36219 21471
rect 36369 21437 36403 21471
rect 38025 21437 38059 21471
rect 38301 21437 38335 21471
rect 40693 21437 40727 21471
rect 40785 21437 40819 21471
rect 5457 21369 5491 21403
rect 14289 21369 14323 21403
rect 20269 21369 20303 21403
rect 24225 21369 24259 21403
rect 29561 21369 29595 21403
rect 32781 21369 32815 21403
rect 33241 21369 33275 21403
rect 37473 21369 37507 21403
rect 48605 21369 48639 21403
rect 10149 21301 10183 21335
rect 16865 21301 16899 21335
rect 19809 21301 19843 21335
rect 20361 21301 20395 21335
rect 20729 21301 20763 21335
rect 22109 21301 22143 21335
rect 24777 21301 24811 21335
rect 30757 21301 30791 21335
rect 34437 21301 34471 21335
rect 35725 21301 35759 21335
rect 36829 21301 36863 21335
rect 37381 21301 37415 21335
rect 39773 21301 39807 21335
rect 42073 21301 42107 21335
rect 43269 21301 43303 21335
rect 43729 21301 43763 21335
rect 44373 21301 44407 21335
rect 45017 21301 45051 21335
rect 45661 21301 45695 21335
rect 46949 21301 46983 21335
rect 49249 21301 49283 21335
rect 7665 21097 7699 21131
rect 8493 21097 8527 21131
rect 10333 21097 10367 21131
rect 16957 21097 16991 21131
rect 18153 21097 18187 21131
rect 22017 21097 22051 21131
rect 27905 21097 27939 21131
rect 28365 21097 28399 21131
rect 30757 21097 30791 21131
rect 36921 21097 36955 21131
rect 37105 21097 37139 21131
rect 39405 21097 39439 21131
rect 40049 21097 40083 21131
rect 44373 21097 44407 21131
rect 45845 21097 45879 21131
rect 46029 21097 46063 21131
rect 47041 21097 47075 21131
rect 47777 21097 47811 21131
rect 48421 21097 48455 21131
rect 9045 21029 9079 21063
rect 9229 21029 9263 21063
rect 9413 21029 9447 21063
rect 13001 21029 13035 21063
rect 19809 21029 19843 21063
rect 22845 21029 22879 21063
rect 23305 21029 23339 21063
rect 29745 21029 29779 21063
rect 31861 21029 31895 21063
rect 45201 21029 45235 21063
rect 4445 20961 4479 20995
rect 6285 20961 6319 20995
rect 13645 20961 13679 20995
rect 14381 20961 14415 20995
rect 17417 20961 17451 20995
rect 17509 20961 17543 20995
rect 18705 20961 18739 20995
rect 20269 20961 20303 20995
rect 23765 20961 23799 20995
rect 23857 20961 23891 20995
rect 26341 20961 26375 20995
rect 27537 20961 27571 20995
rect 28825 20961 28859 20995
rect 28917 20961 28951 20995
rect 31217 20961 31251 20995
rect 31401 20961 31435 20995
rect 32781 20961 32815 20995
rect 34897 20961 34931 20995
rect 35173 20961 35207 20995
rect 37933 20961 37967 20995
rect 40509 20961 40543 20995
rect 40601 20961 40635 20995
rect 41797 20961 41831 20995
rect 42441 20961 42475 20995
rect 42717 20961 42751 20995
rect 1777 20893 1811 20927
rect 4077 20893 4111 20927
rect 6009 20893 6043 20927
rect 7849 20893 7883 20927
rect 9733 20893 9767 20927
rect 10793 20893 10827 20927
rect 11897 20893 11931 20927
rect 13369 20893 13403 20927
rect 14657 20893 14691 20927
rect 22661 20893 22695 20927
rect 24593 20893 24627 20927
rect 27261 20893 27295 20927
rect 29929 20893 29963 20927
rect 31953 20893 31987 20927
rect 32505 20893 32539 20927
rect 37657 20893 37691 20927
rect 41613 20893 41647 20927
rect 43913 20893 43947 20927
rect 44557 20893 44591 20927
rect 45385 20893 45419 20927
rect 45661 20893 45695 20927
rect 46581 20893 46615 20927
rect 47225 20893 47259 20927
rect 47961 20893 47995 20927
rect 48605 20893 48639 20927
rect 49065 20893 49099 20927
rect 2789 20825 2823 20859
rect 8401 20825 8435 20859
rect 11437 20825 11471 20859
rect 14933 20825 14967 20859
rect 17969 20825 18003 20859
rect 18521 20825 18555 20859
rect 19625 20825 19659 20859
rect 20545 20825 20579 20859
rect 27353 20825 27387 20859
rect 30481 20825 30515 20859
rect 40417 20825 40451 20859
rect 41705 20825 41739 20859
rect 12541 20757 12575 20791
rect 13461 20757 13495 20791
rect 14197 20757 14231 20791
rect 16405 20757 16439 20791
rect 17325 20757 17359 20791
rect 18613 20757 18647 20791
rect 23673 20757 23707 20791
rect 25237 20757 25271 20791
rect 25697 20757 25731 20791
rect 26065 20757 26099 20791
rect 26157 20757 26191 20791
rect 26893 20757 26927 20791
rect 28733 20757 28767 20791
rect 30205 20757 30239 20791
rect 31125 20757 31159 20791
rect 32137 20757 32171 20791
rect 34253 20757 34287 20791
rect 36645 20757 36679 20791
rect 37289 20757 37323 20791
rect 41245 20757 41279 20791
rect 43729 20757 43763 20791
rect 46397 20757 46431 20791
rect 49249 20757 49283 20791
rect 8309 20553 8343 20587
rect 8401 20553 8435 20587
rect 13369 20553 13403 20587
rect 20729 20553 20763 20587
rect 22017 20553 22051 20587
rect 22753 20553 22787 20587
rect 26709 20553 26743 20587
rect 29009 20553 29043 20587
rect 29929 20553 29963 20587
rect 34069 20553 34103 20587
rect 34621 20553 34655 20587
rect 36093 20553 36127 20587
rect 36553 20553 36587 20587
rect 42165 20553 42199 20587
rect 43085 20553 43119 20587
rect 43821 20553 43855 20587
rect 44281 20553 44315 20587
rect 44649 20553 44683 20587
rect 44833 20553 44867 20587
rect 46581 20553 46615 20587
rect 47041 20553 47075 20587
rect 48053 20553 48087 20587
rect 5549 20485 5583 20519
rect 6193 20485 6227 20519
rect 11713 20485 11747 20519
rect 12265 20485 12299 20519
rect 26617 20485 26651 20519
rect 31125 20485 31159 20519
rect 31861 20485 31895 20519
rect 34345 20485 34379 20519
rect 38025 20485 38059 20519
rect 40325 20485 40359 20519
rect 42625 20485 42659 20519
rect 44373 20485 44407 20519
rect 46673 20485 46707 20519
rect 47225 20485 47259 20519
rect 1777 20417 1811 20451
rect 3617 20417 3651 20451
rect 5365 20417 5399 20451
rect 6561 20417 6595 20451
rect 9137 20417 9171 20451
rect 9873 20417 9907 20451
rect 10517 20417 10551 20451
rect 12081 20417 12115 20451
rect 12725 20417 12759 20451
rect 16129 20417 16163 20451
rect 17325 20417 17359 20451
rect 17417 20417 17451 20451
rect 18061 20417 18095 20451
rect 18153 20417 18187 20451
rect 21097 20417 21131 20451
rect 22661 20417 22695 20451
rect 23305 20417 23339 20451
rect 23489 20417 23523 20451
rect 26249 20417 26283 20451
rect 27261 20417 27295 20451
rect 29837 20417 29871 20451
rect 31033 20417 31067 20451
rect 35265 20417 35299 20451
rect 35357 20417 35391 20451
rect 36461 20417 36495 20451
rect 37289 20417 37323 20451
rect 41153 20417 41187 20451
rect 43545 20417 43579 20451
rect 47317 20417 47351 20451
rect 47961 20417 47995 20451
rect 48605 20417 48639 20451
rect 49065 20417 49099 20451
rect 2789 20349 2823 20383
rect 3893 20349 3927 20383
rect 7205 20349 7239 20383
rect 9321 20349 9355 20383
rect 10057 20349 10091 20383
rect 13829 20349 13863 20383
rect 14105 20349 14139 20383
rect 15577 20349 15611 20383
rect 17509 20349 17543 20383
rect 18521 20349 18555 20383
rect 18797 20349 18831 20383
rect 21189 20349 21223 20383
rect 21373 20349 21407 20383
rect 22937 20349 22971 20383
rect 23857 20349 23891 20383
rect 24133 20349 24167 20383
rect 25605 20349 25639 20383
rect 27537 20349 27571 20383
rect 30113 20349 30147 20383
rect 31217 20349 31251 20383
rect 32321 20349 32355 20383
rect 32597 20349 32631 20383
rect 35541 20349 35575 20383
rect 36737 20349 36771 20383
rect 37749 20349 37783 20383
rect 40417 20349 40451 20383
rect 40601 20349 40635 20383
rect 43729 20349 43763 20383
rect 47777 20349 47811 20383
rect 6009 20281 6043 20315
rect 22293 20281 22327 20315
rect 26065 20281 26099 20315
rect 29469 20281 29503 20315
rect 43361 20281 43395 20315
rect 49249 20281 49283 20315
rect 11161 20213 11195 20247
rect 16221 20213 16255 20247
rect 16773 20213 16807 20247
rect 16957 20213 16991 20247
rect 20269 20213 20303 20247
rect 30665 20213 30699 20247
rect 31677 20213 31711 20247
rect 34897 20213 34931 20247
rect 39497 20213 39531 20247
rect 39957 20213 39991 20247
rect 41797 20213 41831 20247
rect 48421 20213 48455 20247
rect 10333 20009 10367 20043
rect 12246 20009 12280 20043
rect 15485 20009 15519 20043
rect 18797 20009 18831 20043
rect 19901 20009 19935 20043
rect 26801 20009 26835 20043
rect 29285 20009 29319 20043
rect 30941 20009 30975 20043
rect 37289 20009 37323 20043
rect 42625 20009 42659 20043
rect 43361 20009 43395 20043
rect 47225 20009 47259 20043
rect 47501 20009 47535 20043
rect 47777 20009 47811 20043
rect 14197 19941 14231 19975
rect 14381 19941 14415 19975
rect 19441 19941 19475 19975
rect 23213 19941 23247 19975
rect 29745 19941 29779 19975
rect 33425 19941 33459 19975
rect 39497 19941 39531 19975
rect 42349 19941 42383 19975
rect 48421 19941 48455 19975
rect 4537 19873 4571 19907
rect 6285 19873 6319 19907
rect 11989 19873 12023 19907
rect 17049 19873 17083 19907
rect 20729 19873 20763 19907
rect 23765 19873 23799 19907
rect 26157 19873 26191 19907
rect 27353 19873 27387 19907
rect 28641 19873 28675 19907
rect 30297 19873 30331 19907
rect 31401 19873 31435 19907
rect 31493 19873 31527 19907
rect 32597 19873 32631 19907
rect 32689 19873 32723 19907
rect 33885 19873 33919 19907
rect 34069 19873 34103 19907
rect 35541 19873 35575 19907
rect 36737 19873 36771 19907
rect 37841 19873 37875 19907
rect 38945 19873 38979 19907
rect 39129 19873 39163 19907
rect 40601 19873 40635 19907
rect 42257 19873 42291 19907
rect 49341 19873 49375 19907
rect 1777 19805 1811 19839
rect 4077 19805 4111 19839
rect 6009 19805 6043 19839
rect 7849 19805 7883 19839
rect 8401 19805 8435 19839
rect 10885 19805 10919 19839
rect 14841 19805 14875 19839
rect 15945 19805 15979 19839
rect 20453 19805 20487 19839
rect 24685 19805 24719 19839
rect 25145 19805 25179 19839
rect 27905 19805 27939 19839
rect 28457 19805 28491 19839
rect 30205 19805 30239 19839
rect 31309 19805 31343 19839
rect 32505 19805 32539 19839
rect 33793 19805 33827 19839
rect 38853 19805 38887 19839
rect 40417 19805 40451 19839
rect 40509 19805 40543 19839
rect 41245 19805 41279 19839
rect 43177 19805 43211 19839
rect 48145 19805 48179 19839
rect 48605 19805 48639 19839
rect 2789 19737 2823 19771
rect 9873 19737 9907 19771
rect 10241 19737 10275 19771
rect 17325 19737 17359 19771
rect 19809 19737 19843 19771
rect 22661 19737 22695 19771
rect 22937 19737 22971 19771
rect 23673 19737 23707 19771
rect 28365 19737 28399 19771
rect 34529 19737 34563 19771
rect 36553 19737 36587 19771
rect 42809 19737 42843 19771
rect 42993 19737 43027 19771
rect 47961 19737 47995 19771
rect 49157 19737 49191 19771
rect 7665 19669 7699 19703
rect 8493 19669 8527 19703
rect 9137 19669 9171 19703
rect 9229 19669 9263 19703
rect 11529 19669 11563 19703
rect 13737 19669 13771 19703
rect 14565 19669 14599 19703
rect 16589 19669 16623 19703
rect 22201 19669 22235 19703
rect 22477 19669 22511 19703
rect 23581 19669 23615 19703
rect 24501 19669 24535 19703
rect 24961 19669 24995 19703
rect 25605 19669 25639 19703
rect 25973 19669 26007 19703
rect 26065 19669 26099 19703
rect 27169 19669 27203 19703
rect 27261 19669 27295 19703
rect 27997 19669 28031 19703
rect 29101 19669 29135 19703
rect 30113 19669 30147 19703
rect 32137 19669 32171 19703
rect 34897 19669 34931 19703
rect 35265 19669 35299 19703
rect 35357 19669 35391 19703
rect 36093 19669 36127 19703
rect 36461 19669 36495 19703
rect 37657 19669 37691 19703
rect 37749 19669 37783 19703
rect 38485 19669 38519 19703
rect 40049 19669 40083 19703
rect 41889 19669 41923 19703
rect 47041 19669 47075 19703
rect 7113 19465 7147 19499
rect 8585 19465 8619 19499
rect 9873 19465 9907 19499
rect 12817 19465 12851 19499
rect 15209 19465 15243 19499
rect 16313 19465 16347 19499
rect 16865 19465 16899 19499
rect 17325 19465 17359 19499
rect 20729 19465 20763 19499
rect 21189 19465 21223 19499
rect 22017 19465 22051 19499
rect 25881 19465 25915 19499
rect 26249 19465 26283 19499
rect 27629 19465 27663 19499
rect 28457 19465 28491 19499
rect 28825 19465 28859 19499
rect 32321 19465 32355 19499
rect 32689 19465 32723 19499
rect 33517 19465 33551 19499
rect 34713 19465 34747 19499
rect 35173 19465 35207 19499
rect 40141 19465 40175 19499
rect 40509 19465 40543 19499
rect 42717 19465 42751 19499
rect 4629 19397 4663 19431
rect 11161 19397 11195 19431
rect 13737 19397 13771 19431
rect 20085 19397 20119 19431
rect 21097 19397 21131 19431
rect 30757 19397 30791 19431
rect 31585 19397 31619 19431
rect 36369 19397 36403 19431
rect 40601 19397 40635 19431
rect 1777 19329 1811 19363
rect 2789 19329 2823 19363
rect 3617 19329 3651 19363
rect 5365 19329 5399 19363
rect 6009 19329 6043 19363
rect 7297 19329 7331 19363
rect 7849 19329 7883 19363
rect 8769 19329 8803 19363
rect 9413 19329 9447 19363
rect 10057 19329 10091 19363
rect 10517 19329 10551 19363
rect 11805 19329 11839 19363
rect 12909 19329 12943 19363
rect 14565 19329 14599 19363
rect 15669 19329 15703 19363
rect 17233 19329 17267 19363
rect 18061 19329 18095 19363
rect 22385 19329 22419 19363
rect 22477 19329 22511 19363
rect 23489 19329 23523 19363
rect 29653 19329 29687 19363
rect 30297 19329 30331 19363
rect 32781 19329 32815 19363
rect 33885 19329 33919 19363
rect 33977 19329 34011 19363
rect 35081 19329 35115 19363
rect 36277 19329 36311 19363
rect 37933 19329 37967 19363
rect 41337 19329 41371 19363
rect 41981 19329 42015 19363
rect 48605 19329 48639 19363
rect 49157 19329 49191 19363
rect 6837 19261 6871 19295
rect 8033 19261 8067 19295
rect 13093 19261 13127 19295
rect 13921 19261 13955 19295
rect 17417 19261 17451 19295
rect 18337 19261 18371 19295
rect 20361 19261 20395 19295
rect 21281 19261 21315 19295
rect 22661 19261 22695 19295
rect 23765 19261 23799 19295
rect 26341 19261 26375 19295
rect 26525 19261 26559 19295
rect 27721 19261 27755 19295
rect 27813 19261 27847 19295
rect 28917 19261 28951 19295
rect 29009 19261 29043 19295
rect 32873 19261 32907 19295
rect 34161 19261 34195 19295
rect 35265 19261 35299 19295
rect 36553 19261 36587 19295
rect 37289 19261 37323 19295
rect 37473 19261 37507 19295
rect 38209 19261 38243 19295
rect 40785 19261 40819 19295
rect 48145 19261 48179 19295
rect 48421 19261 48455 19295
rect 9229 19193 9263 19227
rect 11989 19193 12023 19227
rect 25237 19193 25271 19227
rect 25513 19193 25547 19227
rect 35909 19193 35943 19227
rect 42809 19193 42843 19227
rect 47961 19193 47995 19227
rect 5457 19125 5491 19159
rect 6193 19125 6227 19159
rect 6469 19125 6503 19159
rect 6653 19125 6687 19159
rect 12449 19125 12483 19159
rect 14289 19125 14323 19159
rect 23213 19125 23247 19159
rect 27261 19125 27295 19159
rect 36921 19125 36955 19159
rect 39681 19125 39715 19159
rect 42441 19125 42475 19159
rect 47869 19125 47903 19159
rect 48789 19125 48823 19159
rect 49249 19125 49283 19159
rect 6193 18921 6227 18955
rect 12725 18921 12759 18955
rect 16037 18921 16071 18955
rect 16497 18921 16531 18955
rect 19809 18921 19843 18955
rect 22556 18921 22590 18955
rect 24593 18921 24627 18955
rect 28733 18921 28767 18955
rect 30757 18921 30791 18955
rect 32137 18921 32171 18955
rect 33333 18921 33367 18955
rect 37381 18921 37415 18955
rect 41797 18921 41831 18955
rect 9873 18853 9907 18887
rect 12265 18853 12299 18887
rect 12633 18853 12667 18887
rect 17693 18853 17727 18887
rect 18889 18853 18923 18887
rect 38025 18853 38059 18887
rect 43177 18853 43211 18887
rect 4445 18785 4479 18819
rect 9137 18785 9171 18819
rect 9229 18785 9263 18819
rect 10517 18785 10551 18819
rect 17049 18785 17083 18819
rect 18245 18785 18279 18819
rect 20453 18785 20487 18819
rect 21741 18785 21775 18819
rect 25237 18785 25271 18819
rect 26157 18785 26191 18819
rect 27629 18785 27663 18819
rect 30297 18785 30331 18819
rect 31401 18785 31435 18819
rect 31585 18785 31619 18819
rect 32781 18785 32815 18819
rect 33977 18785 34011 18819
rect 35633 18785 35667 18819
rect 35909 18785 35943 18819
rect 38577 18785 38611 18819
rect 40325 18785 40359 18819
rect 1777 18717 1811 18751
rect 4077 18717 4111 18751
rect 6377 18717 6411 18751
rect 7021 18717 7055 18751
rect 7481 18717 7515 18751
rect 10057 18717 10091 18751
rect 13093 18717 13127 18751
rect 14289 18717 14323 18751
rect 18153 18717 18187 18751
rect 19441 18717 19475 18751
rect 19625 18717 19659 18751
rect 20177 18717 20211 18751
rect 21557 18717 21591 18751
rect 22293 18717 22327 18751
rect 25881 18717 25915 18751
rect 28089 18717 28123 18751
rect 29193 18717 29227 18751
rect 30205 18717 30239 18751
rect 31309 18717 31343 18751
rect 34345 18717 34379 18751
rect 39405 18717 39439 18751
rect 40049 18717 40083 18751
rect 42257 18717 42291 18751
rect 48605 18717 48639 18751
rect 49065 18717 49099 18751
rect 2789 18649 2823 18683
rect 8217 18649 8251 18683
rect 8401 18649 8435 18683
rect 10793 18649 10827 18683
rect 13737 18649 13771 18683
rect 14565 18649 14599 18683
rect 32597 18649 32631 18683
rect 5641 18581 5675 18615
rect 6837 18581 6871 18615
rect 8769 18581 8803 18615
rect 16865 18581 16899 18615
rect 16957 18581 16991 18615
rect 18061 18581 18095 18615
rect 19073 18581 19107 18615
rect 19349 18581 19383 18615
rect 20269 18581 20303 18615
rect 21097 18581 21131 18615
rect 21465 18581 21499 18615
rect 24041 18581 24075 18615
rect 24961 18581 24995 18615
rect 25053 18581 25087 18615
rect 29101 18581 29135 18615
rect 29745 18581 29779 18615
rect 30113 18581 30147 18615
rect 30941 18581 30975 18615
rect 32505 18581 32539 18615
rect 33701 18581 33735 18615
rect 33793 18581 33827 18615
rect 34897 18581 34931 18615
rect 37657 18581 37691 18615
rect 38393 18581 38427 18615
rect 38485 18581 38519 18615
rect 39221 18581 39255 18615
rect 42901 18581 42935 18615
rect 48421 18581 48455 18615
rect 49249 18581 49283 18615
rect 14841 18377 14875 18411
rect 15209 18377 15243 18411
rect 16221 18377 16255 18411
rect 17141 18377 17175 18411
rect 17877 18377 17911 18411
rect 24685 18377 24719 18411
rect 25145 18377 25179 18411
rect 26249 18377 26283 18411
rect 29469 18377 29503 18411
rect 30205 18377 30239 18411
rect 30941 18377 30975 18411
rect 31309 18377 31343 18411
rect 35909 18377 35943 18411
rect 36369 18377 36403 18411
rect 39773 18377 39807 18411
rect 40877 18377 40911 18411
rect 42165 18377 42199 18411
rect 48789 18377 48823 18411
rect 3709 18309 3743 18343
rect 5825 18309 5859 18343
rect 7757 18309 7791 18343
rect 8401 18309 8435 18343
rect 18705 18309 18739 18343
rect 23397 18309 23431 18343
rect 24041 18309 24075 18343
rect 27537 18309 27571 18343
rect 28825 18309 28859 18343
rect 40785 18309 40819 18343
rect 1777 18241 1811 18275
rect 3525 18241 3559 18275
rect 4721 18241 4755 18275
rect 5365 18241 5399 18275
rect 7205 18241 7239 18275
rect 7941 18241 7975 18275
rect 11621 18241 11655 18275
rect 12173 18241 12207 18275
rect 16129 18241 16163 18275
rect 17785 18241 17819 18275
rect 19257 18241 19291 18275
rect 22201 18241 22235 18275
rect 22661 18241 22695 18275
rect 25053 18241 25087 18275
rect 27629 18241 27663 18275
rect 28733 18241 28767 18275
rect 30113 18241 30147 18275
rect 32689 18241 32723 18275
rect 32781 18241 32815 18275
rect 36277 18241 36311 18275
rect 37565 18241 37599 18275
rect 41797 18241 41831 18275
rect 42625 18241 42659 18275
rect 48605 18241 48639 18275
rect 49065 18241 49099 18275
rect 2789 18173 2823 18207
rect 8677 18173 8711 18207
rect 8953 18173 8987 18207
rect 10977 18173 11011 18207
rect 12633 18173 12667 18207
rect 12909 18173 12943 18207
rect 14381 18173 14415 18207
rect 15301 18173 15335 18207
rect 15393 18173 15427 18207
rect 17969 18173 18003 18207
rect 19625 18173 19659 18207
rect 19901 18173 19935 18207
rect 25237 18173 25271 18207
rect 26341 18173 26375 18207
rect 26433 18173 26467 18207
rect 27721 18173 27755 18207
rect 28917 18173 28951 18207
rect 30297 18173 30331 18207
rect 31401 18173 31435 18207
rect 31585 18173 31619 18207
rect 32873 18173 32907 18207
rect 33609 18173 33643 18207
rect 33885 18173 33919 18207
rect 36553 18173 36587 18207
rect 36921 18173 36955 18207
rect 37381 18173 37415 18207
rect 38025 18173 38059 18207
rect 38301 18173 38335 18207
rect 40969 18173 41003 18207
rect 5181 18105 5215 18139
rect 6745 18105 6779 18139
rect 10425 18105 10459 18139
rect 11989 18105 12023 18139
rect 16865 18105 16899 18139
rect 18889 18105 18923 18139
rect 40417 18105 40451 18139
rect 41613 18105 41647 18139
rect 4537 18037 4571 18071
rect 7021 18037 7055 18071
rect 10885 18037 10919 18071
rect 16681 18037 16715 18071
rect 17417 18037 17451 18071
rect 21373 18037 21407 18071
rect 22017 18037 22051 18071
rect 25881 18037 25915 18071
rect 27169 18037 27203 18071
rect 28365 18037 28399 18071
rect 29745 18037 29779 18071
rect 32321 18037 32355 18071
rect 35357 18037 35391 18071
rect 37749 18037 37783 18071
rect 40049 18037 40083 18071
rect 43269 18037 43303 18071
rect 49249 18037 49283 18071
rect 8401 17833 8435 17867
rect 9229 17833 9263 17867
rect 13645 17833 13679 17867
rect 16037 17833 16071 17867
rect 17509 17833 17543 17867
rect 24593 17833 24627 17867
rect 25789 17833 25823 17867
rect 27340 17833 27374 17867
rect 33793 17833 33827 17867
rect 40509 17833 40543 17867
rect 42349 17833 42383 17867
rect 42625 17833 42659 17867
rect 13185 17765 13219 17799
rect 19441 17765 19475 17799
rect 31309 17765 31343 17799
rect 37565 17765 37599 17799
rect 38025 17765 38059 17799
rect 42809 17765 42843 17799
rect 2053 17697 2087 17731
rect 4445 17697 4479 17731
rect 5825 17697 5859 17731
rect 10517 17697 10551 17731
rect 14289 17697 14323 17731
rect 18705 17697 18739 17731
rect 20177 17697 20211 17731
rect 23213 17697 23247 17731
rect 25053 17697 25087 17731
rect 25145 17697 25179 17731
rect 26341 17697 26375 17731
rect 27077 17697 27111 17731
rect 31861 17697 31895 17731
rect 33241 17697 33275 17731
rect 33425 17697 33459 17731
rect 35817 17697 35851 17731
rect 36093 17697 36127 17731
rect 38485 17697 38519 17731
rect 38577 17697 38611 17731
rect 39221 17697 39255 17731
rect 40969 17697 41003 17731
rect 41061 17697 41095 17731
rect 1777 17629 1811 17663
rect 4169 17629 4203 17663
rect 6101 17629 6135 17663
rect 7297 17629 7331 17663
rect 8585 17629 8619 17663
rect 9413 17629 9447 17663
rect 11069 17629 11103 17663
rect 13553 17629 13587 17663
rect 16865 17629 16899 17663
rect 19625 17629 19659 17663
rect 29101 17629 29135 17663
rect 29837 17629 29871 17663
rect 31769 17629 31803 17663
rect 32413 17629 32447 17663
rect 41705 17629 41739 17663
rect 48605 17629 48639 17663
rect 49065 17629 49099 17663
rect 7757 17561 7791 17595
rect 10241 17561 10275 17595
rect 11345 17561 11379 17595
rect 14565 17561 14599 17595
rect 17969 17561 18003 17595
rect 20453 17561 20487 17595
rect 22477 17561 22511 17595
rect 23857 17561 23891 17595
rect 26157 17561 26191 17595
rect 30665 17561 30699 17595
rect 34897 17561 34931 17595
rect 40877 17561 40911 17595
rect 7113 17493 7147 17527
rect 9873 17493 9907 17527
rect 10333 17493 10367 17527
rect 12817 17493 12851 17527
rect 16405 17493 16439 17527
rect 21925 17493 21959 17527
rect 24961 17493 24995 17527
rect 26249 17493 26283 17527
rect 28825 17493 28859 17527
rect 29285 17493 29319 17527
rect 31677 17493 31711 17527
rect 32781 17493 32815 17527
rect 33149 17493 33183 17527
rect 34161 17493 34195 17527
rect 35357 17493 35391 17527
rect 38393 17493 38427 17527
rect 39865 17493 39899 17527
rect 40141 17493 40175 17527
rect 48789 17493 48823 17527
rect 49249 17493 49283 17527
rect 3985 17289 4019 17323
rect 4813 17289 4847 17323
rect 5457 17289 5491 17323
rect 9781 17289 9815 17323
rect 10793 17289 10827 17323
rect 13185 17289 13219 17323
rect 14013 17289 14047 17323
rect 18889 17289 18923 17323
rect 24409 17289 24443 17323
rect 24869 17289 24903 17323
rect 25329 17289 25363 17323
rect 27353 17289 27387 17323
rect 27813 17289 27847 17323
rect 29101 17289 29135 17323
rect 29837 17289 29871 17323
rect 30205 17289 30239 17323
rect 37473 17289 37507 17323
rect 37933 17289 37967 17323
rect 42073 17289 42107 17323
rect 48421 17289 48455 17323
rect 21373 17221 21407 17255
rect 26525 17221 26559 17255
rect 26801 17221 26835 17255
rect 31861 17221 31895 17255
rect 32597 17221 32631 17255
rect 1777 17153 1811 17187
rect 4169 17153 4203 17187
rect 4997 17153 5031 17187
rect 5641 17153 5675 17187
rect 6561 17153 6595 17187
rect 6837 17153 6871 17187
rect 8033 17153 8067 17187
rect 8677 17153 8711 17187
rect 9321 17153 9355 17187
rect 9965 17153 9999 17187
rect 11805 17153 11839 17187
rect 13093 17153 13127 17187
rect 14473 17153 14507 17187
rect 15945 17153 15979 17187
rect 16037 17153 16071 17187
rect 19349 17153 19383 17187
rect 21649 17153 21683 17187
rect 22201 17153 22235 17187
rect 22661 17153 22695 17187
rect 25237 17153 25271 17187
rect 26249 17153 26283 17187
rect 27721 17153 27755 17187
rect 29009 17153 29043 17187
rect 30573 17153 30607 17187
rect 31401 17153 31435 17187
rect 32321 17153 32355 17187
rect 34621 17153 34655 17187
rect 36369 17153 36403 17187
rect 37841 17153 37875 17187
rect 41061 17153 41095 17187
rect 48605 17153 48639 17187
rect 49157 17153 49191 17187
rect 2053 17085 2087 17119
rect 10885 17085 10919 17119
rect 10977 17085 11011 17119
rect 13277 17085 13311 17119
rect 13829 17085 13863 17119
rect 16129 17085 16163 17119
rect 17141 17085 17175 17119
rect 17417 17085 17451 17119
rect 19625 17085 19659 17119
rect 22937 17085 22971 17119
rect 25513 17085 25547 17119
rect 27997 17085 28031 17119
rect 29285 17085 29319 17119
rect 30665 17085 30699 17119
rect 30849 17085 30883 17119
rect 35357 17085 35391 17119
rect 36461 17085 36495 17119
rect 36553 17085 36587 17119
rect 38117 17085 38151 17119
rect 38853 17085 38887 17119
rect 39129 17085 39163 17119
rect 7849 17017 7883 17051
rect 9137 17017 9171 17051
rect 10425 17017 10459 17051
rect 12449 17017 12483 17051
rect 14197 17017 14231 17051
rect 15577 17017 15611 17051
rect 22017 17017 22051 17051
rect 26065 17017 26099 17051
rect 28641 17017 28675 17051
rect 34069 17017 34103 17051
rect 37013 17017 37047 17051
rect 41705 17017 41739 17051
rect 8493 16949 8527 16983
rect 11897 16949 11931 16983
rect 12725 16949 12759 16983
rect 15117 16949 15151 16983
rect 16773 16949 16807 16983
rect 21097 16949 21131 16983
rect 26985 16949 27019 16983
rect 29745 16949 29779 16983
rect 36001 16949 36035 16983
rect 38485 16949 38519 16983
rect 40601 16949 40635 16983
rect 49249 16949 49283 16983
rect 4629 16745 4663 16779
rect 7481 16745 7515 16779
rect 8953 16745 8987 16779
rect 16405 16745 16439 16779
rect 20453 16745 20487 16779
rect 25329 16745 25363 16779
rect 31125 16745 31159 16779
rect 34529 16745 34563 16779
rect 36277 16745 36311 16779
rect 39497 16745 39531 16779
rect 48789 16745 48823 16779
rect 9597 16677 9631 16711
rect 20821 16677 20855 16711
rect 25053 16677 25087 16711
rect 30941 16677 30975 16711
rect 33241 16677 33275 16711
rect 8217 16609 8251 16643
rect 8309 16609 8343 16643
rect 11713 16609 11747 16643
rect 13461 16609 13495 16643
rect 13553 16609 13587 16643
rect 14105 16609 14139 16643
rect 14933 16609 14967 16643
rect 15025 16609 15059 16643
rect 18705 16609 18739 16643
rect 20085 16609 20119 16643
rect 21097 16609 21131 16643
rect 21373 16609 21407 16643
rect 23765 16609 23799 16643
rect 23857 16609 23891 16643
rect 25605 16609 25639 16643
rect 30297 16609 30331 16643
rect 31493 16609 31527 16643
rect 34345 16609 34379 16643
rect 35725 16609 35759 16643
rect 36921 16609 36955 16643
rect 38025 16609 38059 16643
rect 1777 16541 1811 16575
rect 4169 16541 4203 16575
rect 4813 16541 4847 16575
rect 5457 16541 5491 16575
rect 6745 16541 6779 16575
rect 10057 16541 10091 16575
rect 12541 16541 12575 16575
rect 14841 16541 14875 16575
rect 15761 16541 15795 16575
rect 16865 16541 16899 16575
rect 17509 16541 17543 16575
rect 28089 16541 28123 16575
rect 28549 16541 28583 16575
rect 30205 16541 30239 16575
rect 33793 16541 33827 16575
rect 34897 16541 34931 16575
rect 36737 16541 36771 16575
rect 37289 16541 37323 16575
rect 37749 16541 37783 16575
rect 40049 16541 40083 16575
rect 41153 16541 41187 16575
rect 42257 16541 42291 16575
rect 48605 16541 48639 16575
rect 49065 16541 49099 16575
rect 2513 16473 2547 16507
rect 8125 16473 8159 16507
rect 9413 16473 9447 16507
rect 10701 16473 10735 16507
rect 13369 16473 13403 16507
rect 17969 16473 18003 16507
rect 19901 16473 19935 16507
rect 25881 16473 25915 16507
rect 31769 16473 31803 16507
rect 40693 16473 40727 16507
rect 3985 16405 4019 16439
rect 5273 16405 5307 16439
rect 6561 16405 6595 16439
rect 7757 16405 7791 16439
rect 11161 16405 11195 16439
rect 11529 16405 11563 16439
rect 11621 16405 11655 16439
rect 12357 16405 12391 16439
rect 13001 16405 13035 16439
rect 14473 16405 14507 16439
rect 19441 16405 19475 16439
rect 19809 16405 19843 16439
rect 22845 16405 22879 16439
rect 23305 16405 23339 16439
rect 23673 16405 23707 16439
rect 24593 16405 24627 16439
rect 27353 16405 27387 16439
rect 27905 16405 27939 16439
rect 29193 16405 29227 16439
rect 29745 16405 29779 16439
rect 30113 16405 30147 16439
rect 30757 16405 30791 16439
rect 36645 16405 36679 16439
rect 41797 16405 41831 16439
rect 42901 16405 42935 16439
rect 49249 16405 49283 16439
rect 8401 16201 8435 16235
rect 10149 16201 10183 16235
rect 11989 16201 12023 16235
rect 12449 16201 12483 16235
rect 13185 16201 13219 16235
rect 13553 16201 13587 16235
rect 14381 16201 14415 16235
rect 16037 16201 16071 16235
rect 17877 16201 17911 16235
rect 18337 16201 18371 16235
rect 23121 16201 23155 16235
rect 26341 16201 26375 16235
rect 26617 16201 26651 16235
rect 27629 16201 27663 16235
rect 30113 16201 30147 16235
rect 31033 16201 31067 16235
rect 31861 16201 31895 16235
rect 32781 16201 32815 16235
rect 33977 16201 34011 16235
rect 34621 16201 34655 16235
rect 37473 16201 37507 16235
rect 40969 16201 41003 16235
rect 41613 16201 41647 16235
rect 41705 16201 41739 16235
rect 41889 16201 41923 16235
rect 9873 16133 9907 16167
rect 10057 16133 10091 16167
rect 10609 16133 10643 16167
rect 11253 16133 11287 16167
rect 13645 16133 13679 16167
rect 19349 16133 19383 16167
rect 21189 16133 21223 16167
rect 21557 16133 21591 16167
rect 23489 16133 23523 16167
rect 24869 16133 24903 16167
rect 28641 16133 28675 16167
rect 30941 16133 30975 16167
rect 34805 16133 34839 16167
rect 37657 16133 37691 16167
rect 38485 16133 38519 16167
rect 40877 16133 40911 16167
rect 1777 16065 1811 16099
rect 9321 16065 9355 16099
rect 12357 16065 12391 16099
rect 14749 16065 14783 16099
rect 14841 16065 14875 16099
rect 15945 16065 15979 16099
rect 16957 16065 16991 16099
rect 17693 16065 17727 16099
rect 18245 16065 18279 16099
rect 19073 16065 19107 16099
rect 22017 16065 22051 16099
rect 24593 16065 24627 16099
rect 27537 16065 27571 16099
rect 28365 16065 28399 16099
rect 31585 16065 31619 16099
rect 32689 16065 32723 16099
rect 33885 16065 33919 16099
rect 37841 16065 37875 16099
rect 42625 16065 42659 16099
rect 48789 16065 48823 16099
rect 49065 16065 49099 16099
rect 2053 15997 2087 16031
rect 8493 15997 8527 16031
rect 8677 15997 8711 16031
rect 12633 15997 12667 16031
rect 13737 15997 13771 16031
rect 15025 15997 15059 16031
rect 16221 15997 16255 16031
rect 18521 15997 18555 16031
rect 23581 15997 23615 16031
rect 23765 15997 23799 16031
rect 27721 15997 27755 16031
rect 31217 15997 31251 16031
rect 32965 15997 32999 16031
rect 34161 15997 34195 16031
rect 35081 15997 35115 16031
rect 35357 15997 35391 16031
rect 36829 15997 36863 16031
rect 38209 15997 38243 16031
rect 41061 15997 41095 16031
rect 8033 15929 8067 15963
rect 10793 15929 10827 15963
rect 20821 15929 20855 15963
rect 27169 15929 27203 15963
rect 30573 15929 30607 15963
rect 37289 15929 37323 15963
rect 40509 15929 40543 15963
rect 9413 15861 9447 15895
rect 11161 15861 11195 15895
rect 11713 15861 11747 15895
rect 15577 15861 15611 15895
rect 17049 15861 17083 15895
rect 17601 15861 17635 15895
rect 22661 15861 22695 15895
rect 24133 15861 24167 15895
rect 32321 15861 32355 15895
rect 33517 15861 33551 15895
rect 39957 15861 39991 15895
rect 43269 15861 43303 15895
rect 49249 15861 49283 15895
rect 9873 15657 9907 15691
rect 13001 15657 13035 15691
rect 14933 15657 14967 15691
rect 18153 15657 18187 15691
rect 19809 15657 19843 15691
rect 21189 15657 21223 15691
rect 26985 15657 27019 15691
rect 28825 15657 28859 15691
rect 32229 15657 32263 15691
rect 34345 15657 34379 15691
rect 38012 15657 38046 15691
rect 49157 15657 49191 15691
rect 15393 15589 15427 15623
rect 16865 15589 16899 15623
rect 22385 15589 22419 15623
rect 24685 15589 24719 15623
rect 28457 15589 28491 15623
rect 28733 15589 28767 15623
rect 37197 15589 37231 15623
rect 39497 15589 39531 15623
rect 41797 15589 41831 15623
rect 2053 15521 2087 15555
rect 10793 15521 10827 15555
rect 11069 15521 11103 15555
rect 12541 15521 12575 15555
rect 13553 15521 13587 15555
rect 15853 15521 15887 15555
rect 15945 15521 15979 15555
rect 17509 15521 17543 15555
rect 18705 15521 18739 15555
rect 19349 15521 19383 15555
rect 20361 15521 20395 15555
rect 20913 15521 20947 15555
rect 21741 15521 21775 15555
rect 23581 15521 23615 15555
rect 25145 15521 25179 15555
rect 25329 15521 25363 15555
rect 26341 15521 26375 15555
rect 26433 15521 26467 15555
rect 27997 15521 28031 15555
rect 30757 15521 30791 15555
rect 33149 15521 33183 15555
rect 33333 15521 33367 15555
rect 35173 15521 35207 15555
rect 40049 15521 40083 15555
rect 40325 15521 40359 15555
rect 1777 15453 1811 15487
rect 10057 15453 10091 15487
rect 14289 15453 14323 15487
rect 17233 15453 17267 15487
rect 18521 15453 18555 15487
rect 18613 15453 18647 15487
rect 22569 15453 22603 15487
rect 23489 15453 23523 15487
rect 27905 15453 27939 15487
rect 29285 15453 29319 15487
rect 30481 15453 30515 15487
rect 33885 15453 33919 15487
rect 34897 15453 34931 15487
rect 37289 15453 37323 15487
rect 37749 15453 37783 15487
rect 42257 15453 42291 15487
rect 48881 15453 48915 15487
rect 49341 15453 49375 15487
rect 6561 15385 6595 15419
rect 9413 15385 9447 15419
rect 13369 15385 13403 15419
rect 15761 15385 15795 15419
rect 19441 15385 19475 15419
rect 20269 15385 20303 15419
rect 23397 15385 23431 15419
rect 27813 15385 27847 15419
rect 29009 15385 29043 15419
rect 42901 15385 42935 15419
rect 6653 15317 6687 15351
rect 8677 15317 8711 15351
rect 9045 15317 9079 15351
rect 9505 15317 9539 15351
rect 10517 15317 10551 15351
rect 13461 15317 13495 15351
rect 16589 15317 16623 15351
rect 17325 15317 17359 15351
rect 20177 15317 20211 15351
rect 21557 15317 21591 15351
rect 21649 15317 21683 15351
rect 23029 15317 23063 15351
rect 25053 15317 25087 15351
rect 25881 15317 25915 15351
rect 26249 15317 26283 15351
rect 27077 15317 27111 15351
rect 27445 15317 27479 15351
rect 29837 15317 29871 15351
rect 32689 15317 32723 15351
rect 33057 15317 33091 15351
rect 36645 15317 36679 15351
rect 36921 15317 36955 15351
rect 9873 15113 9907 15147
rect 11805 15113 11839 15147
rect 12265 15113 12299 15147
rect 15117 15113 15151 15147
rect 16865 15113 16899 15147
rect 18061 15113 18095 15147
rect 18705 15113 18739 15147
rect 19533 15113 19567 15147
rect 20729 15113 20763 15147
rect 21925 15113 21959 15147
rect 22937 15113 22971 15147
rect 24133 15113 24167 15147
rect 27077 15113 27111 15147
rect 27353 15113 27387 15147
rect 27629 15113 27663 15147
rect 32321 15113 32355 15147
rect 33885 15113 33919 15147
rect 35081 15113 35115 15147
rect 36277 15113 36311 15147
rect 39681 15113 39715 15147
rect 41521 15113 41555 15147
rect 41797 15113 41831 15147
rect 41981 15113 42015 15147
rect 9965 15045 9999 15079
rect 17233 15045 17267 15079
rect 17325 15045 17359 15079
rect 26341 15045 26375 15079
rect 31585 15045 31619 15079
rect 32781 15045 32815 15079
rect 40049 15045 40083 15079
rect 1777 14977 1811 15011
rect 9229 14977 9263 15011
rect 10977 14977 11011 15011
rect 12173 14977 12207 15011
rect 13001 14977 13035 15011
rect 15669 14977 15703 15011
rect 19901 14977 19935 15011
rect 21097 14977 21131 15011
rect 22293 14977 22327 15011
rect 23305 14977 23339 15011
rect 24501 14977 24535 15011
rect 25145 14977 25179 15011
rect 26249 14977 26283 15011
rect 27261 14977 27295 15011
rect 28089 14977 28123 15011
rect 30665 14977 30699 15011
rect 32689 14977 32723 15011
rect 40141 14977 40175 15011
rect 40877 14977 40911 15011
rect 42809 14977 42843 15011
rect 48789 14977 48823 15011
rect 49065 14977 49099 15011
rect 2053 14909 2087 14943
rect 10057 14909 10091 14943
rect 12357 14909 12391 14943
rect 13277 14909 13311 14943
rect 17417 14909 17451 14943
rect 18797 14909 18831 14943
rect 18889 14909 18923 14943
rect 19993 14909 20027 14943
rect 20085 14909 20119 14943
rect 21189 14909 21223 14943
rect 21281 14909 21315 14943
rect 23397 14909 23431 14943
rect 23581 14909 23615 14943
rect 24593 14909 24627 14943
rect 24685 14909 24719 14943
rect 26433 14909 26467 14943
rect 28365 14909 28399 14943
rect 29837 14909 29871 14943
rect 30757 14909 30791 14943
rect 30849 14909 30883 14943
rect 32965 14909 32999 14943
rect 33977 14909 34011 14943
rect 34161 14909 34195 14943
rect 35173 14909 35207 14943
rect 35357 14909 35391 14943
rect 36369 14909 36403 14943
rect 36553 14909 36587 14943
rect 37473 14909 37507 14943
rect 37749 14909 37783 14943
rect 40233 14909 40267 14943
rect 14749 14841 14783 14875
rect 18337 14841 18371 14875
rect 27721 14841 27755 14875
rect 34713 14841 34747 14875
rect 35909 14841 35943 14875
rect 49249 14841 49283 14875
rect 9505 14773 9539 14807
rect 10609 14773 10643 14807
rect 11069 14773 11103 14807
rect 15301 14773 15335 14807
rect 16313 14773 16347 14807
rect 25329 14773 25363 14807
rect 25513 14773 25547 14807
rect 25881 14773 25915 14807
rect 30297 14773 30331 14807
rect 33517 14773 33551 14807
rect 36921 14773 36955 14807
rect 39221 14773 39255 14807
rect 42625 14773 42659 14807
rect 10425 14569 10459 14603
rect 14197 14569 14231 14603
rect 23765 14569 23799 14603
rect 24225 14569 24259 14603
rect 25960 14569 25994 14603
rect 29745 14569 29779 14603
rect 30941 14569 30975 14603
rect 42073 14569 42107 14603
rect 11805 14501 11839 14535
rect 18153 14501 18187 14535
rect 19625 14501 19659 14535
rect 27905 14501 27939 14535
rect 32137 14501 32171 14535
rect 33333 14501 33367 14535
rect 36645 14501 36679 14535
rect 2053 14433 2087 14467
rect 9045 14433 9079 14467
rect 12449 14433 12483 14467
rect 13461 14433 13495 14467
rect 13553 14433 13587 14467
rect 15117 14433 15151 14467
rect 16221 14433 16255 14467
rect 17417 14433 17451 14467
rect 18613 14433 18647 14467
rect 18705 14433 18739 14467
rect 20177 14433 20211 14467
rect 21097 14433 21131 14467
rect 23121 14433 23155 14467
rect 25697 14433 25731 14467
rect 28365 14433 28399 14467
rect 28549 14433 28583 14467
rect 29101 14433 29135 14467
rect 30297 14433 30331 14467
rect 31585 14433 31619 14467
rect 32781 14433 32815 14467
rect 33793 14433 33827 14467
rect 33977 14433 34011 14467
rect 34897 14433 34931 14467
rect 37105 14433 37139 14467
rect 1777 14365 1811 14399
rect 9781 14365 9815 14399
rect 12173 14365 12207 14399
rect 17233 14365 17267 14399
rect 23949 14365 23983 14399
rect 24593 14365 24627 14399
rect 31309 14365 31343 14399
rect 32597 14365 32631 14399
rect 33701 14365 33735 14399
rect 39497 14365 39531 14399
rect 40049 14365 40083 14399
rect 41153 14365 41187 14399
rect 48605 14365 48639 14399
rect 49065 14365 49099 14399
rect 9597 14297 9631 14331
rect 10333 14297 10367 14331
rect 11161 14297 11195 14331
rect 12265 14297 12299 14331
rect 13369 14297 13403 14331
rect 14841 14297 14875 14331
rect 21373 14297 21407 14331
rect 23397 14297 23431 14331
rect 28273 14297 28307 14331
rect 31401 14297 31435 14331
rect 34345 14297 34379 14331
rect 35173 14297 35207 14331
rect 37381 14297 37415 14331
rect 41797 14297 41831 14331
rect 9229 14229 9263 14263
rect 11253 14229 11287 14263
rect 13001 14229 13035 14263
rect 14473 14229 14507 14263
rect 14933 14229 14967 14263
rect 15669 14229 15703 14263
rect 16037 14229 16071 14263
rect 16129 14229 16163 14263
rect 16865 14229 16899 14263
rect 17325 14229 17359 14263
rect 18521 14229 18555 14263
rect 19349 14229 19383 14263
rect 19993 14229 20027 14263
rect 20085 14229 20119 14263
rect 20729 14229 20763 14263
rect 23673 14229 23707 14263
rect 25237 14229 25271 14263
rect 27445 14229 27479 14263
rect 28917 14229 28951 14263
rect 29285 14229 29319 14263
rect 30113 14229 30147 14263
rect 30205 14229 30239 14263
rect 32505 14229 32539 14263
rect 38853 14229 38887 14263
rect 39313 14229 39347 14263
rect 40693 14229 40727 14263
rect 48697 14229 48731 14263
rect 49249 14229 49283 14263
rect 3617 14025 3651 14059
rect 9873 14025 9907 14059
rect 11161 14025 11195 14059
rect 11621 14025 11655 14059
rect 15117 14025 15151 14059
rect 16313 14025 16347 14059
rect 17877 14025 17911 14059
rect 18245 14025 18279 14059
rect 21465 14025 21499 14059
rect 26617 14025 26651 14059
rect 31585 14025 31619 14059
rect 34897 14025 34931 14059
rect 35725 14025 35759 14059
rect 36093 14025 36127 14059
rect 36829 14025 36863 14059
rect 37473 14025 37507 14059
rect 37841 14025 37875 14059
rect 38669 14025 38703 14059
rect 40509 14025 40543 14059
rect 41337 14025 41371 14059
rect 41797 14025 41831 14059
rect 45661 14025 45695 14059
rect 48421 14025 48455 14059
rect 49249 14025 49283 14059
rect 18337 13957 18371 13991
rect 22293 13957 22327 13991
rect 24225 13957 24259 13991
rect 27169 13957 27203 13991
rect 34989 13957 35023 13991
rect 36185 13957 36219 13991
rect 45017 13957 45051 13991
rect 48145 13957 48179 13991
rect 49157 13957 49191 13991
rect 1777 13889 1811 13923
rect 3525 13889 3559 13923
rect 3985 13889 4019 13923
rect 10517 13889 10551 13923
rect 12357 13889 12391 13923
rect 15669 13889 15703 13923
rect 16773 13889 16807 13923
rect 17417 13889 17451 13923
rect 22017 13889 22051 13923
rect 24869 13889 24903 13923
rect 28917 13889 28951 13923
rect 39037 13889 39071 13923
rect 39865 13889 39899 13923
rect 40877 13889 40911 13923
rect 40969 13889 41003 13923
rect 41521 13889 41555 13923
rect 45845 13889 45879 13923
rect 48605 13889 48639 13923
rect 2053 13821 2087 13855
rect 9597 13821 9631 13855
rect 12449 13821 12483 13855
rect 12541 13821 12575 13855
rect 13001 13821 13035 13855
rect 13369 13821 13403 13855
rect 18429 13821 18463 13855
rect 19073 13821 19107 13855
rect 19717 13821 19751 13855
rect 23765 13821 23799 13855
rect 25145 13821 25179 13855
rect 29377 13821 29411 13855
rect 29653 13821 29687 13855
rect 31125 13821 31159 13855
rect 32321 13821 32355 13855
rect 32597 13821 32631 13855
rect 34069 13821 34103 13855
rect 35081 13821 35115 13855
rect 36277 13821 36311 13855
rect 37933 13821 37967 13855
rect 38117 13821 38151 13855
rect 39129 13821 39163 13855
rect 39313 13821 39347 13855
rect 45201 13821 45235 13855
rect 17233 13753 17267 13787
rect 11989 13685 12023 13719
rect 13632 13685 13666 13719
rect 16957 13685 16991 13719
rect 19974 13685 20008 13719
rect 34529 13685 34563 13719
rect 36921 13685 36955 13719
rect 9597 13481 9631 13515
rect 11148 13481 11182 13515
rect 13093 13481 13127 13515
rect 14473 13481 14507 13515
rect 15209 13481 15243 13515
rect 16405 13481 16439 13515
rect 18705 13481 18739 13515
rect 19533 13481 19567 13515
rect 20729 13481 20763 13515
rect 21925 13481 21959 13515
rect 24133 13481 24167 13515
rect 24869 13481 24903 13515
rect 26709 13481 26743 13515
rect 29009 13481 29043 13515
rect 29377 13481 29411 13515
rect 38209 13481 38243 13515
rect 13277 13413 13311 13447
rect 18889 13413 18923 13447
rect 23121 13413 23155 13447
rect 36185 13413 36219 13447
rect 2789 13345 2823 13379
rect 9781 13345 9815 13379
rect 12633 13345 12667 13379
rect 15669 13345 15703 13379
rect 15853 13345 15887 13379
rect 16865 13345 16899 13379
rect 17049 13345 17083 13379
rect 18245 13345 18279 13379
rect 20085 13345 20119 13379
rect 21373 13345 21407 13379
rect 22385 13345 22419 13379
rect 22569 13345 22603 13379
rect 23765 13345 23799 13379
rect 25421 13345 25455 13379
rect 30297 13345 30331 13379
rect 31217 13345 31251 13379
rect 33977 13345 34011 13379
rect 34069 13345 34103 13379
rect 36737 13345 36771 13379
rect 1777 13277 1811 13311
rect 10885 13277 10919 13311
rect 15577 13277 15611 13311
rect 17969 13277 18003 13311
rect 18061 13277 18095 13311
rect 19901 13277 19935 13311
rect 21097 13277 21131 13311
rect 25237 13277 25271 13311
rect 26065 13277 26099 13311
rect 27169 13277 27203 13311
rect 28365 13277 28399 13311
rect 30113 13277 30147 13311
rect 33885 13277 33919 13311
rect 34897 13277 34931 13311
rect 35725 13277 35759 13311
rect 36461 13277 36495 13311
rect 38669 13277 38703 13311
rect 40049 13277 40083 13311
rect 41153 13277 41187 13311
rect 47961 13277 47995 13311
rect 49157 13277 49191 13311
rect 9965 13209 9999 13243
rect 13553 13209 13587 13243
rect 14381 13209 14415 13243
rect 16773 13209 16807 13243
rect 18981 13209 19015 13243
rect 19993 13209 20027 13243
rect 23581 13209 23615 13243
rect 31493 13209 31527 13243
rect 40693 13209 40727 13243
rect 10241 13141 10275 13175
rect 14841 13141 14875 13175
rect 17601 13141 17635 13175
rect 21189 13141 21223 13175
rect 22293 13141 22327 13175
rect 23489 13141 23523 13175
rect 24501 13141 24535 13175
rect 25329 13141 25363 13175
rect 27813 13141 27847 13175
rect 29745 13141 29779 13175
rect 30205 13141 30239 13175
rect 30757 13141 30791 13175
rect 32965 13141 32999 13175
rect 33517 13141 33551 13175
rect 39313 13141 39347 13175
rect 39589 13141 39623 13175
rect 41797 13141 41831 13175
rect 2881 12937 2915 12971
rect 9873 12937 9907 12971
rect 10885 12937 10919 12971
rect 12081 12937 12115 12971
rect 14841 12937 14875 12971
rect 15945 12937 15979 12971
rect 21097 12937 21131 12971
rect 22753 12937 22787 12971
rect 25697 12937 25731 12971
rect 36921 12937 36955 12971
rect 17141 12869 17175 12903
rect 23121 12869 23155 12903
rect 24225 12869 24259 12903
rect 26801 12869 26835 12903
rect 27445 12869 27479 12903
rect 29653 12869 29687 12903
rect 30389 12869 30423 12903
rect 32597 12869 32631 12903
rect 34529 12869 34563 12903
rect 36369 12869 36403 12903
rect 37749 12869 37783 12903
rect 41153 12869 41187 12903
rect 41889 12869 41923 12903
rect 3065 12801 3099 12835
rect 3341 12801 3375 12835
rect 10793 12801 10827 12835
rect 12173 12801 12207 12835
rect 13093 12801 13127 12835
rect 16037 12801 16071 12835
rect 16865 12801 16899 12835
rect 19533 12801 19567 12835
rect 21005 12801 21039 12835
rect 23213 12801 23247 12835
rect 23949 12801 23983 12835
rect 27169 12801 27203 12835
rect 31401 12801 31435 12835
rect 32321 12801 32355 12835
rect 36277 12801 36311 12835
rect 37473 12801 37507 12835
rect 39957 12801 39991 12835
rect 41613 12801 41647 12835
rect 46213 12801 46247 12835
rect 47961 12801 47995 12835
rect 49157 12801 49191 12835
rect 1593 12733 1627 12767
rect 1869 12733 1903 12767
rect 10977 12733 11011 12767
rect 12357 12733 12391 12767
rect 13369 12733 13403 12767
rect 15209 12733 15243 12767
rect 16221 12733 16255 12767
rect 18613 12733 18647 12767
rect 19625 12733 19659 12767
rect 19809 12733 19843 12767
rect 21189 12733 21223 12767
rect 22017 12733 22051 12767
rect 23305 12733 23339 12767
rect 26157 12733 26191 12767
rect 29193 12733 29227 12767
rect 31493 12733 31527 12767
rect 31677 12733 31711 12767
rect 35265 12733 35299 12767
rect 36461 12733 36495 12767
rect 39497 12733 39531 12767
rect 10149 12665 10183 12699
rect 19165 12665 19199 12699
rect 20637 12665 20671 12699
rect 34069 12665 34103 12699
rect 41337 12665 41371 12699
rect 10425 12597 10459 12631
rect 11713 12597 11747 12631
rect 12817 12597 12851 12631
rect 15577 12597 15611 12631
rect 20269 12597 20303 12631
rect 31033 12597 31067 12631
rect 35909 12597 35943 12631
rect 40601 12597 40635 12631
rect 46029 12597 46063 12631
rect 2789 12393 2823 12427
rect 16773 12393 16807 12427
rect 23305 12393 23339 12427
rect 31769 12393 31803 12427
rect 33977 12393 34011 12427
rect 36645 12393 36679 12427
rect 37105 12393 37139 12427
rect 39221 12393 39255 12427
rect 39405 12393 39439 12427
rect 39589 12393 39623 12427
rect 20913 12325 20947 12359
rect 26341 12325 26375 12359
rect 34253 12325 34287 12359
rect 41429 12325 41463 12359
rect 1869 12257 1903 12291
rect 10977 12257 11011 12291
rect 13461 12257 13495 12291
rect 13645 12257 13679 12291
rect 14657 12257 14691 12291
rect 17417 12257 17451 12291
rect 20177 12257 20211 12291
rect 21465 12257 21499 12291
rect 22753 12257 22787 12291
rect 23949 12257 23983 12291
rect 24869 12257 24903 12291
rect 27537 12257 27571 12291
rect 29009 12257 29043 12291
rect 30021 12257 30055 12291
rect 32229 12257 32263 12291
rect 32505 12257 32539 12291
rect 34529 12257 34563 12291
rect 34897 12257 34931 12291
rect 37565 12257 37599 12291
rect 37749 12257 37783 12291
rect 49157 12257 49191 12291
rect 1593 12189 1627 12223
rect 9597 12189 9631 12223
rect 10701 12189 10735 12223
rect 14381 12189 14415 12223
rect 17969 12189 18003 12223
rect 21281 12189 21315 12223
rect 23673 12189 23707 12223
rect 24593 12189 24627 12223
rect 26709 12189 26743 12223
rect 28917 12189 28951 12223
rect 29745 12189 29779 12223
rect 37473 12189 37507 12223
rect 38301 12189 38335 12223
rect 40969 12189 41003 12223
rect 41613 12189 41647 12223
rect 46121 12189 46155 12223
rect 47961 12189 47995 12223
rect 2881 12121 2915 12155
rect 13369 12121 13403 12155
rect 18705 12121 18739 12155
rect 19441 12121 19475 12155
rect 35173 12121 35207 12155
rect 40141 12121 40175 12155
rect 40325 12121 40359 12155
rect 9229 12053 9263 12087
rect 10241 12053 10275 12087
rect 12449 12053 12483 12087
rect 13001 12053 13035 12087
rect 16129 12053 16163 12087
rect 17141 12053 17175 12087
rect 17233 12053 17267 12087
rect 21373 12053 21407 12087
rect 22109 12053 22143 12087
rect 22477 12053 22511 12087
rect 22569 12053 22603 12087
rect 23765 12053 23799 12087
rect 26985 12053 27019 12087
rect 27353 12053 27387 12087
rect 27445 12053 27479 12087
rect 28089 12053 28123 12087
rect 28457 12053 28491 12087
rect 28825 12053 28859 12087
rect 31493 12053 31527 12087
rect 38945 12053 38979 12087
rect 40785 12053 40819 12087
rect 45937 12053 45971 12087
rect 2329 11849 2363 11883
rect 9965 11849 9999 11883
rect 10149 11849 10183 11883
rect 15577 11849 15611 11883
rect 16497 11849 16531 11883
rect 19073 11849 19107 11883
rect 19901 11849 19935 11883
rect 20729 11849 20763 11883
rect 21097 11849 21131 11883
rect 22293 11849 22327 11883
rect 25697 11849 25731 11883
rect 25973 11849 26007 11883
rect 26433 11849 26467 11883
rect 31217 11849 31251 11883
rect 31309 11849 31343 11883
rect 32321 11849 32355 11883
rect 37841 11849 37875 11883
rect 38669 11849 38703 11883
rect 18981 11781 19015 11815
rect 22109 11781 22143 11815
rect 23397 11781 23431 11815
rect 33885 11781 33919 11815
rect 34621 11781 34655 11815
rect 37933 11781 37967 11815
rect 45109 11781 45143 11815
rect 49157 11781 49191 11815
rect 1593 11713 1627 11747
rect 2513 11713 2547 11747
rect 10517 11713 10551 11747
rect 12357 11713 12391 11747
rect 14381 11713 14415 11747
rect 15485 11713 15519 11747
rect 16865 11713 16899 11747
rect 19809 11713 19843 11747
rect 21925 11713 21959 11747
rect 22569 11713 22603 11747
rect 23949 11713 23983 11747
rect 27537 11713 27571 11747
rect 28181 11713 28215 11747
rect 28549 11713 28583 11747
rect 32689 11713 32723 11747
rect 39037 11713 39071 11747
rect 39865 11713 39899 11747
rect 47961 11713 47995 11747
rect 2789 11645 2823 11679
rect 11713 11645 11747 11679
rect 12633 11645 12667 11679
rect 15669 11645 15703 11679
rect 17141 11645 17175 11679
rect 19993 11645 20027 11679
rect 21189 11645 21223 11679
rect 21373 11645 21407 11679
rect 24225 11645 24259 11679
rect 27629 11645 27663 11679
rect 27813 11645 27847 11679
rect 28825 11645 28859 11679
rect 31401 11645 31435 11679
rect 32781 11645 32815 11679
rect 32873 11645 32907 11679
rect 33977 11645 34011 11679
rect 34161 11645 34195 11679
rect 35173 11645 35207 11679
rect 35449 11645 35483 11679
rect 36921 11645 36955 11679
rect 38117 11645 38151 11679
rect 39129 11645 39163 11679
rect 39221 11645 39255 11679
rect 40785 11645 40819 11679
rect 1777 11577 1811 11611
rect 27169 11577 27203 11611
rect 30297 11577 30331 11611
rect 33517 11577 33551 11611
rect 37473 11577 37507 11611
rect 45293 11577 45327 11611
rect 11161 11509 11195 11543
rect 14841 11509 14875 11543
rect 15117 11509 15151 11543
rect 16221 11509 16255 11543
rect 18613 11509 18647 11543
rect 19441 11509 19475 11543
rect 30849 11509 30883 11543
rect 31953 11509 31987 11543
rect 34805 11509 34839 11543
rect 40509 11509 40543 11543
rect 2145 11305 2179 11339
rect 10425 11305 10459 11339
rect 10885 11305 10919 11339
rect 14565 11305 14599 11339
rect 16957 11305 16991 11339
rect 18153 11305 18187 11339
rect 19441 11305 19475 11339
rect 20624 11305 20658 11339
rect 23305 11305 23339 11339
rect 26341 11305 26375 11339
rect 29009 11305 29043 11339
rect 34713 11305 34747 11339
rect 40233 11305 40267 11339
rect 1777 11237 1811 11271
rect 13921 11237 13955 11271
rect 28641 11237 28675 11271
rect 33517 11237 33551 11271
rect 38853 11237 38887 11271
rect 41521 11237 41555 11271
rect 11161 11169 11195 11203
rect 11437 11169 11471 11203
rect 13369 11169 13403 11203
rect 15025 11169 15059 11203
rect 15117 11169 15151 11203
rect 16221 11169 16255 11203
rect 16313 11169 16347 11203
rect 17601 11169 17635 11203
rect 18613 11169 18647 11203
rect 18797 11169 18831 11203
rect 20361 11169 20395 11203
rect 22569 11169 22603 11203
rect 23949 11169 23983 11203
rect 24593 11169 24627 11203
rect 27169 11169 27203 11203
rect 31401 11169 31435 11203
rect 32873 11169 32907 11203
rect 34069 11169 34103 11203
rect 49157 11169 49191 11203
rect 1593 11101 1627 11135
rect 2329 11101 2363 11135
rect 17325 11101 17359 11135
rect 18521 11101 18555 11135
rect 23673 11101 23707 11135
rect 26893 11101 26927 11135
rect 31125 11101 31159 11135
rect 33977 11101 34011 11135
rect 35725 11101 35759 11135
rect 38209 11101 38243 11135
rect 39497 11101 39531 11135
rect 41705 11101 41739 11135
rect 45661 11101 45695 11135
rect 47961 11101 47995 11135
rect 10609 11033 10643 11067
rect 14289 11033 14323 11067
rect 16129 11033 16163 11067
rect 17417 11033 17451 11067
rect 19717 11033 19751 11067
rect 23765 11033 23799 11067
rect 24869 11033 24903 11067
rect 29745 11033 29779 11067
rect 30481 11033 30515 11067
rect 33885 11033 33919 11067
rect 35265 11033 35299 11067
rect 36001 11033 36035 11067
rect 37749 11033 37783 11067
rect 40141 11033 40175 11067
rect 40877 11033 40911 11067
rect 41061 11033 41095 11067
rect 45845 11033 45879 11067
rect 12909 10965 12943 10999
rect 14933 10965 14967 10999
rect 15761 10965 15795 10999
rect 22109 10965 22143 10999
rect 29101 10965 29135 10999
rect 29285 10965 29319 10999
rect 33241 10965 33275 10999
rect 34989 10965 35023 10999
rect 35173 10965 35207 10999
rect 39313 10965 39347 10999
rect 12357 10761 12391 10795
rect 13645 10761 13679 10795
rect 14841 10761 14875 10795
rect 15577 10761 15611 10795
rect 17417 10761 17451 10795
rect 18061 10761 18095 10795
rect 18797 10761 18831 10795
rect 19533 10761 19567 10795
rect 20729 10761 20763 10795
rect 21097 10761 21131 10795
rect 21189 10761 21223 10795
rect 23765 10761 23799 10795
rect 25329 10761 25363 10795
rect 25513 10761 25547 10795
rect 25697 10761 25731 10795
rect 27169 10761 27203 10795
rect 31401 10761 31435 10795
rect 32781 10761 32815 10795
rect 33333 10761 33367 10795
rect 39221 10761 39255 10795
rect 40233 10761 40267 10795
rect 40693 10761 40727 10795
rect 19993 10693 20027 10727
rect 24685 10693 24719 10727
rect 28825 10693 28859 10727
rect 32689 10693 32723 10727
rect 34069 10693 34103 10727
rect 36553 10693 36587 10727
rect 49157 10693 49191 10727
rect 1593 10625 1627 10659
rect 2329 10625 2363 10659
rect 2881 10625 2915 10659
rect 11621 10625 11655 10659
rect 13553 10625 13587 10659
rect 14749 10625 14783 10659
rect 15945 10625 15979 10659
rect 17325 10625 17359 10659
rect 18705 10625 18739 10659
rect 19901 10625 19935 10659
rect 24593 10625 24627 10659
rect 25973 10625 26007 10659
rect 27537 10625 27571 10659
rect 28733 10625 28767 10659
rect 29837 10625 29871 10659
rect 31309 10625 31343 10659
rect 36461 10625 36495 10659
rect 37473 10625 37507 10659
rect 38577 10625 38611 10659
rect 39773 10625 39807 10659
rect 47961 10625 47995 10659
rect 3065 10557 3099 10591
rect 12449 10557 12483 10591
rect 12541 10557 12575 10591
rect 13829 10557 13863 10591
rect 15025 10557 15059 10591
rect 16037 10557 16071 10591
rect 16221 10557 16255 10591
rect 17601 10557 17635 10591
rect 18889 10557 18923 10591
rect 20177 10557 20211 10591
rect 21373 10557 21407 10591
rect 22017 10557 22051 10591
rect 22293 10557 22327 10591
rect 24869 10557 24903 10591
rect 27629 10557 27663 10591
rect 27813 10557 27847 10591
rect 28917 10557 28951 10591
rect 30481 10557 30515 10591
rect 31585 10557 31619 10591
rect 32873 10557 32907 10591
rect 33793 10557 33827 10591
rect 36737 10557 36771 10591
rect 39957 10557 39991 10591
rect 1777 10489 1811 10523
rect 13185 10489 13219 10523
rect 16957 10489 16991 10523
rect 24225 10489 24259 10523
rect 30941 10489 30975 10523
rect 35541 10489 35575 10523
rect 36093 10489 36127 10523
rect 2513 10421 2547 10455
rect 11253 10421 11287 10455
rect 11989 10421 12023 10455
rect 14381 10421 14415 10455
rect 18337 10421 18371 10455
rect 26617 10421 26651 10455
rect 28365 10421 28399 10455
rect 29469 10421 29503 10455
rect 32321 10421 32355 10455
rect 38117 10421 38151 10455
rect 12541 10217 12575 10251
rect 13001 10217 13035 10251
rect 18521 10217 18555 10251
rect 19349 10217 19383 10251
rect 24856 10217 24890 10251
rect 26709 10217 26743 10251
rect 29377 10217 29411 10251
rect 32137 10217 32171 10251
rect 36645 10217 36679 10251
rect 19073 10149 19107 10183
rect 22109 10149 22143 10183
rect 28733 10149 28767 10183
rect 33333 10149 33367 10183
rect 38485 10149 38519 10183
rect 1869 10081 1903 10115
rect 13553 10081 13587 10115
rect 14289 10081 14323 10115
rect 14565 10081 14599 10115
rect 17049 10081 17083 10115
rect 19625 10081 19659 10115
rect 20361 10081 20395 10115
rect 23305 10081 23339 10115
rect 24593 10081 24627 10115
rect 27261 10081 27295 10115
rect 29745 10081 29779 10115
rect 33977 10081 34011 10115
rect 34437 10081 34471 10115
rect 35173 10081 35207 10115
rect 37749 10081 37783 10115
rect 39497 10081 39531 10115
rect 40325 10081 40359 10115
rect 49157 10081 49191 10115
rect 1593 10013 1627 10047
rect 11897 10013 11931 10047
rect 16773 10013 16807 10047
rect 18797 10013 18831 10047
rect 26985 10013 27019 10047
rect 29101 10013 29135 10047
rect 30389 10013 30423 10047
rect 32597 10013 32631 10047
rect 33701 10013 33735 10047
rect 34897 10013 34931 10047
rect 37105 10013 37139 10047
rect 46121 10013 46155 10047
rect 47961 10013 47995 10047
rect 16313 9945 16347 9979
rect 20624 9945 20658 9979
rect 22569 9945 22603 9979
rect 30665 9945 30699 9979
rect 38301 9945 38335 9979
rect 38761 9945 38795 9979
rect 40141 9945 40175 9979
rect 40601 9945 40635 9979
rect 44373 9945 44407 9979
rect 44557 9945 44591 9979
rect 47317 9945 47351 9979
rect 13369 9877 13403 9911
rect 13461 9877 13495 9911
rect 23857 9877 23891 9911
rect 24041 9877 24075 9911
rect 26341 9877 26375 9911
rect 33793 9877 33827 9911
rect 2145 9673 2179 9707
rect 15393 9673 15427 9707
rect 22017 9673 22051 9707
rect 35633 9673 35667 9707
rect 37289 9673 37323 9707
rect 12817 9605 12851 9639
rect 15853 9605 15887 9639
rect 16129 9605 16163 9639
rect 23121 9605 23155 9639
rect 26249 9605 26283 9639
rect 32965 9605 32999 9639
rect 34161 9605 34195 9639
rect 37105 9605 37139 9639
rect 37841 9605 37875 9639
rect 49157 9605 49191 9639
rect 1685 9537 1719 9571
rect 2329 9537 2363 9571
rect 12909 9537 12943 9571
rect 22385 9537 22419 9571
rect 23581 9537 23615 9571
rect 26157 9537 26191 9571
rect 31861 9537 31895 9571
rect 32321 9537 32355 9571
rect 33057 9537 33091 9571
rect 36093 9537 36127 9571
rect 47961 9537 47995 9571
rect 1869 9469 1903 9503
rect 13093 9469 13127 9503
rect 13645 9469 13679 9503
rect 13921 9469 13955 9503
rect 16865 9469 16899 9503
rect 17141 9469 17175 9503
rect 18889 9469 18923 9503
rect 19349 9469 19383 9503
rect 19625 9469 19659 9503
rect 22477 9469 22511 9503
rect 22661 9469 22695 9503
rect 23857 9469 23891 9503
rect 26433 9469 26467 9503
rect 27537 9469 27571 9503
rect 27813 9469 27847 9503
rect 29745 9469 29779 9503
rect 30021 9469 30055 9503
rect 33149 9469 33183 9503
rect 33885 9469 33919 9503
rect 12449 9401 12483 9435
rect 21465 9401 21499 9435
rect 25789 9401 25823 9435
rect 12081 9333 12115 9367
rect 21097 9333 21131 9367
rect 21649 9333 21683 9367
rect 25329 9333 25363 9367
rect 27077 9333 27111 9367
rect 27261 9333 27295 9367
rect 29285 9333 29319 9367
rect 31493 9333 31527 9367
rect 32597 9333 32631 9367
rect 36737 9333 36771 9367
rect 13001 9129 13035 9163
rect 18889 9129 18923 9163
rect 21649 9129 21683 9163
rect 23121 9129 23155 9163
rect 25973 9129 26007 9163
rect 27721 9129 27755 9163
rect 28181 9129 28215 9163
rect 32505 9129 32539 9163
rect 32965 9129 32999 9163
rect 34897 9129 34931 9163
rect 21189 9061 21223 9095
rect 36645 9061 36679 9095
rect 13461 8993 13495 9027
rect 13645 8993 13679 9027
rect 22201 8993 22235 9027
rect 23765 8993 23799 9027
rect 24133 8993 24167 9027
rect 24685 8993 24719 9027
rect 26433 8993 26467 9027
rect 28825 8993 28859 9027
rect 29745 8993 29779 9027
rect 31033 8993 31067 9027
rect 33609 8993 33643 9027
rect 34069 8993 34103 9027
rect 35357 8993 35391 9027
rect 35449 8993 35483 9027
rect 49157 8993 49191 9027
rect 2329 8925 2363 8959
rect 2881 8925 2915 8959
rect 14289 8925 14323 8959
rect 16681 8925 16715 8959
rect 17141 8925 17175 8959
rect 19441 8925 19475 8959
rect 22109 8925 22143 8959
rect 23489 8925 23523 8959
rect 23581 8925 23615 8959
rect 25329 8925 25363 8959
rect 27077 8925 27111 8959
rect 30389 8925 30423 8959
rect 30757 8925 30791 8959
rect 33333 8925 33367 8959
rect 33425 8925 33459 8959
rect 34161 8925 34195 8959
rect 36829 8925 36863 8959
rect 37841 8925 37875 8959
rect 39865 8925 39899 8959
rect 47961 8925 47995 8959
rect 1685 8857 1719 8891
rect 3065 8857 3099 8891
rect 13369 8857 13403 8891
rect 14565 8857 14599 8891
rect 17417 8857 17451 8891
rect 19717 8857 19751 8891
rect 22753 8857 22787 8891
rect 28549 8857 28583 8891
rect 35265 8857 35299 8891
rect 36001 8857 36035 8891
rect 36185 8857 36219 8891
rect 39313 8857 39347 8891
rect 39497 8857 39531 8891
rect 1777 8789 1811 8823
rect 2513 8789 2547 8823
rect 16037 8789 16071 8823
rect 16497 8789 16531 8823
rect 22017 8789 22051 8823
rect 28641 8789 28675 8823
rect 29285 8789 29319 8823
rect 30205 8789 30239 8823
rect 34529 8789 34563 8823
rect 37657 8789 37691 8823
rect 13737 8585 13771 8619
rect 14749 8585 14783 8619
rect 15117 8585 15151 8619
rect 15761 8585 15795 8619
rect 15853 8585 15887 8619
rect 19073 8585 19107 8619
rect 21465 8585 21499 8619
rect 22109 8585 22143 8619
rect 24133 8585 24167 8619
rect 24501 8585 24535 8619
rect 25513 8585 25547 8619
rect 25881 8585 25915 8619
rect 28365 8585 28399 8619
rect 31033 8585 31067 8619
rect 31493 8585 31527 8619
rect 34345 8585 34379 8619
rect 34621 8585 34655 8619
rect 34897 8585 34931 8619
rect 35357 8585 35391 8619
rect 38945 8585 38979 8619
rect 17141 8517 17175 8551
rect 44189 8517 44223 8551
rect 44373 8517 44407 8551
rect 49157 8517 49191 8551
rect 1869 8449 1903 8483
rect 14105 8449 14139 8483
rect 16865 8449 16899 8483
rect 19717 8449 19751 8483
rect 24869 8449 24903 8483
rect 27721 8449 27755 8483
rect 28825 8449 28859 8483
rect 31401 8449 31435 8483
rect 32321 8449 32355 8483
rect 35265 8449 35299 8483
rect 37657 8449 37691 8483
rect 39129 8449 39163 8483
rect 40325 8449 40359 8483
rect 40877 8449 40911 8483
rect 45845 8449 45879 8483
rect 47961 8449 47995 8483
rect 1593 8381 1627 8415
rect 15945 8381 15979 8415
rect 19993 8381 20027 8415
rect 21833 8381 21867 8415
rect 22385 8381 22419 8415
rect 22661 8381 22695 8415
rect 29101 8381 29135 8415
rect 31677 8381 31711 8415
rect 32597 8381 32631 8415
rect 35449 8381 35483 8415
rect 40509 8381 40543 8415
rect 46857 8381 46891 8415
rect 18613 8313 18647 8347
rect 26065 8313 26099 8347
rect 30573 8313 30607 8347
rect 34069 8313 34103 8347
rect 37473 8313 37507 8347
rect 15393 8245 15427 8279
rect 16405 8245 16439 8279
rect 2145 8041 2179 8075
rect 16589 8041 16623 8075
rect 17509 8041 17543 8075
rect 17969 8041 18003 8075
rect 20453 8041 20487 8075
rect 23121 8041 23155 8075
rect 25237 8041 25271 8075
rect 30389 8041 30423 8075
rect 31033 8041 31067 8075
rect 15393 7973 15427 8007
rect 20913 7973 20947 8007
rect 32873 7973 32907 8007
rect 15853 7905 15887 7939
rect 16037 7905 16071 7939
rect 18429 7905 18463 7939
rect 18521 7905 18555 7939
rect 19901 7905 19935 7939
rect 19993 7905 20027 7939
rect 21373 7905 21407 7939
rect 29009 7905 29043 7939
rect 31493 7905 31527 7939
rect 31677 7905 31711 7939
rect 49157 7905 49191 7939
rect 1593 7837 1627 7871
rect 2329 7837 2363 7871
rect 15761 7837 15795 7871
rect 16865 7837 16899 7871
rect 24593 7837 24627 7871
rect 29745 7837 29779 7871
rect 32229 7837 32263 7871
rect 38761 7837 38795 7871
rect 39221 7837 39255 7871
rect 47961 7837 47995 7871
rect 20729 7769 20763 7803
rect 21649 7769 21683 7803
rect 31401 7769 31435 7803
rect 33333 7769 33367 7803
rect 38025 7769 38059 7803
rect 38945 7769 38979 7803
rect 1777 7701 1811 7735
rect 15117 7701 15151 7735
rect 18337 7701 18371 7735
rect 18981 7701 19015 7735
rect 19441 7701 19475 7735
rect 19809 7701 19843 7735
rect 21005 7701 21039 7735
rect 23489 7701 23523 7735
rect 23673 7701 23707 7735
rect 24133 7701 24167 7735
rect 27997 7701 28031 7735
rect 30757 7701 30791 7735
rect 37565 7701 37599 7735
rect 38117 7701 38151 7735
rect 17509 7497 17543 7531
rect 18245 7497 18279 7531
rect 18613 7497 18647 7531
rect 18705 7497 18739 7531
rect 20085 7497 20119 7531
rect 20361 7497 20395 7531
rect 21465 7497 21499 7531
rect 22661 7497 22695 7531
rect 23765 7497 23799 7531
rect 29653 7497 29687 7531
rect 31401 7497 31435 7531
rect 32965 7497 32999 7531
rect 37381 7497 37415 7531
rect 30941 7429 30975 7463
rect 37841 7429 37875 7463
rect 44833 7429 44867 7463
rect 49157 7429 49191 7463
rect 1593 7361 1627 7395
rect 2145 7361 2179 7395
rect 16221 7361 16255 7395
rect 16865 7361 16899 7395
rect 19441 7361 19475 7395
rect 20821 7361 20855 7395
rect 22017 7361 22051 7395
rect 23121 7361 23155 7395
rect 30297 7361 30331 7395
rect 32321 7361 32355 7395
rect 38577 7361 38611 7395
rect 39037 7361 39071 7395
rect 47961 7361 47995 7395
rect 18889 7293 18923 7327
rect 1777 7225 1811 7259
rect 16037 7225 16071 7259
rect 38761 7225 38795 7259
rect 45017 7225 45051 7259
rect 15761 7157 15795 7191
rect 17969 7157 18003 7191
rect 37933 7157 37967 7191
rect 19901 6953 19935 6987
rect 31309 6953 31343 6987
rect 18889 6817 18923 6851
rect 21005 6817 21039 6851
rect 22201 6817 22235 6851
rect 31033 6817 31067 6851
rect 49157 6817 49191 6851
rect 2513 6749 2547 6783
rect 2789 6749 2823 6783
rect 18245 6749 18279 6783
rect 20361 6749 20395 6783
rect 21557 6749 21591 6783
rect 30389 6749 30423 6783
rect 46121 6749 46155 6783
rect 47961 6749 47995 6783
rect 1685 6681 1719 6715
rect 1869 6681 1903 6715
rect 47317 6681 47351 6715
rect 2329 6613 2363 6647
rect 16405 6613 16439 6647
rect 17785 6613 17819 6647
rect 19441 6613 19475 6647
rect 2145 6409 2179 6443
rect 18705 6409 18739 6443
rect 19901 6409 19935 6443
rect 37565 6341 37599 6375
rect 38025 6341 38059 6375
rect 44005 6341 44039 6375
rect 49157 6341 49191 6375
rect 1593 6273 1627 6307
rect 2329 6273 2363 6307
rect 18337 6273 18371 6307
rect 19257 6273 19291 6307
rect 20545 6273 20579 6307
rect 47961 6273 47995 6307
rect 1777 6137 1811 6171
rect 18153 6137 18187 6171
rect 44189 6137 44223 6171
rect 20361 6069 20395 6103
rect 37657 6069 37691 6103
rect 1777 5797 1811 5831
rect 3065 5729 3099 5763
rect 49157 5729 49191 5763
rect 1593 5661 1627 5695
rect 2329 5661 2363 5695
rect 2881 5661 2915 5695
rect 43729 5661 43763 5695
rect 47961 5661 47995 5695
rect 43913 5593 43947 5627
rect 2513 5525 2547 5559
rect 37381 5321 37415 5355
rect 38577 5253 38611 5287
rect 39037 5253 39071 5287
rect 49157 5253 49191 5287
rect 37841 5185 37875 5219
rect 45845 5185 45879 5219
rect 47961 5185 47995 5219
rect 1593 5117 1627 5151
rect 1869 5117 1903 5151
rect 46857 5117 46891 5151
rect 38761 5049 38795 5083
rect 37933 4981 37967 5015
rect 2145 4777 2179 4811
rect 36921 4777 36955 4811
rect 25237 4641 25271 4675
rect 26249 4641 26283 4675
rect 49157 4641 49191 4675
rect 1593 4573 1627 4607
rect 2329 4573 2363 4607
rect 22252 4573 22286 4607
rect 22880 4573 22914 4607
rect 23708 4573 23742 4607
rect 38117 4573 38151 4607
rect 38577 4573 38611 4607
rect 47961 4573 47995 4607
rect 22339 4505 22373 4539
rect 23811 4505 23845 4539
rect 25421 4505 25455 4539
rect 37381 4505 37415 4539
rect 38301 4505 38335 4539
rect 1777 4437 1811 4471
rect 22983 4437 23017 4471
rect 24225 4437 24259 4471
rect 37473 4437 37507 4471
rect 1685 4165 1719 4199
rect 24501 4165 24535 4199
rect 27353 4165 27387 4199
rect 2329 4097 2363 4131
rect 3065 4097 3099 4131
rect 18337 4097 18371 4131
rect 27169 4097 27203 4131
rect 45845 4097 45879 4131
rect 47961 4097 47995 4131
rect 49157 4097 49191 4131
rect 2881 4029 2915 4063
rect 18521 4029 18555 4063
rect 20177 4029 20211 4063
rect 22017 4029 22051 4063
rect 22293 4029 22327 4063
rect 24317 4029 24351 4063
rect 25697 4029 25731 4063
rect 27629 4029 27663 4063
rect 46673 4029 46707 4063
rect 2513 3961 2547 3995
rect 1777 3893 1811 3927
rect 23765 3893 23799 3927
rect 20085 3689 20119 3723
rect 23995 3689 24029 3723
rect 36553 3689 36587 3723
rect 17601 3621 17635 3655
rect 21189 3553 21223 3587
rect 21373 3553 21407 3587
rect 24777 3553 24811 3587
rect 25053 3553 25087 3587
rect 49157 3553 49191 3587
rect 1593 3485 1627 3519
rect 1869 3485 1903 3519
rect 16497 3485 16531 3519
rect 17785 3485 17819 3519
rect 19441 3485 19475 3519
rect 23892 3485 23926 3519
rect 24593 3485 24627 3519
rect 36461 3485 36495 3519
rect 36921 3485 36955 3519
rect 46121 3485 46155 3519
rect 47961 3485 47995 3519
rect 23029 3417 23063 3451
rect 47317 3417 47351 3451
rect 16589 3349 16623 3383
rect 2145 3145 2179 3179
rect 31217 3145 31251 3179
rect 22937 3077 22971 3111
rect 49157 3077 49191 3111
rect 1593 3009 1627 3043
rect 2513 3009 2547 3043
rect 14565 3009 14599 3043
rect 17049 3009 17083 3043
rect 19073 3009 19107 3043
rect 19625 3009 19659 3043
rect 22753 3009 22787 3043
rect 25053 3009 25087 3043
rect 27905 3009 27939 3043
rect 29101 3009 29135 3043
rect 44005 3009 44039 3043
rect 45845 3009 45879 3043
rect 47961 3009 47995 3043
rect 14841 2941 14875 2975
rect 17325 2941 17359 2975
rect 19809 2941 19843 2975
rect 21465 2941 21499 2975
rect 24593 2941 24627 2975
rect 28549 2941 28583 2975
rect 29377 2941 29411 2975
rect 45201 2941 45235 2975
rect 46857 2941 46891 2975
rect 1777 2873 1811 2907
rect 18889 2873 18923 2907
rect 2329 2805 2363 2839
rect 2789 2805 2823 2839
rect 16313 2805 16347 2839
rect 25697 2805 25731 2839
rect 30849 2805 30883 2839
rect 3065 2601 3099 2635
rect 9689 2601 9723 2635
rect 16405 2601 16439 2635
rect 21005 2601 21039 2635
rect 22753 2601 22787 2635
rect 23765 2601 23799 2635
rect 26341 2601 26375 2635
rect 27905 2601 27939 2635
rect 32965 2601 32999 2635
rect 35081 2601 35115 2635
rect 2513 2533 2547 2567
rect 21373 2533 21407 2567
rect 22937 2533 22971 2567
rect 23949 2533 23983 2567
rect 12265 2465 12299 2499
rect 14749 2465 14783 2499
rect 24593 2465 24627 2499
rect 24869 2465 24903 2499
rect 26709 2465 26743 2499
rect 37749 2465 37783 2499
rect 41429 2465 41463 2499
rect 49157 2465 49191 2499
rect 1593 2397 1627 2431
rect 2329 2397 2363 2431
rect 3249 2397 3283 2431
rect 3525 2397 3559 2431
rect 9873 2397 9907 2431
rect 10149 2397 10183 2431
rect 11989 2397 12023 2431
rect 14473 2397 14507 2431
rect 17693 2397 17727 2431
rect 20453 2397 20487 2431
rect 20913 2397 20947 2431
rect 22477 2397 22511 2431
rect 23489 2397 23523 2431
rect 27629 2397 27663 2431
rect 28917 2397 28951 2431
rect 29193 2397 29227 2431
rect 31033 2397 31067 2431
rect 31309 2397 31343 2431
rect 33149 2397 33183 2431
rect 33425 2397 33459 2431
rect 35265 2397 35299 2431
rect 35541 2397 35575 2431
rect 37473 2397 37507 2431
rect 40693 2397 40727 2431
rect 45845 2397 45879 2431
rect 47961 2397 47995 2431
rect 18429 2329 18463 2363
rect 47041 2329 47075 2363
rect 1777 2261 1811 2295
rect 20269 2261 20303 2295
rect 28089 2261 28123 2295
rect 28733 2261 28767 2295
rect 30849 2261 30883 2295
rect 37105 2261 37139 2295
<< metal1 >>
rect 24670 26324 24676 26376
rect 24728 26364 24734 26376
rect 43898 26364 43904 26376
rect 24728 26336 43904 26364
rect 24728 26324 24734 26336
rect 43898 26324 43904 26336
rect 43956 26324 43962 26376
rect 28902 26256 28908 26308
rect 28960 26296 28966 26308
rect 45094 26296 45100 26308
rect 28960 26268 45100 26296
rect 28960 26256 28966 26268
rect 45094 26256 45100 26268
rect 45152 26256 45158 26308
rect 27522 26188 27528 26240
rect 27580 26228 27586 26240
rect 40034 26228 40040 26240
rect 27580 26200 40040 26228
rect 27580 26188 27586 26200
rect 40034 26188 40040 26200
rect 40092 26188 40098 26240
rect 33410 26120 33416 26172
rect 33468 26160 33474 26172
rect 45278 26160 45284 26172
rect 33468 26132 45284 26160
rect 33468 26120 33474 26132
rect 45278 26120 45284 26132
rect 45336 26120 45342 26172
rect 34422 26052 34428 26104
rect 34480 26092 34486 26104
rect 45830 26092 45836 26104
rect 34480 26064 45836 26092
rect 34480 26052 34486 26064
rect 45830 26052 45836 26064
rect 45888 26052 45894 26104
rect 33778 25984 33784 26036
rect 33836 26024 33842 26036
rect 44634 26024 44640 26036
rect 33836 25996 44640 26024
rect 33836 25984 33842 25996
rect 44634 25984 44640 25996
rect 44692 25984 44698 26036
rect 36998 25916 37004 25968
rect 37056 25956 37062 25968
rect 46014 25956 46020 25968
rect 37056 25928 46020 25956
rect 37056 25916 37062 25928
rect 46014 25916 46020 25928
rect 46072 25916 46078 25968
rect 25222 25712 25228 25764
rect 25280 25752 25286 25764
rect 38654 25752 38660 25764
rect 25280 25724 38660 25752
rect 25280 25712 25286 25724
rect 38654 25712 38660 25724
rect 38712 25712 38718 25764
rect 31846 25644 31852 25696
rect 31904 25684 31910 25696
rect 38930 25684 38936 25696
rect 31904 25656 38936 25684
rect 31904 25644 31910 25656
rect 38930 25644 38936 25656
rect 38988 25644 38994 25696
rect 25866 25576 25872 25628
rect 25924 25616 25930 25628
rect 40586 25616 40592 25628
rect 25924 25588 40592 25616
rect 25924 25576 25930 25588
rect 40586 25576 40592 25588
rect 40644 25576 40650 25628
rect 24026 25508 24032 25560
rect 24084 25548 24090 25560
rect 42610 25548 42616 25560
rect 24084 25520 42616 25548
rect 24084 25508 24090 25520
rect 42610 25508 42616 25520
rect 42668 25508 42674 25560
rect 29822 25440 29828 25492
rect 29880 25480 29886 25492
rect 43346 25480 43352 25492
rect 29880 25452 43352 25480
rect 29880 25440 29886 25452
rect 43346 25440 43352 25452
rect 43404 25440 43410 25492
rect 31570 25372 31576 25424
rect 31628 25412 31634 25424
rect 48406 25412 48412 25424
rect 31628 25384 48412 25412
rect 31628 25372 31634 25384
rect 48406 25372 48412 25384
rect 48464 25372 48470 25424
rect 22462 25304 22468 25356
rect 22520 25344 22526 25356
rect 48774 25344 48780 25356
rect 22520 25316 48780 25344
rect 22520 25304 22526 25316
rect 48774 25304 48780 25316
rect 48832 25304 48838 25356
rect 28626 25236 28632 25288
rect 28684 25276 28690 25288
rect 38838 25276 38844 25288
rect 28684 25248 38844 25276
rect 28684 25236 28690 25248
rect 38838 25236 38844 25248
rect 38896 25236 38902 25288
rect 38930 25236 38936 25288
rect 38988 25276 38994 25288
rect 43438 25276 43444 25288
rect 38988 25248 43444 25276
rect 38988 25236 38994 25248
rect 43438 25236 43444 25248
rect 43496 25236 43502 25288
rect 37734 25168 37740 25220
rect 37792 25208 37798 25220
rect 48958 25208 48964 25220
rect 37792 25180 48964 25208
rect 37792 25168 37798 25180
rect 48958 25168 48964 25180
rect 49016 25168 49022 25220
rect 35986 25100 35992 25152
rect 36044 25140 36050 25152
rect 42518 25140 42524 25152
rect 36044 25112 42524 25140
rect 36044 25100 36050 25112
rect 42518 25100 42524 25112
rect 42576 25100 42582 25152
rect 35802 25032 35808 25084
rect 35860 25072 35866 25084
rect 44358 25072 44364 25084
rect 35860 25044 44364 25072
rect 35860 25032 35866 25044
rect 44358 25032 44364 25044
rect 44416 25032 44422 25084
rect 33318 24964 33324 25016
rect 33376 25004 33382 25016
rect 42334 25004 42340 25016
rect 33376 24976 42340 25004
rect 33376 24964 33382 24976
rect 42334 24964 42340 24976
rect 42392 24964 42398 25016
rect 37642 24896 37648 24948
rect 37700 24936 37706 24948
rect 44450 24936 44456 24948
rect 37700 24908 44456 24936
rect 37700 24896 37706 24908
rect 44450 24896 44456 24908
rect 44508 24896 44514 24948
rect 3050 24828 3056 24880
rect 3108 24868 3114 24880
rect 9858 24868 9864 24880
rect 3108 24840 9864 24868
rect 3108 24828 3114 24840
rect 9858 24828 9864 24840
rect 9916 24828 9922 24880
rect 36722 24828 36728 24880
rect 36780 24868 36786 24880
rect 43990 24868 43996 24880
rect 36780 24840 43996 24868
rect 36780 24828 36786 24840
rect 43990 24828 43996 24840
rect 44048 24828 44054 24880
rect 3418 24760 3424 24812
rect 3476 24800 3482 24812
rect 7190 24800 7196 24812
rect 3476 24772 7196 24800
rect 3476 24760 3482 24772
rect 7190 24760 7196 24772
rect 7248 24760 7254 24812
rect 19426 24760 19432 24812
rect 19484 24800 19490 24812
rect 25498 24800 25504 24812
rect 19484 24772 25504 24800
rect 19484 24760 19490 24772
rect 25498 24760 25504 24772
rect 25556 24760 25562 24812
rect 34238 24760 34244 24812
rect 34296 24800 34302 24812
rect 38746 24800 38752 24812
rect 34296 24772 38752 24800
rect 34296 24760 34302 24772
rect 38746 24760 38752 24772
rect 38804 24760 38810 24812
rect 40218 24760 40224 24812
rect 40276 24800 40282 24812
rect 45646 24800 45652 24812
rect 40276 24772 45652 24800
rect 40276 24760 40282 24772
rect 45646 24760 45652 24772
rect 45704 24760 45710 24812
rect 20530 24692 20536 24744
rect 20588 24732 20594 24744
rect 28350 24732 28356 24744
rect 20588 24704 28356 24732
rect 20588 24692 20594 24704
rect 28350 24692 28356 24704
rect 28408 24692 28414 24744
rect 34054 24692 34060 24744
rect 34112 24732 34118 24744
rect 39666 24732 39672 24744
rect 34112 24704 39672 24732
rect 34112 24692 34118 24704
rect 39666 24692 39672 24704
rect 39724 24692 39730 24744
rect 43806 24692 43812 24744
rect 43864 24732 43870 24744
rect 46566 24732 46572 24744
rect 43864 24704 46572 24732
rect 43864 24692 43870 24704
rect 46566 24692 46572 24704
rect 46624 24692 46630 24744
rect 11790 24624 11796 24676
rect 11848 24664 11854 24676
rect 25406 24664 25412 24676
rect 11848 24636 25412 24664
rect 11848 24624 11854 24636
rect 25406 24624 25412 24636
rect 25464 24624 25470 24676
rect 36538 24624 36544 24676
rect 36596 24664 36602 24676
rect 40310 24664 40316 24676
rect 36596 24636 40316 24664
rect 36596 24624 36602 24636
rect 40310 24624 40316 24636
rect 40368 24624 40374 24676
rect 42426 24624 42432 24676
rect 42484 24664 42490 24676
rect 47578 24664 47584 24676
rect 42484 24636 47584 24664
rect 42484 24624 42490 24636
rect 47578 24624 47584 24636
rect 47636 24624 47642 24676
rect 2130 24556 2136 24608
rect 2188 24596 2194 24608
rect 10962 24596 10968 24608
rect 2188 24568 10968 24596
rect 2188 24556 2194 24568
rect 10962 24556 10968 24568
rect 11020 24556 11026 24608
rect 19610 24556 19616 24608
rect 19668 24596 19674 24608
rect 25774 24596 25780 24608
rect 19668 24568 25780 24596
rect 19668 24556 19674 24568
rect 25774 24556 25780 24568
rect 25832 24556 25838 24608
rect 30282 24556 30288 24608
rect 30340 24596 30346 24608
rect 35802 24596 35808 24608
rect 30340 24568 35808 24596
rect 30340 24556 30346 24568
rect 35802 24556 35808 24568
rect 35860 24556 35866 24608
rect 36722 24556 36728 24608
rect 36780 24596 36786 24608
rect 39206 24596 39212 24608
rect 36780 24568 39212 24596
rect 36780 24556 36786 24568
rect 39206 24556 39212 24568
rect 39264 24556 39270 24608
rect 43622 24556 43628 24608
rect 43680 24596 43686 24608
rect 47946 24596 47952 24608
rect 43680 24568 47952 24596
rect 43680 24556 43686 24568
rect 47946 24556 47952 24568
rect 48004 24556 48010 24608
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 2774 24352 2780 24404
rect 2832 24392 2838 24404
rect 6178 24392 6184 24404
rect 2832 24364 6184 24392
rect 2832 24352 2838 24364
rect 6178 24352 6184 24364
rect 6236 24352 6242 24404
rect 13446 24392 13452 24404
rect 6564 24364 13452 24392
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 3510 24256 3516 24268
rect 3283 24228 3516 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 5813 24259 5871 24265
rect 5813 24225 5825 24259
rect 5859 24256 5871 24259
rect 6454 24256 6460 24268
rect 5859 24228 6460 24256
rect 5859 24225 5871 24228
rect 5813 24219 5871 24225
rect 6454 24216 6460 24228
rect 6512 24216 6518 24268
rect 6564 24265 6592 24364
rect 13446 24352 13452 24364
rect 13504 24352 13510 24404
rect 16853 24395 16911 24401
rect 16853 24361 16865 24395
rect 16899 24392 16911 24395
rect 21726 24392 21732 24404
rect 16899 24364 21732 24392
rect 16899 24361 16911 24364
rect 16853 24355 16911 24361
rect 21726 24352 21732 24364
rect 21784 24352 21790 24404
rect 22278 24352 22284 24404
rect 22336 24392 22342 24404
rect 22336 24364 24808 24392
rect 22336 24352 22342 24364
rect 6886 24296 12020 24324
rect 6549 24259 6607 24265
rect 6549 24225 6561 24259
rect 6595 24225 6607 24259
rect 6549 24219 6607 24225
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 2314 24188 2320 24200
rect 2271 24160 2320 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 2314 24148 2320 24160
rect 2372 24148 2378 24200
rect 4157 24191 4215 24197
rect 4157 24157 4169 24191
rect 4203 24157 4215 24191
rect 4157 24151 4215 24157
rect 4801 24191 4859 24197
rect 4801 24157 4813 24191
rect 4847 24188 4859 24191
rect 4890 24188 4896 24200
rect 4847 24160 4896 24188
rect 4847 24157 4859 24160
rect 4801 24151 4859 24157
rect 4172 24120 4200 24151
rect 4890 24148 4896 24160
rect 4948 24148 4954 24200
rect 5258 24148 5264 24200
rect 5316 24188 5322 24200
rect 6886 24188 6914 24296
rect 8205 24259 8263 24265
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 8662 24256 8668 24268
rect 8251 24228 8668 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 8662 24216 8668 24228
rect 8720 24216 8726 24268
rect 5316 24160 6914 24188
rect 5316 24148 5322 24160
rect 7374 24148 7380 24200
rect 7432 24148 7438 24200
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24188 9367 24191
rect 9674 24188 9680 24200
rect 9355 24160 9680 24188
rect 9355 24157 9367 24160
rect 9309 24151 9367 24157
rect 9674 24148 9680 24160
rect 9732 24148 9738 24200
rect 9953 24191 10011 24197
rect 9953 24157 9965 24191
rect 9999 24188 10011 24191
rect 10778 24188 10784 24200
rect 9999 24160 10784 24188
rect 9999 24157 10011 24160
rect 9953 24151 10011 24157
rect 10778 24148 10784 24160
rect 10836 24148 10842 24200
rect 11606 24148 11612 24200
rect 11664 24188 11670 24200
rect 11885 24191 11943 24197
rect 11885 24188 11897 24191
rect 11664 24160 11897 24188
rect 11664 24148 11670 24160
rect 11885 24157 11897 24160
rect 11931 24157 11943 24191
rect 11992 24188 12020 24296
rect 14274 24284 14280 24336
rect 14332 24324 14338 24336
rect 14332 24296 19380 24324
rect 14332 24284 14338 24296
rect 13541 24259 13599 24265
rect 13541 24225 13553 24259
rect 13587 24256 13599 24259
rect 14458 24256 14464 24268
rect 13587 24228 14464 24256
rect 13587 24225 13599 24228
rect 13541 24219 13599 24225
rect 14458 24216 14464 24228
rect 14516 24216 14522 24268
rect 16117 24259 16175 24265
rect 16117 24225 16129 24259
rect 16163 24256 16175 24259
rect 18322 24256 18328 24268
rect 16163 24228 18328 24256
rect 16163 24225 16175 24228
rect 16117 24219 16175 24225
rect 18322 24216 18328 24228
rect 18380 24216 18386 24268
rect 18693 24259 18751 24265
rect 18693 24225 18705 24259
rect 18739 24256 18751 24259
rect 19242 24256 19248 24268
rect 18739 24228 19248 24256
rect 18739 24225 18751 24228
rect 18693 24219 18751 24225
rect 19242 24216 19248 24228
rect 19300 24216 19306 24268
rect 19352 24256 19380 24296
rect 19426 24284 19432 24336
rect 19484 24284 19490 24336
rect 22370 24324 22376 24336
rect 19536 24296 22376 24324
rect 19536 24256 19564 24296
rect 22370 24284 22376 24296
rect 22428 24284 22434 24336
rect 19352 24228 19564 24256
rect 19720 24228 20208 24256
rect 12345 24191 12403 24197
rect 12345 24188 12357 24191
rect 11992 24160 12357 24188
rect 11885 24151 11943 24157
rect 12345 24157 12357 24160
rect 12391 24157 12403 24191
rect 12345 24151 12403 24157
rect 15105 24191 15163 24197
rect 15105 24157 15117 24191
rect 15151 24157 15163 24191
rect 15105 24151 15163 24157
rect 17037 24191 17095 24197
rect 17037 24157 17049 24191
rect 17083 24188 17095 24191
rect 17126 24188 17132 24200
rect 17083 24160 17132 24188
rect 17083 24157 17095 24160
rect 17037 24151 17095 24157
rect 5902 24120 5908 24132
rect 4172 24092 5908 24120
rect 5902 24080 5908 24092
rect 5960 24080 5966 24132
rect 10965 24123 11023 24129
rect 10965 24089 10977 24123
rect 11011 24120 11023 24123
rect 12526 24120 12532 24132
rect 11011 24092 12532 24120
rect 11011 24089 11023 24092
rect 10965 24083 11023 24089
rect 12526 24080 12532 24092
rect 12584 24080 12590 24132
rect 15120 24120 15148 24151
rect 17126 24148 17132 24160
rect 17184 24148 17190 24200
rect 17681 24191 17739 24197
rect 17681 24157 17693 24191
rect 17727 24188 17739 24191
rect 17770 24188 17776 24200
rect 17727 24160 17776 24188
rect 17727 24157 17739 24160
rect 17681 24151 17739 24157
rect 17770 24148 17776 24160
rect 17828 24148 17834 24200
rect 19610 24148 19616 24200
rect 19668 24148 19674 24200
rect 19720 24120 19748 24228
rect 20073 24191 20131 24197
rect 20073 24157 20085 24191
rect 20119 24157 20131 24191
rect 20180 24188 20208 24228
rect 20898 24216 20904 24268
rect 20956 24216 20962 24268
rect 23382 24256 23388 24268
rect 22066 24228 23388 24256
rect 22066 24188 22094 24228
rect 23382 24216 23388 24228
rect 23440 24216 23446 24268
rect 24780 24256 24808 24364
rect 24854 24352 24860 24404
rect 24912 24352 24918 24404
rect 25130 24352 25136 24404
rect 25188 24392 25194 24404
rect 28997 24395 29055 24401
rect 28997 24392 29009 24395
rect 25188 24364 29009 24392
rect 25188 24352 25194 24364
rect 28997 24361 29009 24364
rect 29043 24361 29055 24395
rect 28997 24355 29055 24361
rect 30190 24352 30196 24404
rect 30248 24392 30254 24404
rect 36262 24392 36268 24404
rect 30248 24364 36268 24392
rect 30248 24352 30254 24364
rect 36262 24352 36268 24364
rect 36320 24352 36326 24404
rect 39390 24352 39396 24404
rect 39448 24392 39454 24404
rect 39577 24395 39635 24401
rect 39577 24392 39589 24395
rect 39448 24364 39589 24392
rect 39448 24352 39454 24364
rect 39577 24361 39589 24364
rect 39623 24361 39635 24395
rect 39577 24355 39635 24361
rect 26421 24327 26479 24333
rect 26421 24293 26433 24327
rect 26467 24324 26479 24327
rect 27614 24324 27620 24336
rect 26467 24296 27620 24324
rect 26467 24293 26479 24296
rect 26421 24287 26479 24293
rect 27614 24284 27620 24296
rect 27672 24284 27678 24336
rect 29638 24284 29644 24336
rect 29696 24324 29702 24336
rect 30282 24324 30288 24336
rect 29696 24296 30288 24324
rect 29696 24284 29702 24296
rect 30282 24284 30288 24296
rect 30340 24324 30346 24336
rect 30469 24327 30527 24333
rect 30469 24324 30481 24327
rect 30340 24296 30481 24324
rect 30340 24284 30346 24296
rect 30469 24293 30481 24296
rect 30515 24293 30527 24327
rect 30469 24287 30527 24293
rect 33980 24296 35204 24324
rect 33980 24256 34008 24296
rect 24780 24228 34008 24256
rect 20180 24160 22094 24188
rect 22189 24191 22247 24197
rect 20073 24151 20131 24157
rect 22189 24157 22201 24191
rect 22235 24188 22247 24191
rect 22554 24188 22560 24200
rect 22235 24160 22560 24188
rect 22235 24157 22247 24160
rect 22189 24151 22247 24157
rect 15120 24092 19748 24120
rect 3970 24012 3976 24064
rect 4028 24012 4034 24064
rect 8846 24012 8852 24064
rect 8904 24052 8910 24064
rect 9125 24055 9183 24061
rect 9125 24052 9137 24055
rect 8904 24024 9137 24052
rect 8904 24012 8910 24024
rect 9125 24021 9137 24024
rect 9171 24021 9183 24055
rect 9125 24015 9183 24021
rect 11701 24055 11759 24061
rect 11701 24021 11713 24055
rect 11747 24052 11759 24055
rect 12434 24052 12440 24064
rect 11747 24024 12440 24052
rect 11747 24021 11759 24024
rect 11701 24015 11759 24021
rect 12434 24012 12440 24024
rect 12492 24012 12498 24064
rect 14277 24055 14335 24061
rect 14277 24021 14289 24055
rect 14323 24052 14335 24055
rect 15010 24052 15016 24064
rect 14323 24024 15016 24052
rect 14323 24021 14335 24024
rect 14277 24015 14335 24021
rect 15010 24012 15016 24024
rect 15068 24012 15074 24064
rect 17402 24012 17408 24064
rect 17460 24052 17466 24064
rect 19150 24052 19156 24064
rect 17460 24024 19156 24052
rect 17460 24012 17466 24024
rect 19150 24012 19156 24024
rect 19208 24012 19214 24064
rect 20088 24052 20116 24151
rect 22554 24148 22560 24160
rect 22612 24148 22618 24200
rect 22925 24191 22983 24197
rect 22925 24188 22937 24191
rect 22664 24160 22937 24188
rect 20254 24080 20260 24132
rect 20312 24120 20318 24132
rect 22664 24120 22692 24160
rect 22925 24157 22937 24160
rect 22971 24157 22983 24191
rect 22925 24151 22983 24157
rect 24026 24148 24032 24200
rect 24084 24148 24090 24200
rect 24780 24197 24808 24228
rect 34054 24216 34060 24268
rect 34112 24216 34118 24268
rect 34238 24216 34244 24268
rect 34296 24216 34302 24268
rect 35176 24256 35204 24296
rect 35250 24284 35256 24336
rect 35308 24324 35314 24336
rect 39301 24327 39359 24333
rect 39301 24324 39313 24327
rect 35308 24296 39313 24324
rect 35308 24284 35314 24296
rect 39301 24293 39313 24296
rect 39347 24293 39359 24327
rect 39592 24324 39620 24355
rect 40034 24352 40040 24404
rect 40092 24392 40098 24404
rect 41138 24392 41144 24404
rect 40092 24364 41144 24392
rect 40092 24352 40098 24364
rect 41138 24352 41144 24364
rect 41196 24392 41202 24404
rect 47029 24395 47087 24401
rect 47029 24392 47041 24395
rect 41196 24364 47041 24392
rect 41196 24352 41202 24364
rect 47029 24361 47041 24364
rect 47075 24361 47087 24395
rect 47029 24355 47087 24361
rect 47946 24352 47952 24404
rect 48004 24352 48010 24404
rect 44726 24324 44732 24336
rect 39592 24296 44732 24324
rect 39301 24287 39359 24293
rect 44726 24284 44732 24296
rect 44784 24284 44790 24336
rect 44818 24284 44824 24336
rect 44876 24324 44882 24336
rect 46753 24327 46811 24333
rect 46753 24324 46765 24327
rect 44876 24296 46765 24324
rect 44876 24284 44882 24296
rect 46753 24293 46765 24296
rect 46799 24293 46811 24327
rect 46753 24287 46811 24293
rect 47210 24284 47216 24336
rect 47268 24284 47274 24336
rect 35342 24256 35348 24268
rect 35176 24228 35348 24256
rect 35342 24216 35348 24228
rect 35400 24216 35406 24268
rect 35529 24259 35587 24265
rect 35529 24225 35541 24259
rect 35575 24256 35587 24259
rect 35802 24256 35808 24268
rect 35575 24228 35808 24256
rect 35575 24225 35587 24228
rect 35529 24219 35587 24225
rect 35802 24216 35808 24228
rect 35860 24216 35866 24268
rect 36538 24216 36544 24268
rect 36596 24216 36602 24268
rect 36722 24216 36728 24268
rect 36780 24216 36786 24268
rect 37918 24216 37924 24268
rect 37976 24216 37982 24268
rect 38105 24259 38163 24265
rect 38105 24225 38117 24259
rect 38151 24256 38163 24259
rect 38378 24256 38384 24268
rect 38151 24228 38384 24256
rect 38151 24225 38163 24228
rect 38105 24219 38163 24225
rect 38378 24216 38384 24228
rect 38436 24216 38442 24268
rect 39482 24216 39488 24268
rect 39540 24256 39546 24268
rect 39540 24228 40816 24256
rect 39540 24216 39546 24228
rect 24765 24191 24823 24197
rect 24765 24157 24777 24191
rect 24811 24157 24823 24191
rect 24765 24151 24823 24157
rect 25409 24191 25467 24197
rect 25409 24157 25421 24191
rect 25455 24188 25467 24191
rect 26602 24188 26608 24200
rect 25455 24160 26608 24188
rect 25455 24157 25467 24160
rect 25409 24151 25467 24157
rect 26602 24148 26608 24160
rect 26660 24148 26666 24200
rect 27249 24191 27307 24197
rect 27249 24157 27261 24191
rect 27295 24188 27307 24191
rect 27338 24188 27344 24200
rect 27295 24160 27344 24188
rect 27295 24157 27307 24160
rect 27249 24151 27307 24157
rect 27338 24148 27344 24160
rect 27396 24148 27402 24200
rect 28350 24148 28356 24200
rect 28408 24148 28414 24200
rect 30282 24148 30288 24200
rect 30340 24188 30346 24200
rect 30837 24191 30895 24197
rect 30837 24188 30849 24191
rect 30340 24160 30849 24188
rect 30340 24148 30346 24160
rect 30837 24157 30849 24160
rect 30883 24157 30895 24191
rect 30837 24151 30895 24157
rect 31478 24148 31484 24200
rect 31536 24188 31542 24200
rect 32493 24191 32551 24197
rect 32493 24188 32505 24191
rect 31536 24160 32505 24188
rect 31536 24148 31542 24160
rect 32493 24157 32505 24160
rect 32539 24157 32551 24191
rect 32493 24151 32551 24157
rect 35066 24148 35072 24200
rect 35124 24188 35130 24200
rect 35253 24191 35311 24197
rect 35253 24188 35265 24191
rect 35124 24160 35265 24188
rect 35124 24148 35130 24160
rect 35253 24157 35265 24160
rect 35299 24188 35311 24191
rect 37826 24188 37832 24200
rect 35299 24160 37832 24188
rect 35299 24157 35311 24160
rect 35253 24151 35311 24157
rect 37826 24148 37832 24160
rect 37884 24148 37890 24200
rect 38657 24191 38715 24197
rect 38657 24188 38669 24191
rect 37936 24160 38669 24188
rect 20312 24092 22692 24120
rect 20312 24080 20318 24092
rect 22738 24080 22744 24132
rect 22796 24120 22802 24132
rect 26878 24120 26884 24132
rect 22796 24092 26884 24120
rect 22796 24080 22802 24092
rect 26878 24080 26884 24092
rect 26936 24080 26942 24132
rect 29362 24080 29368 24132
rect 29420 24120 29426 24132
rect 29825 24123 29883 24129
rect 29825 24120 29837 24123
rect 29420 24092 29837 24120
rect 29420 24080 29426 24092
rect 29825 24089 29837 24092
rect 29871 24089 29883 24123
rect 29825 24083 29883 24089
rect 30377 24123 30435 24129
rect 30377 24089 30389 24123
rect 30423 24120 30435 24123
rect 31110 24120 31116 24132
rect 30423 24092 31116 24120
rect 30423 24089 30435 24092
rect 30377 24083 30435 24089
rect 31110 24080 31116 24092
rect 31168 24080 31174 24132
rect 31294 24080 31300 24132
rect 31352 24120 31358 24132
rect 31757 24123 31815 24129
rect 31757 24120 31769 24123
rect 31352 24092 31769 24120
rect 31352 24080 31358 24092
rect 31757 24089 31769 24092
rect 31803 24089 31815 24123
rect 31757 24083 31815 24089
rect 33137 24123 33195 24129
rect 33137 24089 33149 24123
rect 33183 24120 33195 24123
rect 33870 24120 33876 24132
rect 33183 24092 33876 24120
rect 33183 24089 33195 24092
rect 33137 24083 33195 24089
rect 33870 24080 33876 24092
rect 33928 24080 33934 24132
rect 33965 24123 34023 24129
rect 33965 24089 33977 24123
rect 34011 24120 34023 24123
rect 34011 24092 35296 24120
rect 34011 24089 34023 24092
rect 33965 24083 34023 24089
rect 23845 24055 23903 24061
rect 23845 24052 23857 24055
rect 20088 24024 23857 24052
rect 23845 24021 23857 24024
rect 23891 24021 23903 24055
rect 23845 24015 23903 24021
rect 25958 24012 25964 24064
rect 26016 24052 26022 24064
rect 26053 24055 26111 24061
rect 26053 24052 26065 24055
rect 26016 24024 26065 24052
rect 26016 24012 26022 24024
rect 26053 24021 26065 24024
rect 26099 24021 26111 24055
rect 26053 24015 26111 24021
rect 26510 24012 26516 24064
rect 26568 24052 26574 24064
rect 26697 24055 26755 24061
rect 26697 24052 26709 24055
rect 26568 24024 26709 24052
rect 26568 24012 26574 24024
rect 26697 24021 26709 24024
rect 26743 24021 26755 24055
rect 26697 24015 26755 24021
rect 26786 24012 26792 24064
rect 26844 24052 26850 24064
rect 27893 24055 27951 24061
rect 27893 24052 27905 24055
rect 26844 24024 27905 24052
rect 26844 24012 26850 24024
rect 27893 24021 27905 24024
rect 27939 24021 27951 24055
rect 27893 24015 27951 24021
rect 29273 24055 29331 24061
rect 29273 24021 29285 24055
rect 29319 24052 29331 24055
rect 29638 24052 29644 24064
rect 29319 24024 29644 24052
rect 29319 24021 29331 24024
rect 29273 24015 29331 24021
rect 29638 24012 29644 24024
rect 29696 24012 29702 24064
rect 29914 24012 29920 24064
rect 29972 24012 29978 24064
rect 31481 24055 31539 24061
rect 31481 24021 31493 24055
rect 31527 24052 31539 24055
rect 31662 24052 31668 24064
rect 31527 24024 31668 24052
rect 31527 24021 31539 24024
rect 31481 24015 31539 24021
rect 31662 24012 31668 24024
rect 31720 24012 31726 24064
rect 32122 24012 32128 24064
rect 32180 24012 32186 24064
rect 33594 24012 33600 24064
rect 33652 24012 33658 24064
rect 34885 24055 34943 24061
rect 34885 24021 34897 24055
rect 34931 24052 34943 24055
rect 35158 24052 35164 24064
rect 34931 24024 35164 24052
rect 34931 24021 34943 24024
rect 34885 24015 34943 24021
rect 35158 24012 35164 24024
rect 35216 24012 35222 24064
rect 35268 24052 35296 24092
rect 35526 24080 35532 24132
rect 35584 24120 35590 24132
rect 37936 24120 37964 24160
rect 38657 24157 38669 24160
rect 38703 24157 38715 24191
rect 38657 24151 38715 24157
rect 39114 24148 39120 24200
rect 39172 24188 39178 24200
rect 39390 24188 39396 24200
rect 39172 24160 39396 24188
rect 39172 24148 39178 24160
rect 39390 24148 39396 24160
rect 39448 24148 39454 24200
rect 40037 24191 40095 24197
rect 40037 24157 40049 24191
rect 40083 24188 40095 24191
rect 40218 24188 40224 24200
rect 40083 24160 40224 24188
rect 40083 24157 40095 24160
rect 40037 24151 40095 24157
rect 40218 24148 40224 24160
rect 40276 24148 40282 24200
rect 35584 24092 37964 24120
rect 35584 24080 35590 24092
rect 38286 24080 38292 24132
rect 38344 24120 38350 24132
rect 40681 24123 40739 24129
rect 40681 24120 40693 24123
rect 38344 24092 40693 24120
rect 38344 24080 38350 24092
rect 40681 24089 40693 24092
rect 40727 24089 40739 24123
rect 40681 24083 40739 24089
rect 35342 24052 35348 24064
rect 35268 24024 35348 24052
rect 35342 24012 35348 24024
rect 35400 24012 35406 24064
rect 36078 24012 36084 24064
rect 36136 24012 36142 24064
rect 36170 24012 36176 24064
rect 36228 24052 36234 24064
rect 36449 24055 36507 24061
rect 36449 24052 36461 24055
rect 36228 24024 36461 24052
rect 36228 24012 36234 24024
rect 36449 24021 36461 24024
rect 36495 24021 36507 24055
rect 36449 24015 36507 24021
rect 37461 24055 37519 24061
rect 37461 24021 37473 24055
rect 37507 24052 37519 24055
rect 39942 24052 39948 24064
rect 37507 24024 39948 24052
rect 37507 24021 37519 24024
rect 37461 24015 37519 24021
rect 39942 24012 39948 24024
rect 40000 24012 40006 24064
rect 40788 24052 40816 24228
rect 41138 24216 41144 24268
rect 41196 24216 41202 24268
rect 41414 24216 41420 24268
rect 41472 24216 41478 24268
rect 45462 24216 45468 24268
rect 45520 24216 45526 24268
rect 46290 24216 46296 24268
rect 46348 24256 46354 24268
rect 47228 24256 47256 24284
rect 46348 24228 47900 24256
rect 46348 24216 46354 24228
rect 45186 24148 45192 24200
rect 45244 24148 45250 24200
rect 47872 24197 47900 24228
rect 48222 24216 48228 24268
rect 48280 24256 48286 24268
rect 48501 24259 48559 24265
rect 48501 24256 48513 24259
rect 48280 24228 48513 24256
rect 48280 24216 48286 24228
rect 48501 24225 48513 24228
rect 48547 24225 48559 24259
rect 48501 24219 48559 24225
rect 48774 24216 48780 24268
rect 48832 24216 48838 24268
rect 47213 24191 47271 24197
rect 47213 24188 47225 24191
rect 45480 24160 47225 24188
rect 42150 24080 42156 24132
rect 42208 24120 42214 24132
rect 42613 24123 42671 24129
rect 42613 24120 42625 24123
rect 42208 24092 42625 24120
rect 42208 24080 42214 24092
rect 42613 24089 42625 24092
rect 42659 24120 42671 24123
rect 45480 24120 45508 24160
rect 47213 24157 47225 24160
rect 47259 24157 47271 24191
rect 47213 24151 47271 24157
rect 47857 24191 47915 24197
rect 47857 24157 47869 24191
rect 47903 24157 47915 24191
rect 47857 24151 47915 24157
rect 42659 24092 45508 24120
rect 46569 24123 46627 24129
rect 42659 24089 42671 24092
rect 42613 24083 42671 24089
rect 46569 24089 46581 24123
rect 46615 24120 46627 24123
rect 46750 24120 46756 24132
rect 46615 24092 46756 24120
rect 46615 24089 46627 24092
rect 46569 24083 46627 24089
rect 41782 24052 41788 24064
rect 40788 24024 41788 24052
rect 41782 24012 41788 24024
rect 41840 24052 41846 24064
rect 42426 24052 42432 24064
rect 41840 24024 42432 24052
rect 41840 24012 41846 24024
rect 42426 24012 42432 24024
rect 42484 24012 42490 24064
rect 44085 24055 44143 24061
rect 44085 24021 44097 24055
rect 44131 24052 44143 24055
rect 44174 24052 44180 24064
rect 44131 24024 44180 24052
rect 44131 24021 44143 24024
rect 44085 24015 44143 24021
rect 44174 24012 44180 24024
rect 44232 24012 44238 24064
rect 44726 24012 44732 24064
rect 44784 24012 44790 24064
rect 45002 24012 45008 24064
rect 45060 24052 45066 24064
rect 46584 24052 46612 24083
rect 46750 24080 46756 24092
rect 46808 24080 46814 24132
rect 47118 24080 47124 24132
rect 47176 24120 47182 24132
rect 48240 24120 48268 24216
rect 47176 24092 48268 24120
rect 47176 24080 47182 24092
rect 45060 24024 46612 24052
rect 45060 24012 45066 24024
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 1854 23808 1860 23860
rect 1912 23848 1918 23860
rect 15562 23848 15568 23860
rect 1912 23820 15568 23848
rect 1912 23808 1918 23820
rect 15562 23808 15568 23820
rect 15620 23808 15626 23860
rect 19702 23848 19708 23860
rect 17144 23820 19708 23848
rect 1765 23783 1823 23789
rect 1765 23749 1777 23783
rect 1811 23780 1823 23783
rect 2130 23780 2136 23792
rect 1811 23752 2136 23780
rect 1811 23749 1823 23752
rect 1765 23743 1823 23749
rect 2130 23740 2136 23752
rect 2188 23740 2194 23792
rect 3970 23740 3976 23792
rect 4028 23780 4034 23792
rect 9125 23783 9183 23789
rect 4028 23752 7972 23780
rect 4028 23740 4034 23752
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23712 3019 23715
rect 3326 23712 3332 23724
rect 3007 23684 3332 23712
rect 3007 23681 3019 23684
rect 2961 23675 3019 23681
rect 3326 23672 3332 23684
rect 3384 23672 3390 23724
rect 4798 23672 4804 23724
rect 4856 23672 4862 23724
rect 6822 23672 6828 23724
rect 6880 23672 6886 23724
rect 7944 23721 7972 23752
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 9306 23780 9312 23792
rect 9171 23752 9312 23780
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 9306 23740 9312 23752
rect 9364 23740 9370 23792
rect 10686 23740 10692 23792
rect 10744 23740 10750 23792
rect 10778 23740 10784 23792
rect 10836 23780 10842 23792
rect 14277 23783 14335 23789
rect 10836 23752 11928 23780
rect 10836 23740 10842 23752
rect 7929 23715 7987 23721
rect 7929 23681 7941 23715
rect 7975 23681 7987 23715
rect 7929 23675 7987 23681
rect 9953 23715 10011 23721
rect 9953 23681 9965 23715
rect 9999 23712 10011 23715
rect 10042 23712 10048 23724
rect 9999 23684 10048 23712
rect 9999 23681 10011 23684
rect 9953 23675 10011 23681
rect 10042 23672 10048 23684
rect 10100 23672 10106 23724
rect 11790 23672 11796 23724
rect 11848 23672 11854 23724
rect 3973 23647 4031 23653
rect 3973 23613 3985 23647
rect 4019 23644 4031 23647
rect 4154 23644 4160 23656
rect 4019 23616 4160 23644
rect 4019 23613 4031 23616
rect 3973 23607 4031 23613
rect 4154 23604 4160 23616
rect 4212 23604 4218 23656
rect 5442 23604 5448 23656
rect 5500 23604 5506 23656
rect 9122 23644 9128 23656
rect 5552 23616 9128 23644
rect 2317 23579 2375 23585
rect 2317 23545 2329 23579
rect 2363 23576 2375 23579
rect 5552 23576 5580 23616
rect 9122 23604 9128 23616
rect 9180 23604 9186 23656
rect 11808 23644 11836 23672
rect 9600 23616 11836 23644
rect 11900 23644 11928 23752
rect 14277 23749 14289 23783
rect 14323 23780 14335 23783
rect 14734 23780 14740 23792
rect 14323 23752 14740 23780
rect 14323 23749 14335 23752
rect 14277 23743 14335 23749
rect 14734 23740 14740 23752
rect 14792 23740 14798 23792
rect 15286 23780 15292 23792
rect 14936 23752 15292 23780
rect 12066 23672 12072 23724
rect 12124 23672 12130 23724
rect 14936 23721 14964 23752
rect 15286 23740 15292 23752
rect 15344 23740 15350 23792
rect 16117 23783 16175 23789
rect 16117 23749 16129 23783
rect 16163 23780 16175 23783
rect 17034 23780 17040 23792
rect 16163 23752 17040 23780
rect 16163 23749 16175 23752
rect 16117 23743 16175 23749
rect 17034 23740 17040 23752
rect 17092 23740 17098 23792
rect 17144 23721 17172 23820
rect 19702 23808 19708 23820
rect 19760 23808 19766 23860
rect 20530 23808 20536 23860
rect 20588 23808 20594 23860
rect 20901 23851 20959 23857
rect 20901 23817 20913 23851
rect 20947 23848 20959 23851
rect 22278 23848 22284 23860
rect 20947 23820 22284 23848
rect 20947 23817 20959 23820
rect 20901 23811 20959 23817
rect 22278 23808 22284 23820
rect 22336 23808 22342 23860
rect 22370 23808 22376 23860
rect 22428 23808 22434 23860
rect 22462 23808 22468 23860
rect 22520 23808 22526 23860
rect 23477 23851 23535 23857
rect 23477 23817 23489 23851
rect 23523 23848 23535 23851
rect 23566 23848 23572 23860
rect 23523 23820 23572 23848
rect 23523 23817 23535 23820
rect 23477 23811 23535 23817
rect 23566 23808 23572 23820
rect 23624 23848 23630 23860
rect 24670 23848 24676 23860
rect 23624 23820 24676 23848
rect 23624 23808 23630 23820
rect 24670 23808 24676 23820
rect 24728 23808 24734 23860
rect 26786 23848 26792 23860
rect 25148 23820 26792 23848
rect 18141 23783 18199 23789
rect 18141 23749 18153 23783
rect 18187 23780 18199 23783
rect 18966 23780 18972 23792
rect 18187 23752 18972 23780
rect 18187 23749 18199 23752
rect 18141 23743 18199 23749
rect 18966 23740 18972 23752
rect 19024 23740 19030 23792
rect 20346 23780 20352 23792
rect 20286 23752 20352 23780
rect 20346 23740 20352 23752
rect 20404 23740 20410 23792
rect 20990 23740 20996 23792
rect 21048 23780 21054 23792
rect 21266 23780 21272 23792
rect 21048 23752 21272 23780
rect 21048 23740 21054 23752
rect 21266 23740 21272 23752
rect 21324 23740 21330 23792
rect 21634 23740 21640 23792
rect 21692 23780 21698 23792
rect 25148 23789 25176 23820
rect 26786 23808 26792 23820
rect 26844 23808 26850 23860
rect 29362 23808 29368 23860
rect 29420 23808 29426 23860
rect 32309 23851 32367 23857
rect 32309 23848 32321 23851
rect 29472 23820 32321 23848
rect 24397 23783 24455 23789
rect 24397 23780 24409 23783
rect 21692 23752 24409 23780
rect 21692 23740 21698 23752
rect 24397 23749 24409 23752
rect 24443 23749 24455 23783
rect 24397 23743 24455 23749
rect 25133 23783 25191 23789
rect 25133 23749 25145 23783
rect 25179 23749 25191 23783
rect 26510 23780 26516 23792
rect 26358 23752 26516 23780
rect 25133 23743 25191 23749
rect 26510 23740 26516 23752
rect 26568 23740 26574 23792
rect 28534 23740 28540 23792
rect 28592 23780 28598 23792
rect 29472 23780 29500 23820
rect 32309 23817 32321 23820
rect 32355 23817 32367 23851
rect 35253 23851 35311 23857
rect 35253 23848 35265 23851
rect 32309 23811 32367 23817
rect 32968 23820 35265 23848
rect 30558 23780 30564 23792
rect 28592 23752 29500 23780
rect 29564 23752 30564 23780
rect 28592 23740 28598 23752
rect 13265 23715 13323 23721
rect 13265 23681 13277 23715
rect 13311 23712 13323 23715
rect 14921 23715 14979 23721
rect 13311 23684 14872 23712
rect 13311 23681 13323 23684
rect 13265 23675 13323 23681
rect 14734 23644 14740 23656
rect 11900 23616 14740 23644
rect 2363 23548 5580 23576
rect 6549 23579 6607 23585
rect 2363 23545 2375 23548
rect 2317 23539 2375 23545
rect 6549 23545 6561 23579
rect 6595 23576 6607 23579
rect 9600 23576 9628 23616
rect 14734 23604 14740 23616
rect 14792 23604 14798 23656
rect 14844 23644 14872 23684
rect 14921 23681 14933 23715
rect 14967 23681 14979 23715
rect 17129 23715 17187 23721
rect 14921 23675 14979 23681
rect 15028 23684 16896 23712
rect 15028 23644 15056 23684
rect 16758 23644 16764 23656
rect 14844 23616 15056 23644
rect 15212 23616 16764 23644
rect 6595 23548 9628 23576
rect 6595 23545 6607 23548
rect 6549 23539 6607 23545
rect 9674 23536 9680 23588
rect 9732 23576 9738 23588
rect 15212 23576 15240 23616
rect 16758 23604 16764 23616
rect 16816 23604 16822 23656
rect 16868 23644 16896 23684
rect 17129 23681 17141 23715
rect 17175 23681 17187 23715
rect 17129 23675 17187 23681
rect 17218 23672 17224 23724
rect 17276 23712 17282 23724
rect 17276 23684 18460 23712
rect 17276 23672 17282 23684
rect 18322 23644 18328 23656
rect 16868 23616 18328 23644
rect 18322 23604 18328 23616
rect 18380 23604 18386 23656
rect 18432 23644 18460 23684
rect 18782 23672 18788 23724
rect 18840 23672 18846 23724
rect 23787 23715 23845 23721
rect 23787 23681 23799 23715
rect 23833 23712 23845 23715
rect 24118 23712 24124 23724
rect 23833 23684 24124 23712
rect 23833 23681 23845 23684
rect 23787 23675 23845 23681
rect 24118 23672 24124 23684
rect 24176 23672 24182 23724
rect 27157 23715 27215 23721
rect 27157 23681 27169 23715
rect 27203 23712 27215 23715
rect 27430 23712 27436 23724
rect 27203 23684 27436 23712
rect 27203 23681 27215 23684
rect 27157 23675 27215 23681
rect 27430 23672 27436 23684
rect 27488 23672 27494 23724
rect 28166 23672 28172 23724
rect 28224 23712 28230 23724
rect 29564 23721 29592 23752
rect 30558 23740 30564 23752
rect 30616 23740 30622 23792
rect 30926 23740 30932 23792
rect 30984 23740 30990 23792
rect 28261 23715 28319 23721
rect 28261 23712 28273 23715
rect 28224 23684 28273 23712
rect 28224 23672 28230 23684
rect 28261 23681 28273 23684
rect 28307 23681 28319 23715
rect 28261 23675 28319 23681
rect 29549 23715 29607 23721
rect 29549 23681 29561 23715
rect 29595 23681 29607 23715
rect 29549 23675 29607 23681
rect 32674 23672 32680 23724
rect 32732 23672 32738 23724
rect 19061 23647 19119 23653
rect 19061 23644 19073 23647
rect 18432 23616 19073 23644
rect 19061 23613 19073 23616
rect 19107 23613 19119 23647
rect 19061 23607 19119 23613
rect 19150 23604 19156 23656
rect 19208 23644 19214 23656
rect 19208 23616 22048 23644
rect 19208 23604 19214 23616
rect 9732 23548 15240 23576
rect 9732 23536 9738 23548
rect 15286 23536 15292 23588
rect 15344 23576 15350 23588
rect 22020 23585 22048 23616
rect 22554 23604 22560 23656
rect 22612 23604 22618 23656
rect 23109 23647 23167 23653
rect 23109 23613 23121 23647
rect 23155 23644 23167 23647
rect 23658 23644 23664 23656
rect 23155 23616 23664 23644
rect 23155 23613 23167 23616
rect 23109 23607 23167 23613
rect 23658 23604 23664 23616
rect 23716 23604 23722 23656
rect 24854 23604 24860 23656
rect 24912 23604 24918 23656
rect 29730 23604 29736 23656
rect 29788 23644 29794 23656
rect 30009 23647 30067 23653
rect 30009 23644 30021 23647
rect 29788 23616 30021 23644
rect 29788 23604 29794 23616
rect 30009 23613 30021 23616
rect 30055 23613 30067 23647
rect 30285 23647 30343 23653
rect 30285 23644 30297 23647
rect 30009 23607 30067 23613
rect 30116 23616 30297 23644
rect 21453 23579 21511 23585
rect 21453 23576 21465 23579
rect 15344 23548 18552 23576
rect 15344 23536 15350 23548
rect 3418 23468 3424 23520
rect 3476 23508 3482 23520
rect 6638 23508 6644 23520
rect 3476 23480 6644 23508
rect 3476 23468 3482 23480
rect 6638 23468 6644 23480
rect 6696 23468 6702 23520
rect 7469 23511 7527 23517
rect 7469 23477 7481 23511
rect 7515 23508 7527 23511
rect 17218 23508 17224 23520
rect 7515 23480 17224 23508
rect 7515 23477 7527 23480
rect 7469 23471 7527 23477
rect 17218 23468 17224 23480
rect 17276 23468 17282 23520
rect 18524 23508 18552 23548
rect 20088 23548 21465 23576
rect 20088 23508 20116 23548
rect 21453 23545 21465 23548
rect 21499 23545 21511 23579
rect 21453 23539 21511 23545
rect 22005 23579 22063 23585
rect 22005 23545 22017 23579
rect 22051 23545 22063 23579
rect 28905 23579 28963 23585
rect 28905 23576 28917 23579
rect 22005 23539 22063 23545
rect 22112 23548 23428 23576
rect 18524 23480 20116 23508
rect 20622 23468 20628 23520
rect 20680 23508 20686 23520
rect 22112 23508 22140 23548
rect 20680 23480 22140 23508
rect 20680 23468 20686 23480
rect 23290 23468 23296 23520
rect 23348 23468 23354 23520
rect 23400 23508 23428 23548
rect 26160 23548 28917 23576
rect 26160 23508 26188 23548
rect 28905 23545 28917 23548
rect 28951 23545 28963 23579
rect 28905 23539 28963 23545
rect 28994 23536 29000 23588
rect 29052 23576 29058 23588
rect 30116 23576 30144 23616
rect 30285 23613 30297 23616
rect 30331 23644 30343 23647
rect 32582 23644 32588 23656
rect 30331 23616 32588 23644
rect 30331 23613 30343 23616
rect 30285 23607 30343 23613
rect 32582 23604 32588 23616
rect 32640 23604 32646 23656
rect 32968 23653 32996 23820
rect 35253 23817 35265 23820
rect 35299 23848 35311 23851
rect 35526 23848 35532 23860
rect 35299 23820 35532 23848
rect 35299 23817 35311 23820
rect 35253 23811 35311 23817
rect 35526 23808 35532 23820
rect 35584 23808 35590 23860
rect 35618 23808 35624 23860
rect 35676 23848 35682 23860
rect 35986 23848 35992 23860
rect 35676 23820 35992 23848
rect 35676 23808 35682 23820
rect 35986 23808 35992 23820
rect 36044 23808 36050 23860
rect 36265 23851 36323 23857
rect 36265 23817 36277 23851
rect 36311 23848 36323 23851
rect 38841 23851 38899 23857
rect 38841 23848 38853 23851
rect 36311 23820 38853 23848
rect 36311 23817 36323 23820
rect 36265 23811 36323 23817
rect 38841 23817 38853 23820
rect 38887 23817 38899 23851
rect 38841 23811 38899 23817
rect 38930 23808 38936 23860
rect 38988 23848 38994 23860
rect 38988 23820 42656 23848
rect 38988 23808 38994 23820
rect 33778 23740 33784 23792
rect 33836 23740 33842 23792
rect 34238 23740 34244 23792
rect 34296 23740 34302 23792
rect 35158 23740 35164 23792
rect 35216 23780 35222 23792
rect 37921 23783 37979 23789
rect 37921 23780 37933 23783
rect 35216 23752 37933 23780
rect 35216 23740 35222 23752
rect 37921 23749 37933 23752
rect 37967 23749 37979 23783
rect 37921 23743 37979 23749
rect 38562 23740 38568 23792
rect 38620 23780 38626 23792
rect 40681 23783 40739 23789
rect 40681 23780 40693 23783
rect 38620 23752 40693 23780
rect 38620 23740 38626 23752
rect 40681 23749 40693 23752
rect 40727 23749 40739 23783
rect 40681 23743 40739 23749
rect 40788 23752 41460 23780
rect 35526 23672 35532 23724
rect 35584 23712 35590 23724
rect 37829 23715 37887 23721
rect 35584 23684 36584 23712
rect 35584 23672 35590 23684
rect 32769 23647 32827 23653
rect 32769 23613 32781 23647
rect 32815 23613 32827 23647
rect 32769 23607 32827 23613
rect 32953 23647 33011 23653
rect 32953 23613 32965 23647
rect 32999 23613 33011 23647
rect 32953 23607 33011 23613
rect 29052 23548 30144 23576
rect 29052 23536 29058 23548
rect 23400 23480 26188 23508
rect 26602 23468 26608 23520
rect 26660 23508 26666 23520
rect 27522 23508 27528 23520
rect 26660 23480 27528 23508
rect 26660 23468 26666 23480
rect 27522 23468 27528 23480
rect 27580 23468 27586 23520
rect 27798 23468 27804 23520
rect 27856 23468 27862 23520
rect 30282 23468 30288 23520
rect 30340 23508 30346 23520
rect 31757 23511 31815 23517
rect 31757 23508 31769 23511
rect 30340 23480 31769 23508
rect 30340 23468 30346 23480
rect 31757 23477 31769 23480
rect 31803 23477 31815 23511
rect 32784 23508 32812 23607
rect 33502 23604 33508 23656
rect 33560 23604 33566 23656
rect 35158 23604 35164 23656
rect 35216 23644 35222 23656
rect 36357 23647 36415 23653
rect 36357 23644 36369 23647
rect 35216 23616 36369 23644
rect 35216 23604 35222 23616
rect 36357 23613 36369 23616
rect 36403 23613 36415 23647
rect 36357 23607 36415 23613
rect 36446 23604 36452 23656
rect 36504 23604 36510 23656
rect 36556 23644 36584 23684
rect 37829 23681 37841 23715
rect 37875 23712 37887 23715
rect 39209 23715 39267 23721
rect 37875 23684 39160 23712
rect 37875 23681 37887 23684
rect 37829 23675 37887 23681
rect 38013 23647 38071 23653
rect 38013 23644 38025 23647
rect 36556 23616 38025 23644
rect 38013 23613 38025 23616
rect 38059 23613 38071 23647
rect 38013 23607 38071 23613
rect 37461 23579 37519 23585
rect 37461 23576 37473 23579
rect 35176 23548 36400 23576
rect 35176 23508 35204 23548
rect 32784 23480 35204 23508
rect 31757 23471 31815 23477
rect 35342 23468 35348 23520
rect 35400 23508 35406 23520
rect 35618 23508 35624 23520
rect 35400 23480 35624 23508
rect 35400 23468 35406 23480
rect 35618 23468 35624 23480
rect 35676 23468 35682 23520
rect 35897 23511 35955 23517
rect 35897 23477 35909 23511
rect 35943 23508 35955 23511
rect 36262 23508 36268 23520
rect 35943 23480 36268 23508
rect 35943 23477 35955 23480
rect 35897 23471 35955 23477
rect 36262 23468 36268 23480
rect 36320 23468 36326 23520
rect 36372 23508 36400 23548
rect 36648 23548 37473 23576
rect 36648 23508 36676 23548
rect 37461 23545 37473 23548
rect 37507 23545 37519 23579
rect 37461 23539 37519 23545
rect 36372 23480 36676 23508
rect 36906 23468 36912 23520
rect 36964 23508 36970 23520
rect 38473 23511 38531 23517
rect 38473 23508 38485 23511
rect 36964 23480 38485 23508
rect 36964 23468 36970 23480
rect 38473 23477 38485 23480
rect 38519 23477 38531 23511
rect 39132 23508 39160 23684
rect 39209 23681 39221 23715
rect 39255 23681 39267 23715
rect 39209 23675 39267 23681
rect 39301 23715 39359 23721
rect 39301 23681 39313 23715
rect 39347 23712 39359 23715
rect 39482 23712 39488 23724
rect 39347 23684 39488 23712
rect 39347 23681 39359 23684
rect 39301 23675 39359 23681
rect 39224 23576 39252 23675
rect 39482 23672 39488 23684
rect 39540 23672 39546 23724
rect 39758 23672 39764 23724
rect 39816 23712 39822 23724
rect 40037 23715 40095 23721
rect 40037 23712 40049 23715
rect 39816 23684 40049 23712
rect 39816 23672 39822 23684
rect 40037 23681 40049 23684
rect 40083 23681 40095 23715
rect 40037 23675 40095 23681
rect 39390 23604 39396 23656
rect 39448 23604 39454 23656
rect 39850 23604 39856 23656
rect 39908 23644 39914 23656
rect 40788 23644 40816 23752
rect 41432 23721 41460 23752
rect 42628 23721 42656 23820
rect 44726 23808 44732 23860
rect 44784 23848 44790 23860
rect 47949 23851 48007 23857
rect 47949 23848 47961 23851
rect 44784 23820 47961 23848
rect 44784 23808 44790 23820
rect 47949 23817 47961 23820
rect 47995 23817 48007 23851
rect 47949 23811 48007 23817
rect 45094 23740 45100 23792
rect 45152 23780 45158 23792
rect 45152 23752 46612 23780
rect 45152 23740 45158 23752
rect 41417 23715 41475 23721
rect 41417 23681 41429 23715
rect 41463 23681 41475 23715
rect 41417 23675 41475 23681
rect 42613 23715 42671 23721
rect 42613 23681 42625 23715
rect 42659 23681 42671 23715
rect 42613 23675 42671 23681
rect 42794 23672 42800 23724
rect 42852 23712 42858 23724
rect 44177 23715 44235 23721
rect 44177 23712 44189 23715
rect 42852 23684 44189 23712
rect 42852 23672 42858 23684
rect 44177 23681 44189 23684
rect 44223 23681 44235 23715
rect 44177 23675 44235 23681
rect 44266 23672 44272 23724
rect 44324 23712 44330 23724
rect 45465 23715 45523 23721
rect 45465 23712 45477 23715
rect 44324 23684 45477 23712
rect 44324 23672 44330 23684
rect 45465 23681 45477 23684
rect 45511 23681 45523 23715
rect 45465 23675 45523 23681
rect 45554 23672 45560 23724
rect 45612 23712 45618 23724
rect 46198 23712 46204 23724
rect 45612 23684 46204 23712
rect 45612 23672 45618 23684
rect 46198 23672 46204 23684
rect 46256 23712 46262 23724
rect 46477 23715 46535 23721
rect 46477 23712 46489 23715
rect 46256 23684 46489 23712
rect 46256 23672 46262 23684
rect 46477 23681 46489 23684
rect 46523 23681 46535 23715
rect 46584 23712 46612 23752
rect 46934 23740 46940 23792
rect 46992 23780 46998 23792
rect 47486 23780 47492 23792
rect 46992 23752 47492 23780
rect 46992 23740 46998 23752
rect 47486 23740 47492 23752
rect 47544 23780 47550 23792
rect 47857 23783 47915 23789
rect 47857 23780 47869 23783
rect 47544 23752 47869 23780
rect 47544 23740 47550 23752
rect 47857 23749 47869 23752
rect 47903 23749 47915 23783
rect 47857 23743 47915 23749
rect 46584 23684 47348 23712
rect 46477 23675 46535 23681
rect 39908 23616 40816 23644
rect 39908 23604 39914 23616
rect 41138 23604 41144 23656
rect 41196 23604 41202 23656
rect 42886 23604 42892 23656
rect 42944 23604 42950 23656
rect 43898 23604 43904 23656
rect 43956 23604 43962 23656
rect 45094 23604 45100 23656
rect 45152 23644 45158 23656
rect 45189 23647 45247 23653
rect 45189 23644 45201 23647
rect 45152 23616 45201 23644
rect 45152 23604 45158 23616
rect 45189 23613 45201 23616
rect 45235 23613 45247 23647
rect 47213 23647 47271 23653
rect 47213 23644 47225 23647
rect 45189 23607 45247 23613
rect 45296 23616 47225 23644
rect 43806 23576 43812 23588
rect 39224 23548 43812 23576
rect 43806 23536 43812 23548
rect 43864 23536 43870 23588
rect 43916 23576 43944 23604
rect 45296 23576 45324 23616
rect 47213 23613 47225 23616
rect 47259 23613 47271 23647
rect 47320 23644 47348 23684
rect 47946 23672 47952 23724
rect 48004 23712 48010 23724
rect 48501 23715 48559 23721
rect 48501 23712 48513 23715
rect 48004 23684 48513 23712
rect 48004 23672 48010 23684
rect 48501 23681 48513 23684
rect 48547 23681 48559 23715
rect 48501 23675 48559 23681
rect 49237 23647 49295 23653
rect 49237 23644 49249 23647
rect 47320 23616 49249 23644
rect 47213 23607 47271 23613
rect 49237 23613 49249 23616
rect 49283 23613 49295 23647
rect 49237 23607 49295 23613
rect 43916 23548 45324 23576
rect 45554 23536 45560 23588
rect 45612 23576 45618 23588
rect 49421 23579 49479 23585
rect 49421 23576 49433 23579
rect 45612 23548 49433 23576
rect 45612 23536 45618 23548
rect 49421 23545 49433 23548
rect 49467 23545 49479 23579
rect 49421 23539 49479 23545
rect 40034 23508 40040 23520
rect 39132 23480 40040 23508
rect 38473 23471 38531 23477
rect 40034 23468 40040 23480
rect 40092 23468 40098 23520
rect 40126 23468 40132 23520
rect 40184 23508 40190 23520
rect 41874 23508 41880 23520
rect 40184 23480 41880 23508
rect 40184 23468 40190 23480
rect 41874 23468 41880 23480
rect 41932 23468 41938 23520
rect 41966 23468 41972 23520
rect 42024 23508 42030 23520
rect 46661 23511 46719 23517
rect 46661 23508 46673 23511
rect 42024 23480 46673 23508
rect 42024 23468 42030 23480
rect 46661 23477 46673 23480
rect 46707 23477 46719 23511
rect 46661 23471 46719 23477
rect 47121 23511 47179 23517
rect 47121 23477 47133 23511
rect 47167 23508 47179 23511
rect 47578 23508 47584 23520
rect 47167 23480 47584 23508
rect 47167 23477 47179 23480
rect 47121 23471 47179 23477
rect 47578 23468 47584 23480
rect 47636 23508 47642 23520
rect 48685 23511 48743 23517
rect 48685 23508 48697 23511
rect 47636 23480 48697 23508
rect 47636 23468 47642 23480
rect 48685 23477 48697 23480
rect 48731 23477 48743 23511
rect 48685 23471 48743 23477
rect 49050 23468 49056 23520
rect 49108 23468 49114 23520
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 3605 23307 3663 23313
rect 3605 23273 3617 23307
rect 3651 23304 3663 23307
rect 6822 23304 6828 23316
rect 3651 23276 6828 23304
rect 3651 23273 3663 23276
rect 3605 23267 3663 23273
rect 6822 23264 6828 23276
rect 6880 23264 6886 23316
rect 13262 23264 13268 23316
rect 13320 23304 13326 23316
rect 17126 23304 17132 23316
rect 13320 23276 17132 23304
rect 13320 23264 13326 23276
rect 17126 23264 17132 23276
rect 17184 23264 17190 23316
rect 17586 23264 17592 23316
rect 17644 23304 17650 23316
rect 19610 23304 19616 23316
rect 17644 23276 19616 23304
rect 17644 23264 17650 23276
rect 19610 23264 19616 23276
rect 19668 23264 19674 23316
rect 19702 23264 19708 23316
rect 19760 23264 19766 23316
rect 22554 23304 22560 23316
rect 19812 23276 22560 23304
rect 8570 23196 8576 23248
rect 8628 23236 8634 23248
rect 8628 23208 16528 23236
rect 8628 23196 8634 23208
rect 4249 23171 4307 23177
rect 4249 23137 4261 23171
rect 4295 23168 4307 23171
rect 5258 23168 5264 23180
rect 4295 23140 5264 23168
rect 4295 23137 4307 23140
rect 4249 23131 4307 23137
rect 5258 23128 5264 23140
rect 5316 23128 5322 23180
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 9398 23128 9404 23180
rect 9456 23128 9462 23180
rect 11238 23128 11244 23180
rect 11296 23128 11302 23180
rect 13354 23128 13360 23180
rect 13412 23128 13418 23180
rect 14274 23128 14280 23180
rect 14332 23168 14338 23180
rect 14550 23168 14556 23180
rect 14332 23140 14556 23168
rect 14332 23128 14338 23140
rect 14550 23128 14556 23140
rect 14608 23128 14614 23180
rect 16390 23128 16396 23180
rect 16448 23128 16454 23180
rect 16500 23168 16528 23208
rect 18598 23196 18604 23248
rect 18656 23236 18662 23248
rect 19812 23236 19840 23276
rect 22554 23264 22560 23276
rect 22612 23264 22618 23316
rect 27893 23307 27951 23313
rect 27893 23304 27905 23307
rect 23032 23276 27905 23304
rect 18656 23208 19840 23236
rect 18656 23196 18662 23208
rect 17405 23171 17463 23177
rect 17405 23168 17417 23171
rect 16500 23140 17417 23168
rect 17405 23137 17417 23140
rect 17451 23137 17463 23171
rect 17405 23131 17463 23137
rect 18782 23128 18788 23180
rect 18840 23168 18846 23180
rect 20349 23171 20407 23177
rect 20349 23168 20361 23171
rect 18840 23140 20361 23168
rect 18840 23128 18846 23140
rect 20349 23137 20361 23140
rect 20395 23168 20407 23171
rect 21174 23168 21180 23180
rect 20395 23140 21180 23168
rect 20395 23137 20407 23140
rect 20349 23131 20407 23137
rect 21174 23128 21180 23140
rect 21232 23128 21238 23180
rect 23032 23177 23060 23276
rect 27893 23273 27905 23276
rect 27939 23273 27951 23307
rect 27893 23267 27951 23273
rect 29733 23307 29791 23313
rect 29733 23273 29745 23307
rect 29779 23304 29791 23307
rect 29822 23304 29828 23316
rect 29779 23276 29828 23304
rect 29779 23273 29791 23276
rect 29733 23267 29791 23273
rect 29822 23264 29828 23276
rect 29880 23264 29886 23316
rect 33778 23264 33784 23316
rect 33836 23304 33842 23316
rect 35342 23304 35348 23316
rect 33836 23276 35348 23304
rect 33836 23264 33842 23276
rect 35342 23264 35348 23276
rect 35400 23264 35406 23316
rect 35802 23264 35808 23316
rect 35860 23304 35866 23316
rect 35860 23276 38516 23304
rect 35860 23264 35866 23276
rect 23382 23196 23388 23248
rect 23440 23236 23446 23248
rect 24029 23239 24087 23245
rect 24029 23236 24041 23239
rect 23440 23208 24041 23236
rect 23440 23196 23446 23208
rect 24029 23205 24041 23208
rect 24075 23205 24087 23239
rect 30006 23236 30012 23248
rect 24029 23199 24087 23205
rect 27080 23208 30012 23236
rect 23017 23171 23075 23177
rect 23017 23137 23029 23171
rect 23063 23137 23075 23171
rect 23017 23131 23075 23137
rect 23106 23128 23112 23180
rect 23164 23128 23170 23180
rect 23658 23168 23664 23180
rect 23308 23140 23664 23168
rect 1765 23103 1823 23109
rect 1765 23069 1777 23103
rect 1811 23100 1823 23103
rect 3421 23103 3479 23109
rect 1811 23072 3372 23100
rect 1811 23069 1823 23072
rect 1765 23063 1823 23069
rect 2774 22992 2780 23044
rect 2832 22992 2838 23044
rect 3344 23032 3372 23072
rect 3421 23069 3433 23103
rect 3467 23100 3479 23103
rect 3970 23100 3976 23112
rect 3467 23072 3976 23100
rect 3467 23069 3479 23072
rect 3421 23063 3479 23069
rect 3970 23060 3976 23072
rect 4028 23060 4034 23112
rect 4430 23060 4436 23112
rect 4488 23100 4494 23112
rect 5353 23103 5411 23109
rect 5353 23100 5365 23103
rect 4488 23072 5365 23100
rect 4488 23060 4494 23072
rect 5353 23069 5365 23072
rect 5399 23069 5411 23103
rect 5353 23063 5411 23069
rect 7098 23060 7104 23112
rect 7156 23100 7162 23112
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 7156 23072 7205 23100
rect 7156 23060 7162 23072
rect 7193 23069 7205 23072
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 9125 23103 9183 23109
rect 9125 23069 9137 23103
rect 9171 23100 9183 23103
rect 9214 23100 9220 23112
rect 9171 23072 9220 23100
rect 9171 23069 9183 23072
rect 9125 23063 9183 23069
rect 9214 23060 9220 23072
rect 9272 23060 9278 23112
rect 10689 23103 10747 23109
rect 10689 23069 10701 23103
rect 10735 23069 10747 23103
rect 10689 23063 10747 23069
rect 4338 23032 4344 23044
rect 3344 23004 4344 23032
rect 4338 22992 4344 23004
rect 4396 22992 4402 23044
rect 10704 23032 10732 23063
rect 12434 23060 12440 23112
rect 12492 23060 12498 23112
rect 15473 23103 15531 23109
rect 15473 23069 15485 23103
rect 15519 23100 15531 23103
rect 16666 23100 16672 23112
rect 15519 23072 16672 23100
rect 15519 23069 15531 23072
rect 15473 23063 15531 23069
rect 16666 23060 16672 23072
rect 16724 23060 16730 23112
rect 17126 23060 17132 23112
rect 17184 23060 17190 23112
rect 19886 23060 19892 23112
rect 19944 23060 19950 23112
rect 22002 23060 22008 23112
rect 22060 23100 22066 23112
rect 23308 23100 23336 23140
rect 23658 23128 23664 23140
rect 23716 23168 23722 23180
rect 25685 23171 25743 23177
rect 25685 23168 25697 23171
rect 23716 23140 25697 23168
rect 23716 23128 23722 23140
rect 25685 23137 25697 23140
rect 25731 23137 25743 23171
rect 25685 23131 25743 23137
rect 25958 23128 25964 23180
rect 26016 23128 26022 23180
rect 22060 23072 23336 23100
rect 22060 23060 22066 23072
rect 23842 23060 23848 23112
rect 23900 23060 23906 23112
rect 24581 23103 24639 23109
rect 24581 23069 24593 23103
rect 24627 23100 24639 23103
rect 25590 23100 25596 23112
rect 24627 23072 25596 23100
rect 24627 23069 24639 23072
rect 24581 23063 24639 23069
rect 25590 23060 25596 23072
rect 25648 23060 25654 23112
rect 26970 23060 26976 23112
rect 27028 23100 27034 23112
rect 27080 23100 27108 23208
rect 30006 23196 30012 23208
rect 30064 23236 30070 23248
rect 30926 23236 30932 23248
rect 30064 23208 30932 23236
rect 30064 23196 30070 23208
rect 30926 23196 30932 23208
rect 30984 23196 30990 23248
rect 38488 23236 38516 23276
rect 38746 23264 38752 23316
rect 38804 23304 38810 23316
rect 38933 23307 38991 23313
rect 38933 23304 38945 23307
rect 38804 23276 38945 23304
rect 38804 23264 38810 23276
rect 38933 23273 38945 23276
rect 38979 23304 38991 23307
rect 39758 23304 39764 23316
rect 38979 23276 39764 23304
rect 38979 23273 38991 23276
rect 38933 23267 38991 23273
rect 39758 23264 39764 23276
rect 39816 23264 39822 23316
rect 40034 23264 40040 23316
rect 40092 23264 40098 23316
rect 41046 23264 41052 23316
rect 41104 23264 41110 23316
rect 43254 23264 43260 23316
rect 43312 23304 43318 23316
rect 43530 23304 43536 23316
rect 43312 23276 43536 23304
rect 43312 23264 43318 23276
rect 43530 23264 43536 23276
rect 43588 23264 43594 23316
rect 43898 23304 43904 23316
rect 43732 23276 43904 23304
rect 39390 23236 39396 23248
rect 38488 23208 39396 23236
rect 39390 23196 39396 23208
rect 39448 23196 39454 23248
rect 39482 23196 39488 23248
rect 39540 23236 39546 23248
rect 39669 23239 39727 23245
rect 39669 23236 39681 23239
rect 39540 23208 39681 23236
rect 39540 23196 39546 23208
rect 39669 23205 39681 23208
rect 39715 23236 39727 23239
rect 40126 23236 40132 23248
rect 39715 23208 40132 23236
rect 39715 23205 39727 23208
rect 39669 23199 39727 23205
rect 40126 23196 40132 23208
rect 40184 23196 40190 23248
rect 40402 23196 40408 23248
rect 40460 23196 40466 23248
rect 42886 23196 42892 23248
rect 42944 23236 42950 23248
rect 43622 23236 43628 23248
rect 42944 23208 43628 23236
rect 42944 23196 42950 23208
rect 43622 23196 43628 23208
rect 43680 23196 43686 23248
rect 27614 23128 27620 23180
rect 27672 23168 27678 23180
rect 28350 23168 28356 23180
rect 27672 23140 28356 23168
rect 27672 23128 27678 23140
rect 28350 23128 28356 23140
rect 28408 23128 28414 23180
rect 28445 23171 28503 23177
rect 28445 23137 28457 23171
rect 28491 23137 28503 23171
rect 28445 23131 28503 23137
rect 27028 23086 27108 23100
rect 27028 23072 27094 23086
rect 27028 23060 27034 23072
rect 14090 23032 14096 23044
rect 10704 23004 14096 23032
rect 14090 22992 14096 23004
rect 14148 22992 14154 23044
rect 14642 22992 14648 23044
rect 14700 22992 14706 23044
rect 14829 23035 14887 23041
rect 14829 23001 14841 23035
rect 14875 23032 14887 23035
rect 17494 23032 17500 23044
rect 14875 23004 17500 23032
rect 14875 23001 14887 23004
rect 14829 22995 14887 23001
rect 17494 22992 17500 23004
rect 17552 22992 17558 23044
rect 18414 22992 18420 23044
rect 18472 22992 18478 23044
rect 19429 23035 19487 23041
rect 19429 23001 19441 23035
rect 19475 23032 19487 23035
rect 19475 23004 20576 23032
rect 19475 23001 19487 23004
rect 19429 22995 19487 23001
rect 14274 22924 14280 22976
rect 14332 22964 14338 22976
rect 17586 22964 17592 22976
rect 14332 22936 17592 22964
rect 14332 22924 14338 22936
rect 17586 22924 17592 22936
rect 17644 22924 17650 22976
rect 17770 22924 17776 22976
rect 17828 22964 17834 22976
rect 18877 22967 18935 22973
rect 18877 22964 18889 22967
rect 17828 22936 18889 22964
rect 17828 22924 17834 22936
rect 18877 22933 18889 22936
rect 18923 22933 18935 22967
rect 20548 22964 20576 23004
rect 20622 22992 20628 23044
rect 20680 22992 20686 23044
rect 20714 22992 20720 23044
rect 20772 23032 20778 23044
rect 21082 23032 21088 23044
rect 20772 23004 21088 23032
rect 20772 22992 20778 23004
rect 21082 22992 21088 23004
rect 21140 22992 21146 23044
rect 24026 23032 24032 23044
rect 21928 23004 24032 23032
rect 21928 22964 21956 23004
rect 24026 22992 24032 23004
rect 24084 22992 24090 23044
rect 24210 22992 24216 23044
rect 24268 23032 24274 23044
rect 28166 23032 28172 23044
rect 24268 23004 26372 23032
rect 24268 22992 24274 23004
rect 20548 22936 21956 22964
rect 18877 22927 18935 22933
rect 22094 22924 22100 22976
rect 22152 22924 22158 22976
rect 22462 22924 22468 22976
rect 22520 22964 22526 22976
rect 22557 22967 22615 22973
rect 22557 22964 22569 22967
rect 22520 22936 22569 22964
rect 22520 22924 22526 22936
rect 22557 22933 22569 22936
rect 22603 22933 22615 22967
rect 22557 22927 22615 22933
rect 22925 22967 22983 22973
rect 22925 22933 22937 22967
rect 22971 22964 22983 22967
rect 23750 22964 23756 22976
rect 22971 22936 23756 22964
rect 22971 22933 22983 22936
rect 22925 22927 22983 22933
rect 23750 22924 23756 22936
rect 23808 22924 23814 22976
rect 25225 22967 25283 22973
rect 25225 22933 25237 22967
rect 25271 22964 25283 22967
rect 25314 22964 25320 22976
rect 25271 22936 25320 22964
rect 25271 22933 25283 22936
rect 25225 22927 25283 22933
rect 25314 22924 25320 22936
rect 25372 22924 25378 22976
rect 26344 22964 26372 23004
rect 27356 23004 28172 23032
rect 27356 22964 27384 23004
rect 28166 22992 28172 23004
rect 28224 23032 28230 23044
rect 28460 23032 28488 23131
rect 30190 23128 30196 23180
rect 30248 23128 30254 23180
rect 30282 23128 30288 23180
rect 30340 23128 30346 23180
rect 31662 23128 31668 23180
rect 31720 23128 31726 23180
rect 32858 23128 32864 23180
rect 32916 23168 32922 23180
rect 34333 23171 34391 23177
rect 34333 23168 34345 23171
rect 32916 23140 34345 23168
rect 32916 23128 32922 23140
rect 34333 23137 34345 23140
rect 34379 23137 34391 23171
rect 34333 23131 34391 23137
rect 34882 23128 34888 23180
rect 34940 23168 34946 23180
rect 34977 23171 35035 23177
rect 34977 23168 34989 23171
rect 34940 23140 34989 23168
rect 34940 23128 34946 23140
rect 34977 23137 34989 23140
rect 35023 23168 35035 23171
rect 37185 23171 37243 23177
rect 37185 23168 37197 23171
rect 35023 23140 37197 23168
rect 35023 23137 35035 23140
rect 34977 23131 35035 23137
rect 37185 23137 37197 23140
rect 37231 23168 37243 23171
rect 37458 23168 37464 23180
rect 37231 23140 37464 23168
rect 37231 23137 37243 23140
rect 37185 23131 37243 23137
rect 37458 23128 37464 23140
rect 37516 23168 37522 23180
rect 39022 23168 39028 23180
rect 37516 23140 39028 23168
rect 37516 23128 37522 23140
rect 39022 23128 39028 23140
rect 39080 23128 39086 23180
rect 39298 23128 39304 23180
rect 39356 23168 39362 23180
rect 39758 23168 39764 23180
rect 39356 23140 39764 23168
rect 39356 23128 39362 23140
rect 39758 23128 39764 23140
rect 39816 23128 39822 23180
rect 31018 23100 31024 23112
rect 28224 23004 28488 23032
rect 28644 23072 31024 23100
rect 28224 22992 28230 23004
rect 26344 22936 27384 22964
rect 27430 22924 27436 22976
rect 27488 22924 27494 22976
rect 28261 22967 28319 22973
rect 28261 22933 28273 22967
rect 28307 22964 28319 22967
rect 28644 22964 28672 23072
rect 31018 23060 31024 23072
rect 31076 23060 31082 23112
rect 31202 23060 31208 23112
rect 31260 23100 31266 23112
rect 31389 23103 31447 23109
rect 31389 23100 31401 23103
rect 31260 23072 31401 23100
rect 31260 23060 31266 23072
rect 31389 23069 31401 23072
rect 31435 23069 31447 23103
rect 31389 23063 31447 23069
rect 33689 23103 33747 23109
rect 33689 23069 33701 23103
rect 33735 23100 33747 23103
rect 33962 23100 33968 23112
rect 33735 23072 33968 23100
rect 33735 23069 33747 23072
rect 33689 23063 33747 23069
rect 33962 23060 33968 23072
rect 34020 23060 34026 23112
rect 40420 23109 40448 23196
rect 40681 23171 40739 23177
rect 40681 23137 40693 23171
rect 40727 23137 40739 23171
rect 40681 23131 40739 23137
rect 40405 23103 40463 23109
rect 40405 23069 40417 23103
rect 40451 23069 40463 23103
rect 40696 23100 40724 23131
rect 41506 23128 41512 23180
rect 41564 23128 41570 23180
rect 40770 23100 40776 23112
rect 40696 23072 40776 23100
rect 40405 23063 40463 23069
rect 40770 23060 40776 23072
rect 40828 23060 40834 23112
rect 43070 23100 43076 23112
rect 42918 23072 43076 23100
rect 43070 23060 43076 23072
rect 43128 23100 43134 23112
rect 43732 23100 43760 23276
rect 43898 23264 43904 23276
rect 43956 23264 43962 23316
rect 44174 23264 44180 23316
rect 44232 23304 44238 23316
rect 44818 23304 44824 23316
rect 44232 23276 44824 23304
rect 44232 23264 44238 23276
rect 44818 23264 44824 23276
rect 44876 23264 44882 23316
rect 45094 23264 45100 23316
rect 45152 23304 45158 23316
rect 45278 23304 45284 23316
rect 45152 23276 45284 23304
rect 45152 23264 45158 23276
rect 45278 23264 45284 23276
rect 45336 23264 45342 23316
rect 47578 23264 47584 23316
rect 47636 23264 47642 23316
rect 47762 23264 47768 23316
rect 47820 23304 47826 23316
rect 47949 23307 48007 23313
rect 47949 23304 47961 23307
rect 47820 23276 47961 23304
rect 47820 23264 47826 23276
rect 47949 23273 47961 23276
rect 47995 23273 48007 23307
rect 47949 23267 48007 23273
rect 48498 23264 48504 23316
rect 48556 23264 48562 23316
rect 48958 23264 48964 23316
rect 49016 23304 49022 23316
rect 49237 23307 49295 23313
rect 49237 23304 49249 23307
rect 49016 23276 49249 23304
rect 49016 23264 49022 23276
rect 49237 23273 49249 23276
rect 49283 23273 49295 23307
rect 49237 23267 49295 23273
rect 44082 23196 44088 23248
rect 44140 23236 44146 23248
rect 47857 23239 47915 23245
rect 47857 23236 47869 23239
rect 44140 23208 47869 23236
rect 44140 23196 44146 23208
rect 47857 23205 47869 23208
rect 47903 23205 47915 23239
rect 47857 23199 47915 23205
rect 43898 23128 43904 23180
rect 43956 23168 43962 23180
rect 45189 23171 45247 23177
rect 45189 23168 45201 23171
rect 43956 23140 45201 23168
rect 43956 23128 43962 23140
rect 45189 23137 45201 23140
rect 45235 23168 45247 23171
rect 45554 23168 45560 23180
rect 45235 23140 45560 23168
rect 45235 23137 45247 23140
rect 45189 23131 45247 23137
rect 45554 23128 45560 23140
rect 45612 23128 45618 23180
rect 45664 23140 46796 23168
rect 43128 23072 43760 23100
rect 43128 23060 43134 23072
rect 44082 23060 44088 23112
rect 44140 23100 44146 23112
rect 44269 23103 44327 23109
rect 44269 23100 44281 23103
rect 44140 23072 44281 23100
rect 44140 23060 44146 23072
rect 44269 23069 44281 23072
rect 44315 23069 44327 23103
rect 44269 23063 44327 23069
rect 44542 23060 44548 23112
rect 44600 23100 44606 23112
rect 45465 23103 45523 23109
rect 45465 23100 45477 23103
rect 44600 23072 45477 23100
rect 44600 23060 44606 23072
rect 45465 23069 45477 23072
rect 45511 23069 45523 23103
rect 45465 23063 45523 23069
rect 28718 22992 28724 23044
rect 28776 23032 28782 23044
rect 30834 23032 30840 23044
rect 28776 23004 30840 23032
rect 28776 22992 28782 23004
rect 30834 22992 30840 23004
rect 30892 22992 30898 23044
rect 30926 22992 30932 23044
rect 30984 23032 30990 23044
rect 32122 23032 32128 23044
rect 30984 23004 32128 23032
rect 30984 22992 30990 23004
rect 32122 22992 32128 23004
rect 32180 22992 32186 23044
rect 35250 22992 35256 23044
rect 35308 22992 35314 23044
rect 35986 22992 35992 23044
rect 36044 22992 36050 23044
rect 37461 23035 37519 23041
rect 37461 23001 37473 23035
rect 37507 23001 37519 23035
rect 39482 23032 39488 23044
rect 38686 23004 39488 23032
rect 37461 22995 37519 23001
rect 28307 22936 28672 22964
rect 28997 22967 29055 22973
rect 28307 22933 28319 22936
rect 28261 22927 28319 22933
rect 28997 22933 29009 22967
rect 29043 22964 29055 22967
rect 29086 22964 29092 22976
rect 29043 22936 29092 22964
rect 29043 22933 29055 22936
rect 28997 22927 29055 22933
rect 29086 22924 29092 22936
rect 29144 22924 29150 22976
rect 29181 22967 29239 22973
rect 29181 22933 29193 22967
rect 29227 22964 29239 22967
rect 29270 22964 29276 22976
rect 29227 22936 29276 22964
rect 29227 22933 29239 22936
rect 29181 22927 29239 22933
rect 29270 22924 29276 22936
rect 29328 22924 29334 22976
rect 29362 22924 29368 22976
rect 29420 22924 29426 22976
rect 30098 22924 30104 22976
rect 30156 22924 30162 22976
rect 30650 22924 30656 22976
rect 30708 22964 30714 22976
rect 30745 22967 30803 22973
rect 30745 22964 30757 22967
rect 30708 22936 30757 22964
rect 30708 22924 30714 22936
rect 30745 22933 30757 22936
rect 30791 22933 30803 22967
rect 30745 22927 30803 22933
rect 31478 22924 31484 22976
rect 31536 22964 31542 22976
rect 33137 22967 33195 22973
rect 33137 22964 33149 22967
rect 31536 22936 33149 22964
rect 31536 22924 31542 22936
rect 33137 22933 33149 22936
rect 33183 22964 33195 22967
rect 35894 22964 35900 22976
rect 33183 22936 35900 22964
rect 33183 22933 33195 22936
rect 33137 22927 33195 22933
rect 35894 22924 35900 22936
rect 35952 22924 35958 22976
rect 36722 22924 36728 22976
rect 36780 22924 36786 22976
rect 37476 22964 37504 22995
rect 39482 22992 39488 23004
rect 39540 22992 39546 23044
rect 40494 22992 40500 23044
rect 40552 22992 40558 23044
rect 41690 23032 41696 23044
rect 41340 23004 41696 23032
rect 38286 22964 38292 22976
rect 37476 22936 38292 22964
rect 38286 22924 38292 22936
rect 38344 22924 38350 22976
rect 39298 22924 39304 22976
rect 39356 22924 39362 22976
rect 39758 22924 39764 22976
rect 39816 22964 39822 22976
rect 41340 22964 41368 23004
rect 41690 22992 41696 23004
rect 41748 22992 41754 23044
rect 41785 23035 41843 23041
rect 41785 23001 41797 23035
rect 41831 23001 41843 23035
rect 41785 22995 41843 23001
rect 43533 23035 43591 23041
rect 43533 23001 43545 23035
rect 43579 23032 43591 23035
rect 43622 23032 43628 23044
rect 43579 23004 43628 23032
rect 43579 23001 43591 23004
rect 43533 22995 43591 23001
rect 39816 22936 41368 22964
rect 41800 22964 41828 22995
rect 43622 22992 43628 23004
rect 43680 22992 43686 23044
rect 44453 23035 44511 23041
rect 44453 23001 44465 23035
rect 44499 23032 44511 23035
rect 44634 23032 44640 23044
rect 44499 23004 44640 23032
rect 44499 23001 44511 23004
rect 44453 22995 44511 23001
rect 44634 22992 44640 23004
rect 44692 22992 44698 23044
rect 44818 22992 44824 23044
rect 44876 23032 44882 23044
rect 45664 23032 45692 23140
rect 46768 23109 46796 23140
rect 46477 23103 46535 23109
rect 46477 23069 46489 23103
rect 46523 23069 46535 23103
rect 46477 23063 46535 23069
rect 46753 23103 46811 23109
rect 46753 23069 46765 23103
rect 46799 23069 46811 23103
rect 46753 23063 46811 23069
rect 44876 23004 45692 23032
rect 44876 22992 44882 23004
rect 46492 22976 46520 23063
rect 48314 23060 48320 23112
rect 48372 23060 48378 23112
rect 49053 23103 49111 23109
rect 49053 23069 49065 23103
rect 49099 23069 49111 23103
rect 49053 23063 49111 23069
rect 47302 22992 47308 23044
rect 47360 23032 47366 23044
rect 49068 23032 49096 23063
rect 47360 23004 49096 23032
rect 47360 22992 47366 23004
rect 43714 22964 43720 22976
rect 41800 22936 43720 22964
rect 39816 22924 39822 22936
rect 43714 22924 43720 22936
rect 43772 22924 43778 22976
rect 43990 22924 43996 22976
rect 44048 22964 44054 22976
rect 46474 22964 46480 22976
rect 44048 22936 46480 22964
rect 44048 22924 44054 22936
rect 46474 22924 46480 22936
rect 46532 22924 46538 22976
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 3142 22720 3148 22772
rect 3200 22760 3206 22772
rect 6730 22760 6736 22772
rect 3200 22732 6736 22760
rect 3200 22720 3206 22732
rect 6730 22720 6736 22732
rect 6788 22720 6794 22772
rect 6822 22720 6828 22772
rect 6880 22760 6886 22772
rect 16574 22760 16580 22772
rect 6880 22720 6914 22760
rect 2866 22652 2872 22704
rect 2924 22692 2930 22704
rect 4246 22692 4252 22704
rect 2924 22664 4252 22692
rect 2924 22652 2930 22664
rect 4246 22652 4252 22664
rect 4304 22652 4310 22704
rect 6886 22692 6914 22720
rect 15120 22732 16580 22760
rect 14458 22692 14464 22704
rect 6886 22664 14464 22692
rect 14458 22652 14464 22664
rect 14516 22652 14522 22704
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22624 1823 22627
rect 1854 22624 1860 22636
rect 1811 22596 1860 22624
rect 1811 22593 1823 22596
rect 1765 22587 1823 22593
rect 1854 22584 1860 22596
rect 1912 22584 1918 22636
rect 3605 22627 3663 22633
rect 3605 22593 3617 22627
rect 3651 22624 3663 22627
rect 3878 22624 3884 22636
rect 3651 22596 3884 22624
rect 3651 22593 3663 22596
rect 3605 22587 3663 22593
rect 3878 22584 3884 22596
rect 3936 22624 3942 22636
rect 3973 22627 4031 22633
rect 3973 22624 3985 22627
rect 3936 22596 3985 22624
rect 3936 22584 3942 22596
rect 3973 22593 3985 22596
rect 4019 22593 4031 22627
rect 3973 22587 4031 22593
rect 4062 22584 4068 22636
rect 4120 22624 4126 22636
rect 4617 22627 4675 22633
rect 4617 22624 4629 22627
rect 4120 22596 4629 22624
rect 4120 22584 4126 22596
rect 4617 22593 4629 22596
rect 4663 22593 4675 22627
rect 4617 22587 4675 22593
rect 5810 22584 5816 22636
rect 5868 22624 5874 22636
rect 6825 22627 6883 22633
rect 6825 22624 6837 22627
rect 5868 22596 6837 22624
rect 5868 22584 5874 22596
rect 6825 22593 6837 22596
rect 6871 22593 6883 22627
rect 6825 22587 6883 22593
rect 6914 22584 6920 22636
rect 6972 22624 6978 22636
rect 7469 22627 7527 22633
rect 7469 22624 7481 22627
rect 6972 22596 7481 22624
rect 6972 22584 6978 22596
rect 7469 22593 7481 22596
rect 7515 22593 7527 22627
rect 7469 22587 7527 22593
rect 9766 22584 9772 22636
rect 9824 22584 9830 22636
rect 15120 22633 15148 22732
rect 16574 22720 16580 22732
rect 16632 22720 16638 22772
rect 16666 22720 16672 22772
rect 16724 22760 16730 22772
rect 16724 22732 18552 22760
rect 16724 22720 16730 22732
rect 15838 22652 15844 22704
rect 15896 22652 15902 22704
rect 17129 22695 17187 22701
rect 17129 22692 17141 22695
rect 15948 22664 17141 22692
rect 13081 22627 13139 22633
rect 13081 22624 13093 22627
rect 9876 22596 13093 22624
rect 2777 22559 2835 22565
rect 2777 22525 2789 22559
rect 2823 22556 2835 22559
rect 2866 22556 2872 22568
rect 2823 22528 2872 22556
rect 2823 22525 2835 22528
rect 2777 22519 2835 22525
rect 2866 22516 2872 22528
rect 2924 22516 2930 22568
rect 4154 22516 4160 22568
rect 4212 22516 4218 22568
rect 5074 22516 5080 22568
rect 5132 22516 5138 22568
rect 7650 22516 7656 22568
rect 7708 22556 7714 22568
rect 7929 22559 7987 22565
rect 7929 22556 7941 22559
rect 7708 22528 7941 22556
rect 7708 22516 7714 22528
rect 7929 22525 7941 22528
rect 7975 22525 7987 22559
rect 7929 22519 7987 22525
rect 9674 22516 9680 22568
rect 9732 22556 9738 22568
rect 9876 22556 9904 22596
rect 13081 22593 13093 22596
rect 13127 22593 13139 22627
rect 13081 22587 13139 22593
rect 15105 22627 15163 22633
rect 15105 22593 15117 22627
rect 15151 22593 15163 22627
rect 15105 22587 15163 22593
rect 9732 22528 9904 22556
rect 9732 22516 9738 22528
rect 9950 22516 9956 22568
rect 10008 22556 10014 22568
rect 10229 22559 10287 22565
rect 10229 22556 10241 22559
rect 10008 22528 10241 22556
rect 10008 22516 10014 22528
rect 10229 22525 10241 22528
rect 10275 22525 10287 22559
rect 11606 22556 11612 22568
rect 10229 22519 10287 22525
rect 10336 22528 11612 22556
rect 3418 22448 3424 22500
rect 3476 22488 3482 22500
rect 5626 22488 5632 22500
rect 3476 22460 5632 22488
rect 3476 22448 3482 22460
rect 5626 22448 5632 22460
rect 5684 22448 5690 22500
rect 6457 22491 6515 22497
rect 6457 22457 6469 22491
rect 6503 22488 6515 22491
rect 10336 22488 10364 22528
rect 11606 22516 11612 22528
rect 11664 22516 11670 22568
rect 11701 22559 11759 22565
rect 11701 22525 11713 22559
rect 11747 22556 11759 22559
rect 11790 22556 11796 22568
rect 11747 22528 11796 22556
rect 11747 22525 11759 22528
rect 11701 22519 11759 22525
rect 11790 22516 11796 22528
rect 11848 22516 11854 22568
rect 11974 22516 11980 22568
rect 12032 22516 12038 22568
rect 13814 22516 13820 22568
rect 13872 22516 13878 22568
rect 6503 22460 10364 22488
rect 6503 22457 6515 22460
rect 6457 22451 6515 22457
rect 10410 22448 10416 22500
rect 10468 22488 10474 22500
rect 15948 22488 15976 22664
rect 17129 22661 17141 22664
rect 17175 22661 17187 22695
rect 18414 22692 18420 22704
rect 18354 22664 18420 22692
rect 17129 22655 17187 22661
rect 18414 22652 18420 22664
rect 18472 22652 18478 22704
rect 18524 22692 18552 22732
rect 18598 22720 18604 22772
rect 18656 22720 18662 22772
rect 19058 22720 19064 22772
rect 19116 22720 19122 22772
rect 25130 22760 25136 22772
rect 22664 22732 25136 22760
rect 19518 22692 19524 22704
rect 18524 22664 19524 22692
rect 19518 22652 19524 22664
rect 19576 22652 19582 22704
rect 20346 22652 20352 22704
rect 20404 22652 20410 22704
rect 21082 22652 21088 22704
rect 21140 22692 21146 22704
rect 21818 22692 21824 22704
rect 21140 22664 21824 22692
rect 21140 22652 21146 22664
rect 21818 22652 21824 22664
rect 21876 22652 21882 22704
rect 22281 22695 22339 22701
rect 22281 22661 22293 22695
rect 22327 22692 22339 22695
rect 22664 22692 22692 22732
rect 25130 22720 25136 22732
rect 25188 22720 25194 22772
rect 26418 22760 26424 22772
rect 25516 22732 26424 22760
rect 22327 22664 22692 22692
rect 22327 22661 22339 22664
rect 22281 22655 22339 22661
rect 23290 22652 23296 22704
rect 23348 22652 23354 22704
rect 23566 22652 23572 22704
rect 23624 22692 23630 22704
rect 24394 22692 24400 22704
rect 23624 22664 24400 22692
rect 23624 22652 23630 22664
rect 24394 22652 24400 22664
rect 24452 22652 24458 22704
rect 25516 22692 25544 22732
rect 26418 22720 26424 22732
rect 26476 22720 26482 22772
rect 26878 22720 26884 22772
rect 26936 22760 26942 22772
rect 27341 22763 27399 22769
rect 27341 22760 27353 22763
rect 26936 22732 27353 22760
rect 26936 22720 26942 22732
rect 27341 22729 27353 22732
rect 27387 22729 27399 22763
rect 27341 22723 27399 22729
rect 27430 22720 27436 22772
rect 27488 22760 27494 22772
rect 27488 22732 30512 22760
rect 27488 22720 27494 22732
rect 26510 22692 26516 22704
rect 24780 22664 25544 22692
rect 26358 22664 26516 22692
rect 16850 22584 16856 22636
rect 16908 22584 16914 22636
rect 21174 22584 21180 22636
rect 21232 22624 21238 22636
rect 22002 22624 22008 22636
rect 21232 22596 22008 22624
rect 21232 22584 21238 22596
rect 22002 22584 22008 22596
rect 22060 22584 22066 22636
rect 24780 22624 24808 22664
rect 26510 22652 26516 22664
rect 26568 22692 26574 22704
rect 26970 22692 26976 22704
rect 26568 22664 26976 22692
rect 26568 22652 26574 22664
rect 26970 22652 26976 22664
rect 27028 22652 27034 22704
rect 27706 22652 27712 22704
rect 27764 22692 27770 22704
rect 27801 22695 27859 22701
rect 27801 22692 27813 22695
rect 27764 22664 27813 22692
rect 27764 22652 27770 22664
rect 27801 22661 27813 22664
rect 27847 22692 27859 22695
rect 28626 22692 28632 22704
rect 27847 22664 28632 22692
rect 27847 22661 27859 22664
rect 27801 22655 27859 22661
rect 28626 22652 28632 22664
rect 28684 22652 28690 22704
rect 30006 22692 30012 22704
rect 29578 22664 30012 22692
rect 30006 22652 30012 22664
rect 30064 22652 30070 22704
rect 24412 22596 24808 22624
rect 16960 22528 19380 22556
rect 16960 22488 16988 22528
rect 10468 22460 15976 22488
rect 16040 22460 16988 22488
rect 10468 22448 10474 22460
rect 5718 22380 5724 22432
rect 5776 22420 5782 22432
rect 6917 22423 6975 22429
rect 6917 22420 6929 22423
rect 5776 22392 6929 22420
rect 5776 22380 5782 22392
rect 6917 22389 6929 22392
rect 6963 22389 6975 22423
rect 6917 22383 6975 22389
rect 9309 22423 9367 22429
rect 9309 22389 9321 22423
rect 9355 22420 9367 22423
rect 9398 22420 9404 22432
rect 9355 22392 9404 22420
rect 9355 22389 9367 22392
rect 9309 22383 9367 22389
rect 9398 22380 9404 22392
rect 9456 22380 9462 22432
rect 9493 22423 9551 22429
rect 9493 22389 9505 22423
rect 9539 22420 9551 22423
rect 13262 22420 13268 22432
rect 9539 22392 13268 22420
rect 9539 22389 9551 22392
rect 9493 22383 9551 22389
rect 13262 22380 13268 22392
rect 13320 22380 13326 22432
rect 13354 22380 13360 22432
rect 13412 22420 13418 22432
rect 16040 22420 16068 22460
rect 18782 22448 18788 22500
rect 18840 22488 18846 22500
rect 19352 22488 19380 22528
rect 19426 22516 19432 22568
rect 19484 22556 19490 22568
rect 19521 22559 19579 22565
rect 19521 22556 19533 22559
rect 19484 22528 19533 22556
rect 19484 22516 19490 22528
rect 19521 22525 19533 22528
rect 19567 22525 19579 22559
rect 19797 22559 19855 22565
rect 19797 22556 19809 22559
rect 19521 22519 19579 22525
rect 19628 22528 19809 22556
rect 19628 22488 19656 22528
rect 19797 22525 19809 22528
rect 19843 22525 19855 22559
rect 19797 22519 19855 22525
rect 21269 22559 21327 22565
rect 21269 22525 21281 22559
rect 21315 22556 21327 22559
rect 22646 22556 22652 22568
rect 21315 22528 22652 22556
rect 21315 22525 21327 22528
rect 21269 22519 21327 22525
rect 22646 22516 22652 22528
rect 22704 22516 22710 22568
rect 23753 22559 23811 22565
rect 23753 22525 23765 22559
rect 23799 22556 23811 22559
rect 24118 22556 24124 22568
rect 23799 22528 24124 22556
rect 23799 22525 23811 22528
rect 23753 22519 23811 22525
rect 24118 22516 24124 22528
rect 24176 22516 24182 22568
rect 24213 22559 24271 22565
rect 24213 22525 24225 22559
rect 24259 22556 24271 22559
rect 24302 22556 24308 22568
rect 24259 22528 24308 22556
rect 24259 22525 24271 22528
rect 24213 22519 24271 22525
rect 24302 22516 24308 22528
rect 24360 22516 24366 22568
rect 18840 22460 19288 22488
rect 19352 22460 19656 22488
rect 18840 22448 18846 22460
rect 13412 22392 16068 22420
rect 13412 22380 13418 22392
rect 16850 22380 16856 22432
rect 16908 22420 16914 22432
rect 17126 22420 17132 22432
rect 16908 22392 17132 22420
rect 16908 22380 16914 22392
rect 17126 22380 17132 22392
rect 17184 22420 17190 22432
rect 17862 22420 17868 22432
rect 17184 22392 17868 22420
rect 17184 22380 17190 22392
rect 17862 22380 17868 22392
rect 17920 22380 17926 22432
rect 19260 22429 19288 22460
rect 19245 22423 19303 22429
rect 19245 22389 19257 22423
rect 19291 22420 19303 22423
rect 22094 22420 22100 22432
rect 19291 22392 22100 22420
rect 19291 22389 19303 22392
rect 19245 22383 19303 22389
rect 22094 22380 22100 22392
rect 22152 22380 22158 22432
rect 22738 22380 22744 22432
rect 22796 22420 22802 22432
rect 24305 22423 24363 22429
rect 24305 22420 24317 22423
rect 22796 22392 24317 22420
rect 22796 22380 22802 22392
rect 24305 22389 24317 22392
rect 24351 22420 24363 22423
rect 24412 22420 24440 22596
rect 24854 22584 24860 22636
rect 24912 22584 24918 22636
rect 27249 22627 27307 22633
rect 27249 22593 27261 22627
rect 27295 22624 27307 22627
rect 27430 22624 27436 22636
rect 27295 22596 27436 22624
rect 27295 22593 27307 22596
rect 27249 22587 27307 22593
rect 27430 22584 27436 22596
rect 27488 22584 27494 22636
rect 24578 22516 24584 22568
rect 24636 22556 24642 22568
rect 25133 22559 25191 22565
rect 24636 22528 24992 22556
rect 24636 22516 24642 22528
rect 24351 22392 24440 22420
rect 24351 22389 24363 22392
rect 24305 22383 24363 22389
rect 24578 22380 24584 22432
rect 24636 22380 24642 22432
rect 24964 22420 24992 22528
rect 25133 22525 25145 22559
rect 25179 22556 25191 22559
rect 27798 22556 27804 22568
rect 25179 22528 27804 22556
rect 25179 22525 25191 22528
rect 25133 22519 25191 22525
rect 27798 22516 27804 22528
rect 27856 22516 27862 22568
rect 28077 22559 28135 22565
rect 28077 22525 28089 22559
rect 28123 22525 28135 22559
rect 28077 22519 28135 22525
rect 28353 22559 28411 22565
rect 28353 22525 28365 22559
rect 28399 22556 28411 22559
rect 30374 22556 30380 22568
rect 28399 22528 30380 22556
rect 28399 22525 28411 22528
rect 28353 22519 28411 22525
rect 26142 22448 26148 22500
rect 26200 22488 26206 22500
rect 26510 22488 26516 22500
rect 26200 22460 26516 22488
rect 26200 22448 26206 22460
rect 26510 22448 26516 22460
rect 26568 22448 26574 22500
rect 27246 22448 27252 22500
rect 27304 22488 27310 22500
rect 28092 22488 28120 22519
rect 30374 22516 30380 22528
rect 30432 22516 30438 22568
rect 30484 22556 30512 22732
rect 30834 22720 30840 22772
rect 30892 22760 30898 22772
rect 31573 22763 31631 22769
rect 31573 22760 31585 22763
rect 30892 22732 31585 22760
rect 30892 22720 30898 22732
rect 31573 22729 31585 22732
rect 31619 22729 31631 22763
rect 31573 22723 31631 22729
rect 31754 22720 31760 22772
rect 31812 22760 31818 22772
rect 32309 22763 32367 22769
rect 32309 22760 32321 22763
rect 31812 22732 32321 22760
rect 31812 22720 31818 22732
rect 32309 22729 32321 22732
rect 32355 22729 32367 22763
rect 32309 22723 32367 22729
rect 33410 22720 33416 22772
rect 33468 22720 33474 22772
rect 33502 22720 33508 22772
rect 33560 22760 33566 22772
rect 34882 22760 34888 22772
rect 33560 22732 34888 22760
rect 33560 22720 33566 22732
rect 30653 22695 30711 22701
rect 30653 22661 30665 22695
rect 30699 22692 30711 22695
rect 33594 22692 33600 22704
rect 30699 22664 33600 22692
rect 30699 22661 30711 22664
rect 30653 22655 30711 22661
rect 33594 22652 33600 22664
rect 33652 22652 33658 22704
rect 30745 22627 30803 22633
rect 30745 22593 30757 22627
rect 30791 22624 30803 22627
rect 32490 22624 32496 22636
rect 30791 22596 32496 22624
rect 30791 22593 30803 22596
rect 30745 22587 30803 22593
rect 32490 22584 32496 22596
rect 32548 22584 32554 22636
rect 33704 22633 33732 22732
rect 34882 22720 34888 22732
rect 34940 22720 34946 22772
rect 35618 22720 35624 22772
rect 35676 22760 35682 22772
rect 36081 22763 36139 22769
rect 36081 22760 36093 22763
rect 35676 22732 36093 22760
rect 35676 22720 35682 22732
rect 36081 22729 36093 22732
rect 36127 22729 36139 22763
rect 41509 22763 41567 22769
rect 41509 22760 41521 22763
rect 36081 22723 36139 22729
rect 37752 22732 41521 22760
rect 33870 22652 33876 22704
rect 33928 22692 33934 22704
rect 33965 22695 34023 22701
rect 33965 22692 33977 22695
rect 33928 22664 33977 22692
rect 33928 22652 33934 22664
rect 33965 22661 33977 22664
rect 34011 22661 34023 22695
rect 33965 22655 34023 22661
rect 34238 22652 34244 22704
rect 34296 22692 34302 22704
rect 37752 22701 37780 22732
rect 41509 22729 41521 22732
rect 41555 22729 41567 22763
rect 41509 22723 41567 22729
rect 41690 22720 41696 22772
rect 41748 22760 41754 22772
rect 44266 22760 44272 22772
rect 41748 22732 44272 22760
rect 41748 22720 41754 22732
rect 44266 22720 44272 22732
rect 44324 22720 44330 22772
rect 46934 22720 46940 22772
rect 46992 22720 46998 22772
rect 47302 22720 47308 22772
rect 47360 22760 47366 22772
rect 47765 22763 47823 22769
rect 47765 22760 47777 22763
rect 47360 22732 47777 22760
rect 47360 22720 47366 22732
rect 47765 22729 47777 22732
rect 47811 22729 47823 22763
rect 47765 22723 47823 22729
rect 48498 22720 48504 22772
rect 48556 22720 48562 22772
rect 49142 22720 49148 22772
rect 49200 22760 49206 22772
rect 49237 22763 49295 22769
rect 49237 22760 49249 22763
rect 49200 22732 49249 22760
rect 49200 22720 49206 22732
rect 49237 22729 49249 22732
rect 49283 22729 49295 22763
rect 49237 22723 49295 22729
rect 37737 22695 37795 22701
rect 34296 22664 34454 22692
rect 34296 22652 34302 22664
rect 37737 22661 37749 22695
rect 37783 22661 37795 22695
rect 39482 22692 39488 22704
rect 38962 22664 39488 22692
rect 37737 22655 37795 22661
rect 39482 22652 39488 22664
rect 39540 22652 39546 22704
rect 39574 22652 39580 22704
rect 39632 22692 39638 22704
rect 39632 22664 40448 22692
rect 39632 22652 39638 22664
rect 32677 22627 32735 22633
rect 32677 22593 32689 22627
rect 32723 22624 32735 22627
rect 33689 22627 33747 22633
rect 32723 22596 33640 22624
rect 32723 22593 32735 22596
rect 32677 22587 32735 22593
rect 30837 22559 30895 22565
rect 30837 22556 30849 22559
rect 30484 22528 30849 22556
rect 30837 22525 30849 22528
rect 30883 22525 30895 22559
rect 30837 22519 30895 22525
rect 31662 22516 31668 22568
rect 31720 22556 31726 22568
rect 31720 22528 32352 22556
rect 31720 22516 31726 22528
rect 31202 22488 31208 22500
rect 27304 22460 28120 22488
rect 27304 22448 27310 22460
rect 26234 22420 26240 22432
rect 24964 22392 26240 22420
rect 26234 22380 26240 22392
rect 26292 22380 26298 22432
rect 26602 22380 26608 22432
rect 26660 22380 26666 22432
rect 28092 22420 28120 22460
rect 29748 22460 31208 22488
rect 29748 22432 29776 22460
rect 31202 22448 31208 22460
rect 31260 22448 31266 22500
rect 32324 22488 32352 22528
rect 32766 22516 32772 22568
rect 32824 22516 32830 22568
rect 32861 22559 32919 22565
rect 32861 22525 32873 22559
rect 32907 22525 32919 22559
rect 32861 22519 32919 22525
rect 32876 22488 32904 22519
rect 32324 22460 32904 22488
rect 29730 22420 29736 22432
rect 28092 22392 29736 22420
rect 29730 22380 29736 22392
rect 29788 22380 29794 22432
rect 29825 22423 29883 22429
rect 29825 22389 29837 22423
rect 29871 22420 29883 22423
rect 29914 22420 29920 22432
rect 29871 22392 29920 22420
rect 29871 22389 29883 22392
rect 29825 22383 29883 22389
rect 29914 22380 29920 22392
rect 29972 22380 29978 22432
rect 30282 22380 30288 22432
rect 30340 22380 30346 22432
rect 33612 22420 33640 22596
rect 33689 22593 33701 22627
rect 33735 22593 33747 22627
rect 33689 22587 33747 22593
rect 36449 22627 36507 22633
rect 36449 22593 36461 22627
rect 36495 22624 36507 22627
rect 37090 22624 37096 22636
rect 36495 22596 37096 22624
rect 36495 22593 36507 22596
rect 36449 22587 36507 22593
rect 37090 22584 37096 22596
rect 37148 22584 37154 22636
rect 37458 22584 37464 22636
rect 37516 22584 37522 22636
rect 40034 22584 40040 22636
rect 40092 22584 40098 22636
rect 34422 22556 34428 22568
rect 33704 22528 34428 22556
rect 33704 22500 33732 22528
rect 34422 22516 34428 22528
rect 34480 22516 34486 22568
rect 34606 22516 34612 22568
rect 34664 22556 34670 22568
rect 36541 22559 36599 22565
rect 36541 22556 36553 22559
rect 34664 22528 36553 22556
rect 34664 22516 34670 22528
rect 36541 22525 36553 22528
rect 36587 22525 36599 22559
rect 36541 22519 36599 22525
rect 36725 22559 36783 22565
rect 36725 22525 36737 22559
rect 36771 22556 36783 22559
rect 39209 22559 39267 22565
rect 39209 22556 39221 22559
rect 36771 22528 39221 22556
rect 36771 22525 36783 22528
rect 36725 22519 36783 22525
rect 39209 22525 39221 22528
rect 39255 22525 39267 22559
rect 39209 22519 39267 22525
rect 33686 22448 33692 22500
rect 33744 22448 33750 22500
rect 35437 22491 35495 22497
rect 35437 22457 35449 22491
rect 35483 22488 35495 22491
rect 35526 22488 35532 22500
rect 35483 22460 35532 22488
rect 35483 22457 35495 22460
rect 35437 22451 35495 22457
rect 35526 22448 35532 22460
rect 35584 22448 35590 22500
rect 39224 22488 39252 22519
rect 40126 22516 40132 22568
rect 40184 22516 40190 22568
rect 40218 22516 40224 22568
rect 40276 22516 40282 22568
rect 40420 22556 40448 22664
rect 40494 22652 40500 22704
rect 40552 22692 40558 22704
rect 41322 22692 41328 22704
rect 40552 22664 41328 22692
rect 40552 22652 40558 22664
rect 41322 22652 41328 22664
rect 41380 22652 41386 22704
rect 41874 22652 41880 22704
rect 41932 22692 41938 22704
rect 42061 22695 42119 22701
rect 42061 22692 42073 22695
rect 41932 22664 42073 22692
rect 41932 22652 41938 22664
rect 42061 22661 42073 22664
rect 42107 22692 42119 22695
rect 42150 22692 42156 22704
rect 42107 22664 42156 22692
rect 42107 22661 42119 22664
rect 42061 22655 42119 22661
rect 42150 22652 42156 22664
rect 42208 22692 42214 22704
rect 42245 22695 42303 22701
rect 42245 22692 42257 22695
rect 42208 22664 42257 22692
rect 42208 22652 42214 22664
rect 42245 22661 42257 22664
rect 42291 22692 42303 22695
rect 43070 22692 43076 22704
rect 42291 22664 43076 22692
rect 42291 22661 42303 22664
rect 42245 22655 42303 22661
rect 43070 22652 43076 22664
rect 43128 22652 43134 22704
rect 46474 22652 46480 22704
rect 46532 22692 46538 22704
rect 47581 22695 47639 22701
rect 47581 22692 47593 22695
rect 46532 22664 47593 22692
rect 46532 22652 46538 22664
rect 47581 22661 47593 22664
rect 47627 22661 47639 22695
rect 47581 22655 47639 22661
rect 40865 22627 40923 22633
rect 40865 22593 40877 22627
rect 40911 22624 40923 22627
rect 41046 22624 41052 22636
rect 40911 22596 41052 22624
rect 40911 22593 40923 22596
rect 40865 22587 40923 22593
rect 41046 22584 41052 22596
rect 41104 22584 41110 22636
rect 42797 22627 42855 22633
rect 42797 22593 42809 22627
rect 42843 22624 42855 22627
rect 43346 22624 43352 22636
rect 42843 22596 43352 22624
rect 42843 22593 42855 22596
rect 42797 22587 42855 22593
rect 43346 22584 43352 22596
rect 43404 22584 43410 22636
rect 43530 22584 43536 22636
rect 43588 22584 43594 22636
rect 44358 22584 44364 22636
rect 44416 22624 44422 22636
rect 44821 22627 44879 22633
rect 44821 22624 44833 22627
rect 44416 22596 44833 22624
rect 44416 22584 44422 22596
rect 44821 22593 44833 22596
rect 44867 22593 44879 22627
rect 44821 22587 44879 22593
rect 45830 22584 45836 22636
rect 45888 22624 45894 22636
rect 45888 22596 46244 22624
rect 45888 22584 45894 22596
rect 43257 22559 43315 22565
rect 40420 22528 43208 22556
rect 40236 22488 40264 22516
rect 39224 22460 40264 22488
rect 40402 22448 40408 22500
rect 40460 22488 40466 22500
rect 40460 22460 42564 22488
rect 40460 22448 40466 22460
rect 34698 22420 34704 22432
rect 33612 22392 34704 22420
rect 34698 22380 34704 22392
rect 34756 22380 34762 22432
rect 35805 22423 35863 22429
rect 35805 22389 35817 22423
rect 35851 22420 35863 22423
rect 35894 22420 35900 22432
rect 35851 22392 35900 22420
rect 35851 22389 35863 22392
rect 35805 22383 35863 22389
rect 35894 22380 35900 22392
rect 35952 22380 35958 22432
rect 36722 22380 36728 22432
rect 36780 22420 36786 22432
rect 38746 22420 38752 22432
rect 36780 22392 38752 22420
rect 36780 22380 36786 22392
rect 38746 22380 38752 22392
rect 38804 22380 38810 22432
rect 39666 22380 39672 22432
rect 39724 22380 39730 22432
rect 42536 22420 42564 22460
rect 42610 22448 42616 22500
rect 42668 22448 42674 22500
rect 43180 22488 43208 22528
rect 43257 22525 43269 22559
rect 43303 22556 43315 22559
rect 44082 22556 44088 22568
rect 43303 22528 44088 22556
rect 43303 22525 43315 22528
rect 43257 22519 43315 22525
rect 44082 22516 44088 22528
rect 44140 22516 44146 22568
rect 44545 22559 44603 22565
rect 44545 22525 44557 22559
rect 44591 22556 44603 22559
rect 44726 22556 44732 22568
rect 44591 22528 44732 22556
rect 44591 22525 44603 22528
rect 44545 22519 44603 22525
rect 44726 22516 44732 22528
rect 44784 22556 44790 22568
rect 45002 22556 45008 22568
rect 44784 22528 45008 22556
rect 44784 22516 44790 22528
rect 45002 22516 45008 22528
rect 45060 22516 45066 22568
rect 46106 22516 46112 22568
rect 46164 22516 46170 22568
rect 46216 22556 46244 22596
rect 46842 22584 46848 22636
rect 46900 22624 46906 22636
rect 47121 22627 47179 22633
rect 47121 22624 47133 22627
rect 46900 22596 47133 22624
rect 46900 22584 46906 22596
rect 47121 22593 47133 22596
rect 47167 22593 47179 22627
rect 47121 22587 47179 22593
rect 47762 22584 47768 22636
rect 47820 22624 47826 22636
rect 48317 22627 48375 22633
rect 48317 22624 48329 22627
rect 47820 22596 48329 22624
rect 47820 22584 47826 22596
rect 48317 22593 48329 22596
rect 48363 22593 48375 22627
rect 48317 22587 48375 22593
rect 49053 22627 49111 22633
rect 49053 22593 49065 22627
rect 49099 22624 49111 22627
rect 49326 22624 49332 22636
rect 49099 22596 49332 22624
rect 49099 22593 49111 22596
rect 49053 22587 49111 22593
rect 49326 22584 49332 22596
rect 49384 22584 49390 22636
rect 47305 22559 47363 22565
rect 47305 22556 47317 22559
rect 46216 22528 47317 22556
rect 47305 22525 47317 22528
rect 47351 22525 47363 22559
rect 47305 22519 47363 22525
rect 46842 22488 46848 22500
rect 43180 22460 46848 22488
rect 46842 22448 46848 22460
rect 46900 22448 46906 22500
rect 48041 22491 48099 22497
rect 48041 22457 48053 22491
rect 48087 22488 48099 22491
rect 49142 22488 49148 22500
rect 48087 22460 49148 22488
rect 48087 22457 48099 22460
rect 48041 22451 48099 22457
rect 49142 22448 49148 22460
rect 49200 22448 49206 22500
rect 48314 22420 48320 22432
rect 42536 22392 48320 22420
rect 48314 22380 48320 22392
rect 48372 22380 48378 22432
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 1578 22176 1584 22228
rect 1636 22216 1642 22228
rect 4614 22216 4620 22228
rect 1636 22188 4620 22216
rect 1636 22176 1642 22188
rect 4614 22176 4620 22188
rect 4672 22176 4678 22228
rect 13906 22176 13912 22228
rect 13964 22216 13970 22228
rect 15454 22219 15512 22225
rect 15454 22216 15466 22219
rect 13964 22188 15466 22216
rect 13964 22176 13970 22188
rect 15454 22185 15466 22188
rect 15500 22185 15512 22219
rect 15454 22179 15512 22185
rect 16850 22176 16856 22228
rect 16908 22216 16914 22228
rect 18414 22216 18420 22228
rect 16908 22188 18420 22216
rect 16908 22176 16914 22188
rect 18414 22176 18420 22188
rect 18472 22176 18478 22228
rect 21440 22219 21498 22225
rect 21440 22185 21452 22219
rect 21486 22216 21498 22219
rect 21634 22216 21640 22228
rect 21486 22188 21640 22216
rect 21486 22185 21498 22188
rect 21440 22179 21498 22185
rect 21634 22176 21640 22188
rect 21692 22176 21698 22228
rect 21818 22176 21824 22228
rect 21876 22216 21882 22228
rect 21876 22188 22600 22216
rect 21876 22176 21882 22188
rect 2222 22108 2228 22160
rect 2280 22148 2286 22160
rect 4522 22148 4528 22160
rect 2280 22120 4528 22148
rect 2280 22108 2286 22120
rect 4522 22108 4528 22120
rect 4580 22108 4586 22160
rect 11790 22148 11796 22160
rect 11624 22120 11796 22148
rect 1302 22040 1308 22092
rect 1360 22080 1366 22092
rect 2041 22083 2099 22089
rect 2041 22080 2053 22083
rect 1360 22052 2053 22080
rect 1360 22040 1366 22052
rect 2041 22049 2053 22052
rect 2087 22049 2099 22083
rect 2041 22043 2099 22049
rect 3786 22040 3792 22092
rect 3844 22080 3850 22092
rect 4433 22083 4491 22089
rect 4433 22080 4445 22083
rect 3844 22052 4445 22080
rect 3844 22040 3850 22052
rect 4433 22049 4445 22052
rect 4479 22049 4491 22083
rect 4433 22043 4491 22049
rect 6730 22040 6736 22092
rect 6788 22040 6794 22092
rect 8570 22040 8576 22092
rect 8628 22040 8634 22092
rect 9858 22040 9864 22092
rect 9916 22040 9922 22092
rect 10042 22040 10048 22092
rect 10100 22080 10106 22092
rect 11241 22083 11299 22089
rect 11241 22080 11253 22083
rect 10100 22052 11253 22080
rect 10100 22040 10106 22052
rect 11241 22049 11253 22052
rect 11287 22049 11299 22083
rect 11241 22043 11299 22049
rect 1762 21972 1768 22024
rect 1820 21972 1826 22024
rect 4065 22015 4123 22021
rect 4065 21981 4077 22015
rect 4111 21981 4123 22015
rect 4065 21975 4123 21981
rect 5997 22015 6055 22021
rect 5997 21981 6009 22015
rect 6043 22012 6055 22015
rect 7650 22012 7656 22024
rect 6043 21984 7656 22012
rect 6043 21981 6055 21984
rect 5997 21975 6055 21981
rect 4080 21876 4108 21975
rect 7650 21972 7656 21984
rect 7708 21972 7714 22024
rect 7926 21972 7932 22024
rect 7984 21972 7990 22024
rect 9122 21972 9128 22024
rect 9180 21972 9186 22024
rect 11624 22012 11652 22120
rect 11790 22108 11796 22120
rect 11848 22108 11854 22160
rect 11882 22108 11888 22160
rect 11940 22148 11946 22160
rect 11940 22120 12480 22148
rect 11940 22108 11946 22120
rect 11698 22040 11704 22092
rect 11756 22040 11762 22092
rect 12452 22089 12480 22120
rect 13630 22108 13636 22160
rect 13688 22148 13694 22160
rect 13688 22120 15332 22148
rect 13688 22108 13694 22120
rect 12437 22083 12495 22089
rect 12437 22049 12449 22083
rect 12483 22049 12495 22083
rect 12437 22043 12495 22049
rect 13909 22083 13967 22089
rect 13909 22049 13921 22083
rect 13955 22080 13967 22083
rect 14274 22080 14280 22092
rect 13955 22052 14280 22080
rect 13955 22049 13967 22052
rect 13909 22043 13967 22049
rect 14274 22040 14280 22052
rect 14332 22040 14338 22092
rect 14734 22040 14740 22092
rect 14792 22040 14798 22092
rect 15304 22080 15332 22120
rect 17126 22108 17132 22160
rect 17184 22148 17190 22160
rect 17184 22120 18092 22148
rect 17184 22108 17190 22120
rect 18064 22080 18092 22120
rect 20346 22080 20352 22092
rect 15304 22052 17908 22080
rect 18064 22052 20352 22080
rect 9600 21984 11652 22012
rect 7561 21947 7619 21953
rect 7561 21913 7573 21947
rect 7607 21944 7619 21947
rect 9600 21944 9628 21984
rect 11790 21972 11796 22024
rect 11848 22012 11854 22024
rect 11977 22015 12035 22021
rect 11977 22012 11989 22015
rect 11848 21984 11989 22012
rect 11848 21972 11854 21984
rect 11977 21981 11989 21984
rect 12023 21981 12035 22015
rect 11977 21975 12035 21981
rect 15194 21972 15200 22024
rect 15252 21972 15258 22024
rect 17494 21972 17500 22024
rect 17552 21972 17558 22024
rect 7607 21916 9628 21944
rect 7607 21913 7619 21916
rect 7561 21907 7619 21913
rect 11054 21904 11060 21956
rect 11112 21904 11118 21956
rect 13725 21947 13783 21953
rect 13725 21913 13737 21947
rect 13771 21944 13783 21947
rect 14366 21944 14372 21956
rect 13771 21916 14372 21944
rect 13771 21913 13783 21916
rect 13725 21907 13783 21913
rect 14366 21904 14372 21916
rect 14424 21904 14430 21956
rect 14553 21947 14611 21953
rect 14553 21913 14565 21947
rect 14599 21944 14611 21947
rect 14826 21944 14832 21956
rect 14599 21916 14832 21944
rect 14599 21913 14611 21916
rect 14553 21907 14611 21913
rect 14826 21904 14832 21916
rect 14884 21904 14890 21956
rect 16850 21944 16856 21956
rect 16698 21916 16856 21944
rect 16850 21904 16856 21916
rect 16908 21904 16914 21956
rect 9398 21876 9404 21888
rect 4080 21848 9404 21876
rect 9398 21836 9404 21848
rect 9456 21836 9462 21888
rect 14182 21836 14188 21888
rect 14240 21836 14246 21888
rect 15286 21836 15292 21888
rect 15344 21876 15350 21888
rect 16945 21879 17003 21885
rect 16945 21876 16957 21879
rect 15344 21848 16957 21876
rect 15344 21836 15350 21848
rect 16945 21845 16957 21848
rect 16991 21845 17003 21879
rect 16945 21839 17003 21845
rect 17034 21836 17040 21888
rect 17092 21876 17098 21888
rect 17770 21876 17776 21888
rect 17092 21848 17776 21876
rect 17092 21836 17098 21848
rect 17770 21836 17776 21848
rect 17828 21836 17834 21888
rect 17880 21876 17908 22052
rect 20346 22040 20352 22052
rect 20404 22040 20410 22092
rect 20438 22040 20444 22092
rect 20496 22080 20502 22092
rect 20533 22083 20591 22089
rect 20533 22080 20545 22083
rect 20496 22052 20545 22080
rect 20496 22040 20502 22052
rect 20533 22049 20545 22052
rect 20579 22049 20591 22083
rect 20533 22043 20591 22049
rect 20622 22040 20628 22092
rect 20680 22080 20686 22092
rect 22462 22080 22468 22092
rect 20680 22052 22468 22080
rect 20680 22040 20686 22052
rect 22462 22040 22468 22052
rect 22520 22040 22526 22092
rect 18046 21972 18052 22024
rect 18104 22012 18110 22024
rect 19334 22012 19340 22024
rect 18104 21984 19340 22012
rect 18104 21972 18110 21984
rect 19334 21972 19340 21984
rect 19392 21972 19398 22024
rect 19426 21972 19432 22024
rect 19484 22012 19490 22024
rect 19521 22015 19579 22021
rect 19521 22012 19533 22015
rect 19484 21984 19533 22012
rect 19484 21972 19490 21984
rect 19521 21981 19533 21984
rect 19567 22012 19579 22015
rect 19705 22015 19763 22021
rect 19705 22012 19717 22015
rect 19567 21984 19717 22012
rect 19567 21981 19579 21984
rect 19521 21975 19579 21981
rect 19705 21981 19717 21984
rect 19751 22012 19763 22015
rect 20070 22012 20076 22024
rect 19751 21984 20076 22012
rect 19751 21981 19763 21984
rect 19705 21975 19763 21981
rect 20070 21972 20076 21984
rect 20128 21972 20134 22024
rect 21174 21972 21180 22024
rect 21232 21972 21238 22024
rect 22572 22012 22600 22188
rect 23750 22176 23756 22228
rect 23808 22216 23814 22228
rect 24581 22219 24639 22225
rect 24581 22216 24593 22219
rect 23808 22188 24593 22216
rect 23808 22176 23814 22188
rect 24581 22185 24593 22188
rect 24627 22185 24639 22219
rect 24581 22179 24639 22185
rect 25130 22176 25136 22228
rect 25188 22216 25194 22228
rect 27246 22216 27252 22228
rect 25188 22188 27252 22216
rect 25188 22176 25194 22188
rect 27246 22176 27252 22188
rect 27304 22176 27310 22228
rect 27338 22176 27344 22228
rect 27396 22216 27402 22228
rect 27396 22188 28994 22216
rect 27396 22176 27402 22188
rect 22646 22108 22652 22160
rect 22704 22148 22710 22160
rect 22704 22120 23612 22148
rect 22704 22108 22710 22120
rect 22738 22040 22744 22092
rect 22796 22080 22802 22092
rect 23584 22080 23612 22120
rect 25774 22108 25780 22160
rect 25832 22148 25838 22160
rect 26602 22148 26608 22160
rect 25832 22120 26608 22148
rect 25832 22108 25838 22120
rect 24210 22080 24216 22092
rect 22796 22052 23520 22080
rect 23584 22052 24216 22080
rect 22796 22040 22802 22052
rect 23198 22012 23204 22024
rect 22572 21998 23204 22012
rect 22586 21984 23204 21998
rect 23198 21972 23204 21984
rect 23256 21972 23262 22024
rect 23290 21972 23296 22024
rect 23348 22012 23354 22024
rect 23385 22015 23443 22021
rect 23385 22012 23397 22015
rect 23348 21984 23397 22012
rect 23348 21972 23354 21984
rect 23385 21981 23397 21984
rect 23431 21981 23443 22015
rect 23492 22012 23520 22052
rect 24210 22040 24216 22052
rect 24268 22080 24274 22092
rect 25133 22083 25191 22089
rect 25133 22080 25145 22083
rect 24268 22052 25145 22080
rect 24268 22040 24274 22052
rect 25133 22049 25145 22052
rect 25179 22049 25191 22083
rect 25133 22043 25191 22049
rect 25406 22040 25412 22092
rect 25464 22080 25470 22092
rect 26142 22080 26148 22092
rect 25464 22052 26148 22080
rect 25464 22040 25470 22052
rect 26142 22040 26148 22052
rect 26200 22040 26206 22092
rect 26528 22089 26556 22120
rect 26602 22108 26608 22120
rect 26660 22108 26666 22160
rect 26694 22108 26700 22160
rect 26752 22148 26758 22160
rect 26752 22120 27568 22148
rect 26752 22108 26758 22120
rect 26513 22083 26571 22089
rect 26513 22049 26525 22083
rect 26559 22049 26571 22083
rect 27540 22080 27568 22120
rect 27614 22108 27620 22160
rect 27672 22148 27678 22160
rect 28353 22151 28411 22157
rect 28353 22148 28365 22151
rect 27672 22120 28365 22148
rect 27672 22108 27678 22120
rect 28353 22117 28365 22120
rect 28399 22117 28411 22151
rect 28353 22111 28411 22117
rect 28966 22148 28994 22188
rect 29362 22176 29368 22228
rect 29420 22216 29426 22228
rect 30282 22216 30288 22228
rect 29420 22188 30288 22216
rect 29420 22176 29426 22188
rect 30282 22176 30288 22188
rect 30340 22176 30346 22228
rect 30374 22176 30380 22228
rect 30432 22176 30438 22228
rect 31662 22216 31668 22228
rect 30576 22188 31668 22216
rect 29914 22148 29920 22160
rect 28966 22120 29920 22148
rect 28966 22092 28994 22120
rect 29914 22108 29920 22120
rect 29972 22108 29978 22160
rect 27709 22083 27767 22089
rect 27709 22080 27721 22083
rect 26513 22043 26571 22049
rect 27080 22052 27476 22080
rect 27540 22052 27721 22080
rect 24029 22015 24087 22021
rect 24029 22012 24041 22015
rect 23492 21984 24041 22012
rect 23385 21975 23443 21981
rect 24029 21981 24041 21984
rect 24075 21981 24087 22015
rect 24029 21975 24087 21981
rect 25038 21972 25044 22024
rect 25096 22012 25102 22024
rect 26878 22012 26884 22024
rect 25096 21984 26884 22012
rect 25096 21972 25102 21984
rect 26878 21972 26884 21984
rect 26936 21972 26942 22024
rect 18138 21904 18144 21956
rect 18196 21944 18202 21956
rect 18417 21947 18475 21953
rect 18417 21944 18429 21947
rect 18196 21916 18429 21944
rect 18196 21904 18202 21916
rect 18417 21913 18429 21916
rect 18463 21913 18475 21947
rect 20162 21944 20168 21956
rect 18417 21907 18475 21913
rect 18524 21916 20168 21944
rect 18524 21876 18552 21916
rect 20162 21904 20168 21916
rect 20220 21904 20226 21956
rect 20349 21947 20407 21953
rect 20349 21913 20361 21947
rect 20395 21944 20407 21947
rect 20714 21944 20720 21956
rect 20395 21916 20720 21944
rect 20395 21913 20407 21916
rect 20349 21907 20407 21913
rect 20714 21904 20720 21916
rect 20772 21904 20778 21956
rect 26421 21947 26479 21953
rect 22756 21916 26004 21944
rect 17880 21848 18552 21876
rect 19337 21879 19395 21885
rect 19337 21845 19349 21879
rect 19383 21876 19395 21879
rect 19426 21876 19432 21888
rect 19383 21848 19432 21876
rect 19383 21845 19395 21848
rect 19337 21839 19395 21845
rect 19426 21836 19432 21848
rect 19484 21836 19490 21888
rect 19978 21836 19984 21888
rect 20036 21836 20042 21888
rect 20441 21879 20499 21885
rect 20441 21845 20453 21879
rect 20487 21876 20499 21879
rect 22756 21876 22784 21916
rect 20487 21848 22784 21876
rect 22925 21879 22983 21885
rect 20487 21845 20499 21848
rect 20441 21839 20499 21845
rect 22925 21845 22937 21879
rect 22971 21876 22983 21879
rect 23014 21876 23020 21888
rect 22971 21848 23020 21876
rect 22971 21845 22983 21848
rect 22925 21839 22983 21845
rect 23014 21836 23020 21848
rect 23072 21836 23078 21888
rect 24302 21836 24308 21888
rect 24360 21876 24366 21888
rect 24949 21879 25007 21885
rect 24949 21876 24961 21879
rect 24360 21848 24961 21876
rect 24360 21836 24366 21848
rect 24949 21845 24961 21848
rect 24995 21845 25007 21879
rect 24949 21839 25007 21845
rect 25406 21836 25412 21888
rect 25464 21876 25470 21888
rect 25976 21885 26004 21916
rect 26421 21913 26433 21947
rect 26467 21944 26479 21947
rect 27080 21944 27108 22052
rect 26467 21916 27108 21944
rect 27448 21944 27476 22052
rect 27709 22049 27721 22052
rect 27755 22049 27767 22083
rect 27709 22043 27767 22049
rect 28902 22040 28908 22092
rect 28960 22089 28994 22092
rect 28960 22083 29009 22089
rect 28960 22049 28963 22083
rect 28997 22049 29009 22083
rect 28960 22043 29009 22049
rect 28960 22040 28966 22043
rect 28721 22015 28779 22021
rect 28721 21981 28733 22015
rect 28767 22012 28779 22015
rect 28810 22012 28816 22024
rect 28767 21984 28816 22012
rect 28767 21981 28779 21984
rect 28721 21975 28779 21981
rect 28810 21972 28816 21984
rect 28868 21972 28874 22024
rect 29638 21972 29644 22024
rect 29696 22012 29702 22024
rect 29733 22015 29791 22021
rect 29733 22012 29745 22015
rect 29696 21984 29745 22012
rect 29696 21972 29702 21984
rect 29733 21981 29745 21984
rect 29779 22012 29791 22015
rect 30576 22012 30604 22188
rect 31662 22176 31668 22188
rect 31720 22176 31726 22228
rect 32490 22176 32496 22228
rect 32548 22216 32554 22228
rect 34238 22216 34244 22228
rect 32548 22188 34244 22216
rect 32548 22176 32554 22188
rect 34238 22176 34244 22188
rect 34296 22176 34302 22228
rect 37540 22219 37598 22225
rect 35544 22188 35848 22216
rect 32582 22108 32588 22160
rect 32640 22108 32646 22160
rect 33778 22148 33784 22160
rect 33612 22120 33784 22148
rect 30837 22083 30895 22089
rect 30837 22049 30849 22083
rect 30883 22080 30895 22083
rect 31202 22080 31208 22092
rect 30883 22052 31208 22080
rect 30883 22049 30895 22052
rect 30837 22043 30895 22049
rect 31202 22040 31208 22052
rect 31260 22080 31266 22092
rect 32306 22080 32312 22092
rect 31260 22052 32312 22080
rect 31260 22040 31266 22052
rect 32306 22040 32312 22052
rect 32364 22040 32370 22092
rect 33318 22040 33324 22092
rect 33376 22080 33382 22092
rect 33376 22052 33456 22080
rect 33376 22040 33382 22052
rect 29779 21984 30604 22012
rect 29779 21981 29791 21984
rect 29733 21975 29791 21981
rect 29362 21944 29368 21956
rect 27448 21916 29368 21944
rect 26467 21913 26479 21916
rect 26421 21907 26479 21913
rect 29362 21904 29368 21916
rect 29420 21904 29426 21956
rect 31113 21947 31171 21953
rect 31113 21913 31125 21947
rect 31159 21944 31171 21947
rect 31202 21944 31208 21956
rect 31159 21916 31208 21944
rect 31159 21913 31171 21916
rect 31113 21907 31171 21913
rect 31202 21904 31208 21916
rect 31260 21944 31266 21956
rect 31386 21944 31392 21956
rect 31260 21916 31392 21944
rect 31260 21904 31266 21916
rect 31386 21904 31392 21916
rect 31444 21904 31450 21956
rect 32122 21904 32128 21956
rect 32180 21904 32186 21956
rect 33428 21953 33456 22052
rect 33502 22040 33508 22092
rect 33560 22040 33566 22092
rect 33612 22089 33640 22120
rect 33778 22108 33784 22120
rect 33836 22108 33842 22160
rect 34330 22108 34336 22160
rect 34388 22148 34394 22160
rect 35544 22148 35572 22188
rect 34388 22120 34560 22148
rect 34388 22108 34394 22120
rect 34532 22094 34560 22120
rect 35452 22120 35572 22148
rect 33597 22083 33655 22089
rect 33597 22049 33609 22083
rect 33643 22049 33655 22083
rect 33597 22043 33655 22049
rect 33870 22040 33876 22092
rect 33928 22080 33934 22092
rect 34057 22083 34115 22089
rect 34057 22080 34069 22083
rect 33928 22052 34069 22080
rect 33928 22040 33934 22052
rect 34057 22049 34069 22052
rect 34103 22049 34115 22083
rect 34532 22080 34652 22094
rect 35345 22083 35403 22089
rect 35345 22080 35357 22083
rect 34532 22066 35357 22080
rect 34624 22052 35357 22066
rect 34057 22043 34115 22049
rect 35345 22049 35357 22052
rect 35391 22080 35403 22083
rect 35452 22080 35480 22120
rect 35391 22052 35480 22080
rect 35529 22083 35587 22089
rect 35391 22049 35403 22052
rect 35345 22043 35403 22049
rect 35529 22049 35541 22083
rect 35575 22049 35587 22083
rect 35820 22080 35848 22188
rect 37540 22185 37552 22219
rect 37586 22216 37598 22219
rect 38562 22216 38568 22228
rect 37586 22188 38568 22216
rect 37586 22185 37598 22188
rect 37540 22179 37598 22185
rect 38562 22176 38568 22188
rect 38620 22176 38626 22228
rect 38838 22176 38844 22228
rect 38896 22216 38902 22228
rect 39758 22216 39764 22228
rect 38896 22188 39764 22216
rect 38896 22176 38902 22188
rect 39758 22176 39764 22188
rect 39816 22176 39822 22228
rect 40034 22176 40040 22228
rect 40092 22216 40098 22228
rect 41233 22219 41291 22225
rect 41233 22216 41245 22219
rect 40092 22188 41245 22216
rect 40092 22176 40098 22188
rect 41233 22185 41245 22188
rect 41279 22185 41291 22219
rect 43622 22216 43628 22228
rect 41233 22179 41291 22185
rect 42812 22188 43628 22216
rect 36740 22120 37412 22148
rect 36740 22089 36768 22120
rect 36725 22083 36783 22089
rect 35820 22052 36676 22080
rect 35529 22043 35587 22049
rect 35544 22012 35572 22043
rect 35894 22012 35900 22024
rect 35544 21984 35900 22012
rect 35894 21972 35900 21984
rect 35952 21972 35958 22024
rect 36648 22012 36676 22052
rect 36725 22049 36737 22083
rect 36771 22080 36783 22083
rect 37384 22080 37412 22120
rect 38746 22108 38752 22160
rect 38804 22148 38810 22160
rect 38804 22120 40632 22148
rect 38804 22108 38810 22120
rect 38286 22080 38292 22092
rect 36771 22052 36805 22080
rect 37384 22052 38292 22080
rect 36771 22049 36783 22052
rect 36725 22043 36783 22049
rect 38286 22040 38292 22052
rect 38344 22040 38350 22092
rect 38562 22040 38568 22092
rect 38620 22080 38626 22092
rect 40604 22089 40632 22120
rect 40770 22108 40776 22160
rect 40828 22148 40834 22160
rect 41046 22148 41052 22160
rect 40828 22120 41052 22148
rect 40828 22108 40834 22120
rect 41046 22108 41052 22120
rect 41104 22148 41110 22160
rect 42812 22148 42840 22188
rect 43622 22176 43628 22188
rect 43680 22216 43686 22228
rect 44545 22219 44603 22225
rect 44545 22216 44557 22219
rect 43680 22188 44557 22216
rect 43680 22176 43686 22188
rect 44545 22185 44557 22188
rect 44591 22185 44603 22219
rect 44545 22179 44603 22185
rect 44821 22219 44879 22225
rect 44821 22185 44833 22219
rect 44867 22216 44879 22219
rect 45554 22216 45560 22228
rect 44867 22188 45560 22216
rect 44867 22185 44879 22188
rect 44821 22179 44879 22185
rect 45554 22176 45560 22188
rect 45612 22176 45618 22228
rect 45646 22176 45652 22228
rect 45704 22216 45710 22228
rect 45704 22188 46152 22216
rect 45704 22176 45710 22188
rect 41104 22120 41828 22148
rect 41104 22108 41110 22120
rect 39025 22083 39083 22089
rect 39025 22080 39037 22083
rect 38620 22052 39037 22080
rect 38620 22040 38626 22052
rect 39025 22049 39037 22052
rect 39071 22049 39083 22083
rect 39025 22043 39083 22049
rect 40589 22083 40647 22089
rect 40589 22049 40601 22083
rect 40635 22049 40647 22083
rect 40589 22043 40647 22049
rect 40862 22040 40868 22092
rect 40920 22080 40926 22092
rect 41414 22080 41420 22092
rect 40920 22052 41420 22080
rect 40920 22040 40926 22052
rect 41414 22040 41420 22052
rect 41472 22040 41478 22092
rect 41800 22089 41828 22120
rect 42720 22120 42840 22148
rect 41785 22083 41843 22089
rect 41785 22049 41797 22083
rect 41831 22049 41843 22083
rect 41785 22043 41843 22049
rect 42334 22040 42340 22092
rect 42392 22080 42398 22092
rect 42429 22083 42487 22089
rect 42429 22080 42441 22083
rect 42392 22052 42441 22080
rect 42392 22040 42398 22052
rect 42429 22049 42441 22052
rect 42475 22049 42487 22083
rect 42429 22043 42487 22049
rect 37182 22012 37188 22024
rect 36648 21984 37188 22012
rect 37182 21972 37188 21984
rect 37240 21972 37246 22024
rect 37277 22015 37335 22021
rect 37277 21981 37289 22015
rect 37323 21981 37335 22015
rect 37277 21975 37335 21981
rect 33413 21947 33471 21953
rect 33413 21913 33425 21947
rect 33459 21913 33471 21947
rect 33413 21907 33471 21913
rect 34333 21947 34391 21953
rect 34333 21913 34345 21947
rect 34379 21944 34391 21947
rect 37292 21944 37320 21975
rect 39390 21972 39396 22024
rect 39448 22012 39454 22024
rect 39485 22015 39543 22021
rect 39485 22012 39497 22015
rect 39448 21984 39497 22012
rect 39448 21972 39454 21984
rect 39485 21981 39497 21984
rect 39531 22012 39543 22015
rect 42720 22012 42748 22120
rect 42886 22108 42892 22160
rect 42944 22108 42950 22160
rect 45189 22151 45247 22157
rect 45189 22117 45201 22151
rect 45235 22117 45247 22151
rect 46014 22148 46020 22160
rect 45189 22111 45247 22117
rect 45848 22120 46020 22148
rect 43530 22040 43536 22092
rect 43588 22040 43594 22092
rect 39531 21984 42748 22012
rect 43257 22015 43315 22021
rect 39531 21981 39543 21984
rect 39485 21975 39543 21981
rect 43257 21981 43269 22015
rect 43303 22012 43315 22015
rect 43346 22012 43352 22024
rect 43303 21984 43352 22012
rect 43303 21981 43315 21984
rect 43257 21975 43315 21981
rect 43346 21972 43352 21984
rect 43404 21972 43410 22024
rect 43714 21972 43720 22024
rect 43772 22012 43778 22024
rect 43772 21984 44680 22012
rect 43772 21972 43778 21984
rect 37458 21944 37464 21956
rect 34379 21916 36676 21944
rect 37292 21916 37464 21944
rect 34379 21913 34391 21916
rect 34333 21907 34391 21913
rect 25593 21879 25651 21885
rect 25593 21876 25605 21879
rect 25464 21848 25605 21876
rect 25464 21836 25470 21848
rect 25593 21845 25605 21848
rect 25639 21845 25651 21879
rect 25593 21839 25651 21845
rect 25961 21879 26019 21885
rect 25961 21845 25973 21879
rect 26007 21845 26019 21879
rect 25961 21839 26019 21845
rect 26326 21836 26332 21888
rect 26384 21836 26390 21888
rect 26694 21836 26700 21888
rect 26752 21876 26758 21888
rect 27157 21879 27215 21885
rect 27157 21876 27169 21879
rect 26752 21848 27169 21876
rect 26752 21836 26758 21848
rect 27157 21845 27169 21848
rect 27203 21845 27215 21879
rect 27157 21839 27215 21845
rect 27338 21836 27344 21888
rect 27396 21876 27402 21888
rect 27525 21879 27583 21885
rect 27525 21876 27537 21879
rect 27396 21848 27537 21876
rect 27396 21836 27402 21848
rect 27525 21845 27537 21848
rect 27571 21845 27583 21879
rect 27525 21839 27583 21845
rect 27617 21879 27675 21885
rect 27617 21845 27629 21879
rect 27663 21876 27675 21879
rect 28626 21876 28632 21888
rect 27663 21848 28632 21876
rect 27663 21845 27675 21848
rect 27617 21839 27675 21845
rect 28626 21836 28632 21848
rect 28684 21836 28690 21888
rect 28813 21879 28871 21885
rect 28813 21845 28825 21879
rect 28859 21876 28871 21879
rect 31754 21876 31760 21888
rect 28859 21848 31760 21876
rect 28859 21845 28871 21848
rect 28813 21839 28871 21845
rect 31754 21836 31760 21848
rect 31812 21836 31818 21888
rect 32674 21836 32680 21888
rect 32732 21876 32738 21888
rect 33045 21879 33103 21885
rect 33045 21876 33057 21879
rect 32732 21848 33057 21876
rect 32732 21836 32738 21848
rect 33045 21845 33057 21848
rect 33091 21845 33103 21879
rect 33045 21839 33103 21845
rect 33134 21836 33140 21888
rect 33192 21876 33198 21888
rect 34348 21876 34376 21907
rect 33192 21848 34376 21876
rect 33192 21836 33198 21848
rect 34514 21836 34520 21888
rect 34572 21836 34578 21888
rect 34885 21879 34943 21885
rect 34885 21845 34897 21879
rect 34931 21876 34943 21879
rect 35158 21876 35164 21888
rect 34931 21848 35164 21876
rect 34931 21845 34943 21848
rect 34885 21839 34943 21845
rect 35158 21836 35164 21848
rect 35216 21836 35222 21888
rect 35250 21836 35256 21888
rect 35308 21836 35314 21888
rect 36081 21879 36139 21885
rect 36081 21845 36093 21879
rect 36127 21876 36139 21879
rect 36170 21876 36176 21888
rect 36127 21848 36176 21876
rect 36127 21845 36139 21848
rect 36081 21839 36139 21845
rect 36170 21836 36176 21848
rect 36228 21836 36234 21888
rect 36446 21836 36452 21888
rect 36504 21836 36510 21888
rect 36538 21836 36544 21888
rect 36596 21836 36602 21888
rect 36648 21876 36676 21916
rect 37458 21904 37464 21916
rect 37516 21904 37522 21956
rect 37550 21904 37556 21956
rect 37608 21944 37614 21956
rect 37608 21916 38042 21944
rect 37608 21904 37614 21916
rect 39574 21904 39580 21956
rect 39632 21904 39638 21956
rect 40405 21947 40463 21953
rect 40405 21913 40417 21947
rect 40451 21944 40463 21947
rect 40586 21944 40592 21956
rect 40451 21916 40592 21944
rect 40451 21913 40463 21916
rect 40405 21907 40463 21913
rect 40586 21904 40592 21916
rect 40644 21944 40650 21956
rect 44453 21947 44511 21953
rect 44453 21944 44465 21947
rect 40644 21916 44465 21944
rect 40644 21904 40650 21916
rect 44453 21913 44465 21916
rect 44499 21944 44511 21947
rect 44542 21944 44548 21956
rect 44499 21916 44548 21944
rect 44499 21913 44511 21916
rect 44453 21907 44511 21913
rect 44542 21904 44548 21916
rect 44600 21904 44606 21956
rect 44652 21944 44680 21984
rect 45204 22008 45232 22111
rect 45848 22089 45876 22120
rect 46014 22108 46020 22120
rect 46072 22108 46078 22160
rect 46124 22148 46152 22188
rect 47302 22176 47308 22228
rect 47360 22216 47366 22228
rect 47857 22219 47915 22225
rect 47857 22216 47869 22219
rect 47360 22188 47869 22216
rect 47360 22176 47366 22188
rect 47857 22185 47869 22188
rect 47903 22216 47915 22219
rect 49234 22216 49240 22228
rect 47903 22188 49240 22216
rect 47903 22185 47915 22188
rect 47857 22179 47915 22185
rect 49234 22176 49240 22188
rect 49292 22176 49298 22228
rect 47581 22151 47639 22157
rect 47581 22148 47593 22151
rect 46124 22120 47593 22148
rect 47581 22117 47593 22120
rect 47627 22117 47639 22151
rect 47581 22111 47639 22117
rect 45833 22083 45891 22089
rect 45833 22049 45845 22083
rect 45879 22049 45891 22083
rect 45833 22043 45891 22049
rect 48041 22083 48099 22089
rect 48041 22049 48053 22083
rect 48087 22080 48099 22083
rect 48590 22080 48596 22092
rect 48087 22052 48596 22080
rect 48087 22049 48099 22052
rect 48041 22043 48099 22049
rect 48590 22040 48596 22052
rect 48648 22040 48654 22092
rect 45278 22008 45284 22024
rect 45204 21980 45284 22008
rect 45278 21972 45284 21980
rect 45336 21972 45342 22024
rect 45373 22015 45431 22021
rect 45373 21981 45385 22015
rect 45419 22012 45431 22015
rect 45646 22012 45652 22024
rect 45419 21984 45652 22012
rect 45419 21981 45431 21984
rect 45373 21975 45431 21981
rect 45646 21972 45652 21984
rect 45704 21972 45710 22024
rect 45738 21972 45744 22024
rect 45796 22012 45802 22024
rect 46109 22015 46167 22021
rect 46109 22012 46121 22015
rect 45796 21984 46121 22012
rect 45796 21972 45802 21984
rect 46109 21981 46121 21984
rect 46155 21981 46167 22015
rect 46109 21975 46167 21981
rect 47302 21972 47308 22024
rect 47360 21972 47366 22024
rect 48317 22015 48375 22021
rect 48317 21981 48329 22015
rect 48363 22012 48375 22015
rect 49050 22012 49056 22024
rect 48363 21984 49056 22012
rect 48363 21981 48375 21984
rect 48317 21975 48375 21981
rect 49050 21972 49056 21984
rect 49108 21972 49114 22024
rect 44652 21916 45232 21944
rect 37274 21876 37280 21888
rect 36648 21848 37280 21876
rect 37274 21836 37280 21848
rect 37332 21836 37338 21888
rect 40034 21836 40040 21888
rect 40092 21836 40098 21888
rect 40494 21836 40500 21888
rect 40552 21836 40558 21888
rect 41506 21836 41512 21888
rect 41564 21876 41570 21888
rect 41601 21879 41659 21885
rect 41601 21876 41613 21879
rect 41564 21848 41613 21876
rect 41564 21836 41570 21848
rect 41601 21845 41613 21848
rect 41647 21845 41659 21879
rect 41601 21839 41659 21845
rect 41690 21836 41696 21888
rect 41748 21876 41754 21888
rect 43438 21876 43444 21888
rect 41748 21848 43444 21876
rect 41748 21836 41754 21848
rect 43438 21836 43444 21848
rect 43496 21836 43502 21888
rect 45204 21876 45232 21916
rect 45462 21904 45468 21956
rect 45520 21944 45526 21956
rect 45520 21916 48544 21944
rect 45520 21904 45526 21916
rect 48516 21885 48544 21916
rect 49142 21904 49148 21956
rect 49200 21904 49206 21956
rect 49329 21947 49387 21953
rect 49329 21913 49341 21947
rect 49375 21944 49387 21947
rect 49418 21944 49424 21956
rect 49375 21916 49424 21944
rect 49375 21913 49387 21916
rect 49329 21907 49387 21913
rect 49418 21904 49424 21916
rect 49476 21904 49482 21956
rect 47121 21879 47179 21885
rect 47121 21876 47133 21879
rect 45204 21848 47133 21876
rect 47121 21845 47133 21848
rect 47167 21845 47179 21879
rect 47121 21839 47179 21845
rect 48501 21879 48559 21885
rect 48501 21845 48513 21879
rect 48547 21845 48559 21879
rect 48501 21839 48559 21845
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 5261 21675 5319 21681
rect 5261 21641 5273 21675
rect 5307 21672 5319 21675
rect 9214 21672 9220 21684
rect 5307 21644 9220 21672
rect 5307 21641 5319 21644
rect 5261 21635 5319 21641
rect 9214 21632 9220 21644
rect 9272 21632 9278 21684
rect 11790 21632 11796 21684
rect 11848 21632 11854 21684
rect 13173 21675 13231 21681
rect 13173 21641 13185 21675
rect 13219 21672 13231 21675
rect 13354 21672 13360 21684
rect 13219 21644 13360 21672
rect 13219 21641 13231 21644
rect 13173 21635 13231 21641
rect 13354 21632 13360 21644
rect 13412 21632 13418 21684
rect 14734 21632 14740 21684
rect 14792 21632 14798 21684
rect 15102 21632 15108 21684
rect 15160 21632 15166 21684
rect 15562 21632 15568 21684
rect 15620 21672 15626 21684
rect 16209 21675 16267 21681
rect 16209 21672 16221 21675
rect 15620 21644 16221 21672
rect 15620 21632 15626 21644
rect 16209 21641 16221 21644
rect 16255 21641 16267 21675
rect 16209 21635 16267 21641
rect 17313 21675 17371 21681
rect 17313 21641 17325 21675
rect 17359 21672 17371 21675
rect 20622 21672 20628 21684
rect 17359 21644 20628 21672
rect 17359 21641 17371 21644
rect 17313 21635 17371 21641
rect 20622 21632 20628 21644
rect 20680 21632 20686 21684
rect 21085 21675 21143 21681
rect 21085 21641 21097 21675
rect 21131 21672 21143 21675
rect 22278 21672 22284 21684
rect 21131 21644 22284 21672
rect 21131 21641 21143 21644
rect 21085 21635 21143 21641
rect 22278 21632 22284 21644
rect 22336 21632 22342 21684
rect 25130 21632 25136 21684
rect 25188 21632 25194 21684
rect 27154 21632 27160 21684
rect 27212 21632 27218 21684
rect 28353 21675 28411 21681
rect 28353 21641 28365 21675
rect 28399 21672 28411 21675
rect 28534 21672 28540 21684
rect 28399 21644 28540 21672
rect 28399 21641 28411 21644
rect 28353 21635 28411 21641
rect 28534 21632 28540 21644
rect 28592 21632 28598 21684
rect 28718 21632 28724 21684
rect 28776 21632 28782 21684
rect 29917 21675 29975 21681
rect 29917 21641 29929 21675
rect 29963 21672 29975 21675
rect 31754 21672 31760 21684
rect 29963 21644 31760 21672
rect 29963 21641 29975 21644
rect 29917 21635 29975 21641
rect 31754 21632 31760 21644
rect 31812 21632 31818 21684
rect 31849 21675 31907 21681
rect 31849 21641 31861 21675
rect 31895 21672 31907 21675
rect 32122 21672 32128 21684
rect 31895 21644 32128 21672
rect 31895 21641 31907 21644
rect 31849 21635 31907 21641
rect 32122 21632 32128 21644
rect 32180 21632 32186 21684
rect 32398 21632 32404 21684
rect 32456 21672 32462 21684
rect 35802 21672 35808 21684
rect 32456 21644 35808 21672
rect 32456 21632 32462 21644
rect 35802 21632 35808 21644
rect 35860 21632 35866 21684
rect 36081 21675 36139 21681
rect 36081 21641 36093 21675
rect 36127 21672 36139 21675
rect 40034 21672 40040 21684
rect 36127 21644 40040 21672
rect 36127 21641 36139 21644
rect 36081 21635 36139 21641
rect 40034 21632 40040 21644
rect 40092 21632 40098 21684
rect 40126 21632 40132 21684
rect 40184 21672 40190 21684
rect 40221 21675 40279 21681
rect 40221 21672 40233 21675
rect 40184 21644 40233 21672
rect 40184 21632 40190 21644
rect 40221 21641 40233 21644
rect 40267 21641 40279 21675
rect 40221 21635 40279 21641
rect 40328 21644 41460 21672
rect 1762 21564 1768 21616
rect 1820 21604 1826 21616
rect 3970 21604 3976 21616
rect 1820 21576 3976 21604
rect 1820 21564 1826 21576
rect 3970 21564 3976 21576
rect 4028 21564 4034 21616
rect 4246 21564 4252 21616
rect 4304 21604 4310 21616
rect 4341 21607 4399 21613
rect 4341 21604 4353 21607
rect 4304 21576 4353 21604
rect 4304 21564 4310 21576
rect 4341 21573 4353 21576
rect 4387 21573 4399 21607
rect 4341 21567 4399 21573
rect 5350 21564 5356 21616
rect 5408 21604 5414 21616
rect 5408 21576 6592 21604
rect 5408 21564 5414 21576
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 3418 21536 3424 21548
rect 1719 21508 3424 21536
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 3418 21496 3424 21508
rect 3476 21496 3482 21548
rect 3605 21539 3663 21545
rect 3605 21505 3617 21539
rect 3651 21536 3663 21539
rect 5074 21536 5080 21548
rect 3651 21508 5080 21536
rect 3651 21505 3663 21508
rect 3605 21499 3663 21505
rect 5074 21496 5080 21508
rect 5132 21496 5138 21548
rect 5166 21496 5172 21548
rect 5224 21536 5230 21548
rect 6564 21545 6592 21576
rect 7742 21564 7748 21616
rect 7800 21604 7806 21616
rect 10318 21604 10324 21616
rect 7800 21576 10324 21604
rect 7800 21564 7806 21576
rect 10318 21564 10324 21576
rect 10376 21564 10382 21616
rect 17034 21604 17040 21616
rect 10520 21576 17040 21604
rect 5813 21539 5871 21545
rect 5813 21536 5825 21539
rect 5224 21508 5825 21536
rect 5224 21496 5230 21508
rect 5813 21505 5825 21508
rect 5859 21505 5871 21539
rect 5813 21499 5871 21505
rect 6549 21539 6607 21545
rect 6549 21505 6561 21539
rect 6595 21505 6607 21539
rect 6549 21499 6607 21505
rect 7282 21496 7288 21548
rect 7340 21536 7346 21548
rect 10520 21545 10548 21576
rect 17034 21564 17040 21576
rect 17092 21564 17098 21616
rect 17126 21564 17132 21616
rect 17184 21604 17190 21616
rect 20070 21604 20076 21616
rect 17184 21576 17448 21604
rect 19550 21576 20076 21604
rect 17184 21564 17190 21576
rect 8389 21539 8447 21545
rect 8389 21536 8401 21539
rect 7340 21508 8401 21536
rect 7340 21496 7346 21508
rect 8389 21505 8401 21508
rect 8435 21505 8447 21539
rect 10505 21539 10563 21545
rect 8389 21499 8447 21505
rect 8496 21508 8984 21536
rect 1394 21428 1400 21480
rect 1452 21468 1458 21480
rect 2041 21471 2099 21477
rect 2041 21468 2053 21471
rect 1452 21440 2053 21468
rect 1452 21428 1458 21440
rect 2041 21437 2053 21440
rect 2087 21437 2099 21471
rect 2041 21431 2099 21437
rect 4338 21428 4344 21480
rect 4396 21468 4402 21480
rect 5997 21471 6055 21477
rect 5997 21468 6009 21471
rect 4396 21440 6009 21468
rect 4396 21428 4402 21440
rect 5997 21437 6009 21440
rect 6043 21437 6055 21471
rect 5997 21431 6055 21437
rect 6638 21428 6644 21480
rect 6696 21468 6702 21480
rect 7009 21471 7067 21477
rect 7009 21468 7021 21471
rect 6696 21440 7021 21468
rect 6696 21428 6702 21440
rect 7009 21437 7021 21440
rect 7055 21437 7067 21471
rect 7009 21431 7067 21437
rect 7834 21428 7840 21480
rect 7892 21468 7898 21480
rect 8496 21468 8524 21508
rect 8849 21471 8907 21477
rect 8849 21468 8861 21471
rect 7892 21440 8524 21468
rect 8588 21440 8861 21468
rect 7892 21428 7898 21440
rect 5442 21360 5448 21412
rect 5500 21360 5506 21412
rect 3602 21292 3608 21344
rect 3660 21332 3666 21344
rect 8588 21332 8616 21440
rect 8849 21437 8861 21440
rect 8895 21437 8907 21471
rect 8849 21431 8907 21437
rect 8956 21400 8984 21508
rect 10505 21505 10517 21539
rect 10551 21505 10563 21539
rect 10505 21499 10563 21505
rect 11974 21496 11980 21548
rect 12032 21496 12038 21548
rect 12529 21539 12587 21545
rect 12529 21505 12541 21539
rect 12575 21505 12587 21539
rect 12529 21499 12587 21505
rect 9766 21428 9772 21480
rect 9824 21468 9830 21480
rect 10318 21468 10324 21480
rect 9824 21440 10324 21468
rect 9824 21428 9830 21440
rect 10318 21428 10324 21440
rect 10376 21428 10382 21480
rect 11146 21428 11152 21480
rect 11204 21428 11210 21480
rect 12544 21468 12572 21499
rect 13630 21496 13636 21548
rect 13688 21496 13694 21548
rect 14918 21496 14924 21548
rect 14976 21536 14982 21548
rect 15197 21539 15255 21545
rect 15197 21536 15209 21539
rect 14976 21508 15209 21536
rect 14976 21496 14982 21508
rect 15197 21505 15209 21508
rect 15243 21505 15255 21539
rect 15197 21499 15255 21505
rect 16114 21496 16120 21548
rect 16172 21496 16178 21548
rect 17218 21496 17224 21548
rect 17276 21496 17282 21548
rect 15010 21468 15016 21480
rect 12544 21440 15016 21468
rect 15010 21428 15016 21440
rect 15068 21428 15074 21480
rect 15286 21428 15292 21480
rect 15344 21428 15350 21480
rect 17420 21477 17448 21576
rect 20070 21564 20076 21576
rect 20128 21564 20134 21616
rect 20438 21564 20444 21616
rect 20496 21604 20502 21616
rect 23014 21604 23020 21616
rect 20496 21576 23020 21604
rect 20496 21564 20502 21576
rect 23014 21564 23020 21576
rect 23072 21564 23078 21616
rect 23382 21564 23388 21616
rect 23440 21564 23446 21616
rect 27617 21607 27675 21613
rect 27617 21573 27629 21607
rect 27663 21604 27675 21607
rect 28166 21604 28172 21616
rect 27663 21576 28172 21604
rect 27663 21573 27675 21576
rect 27617 21567 27675 21573
rect 28166 21564 28172 21576
rect 28224 21564 28230 21616
rect 28626 21564 28632 21616
rect 28684 21604 28690 21616
rect 29270 21604 29276 21616
rect 28684 21576 29276 21604
rect 28684 21564 28690 21576
rect 29270 21564 29276 21576
rect 29328 21564 29334 21616
rect 30009 21607 30067 21613
rect 30009 21573 30021 21607
rect 30055 21604 30067 21607
rect 30190 21604 30196 21616
rect 30055 21576 30196 21604
rect 30055 21573 30067 21576
rect 30009 21567 30067 21573
rect 30190 21564 30196 21576
rect 30248 21564 30254 21616
rect 31113 21607 31171 21613
rect 31113 21573 31125 21607
rect 31159 21604 31171 21607
rect 31159 21576 33640 21604
rect 31159 21573 31171 21576
rect 31113 21567 31171 21573
rect 33612 21548 33640 21576
rect 34238 21564 34244 21616
rect 34296 21604 34302 21616
rect 34885 21607 34943 21613
rect 34885 21604 34897 21607
rect 34296 21576 34897 21604
rect 34296 21564 34302 21576
rect 34885 21573 34897 21576
rect 34931 21604 34943 21607
rect 34974 21604 34980 21616
rect 34931 21576 34980 21604
rect 34931 21573 34943 21576
rect 34885 21567 34943 21573
rect 34974 21564 34980 21576
rect 35032 21564 35038 21616
rect 35986 21564 35992 21616
rect 36044 21604 36050 21616
rect 36906 21604 36912 21616
rect 36044 21576 36912 21604
rect 36044 21564 36050 21576
rect 36906 21564 36912 21576
rect 36964 21604 36970 21616
rect 37550 21604 37556 21616
rect 36964 21576 37556 21604
rect 36964 21564 36970 21576
rect 37550 21564 37556 21576
rect 37608 21604 37614 21616
rect 37645 21607 37703 21613
rect 37645 21604 37657 21607
rect 37608 21576 37657 21604
rect 37608 21564 37614 21576
rect 37645 21573 37657 21576
rect 37691 21604 37703 21607
rect 38562 21604 38568 21616
rect 37691 21576 38568 21604
rect 37691 21573 37703 21576
rect 37645 21567 37703 21573
rect 38562 21564 38568 21576
rect 38620 21564 38626 21616
rect 38746 21564 38752 21616
rect 38804 21564 38810 21616
rect 21177 21539 21235 21545
rect 21177 21505 21189 21539
rect 21223 21536 21235 21539
rect 21266 21536 21272 21548
rect 21223 21508 21272 21536
rect 21223 21505 21235 21508
rect 21177 21499 21235 21505
rect 21266 21496 21272 21508
rect 21324 21496 21330 21548
rect 21542 21536 21548 21548
rect 21376 21508 21548 21536
rect 17405 21471 17463 21477
rect 17405 21437 17417 21471
rect 17451 21437 17463 21471
rect 17405 21431 17463 21437
rect 17954 21428 17960 21480
rect 18012 21468 18018 21480
rect 18049 21471 18107 21477
rect 18049 21468 18061 21471
rect 18012 21440 18061 21468
rect 18012 21428 18018 21440
rect 18049 21437 18061 21440
rect 18095 21437 18107 21471
rect 18325 21471 18383 21477
rect 18325 21468 18337 21471
rect 18049 21431 18107 21437
rect 18156 21440 18337 21468
rect 14277 21403 14335 21409
rect 8956 21372 12434 21400
rect 3660 21304 8616 21332
rect 3660 21292 3666 21304
rect 9582 21292 9588 21344
rect 9640 21332 9646 21344
rect 10137 21335 10195 21341
rect 10137 21332 10149 21335
rect 9640 21304 10149 21332
rect 9640 21292 9646 21304
rect 10137 21301 10149 21304
rect 10183 21301 10195 21335
rect 12406 21332 12434 21372
rect 14277 21369 14289 21403
rect 14323 21400 14335 21403
rect 18156 21400 18184 21440
rect 18325 21437 18337 21440
rect 18371 21437 18383 21471
rect 18325 21431 18383 21437
rect 20162 21428 20168 21480
rect 20220 21468 20226 21480
rect 20622 21468 20628 21480
rect 20220 21440 20628 21468
rect 20220 21428 20226 21440
rect 20622 21428 20628 21440
rect 20680 21428 20686 21480
rect 21376 21477 21404 21508
rect 21542 21496 21548 21508
rect 21600 21496 21606 21548
rect 21910 21496 21916 21548
rect 21968 21496 21974 21548
rect 22002 21496 22008 21548
rect 22060 21536 22066 21548
rect 22465 21539 22523 21545
rect 22465 21536 22477 21539
rect 22060 21508 22477 21536
rect 22060 21496 22066 21508
rect 22465 21505 22477 21508
rect 22511 21505 22523 21539
rect 22465 21499 22523 21505
rect 25148 21508 25360 21536
rect 21361 21471 21419 21477
rect 21361 21437 21373 21471
rect 21407 21437 21419 21471
rect 22741 21471 22799 21477
rect 22741 21468 22753 21471
rect 21361 21431 21419 21437
rect 22388 21440 22753 21468
rect 22388 21412 22416 21440
rect 22741 21437 22753 21440
rect 22787 21437 22799 21471
rect 22741 21431 22799 21437
rect 23290 21428 23296 21480
rect 23348 21468 23354 21480
rect 25148 21468 25176 21508
rect 23348 21440 25176 21468
rect 23348 21428 23354 21440
rect 25222 21428 25228 21480
rect 25280 21428 25286 21480
rect 25332 21477 25360 21508
rect 25958 21496 25964 21548
rect 26016 21496 26022 21548
rect 26602 21496 26608 21548
rect 26660 21496 26666 21548
rect 27525 21539 27583 21545
rect 27525 21505 27537 21539
rect 27571 21536 27583 21539
rect 29086 21536 29092 21548
rect 27571 21508 29092 21536
rect 27571 21505 27583 21508
rect 27525 21499 27583 21505
rect 29086 21496 29092 21508
rect 29144 21536 29150 21548
rect 29546 21536 29552 21548
rect 29144 21508 29552 21536
rect 29144 21496 29150 21508
rect 29546 21496 29552 21508
rect 29604 21496 29610 21548
rect 31205 21539 31263 21545
rect 31205 21505 31217 21539
rect 31251 21536 31263 21539
rect 31251 21508 33548 21536
rect 31251 21505 31263 21508
rect 31205 21499 31263 21505
rect 25317 21471 25375 21477
rect 25317 21437 25329 21471
rect 25363 21468 25375 21471
rect 27709 21471 27767 21477
rect 27709 21468 27721 21471
rect 25363 21440 27721 21468
rect 25363 21437 25375 21440
rect 25317 21431 25375 21437
rect 27709 21437 27721 21440
rect 27755 21437 27767 21471
rect 27709 21431 27767 21437
rect 28166 21428 28172 21480
rect 28224 21468 28230 21480
rect 28626 21468 28632 21480
rect 28224 21440 28632 21468
rect 28224 21428 28230 21440
rect 28626 21428 28632 21440
rect 28684 21428 28690 21480
rect 28810 21428 28816 21480
rect 28868 21428 28874 21480
rect 28902 21428 28908 21480
rect 28960 21428 28966 21480
rect 29454 21428 29460 21480
rect 29512 21468 29518 21480
rect 30101 21471 30159 21477
rect 30101 21468 30113 21471
rect 29512 21440 30113 21468
rect 29512 21428 29518 21440
rect 30101 21437 30113 21440
rect 30147 21437 30159 21471
rect 30101 21431 30159 21437
rect 30742 21428 30748 21480
rect 30800 21468 30806 21480
rect 31294 21468 31300 21480
rect 30800 21440 31300 21468
rect 30800 21428 30806 21440
rect 31294 21428 31300 21440
rect 31352 21428 31358 21480
rect 32030 21428 32036 21480
rect 32088 21468 32094 21480
rect 32309 21471 32367 21477
rect 32309 21468 32321 21471
rect 32088 21440 32321 21468
rect 32088 21428 32094 21440
rect 32309 21437 32321 21440
rect 32355 21437 32367 21471
rect 32309 21431 32367 21437
rect 32490 21428 32496 21480
rect 32548 21468 32554 21480
rect 33042 21468 33048 21480
rect 32548 21440 33048 21468
rect 32548 21428 32554 21440
rect 33042 21428 33048 21440
rect 33100 21428 33106 21480
rect 33520 21468 33548 21508
rect 33594 21496 33600 21548
rect 33652 21496 33658 21548
rect 33796 21508 34376 21536
rect 33686 21468 33692 21480
rect 33520 21440 33692 21468
rect 33686 21428 33692 21440
rect 33744 21428 33750 21480
rect 14323 21372 18184 21400
rect 14323 21369 14335 21372
rect 14277 21363 14335 21369
rect 20070 21360 20076 21412
rect 20128 21400 20134 21412
rect 20257 21403 20315 21409
rect 20257 21400 20269 21403
rect 20128 21372 20269 21400
rect 20128 21360 20134 21372
rect 20257 21369 20269 21372
rect 20303 21400 20315 21403
rect 20303 21372 20852 21400
rect 20303 21369 20315 21372
rect 20257 21363 20315 21369
rect 15746 21332 15752 21344
rect 12406 21304 15752 21332
rect 10137 21295 10195 21301
rect 15746 21292 15752 21304
rect 15804 21292 15810 21344
rect 16850 21292 16856 21344
rect 16908 21292 16914 21344
rect 17494 21292 17500 21344
rect 17552 21332 17558 21344
rect 19797 21335 19855 21341
rect 19797 21332 19809 21335
rect 17552 21304 19809 21332
rect 17552 21292 17558 21304
rect 19797 21301 19809 21304
rect 19843 21301 19855 21335
rect 19797 21295 19855 21301
rect 20346 21292 20352 21344
rect 20404 21292 20410 21344
rect 20530 21292 20536 21344
rect 20588 21332 20594 21344
rect 20717 21335 20775 21341
rect 20717 21332 20729 21335
rect 20588 21304 20729 21332
rect 20588 21292 20594 21304
rect 20717 21301 20729 21304
rect 20763 21301 20775 21335
rect 20824 21332 20852 21372
rect 22370 21360 22376 21412
rect 22428 21360 22434 21412
rect 24213 21403 24271 21409
rect 24213 21369 24225 21403
rect 24259 21400 24271 21403
rect 24259 21372 24900 21400
rect 24259 21369 24271 21372
rect 24213 21363 24271 21369
rect 21910 21332 21916 21344
rect 20824 21304 21916 21332
rect 20717 21295 20775 21301
rect 21910 21292 21916 21304
rect 21968 21292 21974 21344
rect 22094 21292 22100 21344
rect 22152 21292 22158 21344
rect 24762 21292 24768 21344
rect 24820 21292 24826 21344
rect 24872 21332 24900 21372
rect 26142 21360 26148 21412
rect 26200 21400 26206 21412
rect 29549 21403 29607 21409
rect 29549 21400 29561 21403
rect 26200 21372 29561 21400
rect 26200 21360 26206 21372
rect 29549 21369 29561 21372
rect 29595 21369 29607 21403
rect 29549 21363 29607 21369
rect 30834 21360 30840 21412
rect 30892 21400 30898 21412
rect 32769 21403 32827 21409
rect 32769 21400 32781 21403
rect 30892 21372 32781 21400
rect 30892 21360 30898 21372
rect 32769 21369 32781 21372
rect 32815 21369 32827 21403
rect 32769 21363 32827 21369
rect 33229 21403 33287 21409
rect 33229 21369 33241 21403
rect 33275 21400 33287 21403
rect 33796 21400 33824 21508
rect 33873 21471 33931 21477
rect 33873 21437 33885 21471
rect 33919 21437 33931 21471
rect 33873 21431 33931 21437
rect 33275 21372 33824 21400
rect 33275 21369 33287 21372
rect 33229 21363 33287 21369
rect 29362 21332 29368 21344
rect 24872 21304 29368 21332
rect 29362 21292 29368 21304
rect 29420 21332 29426 21344
rect 30190 21332 30196 21344
rect 29420 21304 30196 21332
rect 29420 21292 29426 21304
rect 30190 21292 30196 21304
rect 30248 21292 30254 21344
rect 30466 21292 30472 21344
rect 30524 21332 30530 21344
rect 30745 21335 30803 21341
rect 30745 21332 30757 21335
rect 30524 21304 30757 21332
rect 30524 21292 30530 21304
rect 30745 21301 30757 21304
rect 30791 21301 30803 21335
rect 30745 21295 30803 21301
rect 31754 21292 31760 21344
rect 31812 21332 31818 21344
rect 32490 21332 32496 21344
rect 31812 21304 32496 21332
rect 31812 21292 31818 21304
rect 32490 21292 32496 21304
rect 32548 21292 32554 21344
rect 32582 21292 32588 21344
rect 32640 21332 32646 21344
rect 33888 21332 33916 21431
rect 34348 21400 34376 21508
rect 34422 21496 34428 21548
rect 34480 21536 34486 21548
rect 34790 21536 34796 21548
rect 34480 21508 34796 21536
rect 34480 21496 34486 21508
rect 34790 21496 34796 21508
rect 34848 21496 34854 21548
rect 35069 21471 35127 21477
rect 35069 21437 35081 21471
rect 35115 21468 35127 21471
rect 35115 21440 35296 21468
rect 35115 21437 35127 21440
rect 35069 21431 35127 21437
rect 35158 21400 35164 21412
rect 34348 21372 35164 21400
rect 35158 21360 35164 21372
rect 35216 21360 35222 21412
rect 35268 21400 35296 21440
rect 36170 21428 36176 21480
rect 36228 21428 36234 21480
rect 36357 21471 36415 21477
rect 36357 21437 36369 21471
rect 36403 21468 36415 21471
rect 36630 21468 36636 21480
rect 36403 21440 36636 21468
rect 36403 21437 36415 21440
rect 36357 21431 36415 21437
rect 36630 21428 36636 21440
rect 36688 21428 36694 21480
rect 37642 21428 37648 21480
rect 37700 21468 37706 21480
rect 38013 21471 38071 21477
rect 38013 21468 38025 21471
rect 37700 21440 38025 21468
rect 37700 21428 37706 21440
rect 38013 21437 38025 21440
rect 38059 21437 38071 21471
rect 38289 21471 38347 21477
rect 38289 21468 38301 21471
rect 38013 21431 38071 21437
rect 38120 21440 38301 21468
rect 37461 21403 37519 21409
rect 37461 21400 37473 21403
rect 35268 21372 36400 21400
rect 36372 21344 36400 21372
rect 36832 21372 37473 21400
rect 36832 21344 36860 21372
rect 37461 21369 37473 21372
rect 37507 21400 37519 21403
rect 37734 21400 37740 21412
rect 37507 21372 37740 21400
rect 37507 21369 37519 21372
rect 37461 21363 37519 21369
rect 37734 21360 37740 21372
rect 37792 21360 37798 21412
rect 32640 21304 33916 21332
rect 34425 21335 34483 21341
rect 32640 21292 32646 21304
rect 34425 21301 34437 21335
rect 34471 21332 34483 21335
rect 35434 21332 35440 21344
rect 34471 21304 35440 21332
rect 34471 21301 34483 21304
rect 34425 21295 34483 21301
rect 35434 21292 35440 21304
rect 35492 21292 35498 21344
rect 35710 21292 35716 21344
rect 35768 21292 35774 21344
rect 36354 21292 36360 21344
rect 36412 21292 36418 21344
rect 36814 21292 36820 21344
rect 36872 21292 36878 21344
rect 37366 21292 37372 21344
rect 37424 21292 37430 21344
rect 37550 21292 37556 21344
rect 37608 21332 37614 21344
rect 38120 21332 38148 21440
rect 38289 21437 38301 21440
rect 38335 21468 38347 21471
rect 38378 21468 38384 21480
rect 38335 21440 38384 21468
rect 38335 21437 38347 21440
rect 38289 21431 38347 21437
rect 38378 21428 38384 21440
rect 38436 21468 38442 21480
rect 39022 21468 39028 21480
rect 38436 21440 39028 21468
rect 38436 21428 38442 21440
rect 39022 21428 39028 21440
rect 39080 21428 39086 21480
rect 39298 21428 39304 21480
rect 39356 21468 39362 21480
rect 40328 21468 40356 21644
rect 41432 21545 41460 21644
rect 42242 21632 42248 21684
rect 42300 21672 42306 21684
rect 42886 21672 42892 21684
rect 42300 21644 42892 21672
rect 42300 21632 42306 21644
rect 42886 21632 42892 21644
rect 42944 21632 42950 21684
rect 43254 21632 43260 21684
rect 43312 21672 43318 21684
rect 45278 21672 45284 21684
rect 43312 21644 45284 21672
rect 43312 21632 43318 21644
rect 45278 21632 45284 21644
rect 45336 21632 45342 21684
rect 45554 21632 45560 21684
rect 45612 21672 45618 21684
rect 46293 21675 46351 21681
rect 46293 21672 46305 21675
rect 45612 21644 46305 21672
rect 45612 21632 45618 21644
rect 46293 21641 46305 21644
rect 46339 21641 46351 21675
rect 46293 21635 46351 21641
rect 47394 21632 47400 21684
rect 47452 21672 47458 21684
rect 47949 21675 48007 21681
rect 47949 21672 47961 21675
rect 47452 21644 47961 21672
rect 47452 21632 47458 21644
rect 47949 21641 47961 21644
rect 47995 21672 48007 21675
rect 48222 21672 48228 21684
rect 47995 21644 48228 21672
rect 47995 21641 48007 21644
rect 47949 21635 48007 21641
rect 48222 21632 48228 21644
rect 48280 21632 48286 21684
rect 41506 21564 41512 21616
rect 41564 21604 41570 21616
rect 41564 21576 44220 21604
rect 41564 21564 41570 21576
rect 40589 21539 40647 21545
rect 40589 21505 40601 21539
rect 40635 21536 40647 21539
rect 41417 21539 41475 21545
rect 40635 21508 41000 21536
rect 40635 21505 40647 21508
rect 40589 21499 40647 21505
rect 40678 21468 40684 21480
rect 39356 21440 40356 21468
rect 40420 21440 40684 21468
rect 39356 21428 39362 21440
rect 39390 21360 39396 21412
rect 39448 21400 39454 21412
rect 40420 21400 40448 21440
rect 40678 21428 40684 21440
rect 40736 21428 40742 21480
rect 40770 21428 40776 21480
rect 40828 21428 40834 21480
rect 40972 21468 41000 21508
rect 41417 21505 41429 21539
rect 41463 21505 41475 21539
rect 41417 21499 41475 21505
rect 42613 21539 42671 21545
rect 42613 21505 42625 21539
rect 42659 21505 42671 21539
rect 42613 21499 42671 21505
rect 41506 21468 41512 21480
rect 40972 21440 41512 21468
rect 41506 21428 41512 21440
rect 41564 21468 41570 21480
rect 42242 21468 42248 21480
rect 41564 21440 42248 21468
rect 41564 21428 41570 21440
rect 42242 21428 42248 21440
rect 42300 21428 42306 21480
rect 42628 21400 42656 21499
rect 43898 21496 43904 21548
rect 43956 21496 43962 21548
rect 44192 21468 44220 21576
rect 44266 21564 44272 21616
rect 44324 21604 44330 21616
rect 44818 21604 44824 21616
rect 44324 21576 44824 21604
rect 44324 21564 44330 21576
rect 44818 21564 44824 21576
rect 44876 21604 44882 21616
rect 47581 21607 47639 21613
rect 47581 21604 47593 21607
rect 44876 21576 45232 21604
rect 44876 21564 44882 21576
rect 44542 21496 44548 21548
rect 44600 21496 44606 21548
rect 44726 21496 44732 21548
rect 44784 21536 44790 21548
rect 45002 21536 45008 21548
rect 44784 21508 45008 21536
rect 44784 21496 44790 21508
rect 45002 21496 45008 21508
rect 45060 21496 45066 21548
rect 45204 21545 45232 21576
rect 46492 21576 47593 21604
rect 45189 21539 45247 21545
rect 45189 21505 45201 21539
rect 45235 21505 45247 21539
rect 45189 21499 45247 21505
rect 45830 21496 45836 21548
rect 45888 21496 45894 21548
rect 45922 21496 45928 21548
rect 45980 21536 45986 21548
rect 46492 21545 46520 21576
rect 47581 21573 47593 21576
rect 47627 21573 47639 21607
rect 47581 21567 47639 21573
rect 48409 21607 48467 21613
rect 48409 21573 48421 21607
rect 48455 21604 48467 21607
rect 48590 21604 48596 21616
rect 48455 21576 48596 21604
rect 48455 21573 48467 21576
rect 48409 21567 48467 21573
rect 48590 21564 48596 21576
rect 48648 21564 48654 21616
rect 46477 21539 46535 21545
rect 46477 21536 46489 21539
rect 45980 21508 46489 21536
rect 45980 21496 45986 21508
rect 46477 21505 46489 21508
rect 46523 21505 46535 21539
rect 46477 21499 46535 21505
rect 46842 21496 46848 21548
rect 46900 21536 46906 21548
rect 47121 21539 47179 21545
rect 47121 21536 47133 21539
rect 46900 21508 47133 21536
rect 46900 21496 46906 21508
rect 47121 21505 47133 21508
rect 47167 21536 47179 21539
rect 47765 21539 47823 21545
rect 47765 21536 47777 21539
rect 47167 21508 47777 21536
rect 47167 21505 47179 21508
rect 47121 21499 47179 21505
rect 47765 21505 47777 21508
rect 47811 21505 47823 21539
rect 47765 21499 47823 21505
rect 48498 21496 48504 21548
rect 48556 21536 48562 21548
rect 49053 21539 49111 21545
rect 49053 21536 49065 21539
rect 48556 21508 49065 21536
rect 48556 21496 48562 21508
rect 49053 21505 49065 21508
rect 49099 21505 49111 21539
rect 49053 21499 49111 21505
rect 47578 21468 47584 21480
rect 44192 21440 47584 21468
rect 47578 21428 47584 21440
rect 47636 21428 47642 21480
rect 39448 21372 40448 21400
rect 40604 21372 42656 21400
rect 39448 21360 39454 21372
rect 40604 21344 40632 21372
rect 45554 21360 45560 21412
rect 45612 21400 45618 21412
rect 48593 21403 48651 21409
rect 48593 21400 48605 21403
rect 45612 21372 48605 21400
rect 45612 21360 45618 21372
rect 48593 21369 48605 21372
rect 48639 21369 48651 21403
rect 48593 21363 48651 21369
rect 37608 21304 38148 21332
rect 37608 21292 37614 21304
rect 38286 21292 38292 21344
rect 38344 21332 38350 21344
rect 39761 21335 39819 21341
rect 39761 21332 39773 21335
rect 38344 21304 39773 21332
rect 38344 21292 38350 21304
rect 39761 21301 39773 21304
rect 39807 21332 39819 21335
rect 40586 21332 40592 21344
rect 39807 21304 40592 21332
rect 39807 21301 39819 21304
rect 39761 21295 39819 21301
rect 40586 21292 40592 21304
rect 40644 21292 40650 21344
rect 42058 21292 42064 21344
rect 42116 21292 42122 21344
rect 42334 21292 42340 21344
rect 42392 21332 42398 21344
rect 43257 21335 43315 21341
rect 43257 21332 43269 21335
rect 42392 21304 43269 21332
rect 42392 21292 42398 21304
rect 43257 21301 43269 21304
rect 43303 21301 43315 21335
rect 43257 21295 43315 21301
rect 43714 21292 43720 21344
rect 43772 21292 43778 21344
rect 44358 21292 44364 21344
rect 44416 21292 44422 21344
rect 45002 21292 45008 21344
rect 45060 21292 45066 21344
rect 45186 21292 45192 21344
rect 45244 21332 45250 21344
rect 45649 21335 45707 21341
rect 45649 21332 45661 21335
rect 45244 21304 45661 21332
rect 45244 21292 45250 21304
rect 45649 21301 45661 21304
rect 45695 21301 45707 21335
rect 45649 21295 45707 21301
rect 45738 21292 45744 21344
rect 45796 21332 45802 21344
rect 46937 21335 46995 21341
rect 46937 21332 46949 21335
rect 45796 21304 46949 21332
rect 45796 21292 45802 21304
rect 46937 21301 46949 21304
rect 46983 21301 46995 21335
rect 46937 21295 46995 21301
rect 48866 21292 48872 21344
rect 48924 21332 48930 21344
rect 49237 21335 49295 21341
rect 49237 21332 49249 21335
rect 48924 21304 49249 21332
rect 48924 21292 48930 21304
rect 49237 21301 49249 21304
rect 49283 21301 49295 21335
rect 49237 21295 49295 21301
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 3418 21088 3424 21140
rect 3476 21128 3482 21140
rect 6454 21128 6460 21140
rect 3476 21100 6460 21128
rect 3476 21088 3482 21100
rect 6454 21088 6460 21100
rect 6512 21088 6518 21140
rect 7650 21088 7656 21140
rect 7708 21088 7714 21140
rect 8481 21131 8539 21137
rect 8481 21097 8493 21131
rect 8527 21128 8539 21131
rect 9674 21128 9680 21140
rect 8527 21100 9680 21128
rect 8527 21097 8539 21100
rect 8481 21091 8539 21097
rect 9674 21088 9680 21100
rect 9732 21088 9738 21140
rect 10321 21131 10379 21137
rect 10321 21097 10333 21131
rect 10367 21128 10379 21131
rect 10410 21128 10416 21140
rect 10367 21100 10416 21128
rect 10367 21097 10379 21100
rect 10321 21091 10379 21097
rect 10410 21088 10416 21100
rect 10468 21088 10474 21140
rect 15286 21128 15292 21140
rect 10704 21100 15292 21128
rect 3970 21020 3976 21072
rect 4028 21060 4034 21072
rect 8018 21060 8024 21072
rect 4028 21032 8024 21060
rect 4028 21020 4034 21032
rect 8018 21020 8024 21032
rect 8076 21020 8082 21072
rect 9030 21020 9036 21072
rect 9088 21020 9094 21072
rect 9217 21063 9275 21069
rect 9217 21029 9229 21063
rect 9263 21060 9275 21063
rect 9401 21063 9459 21069
rect 9401 21060 9413 21063
rect 9263 21032 9413 21060
rect 9263 21029 9275 21032
rect 9217 21023 9275 21029
rect 9401 21029 9413 21032
rect 9447 21060 9459 21063
rect 9582 21060 9588 21072
rect 9447 21032 9588 21060
rect 9447 21029 9459 21032
rect 9401 21023 9459 21029
rect 9582 21020 9588 21032
rect 9640 21020 9646 21072
rect 1780 20964 4016 20992
rect 1780 20933 1808 20964
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20893 1823 20927
rect 1765 20887 1823 20893
rect 2774 20816 2780 20868
rect 2832 20816 2838 20868
rect 3988 20788 4016 20964
rect 4154 20952 4160 21004
rect 4212 20992 4218 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 4212 20964 4445 20992
rect 4212 20952 4218 20964
rect 4433 20961 4445 20964
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 5626 20952 5632 21004
rect 5684 20992 5690 21004
rect 6273 20995 6331 21001
rect 6273 20992 6285 20995
rect 5684 20964 6285 20992
rect 5684 20952 5690 20964
rect 6273 20961 6285 20964
rect 6319 20961 6331 20995
rect 8294 20992 8300 21004
rect 6273 20955 6331 20961
rect 7116 20964 8300 20992
rect 4065 20927 4123 20933
rect 4065 20893 4077 20927
rect 4111 20893 4123 20927
rect 4065 20887 4123 20893
rect 5997 20927 6055 20933
rect 5997 20893 6009 20927
rect 6043 20924 6055 20927
rect 7006 20924 7012 20936
rect 6043 20896 7012 20924
rect 6043 20893 6055 20896
rect 5997 20887 6055 20893
rect 4080 20856 4108 20887
rect 7006 20884 7012 20896
rect 7064 20884 7070 20936
rect 7116 20856 7144 20964
rect 8294 20952 8300 20964
rect 8352 20952 8358 21004
rect 7834 20884 7840 20936
rect 7892 20884 7898 20936
rect 9490 20924 9496 20936
rect 8036 20896 9496 20924
rect 8036 20856 8064 20896
rect 9490 20884 9496 20896
rect 9548 20884 9554 20936
rect 9721 20927 9779 20933
rect 9721 20893 9733 20927
rect 9767 20924 9779 20927
rect 10704 20924 10732 21100
rect 15286 21088 15292 21100
rect 15344 21088 15350 21140
rect 16942 21088 16948 21140
rect 17000 21088 17006 21140
rect 17218 21088 17224 21140
rect 17276 21128 17282 21140
rect 18141 21131 18199 21137
rect 18141 21128 18153 21131
rect 17276 21100 18153 21128
rect 17276 21088 17282 21100
rect 18141 21097 18153 21100
rect 18187 21097 18199 21131
rect 20530 21128 20536 21140
rect 18141 21091 18199 21097
rect 18248 21100 20536 21128
rect 12989 21063 13047 21069
rect 12989 21029 13001 21063
rect 13035 21029 13047 21063
rect 18248 21060 18276 21100
rect 20530 21088 20536 21100
rect 20588 21088 20594 21140
rect 20622 21088 20628 21140
rect 20680 21128 20686 21140
rect 21542 21128 21548 21140
rect 20680 21100 21548 21128
rect 20680 21088 20686 21100
rect 21542 21088 21548 21100
rect 21600 21128 21606 21140
rect 22005 21131 22063 21137
rect 22005 21128 22017 21131
rect 21600 21100 22017 21128
rect 21600 21088 21606 21100
rect 22005 21097 22017 21100
rect 22051 21097 22063 21131
rect 22005 21091 22063 21097
rect 22278 21088 22284 21140
rect 22336 21128 22342 21140
rect 24762 21128 24768 21140
rect 22336 21100 24768 21128
rect 22336 21088 22342 21100
rect 24762 21088 24768 21100
rect 24820 21088 24826 21140
rect 26234 21088 26240 21140
rect 26292 21128 26298 21140
rect 27893 21131 27951 21137
rect 27893 21128 27905 21131
rect 26292 21100 27905 21128
rect 26292 21088 26298 21100
rect 27893 21097 27905 21100
rect 27939 21097 27951 21131
rect 27893 21091 27951 21097
rect 28353 21131 28411 21137
rect 28353 21097 28365 21131
rect 28399 21128 28411 21131
rect 30098 21128 30104 21140
rect 28399 21100 30104 21128
rect 28399 21097 28411 21100
rect 28353 21091 28411 21097
rect 30098 21088 30104 21100
rect 30156 21088 30162 21140
rect 30558 21088 30564 21140
rect 30616 21128 30622 21140
rect 30745 21131 30803 21137
rect 30745 21128 30757 21131
rect 30616 21100 30757 21128
rect 30616 21088 30622 21100
rect 30745 21097 30757 21100
rect 30791 21097 30803 21131
rect 35710 21128 35716 21140
rect 30745 21091 30803 21097
rect 31220 21100 35716 21128
rect 12989 21023 13047 21029
rect 17420 21032 18276 21060
rect 12894 20992 12900 21004
rect 10796 20964 12900 20992
rect 10796 20933 10824 20964
rect 12894 20952 12900 20964
rect 12952 20952 12958 21004
rect 13004 20992 13032 21023
rect 13004 20964 13124 20992
rect 9767 20896 10732 20924
rect 10781 20927 10839 20933
rect 9767 20893 9779 20896
rect 9721 20887 9779 20893
rect 10781 20893 10793 20927
rect 10827 20893 10839 20927
rect 10781 20887 10839 20893
rect 11885 20927 11943 20933
rect 11885 20893 11897 20927
rect 11931 20924 11943 20927
rect 12526 20924 12532 20936
rect 11931 20896 12532 20924
rect 11931 20893 11943 20896
rect 11885 20887 11943 20893
rect 12526 20884 12532 20896
rect 12584 20884 12590 20936
rect 13096 20868 13124 20964
rect 13262 20952 13268 21004
rect 13320 20992 13326 21004
rect 13633 20995 13691 21001
rect 13633 20992 13645 20995
rect 13320 20964 13645 20992
rect 13320 20952 13326 20964
rect 13633 20961 13645 20964
rect 13679 20992 13691 20995
rect 14182 20992 14188 21004
rect 13679 20964 14188 20992
rect 13679 20961 13691 20964
rect 13633 20955 13691 20961
rect 14182 20952 14188 20964
rect 14240 20952 14246 21004
rect 14366 20952 14372 21004
rect 14424 20952 14430 21004
rect 15010 20952 15016 21004
rect 15068 20992 15074 21004
rect 17420 21001 17448 21032
rect 18322 21020 18328 21072
rect 18380 21060 18386 21072
rect 19797 21063 19855 21069
rect 19797 21060 19809 21063
rect 18380 21032 19809 21060
rect 18380 21020 18386 21032
rect 19797 21029 19809 21032
rect 19843 21029 19855 21063
rect 19797 21023 19855 21029
rect 22830 21020 22836 21072
rect 22888 21020 22894 21072
rect 23293 21063 23351 21069
rect 23293 21029 23305 21063
rect 23339 21060 23351 21063
rect 23339 21032 28856 21060
rect 23339 21029 23351 21032
rect 23293 21023 23351 21029
rect 17405 20995 17463 21001
rect 15068 20964 17356 20992
rect 15068 20952 15074 20964
rect 13357 20927 13415 20933
rect 13357 20893 13369 20927
rect 13403 20924 13415 20927
rect 13446 20924 13452 20936
rect 13403 20896 13452 20924
rect 13403 20893 13415 20896
rect 13357 20887 13415 20893
rect 13446 20884 13452 20896
rect 13504 20884 13510 20936
rect 13814 20884 13820 20936
rect 13872 20924 13878 20936
rect 14645 20927 14703 20933
rect 14645 20924 14657 20927
rect 13872 20896 14657 20924
rect 13872 20884 13878 20896
rect 14645 20893 14657 20896
rect 14691 20893 14703 20927
rect 14645 20887 14703 20893
rect 15930 20884 15936 20936
rect 15988 20924 15994 20936
rect 16758 20924 16764 20936
rect 15988 20896 16764 20924
rect 15988 20884 15994 20896
rect 16758 20884 16764 20896
rect 16816 20884 16822 20936
rect 17328 20924 17356 20964
rect 17405 20961 17417 20995
rect 17451 20961 17463 20995
rect 17405 20955 17463 20961
rect 17494 20952 17500 21004
rect 17552 20952 17558 21004
rect 18693 20995 18751 21001
rect 18693 20992 18705 20995
rect 17604 20964 18705 20992
rect 17512 20924 17540 20952
rect 17328 20896 17540 20924
rect 4080 20828 7144 20856
rect 7208 20828 8064 20856
rect 8389 20859 8447 20865
rect 7208 20788 7236 20828
rect 8389 20825 8401 20859
rect 8435 20856 8447 20859
rect 9950 20856 9956 20868
rect 8435 20828 9956 20856
rect 8435 20825 8447 20828
rect 8389 20819 8447 20825
rect 9950 20816 9956 20828
rect 10008 20816 10014 20868
rect 11425 20859 11483 20865
rect 11425 20825 11437 20859
rect 11471 20856 11483 20859
rect 12802 20856 12808 20868
rect 11471 20828 12808 20856
rect 11471 20825 11483 20828
rect 11425 20819 11483 20825
rect 12802 20816 12808 20828
rect 12860 20816 12866 20868
rect 13078 20816 13084 20868
rect 13136 20816 13142 20868
rect 13170 20816 13176 20868
rect 13228 20856 13234 20868
rect 14921 20859 14979 20865
rect 14921 20856 14933 20859
rect 13228 20828 14933 20856
rect 13228 20816 13234 20828
rect 14921 20825 14933 20828
rect 14967 20825 14979 20859
rect 17604 20856 17632 20964
rect 18693 20961 18705 20964
rect 18739 20992 18751 20995
rect 18782 20992 18788 21004
rect 18739 20964 18788 20992
rect 18739 20961 18751 20964
rect 18693 20955 18751 20961
rect 18782 20952 18788 20964
rect 18840 20952 18846 21004
rect 20257 20995 20315 21001
rect 20257 20961 20269 20995
rect 20303 20992 20315 20995
rect 21174 20992 21180 21004
rect 20303 20964 21180 20992
rect 20303 20961 20315 20964
rect 20257 20955 20315 20961
rect 21174 20952 21180 20964
rect 21232 20952 21238 21004
rect 21726 20992 21732 21004
rect 21652 20964 21732 20992
rect 21652 20910 21680 20964
rect 21726 20952 21732 20964
rect 21784 20992 21790 21004
rect 21910 20992 21916 21004
rect 21784 20964 21916 20992
rect 21784 20952 21790 20964
rect 21910 20952 21916 20964
rect 21968 20952 21974 21004
rect 22738 20992 22744 21004
rect 22066 20964 22744 20992
rect 22066 20924 22094 20964
rect 22738 20952 22744 20964
rect 22796 20952 22802 21004
rect 23750 20952 23756 21004
rect 23808 20952 23814 21004
rect 23842 20952 23848 21004
rect 23900 20952 23906 21004
rect 26326 20952 26332 21004
rect 26384 20952 26390 21004
rect 27522 20952 27528 21004
rect 27580 20952 27586 21004
rect 28828 21001 28856 21032
rect 29730 21020 29736 21072
rect 29788 21020 29794 21072
rect 28813 20995 28871 21001
rect 28813 20961 28825 20995
rect 28859 20961 28871 20995
rect 28813 20955 28871 20961
rect 28905 20995 28963 21001
rect 28905 20961 28917 20995
rect 28951 20992 28963 20995
rect 28994 20992 29000 21004
rect 28951 20964 29000 20992
rect 28951 20961 28963 20964
rect 28905 20955 28963 20961
rect 28994 20952 29000 20964
rect 29052 20952 29058 21004
rect 30098 20952 30104 21004
rect 30156 20992 30162 21004
rect 30742 20992 30748 21004
rect 30156 20964 30748 20992
rect 30156 20952 30162 20964
rect 30742 20952 30748 20964
rect 30800 20952 30806 21004
rect 31220 21001 31248 21100
rect 35710 21088 35716 21100
rect 35768 21088 35774 21140
rect 36906 21088 36912 21140
rect 36964 21128 36970 21140
rect 37093 21131 37151 21137
rect 37093 21128 37105 21131
rect 36964 21100 37105 21128
rect 36964 21088 36970 21100
rect 37093 21097 37105 21100
rect 37139 21097 37151 21131
rect 37093 21091 37151 21097
rect 37182 21088 37188 21140
rect 37240 21128 37246 21140
rect 37240 21100 39160 21128
rect 37240 21088 37246 21100
rect 31754 21020 31760 21072
rect 31812 21060 31818 21072
rect 31849 21063 31907 21069
rect 31849 21060 31861 21063
rect 31812 21032 31861 21060
rect 31812 21020 31818 21032
rect 31849 21029 31861 21032
rect 31895 21060 31907 21063
rect 32398 21060 32404 21072
rect 31895 21032 32404 21060
rect 31895 21029 31907 21032
rect 31849 21023 31907 21029
rect 32398 21020 32404 21032
rect 32456 21020 32462 21072
rect 39132 21060 39160 21100
rect 39206 21088 39212 21140
rect 39264 21128 39270 21140
rect 39393 21131 39451 21137
rect 39393 21128 39405 21131
rect 39264 21100 39405 21128
rect 39264 21088 39270 21100
rect 39393 21097 39405 21100
rect 39439 21097 39451 21131
rect 39393 21091 39451 21097
rect 40037 21131 40095 21137
rect 40037 21097 40049 21131
rect 40083 21128 40095 21131
rect 40310 21128 40316 21140
rect 40083 21100 40316 21128
rect 40083 21097 40095 21100
rect 40037 21091 40095 21097
rect 40310 21088 40316 21100
rect 40368 21088 40374 21140
rect 40494 21088 40500 21140
rect 40552 21128 40558 21140
rect 44266 21128 44272 21140
rect 40552 21100 44272 21128
rect 40552 21088 40558 21100
rect 44266 21088 44272 21100
rect 44324 21088 44330 21140
rect 44361 21131 44419 21137
rect 44361 21097 44373 21131
rect 44407 21128 44419 21131
rect 44910 21128 44916 21140
rect 44407 21100 44916 21128
rect 44407 21097 44419 21100
rect 44361 21091 44419 21097
rect 44910 21088 44916 21100
rect 44968 21088 44974 21140
rect 45830 21088 45836 21140
rect 45888 21088 45894 21140
rect 46014 21088 46020 21140
rect 46072 21088 46078 21140
rect 46566 21088 46572 21140
rect 46624 21128 46630 21140
rect 47029 21131 47087 21137
rect 47029 21128 47041 21131
rect 46624 21100 47041 21128
rect 46624 21088 46630 21100
rect 47029 21097 47041 21100
rect 47075 21097 47087 21131
rect 47029 21091 47087 21097
rect 47578 21088 47584 21140
rect 47636 21128 47642 21140
rect 47765 21131 47823 21137
rect 47765 21128 47777 21131
rect 47636 21100 47777 21128
rect 47636 21088 47642 21100
rect 47765 21097 47777 21100
rect 47811 21097 47823 21131
rect 47765 21091 47823 21097
rect 48314 21088 48320 21140
rect 48372 21128 48378 21140
rect 48409 21131 48467 21137
rect 48409 21128 48421 21131
rect 48372 21100 48421 21128
rect 48372 21088 48378 21100
rect 48409 21097 48421 21100
rect 48455 21097 48467 21131
rect 48409 21091 48467 21097
rect 39298 21060 39304 21072
rect 39132 21032 39304 21060
rect 39298 21020 39304 21032
rect 39356 21020 39362 21072
rect 42334 21060 42340 21072
rect 39684 21032 42340 21060
rect 31205 20995 31263 21001
rect 31205 20961 31217 20995
rect 31251 20961 31263 20995
rect 31205 20955 31263 20961
rect 31389 20995 31447 21001
rect 31389 20961 31401 20995
rect 31435 20992 31447 20995
rect 32769 20995 32827 21001
rect 31435 20964 32260 20992
rect 31435 20961 31447 20964
rect 31389 20955 31447 20961
rect 21836 20896 22094 20924
rect 22649 20927 22707 20933
rect 14921 20819 14979 20825
rect 16316 20828 17632 20856
rect 3988 20760 7236 20788
rect 8018 20748 8024 20800
rect 8076 20788 8082 20800
rect 12250 20788 12256 20800
rect 8076 20760 12256 20788
rect 8076 20748 8082 20760
rect 12250 20748 12256 20760
rect 12308 20748 12314 20800
rect 12529 20791 12587 20797
rect 12529 20757 12541 20791
rect 12575 20788 12587 20791
rect 12618 20788 12624 20800
rect 12575 20760 12624 20788
rect 12575 20757 12587 20760
rect 12529 20751 12587 20757
rect 12618 20748 12624 20760
rect 12676 20748 12682 20800
rect 13449 20791 13507 20797
rect 13449 20757 13461 20791
rect 13495 20788 13507 20791
rect 13722 20788 13728 20800
rect 13495 20760 13728 20788
rect 13495 20757 13507 20760
rect 13449 20751 13507 20757
rect 13722 20748 13728 20760
rect 13780 20748 13786 20800
rect 14185 20791 14243 20797
rect 14185 20757 14197 20791
rect 14231 20788 14243 20791
rect 14458 20788 14464 20800
rect 14231 20760 14464 20788
rect 14231 20757 14243 20760
rect 14185 20751 14243 20757
rect 14458 20748 14464 20760
rect 14516 20788 14522 20800
rect 16316 20788 16344 20828
rect 17954 20816 17960 20868
rect 18012 20856 18018 20868
rect 18509 20859 18567 20865
rect 18509 20856 18521 20859
rect 18012 20828 18521 20856
rect 18012 20816 18018 20828
rect 18509 20825 18521 20828
rect 18555 20825 18567 20859
rect 18509 20819 18567 20825
rect 19613 20859 19671 20865
rect 19613 20825 19625 20859
rect 19659 20856 19671 20859
rect 20254 20856 20260 20868
rect 19659 20828 20260 20856
rect 19659 20825 19671 20828
rect 19613 20819 19671 20825
rect 20254 20816 20260 20828
rect 20312 20816 20318 20868
rect 20533 20859 20591 20865
rect 20533 20825 20545 20859
rect 20579 20825 20591 20859
rect 20533 20819 20591 20825
rect 14516 20760 16344 20788
rect 14516 20748 14522 20760
rect 16390 20748 16396 20800
rect 16448 20748 16454 20800
rect 17310 20748 17316 20800
rect 17368 20748 17374 20800
rect 18598 20748 18604 20800
rect 18656 20748 18662 20800
rect 20548 20788 20576 20819
rect 21836 20788 21864 20896
rect 22649 20893 22661 20927
rect 22695 20924 22707 20927
rect 22830 20924 22836 20936
rect 22695 20896 22836 20924
rect 22695 20893 22707 20896
rect 22649 20887 22707 20893
rect 22830 20884 22836 20896
rect 22888 20884 22894 20936
rect 24581 20927 24639 20933
rect 24581 20893 24593 20927
rect 24627 20924 24639 20927
rect 24762 20924 24768 20936
rect 24627 20896 24768 20924
rect 24627 20893 24639 20896
rect 24581 20887 24639 20893
rect 24762 20884 24768 20896
rect 24820 20884 24826 20936
rect 27249 20927 27307 20933
rect 27249 20893 27261 20927
rect 27295 20924 27307 20927
rect 28534 20924 28540 20936
rect 27295 20896 28540 20924
rect 27295 20893 27307 20896
rect 27249 20887 27307 20893
rect 28534 20884 28540 20896
rect 28592 20884 28598 20936
rect 29914 20884 29920 20936
rect 29972 20884 29978 20936
rect 31294 20924 31300 20936
rect 30392 20896 31300 20924
rect 22738 20816 22744 20868
rect 22796 20856 22802 20868
rect 26786 20856 26792 20868
rect 22796 20828 25728 20856
rect 22796 20816 22802 20828
rect 20548 20760 21864 20788
rect 22554 20748 22560 20800
rect 22612 20788 22618 20800
rect 23290 20788 23296 20800
rect 22612 20760 23296 20788
rect 22612 20748 22618 20760
rect 23290 20748 23296 20760
rect 23348 20748 23354 20800
rect 23658 20748 23664 20800
rect 23716 20748 23722 20800
rect 25130 20748 25136 20800
rect 25188 20788 25194 20800
rect 25700 20797 25728 20828
rect 26068 20828 26792 20856
rect 26068 20797 26096 20828
rect 26786 20816 26792 20828
rect 26844 20816 26850 20868
rect 27341 20859 27399 20865
rect 27341 20825 27353 20859
rect 27387 20856 27399 20859
rect 27614 20856 27620 20868
rect 27387 20828 27620 20856
rect 27387 20825 27399 20828
rect 27341 20819 27399 20825
rect 27614 20816 27620 20828
rect 27672 20816 27678 20868
rect 27798 20816 27804 20868
rect 27856 20856 27862 20868
rect 30392 20856 30420 20896
rect 31294 20884 31300 20896
rect 31352 20884 31358 20936
rect 31846 20884 31852 20936
rect 31904 20924 31910 20936
rect 31941 20927 31999 20933
rect 31941 20924 31953 20927
rect 31904 20896 31953 20924
rect 31904 20884 31910 20896
rect 31941 20893 31953 20896
rect 31987 20893 31999 20927
rect 31941 20887 31999 20893
rect 27856 20828 30420 20856
rect 30469 20859 30527 20865
rect 27856 20816 27862 20828
rect 30469 20825 30481 20859
rect 30515 20856 30527 20859
rect 30558 20856 30564 20868
rect 30515 20828 30564 20856
rect 30515 20825 30527 20828
rect 30469 20819 30527 20825
rect 30558 20816 30564 20828
rect 30616 20856 30622 20868
rect 31570 20856 31576 20868
rect 30616 20828 31576 20856
rect 30616 20816 30622 20828
rect 31570 20816 31576 20828
rect 31628 20816 31634 20868
rect 25225 20791 25283 20797
rect 25225 20788 25237 20791
rect 25188 20760 25237 20788
rect 25188 20748 25194 20760
rect 25225 20757 25237 20760
rect 25271 20757 25283 20791
rect 25225 20751 25283 20757
rect 25685 20791 25743 20797
rect 25685 20757 25697 20791
rect 25731 20757 25743 20791
rect 25685 20751 25743 20757
rect 26053 20791 26111 20797
rect 26053 20757 26065 20791
rect 26099 20757 26111 20791
rect 26053 20751 26111 20757
rect 26142 20748 26148 20800
rect 26200 20748 26206 20800
rect 26326 20748 26332 20800
rect 26384 20788 26390 20800
rect 26881 20791 26939 20797
rect 26881 20788 26893 20791
rect 26384 20760 26893 20788
rect 26384 20748 26390 20760
rect 26881 20757 26893 20760
rect 26927 20757 26939 20791
rect 26881 20751 26939 20757
rect 28718 20748 28724 20800
rect 28776 20748 28782 20800
rect 28902 20748 28908 20800
rect 28960 20788 28966 20800
rect 30098 20788 30104 20800
rect 28960 20760 30104 20788
rect 28960 20748 28966 20760
rect 30098 20748 30104 20760
rect 30156 20788 30162 20800
rect 30193 20791 30251 20797
rect 30193 20788 30205 20791
rect 30156 20760 30205 20788
rect 30156 20748 30162 20760
rect 30193 20757 30205 20760
rect 30239 20757 30251 20791
rect 30193 20751 30251 20757
rect 31113 20791 31171 20797
rect 31113 20757 31125 20791
rect 31159 20788 31171 20791
rect 31294 20788 31300 20800
rect 31159 20760 31300 20788
rect 31159 20757 31171 20760
rect 31113 20751 31171 20757
rect 31294 20748 31300 20760
rect 31352 20748 31358 20800
rect 31846 20748 31852 20800
rect 31904 20788 31910 20800
rect 32125 20791 32183 20797
rect 32125 20788 32137 20791
rect 31904 20760 32137 20788
rect 31904 20748 31910 20760
rect 32125 20757 32137 20760
rect 32171 20757 32183 20791
rect 32232 20788 32260 20964
rect 32769 20961 32781 20995
rect 32815 20992 32827 20995
rect 32858 20992 32864 21004
rect 32815 20964 32864 20992
rect 32815 20961 32827 20964
rect 32769 20955 32827 20961
rect 32858 20952 32864 20964
rect 32916 20952 32922 21004
rect 33134 20952 33140 21004
rect 33192 20992 33198 21004
rect 33192 20964 34100 20992
rect 33192 20952 33198 20964
rect 32306 20884 32312 20936
rect 32364 20924 32370 20936
rect 32493 20927 32551 20933
rect 32493 20924 32505 20927
rect 32364 20896 32505 20924
rect 32364 20884 32370 20896
rect 32493 20893 32505 20896
rect 32539 20893 32551 20927
rect 32493 20887 32551 20893
rect 33042 20816 33048 20868
rect 33100 20856 33106 20868
rect 34072 20856 34100 20964
rect 34882 20952 34888 21004
rect 34940 20952 34946 21004
rect 35161 20995 35219 21001
rect 35161 20961 35173 20995
rect 35207 20992 35219 20995
rect 36722 20992 36728 21004
rect 35207 20964 36728 20992
rect 35207 20961 35219 20964
rect 35161 20955 35219 20961
rect 36722 20952 36728 20964
rect 36780 20952 36786 21004
rect 37921 20995 37979 21001
rect 37921 20961 37933 20995
rect 37967 20992 37979 20995
rect 39684 20992 39712 21032
rect 42334 21020 42340 21032
rect 42392 21020 42398 21072
rect 42794 21020 42800 21072
rect 42852 21060 42858 21072
rect 45189 21063 45247 21069
rect 45189 21060 45201 21063
rect 42852 21032 45201 21060
rect 42852 21020 42858 21032
rect 45189 21029 45201 21032
rect 45235 21029 45247 21063
rect 45189 21023 45247 21029
rect 37967 20964 39712 20992
rect 37967 20961 37979 20964
rect 37921 20955 37979 20961
rect 39942 20952 39948 21004
rect 40000 20992 40006 21004
rect 40497 20995 40555 21001
rect 40497 20992 40509 20995
rect 40000 20964 40509 20992
rect 40000 20952 40006 20964
rect 40497 20961 40509 20964
rect 40543 20961 40555 20995
rect 40497 20955 40555 20961
rect 40586 20952 40592 21004
rect 40644 20952 40650 21004
rect 41785 20995 41843 21001
rect 41785 20992 41797 20995
rect 41386 20964 41797 20992
rect 37642 20884 37648 20936
rect 37700 20884 37706 20936
rect 39206 20884 39212 20936
rect 39264 20924 39270 20936
rect 41386 20924 41414 20964
rect 41785 20961 41797 20964
rect 41831 20961 41843 20995
rect 41785 20955 41843 20961
rect 42426 20952 42432 21004
rect 42484 20952 42490 21004
rect 42702 20952 42708 21004
rect 42760 20952 42766 21004
rect 48774 20992 48780 21004
rect 42812 20964 48780 20992
rect 39264 20896 41414 20924
rect 41601 20927 41659 20933
rect 39264 20884 39270 20896
rect 41601 20893 41613 20927
rect 41647 20924 41659 20927
rect 42812 20924 42840 20964
rect 48774 20952 48780 20964
rect 48832 20952 48838 21004
rect 41647 20896 42840 20924
rect 41647 20893 41659 20896
rect 41601 20887 41659 20893
rect 42886 20884 42892 20936
rect 42944 20924 42950 20936
rect 43806 20924 43812 20936
rect 42944 20896 43812 20924
rect 42944 20884 42950 20896
rect 43806 20884 43812 20896
rect 43864 20924 43870 20936
rect 43901 20927 43959 20933
rect 43901 20924 43913 20927
rect 43864 20896 43913 20924
rect 43864 20884 43870 20896
rect 43901 20893 43913 20896
rect 43947 20893 43959 20927
rect 43901 20887 43959 20893
rect 44450 20884 44456 20936
rect 44508 20924 44514 20936
rect 44545 20927 44603 20933
rect 44545 20924 44557 20927
rect 44508 20896 44557 20924
rect 44508 20884 44514 20896
rect 44545 20893 44557 20896
rect 44591 20893 44603 20927
rect 44545 20887 44603 20893
rect 45094 20884 45100 20936
rect 45152 20924 45158 20936
rect 45373 20927 45431 20933
rect 45373 20924 45385 20927
rect 45152 20896 45385 20924
rect 45152 20884 45158 20896
rect 45373 20893 45385 20896
rect 45419 20924 45431 20927
rect 45649 20927 45707 20933
rect 45649 20924 45661 20927
rect 45419 20896 45661 20924
rect 45419 20893 45431 20896
rect 45373 20887 45431 20893
rect 45649 20893 45661 20896
rect 45695 20893 45707 20927
rect 45649 20887 45707 20893
rect 46382 20884 46388 20936
rect 46440 20924 46446 20936
rect 46569 20927 46627 20933
rect 46569 20924 46581 20927
rect 46440 20896 46581 20924
rect 46440 20884 46446 20896
rect 46569 20893 46581 20896
rect 46615 20893 46627 20927
rect 46569 20887 46627 20893
rect 47026 20884 47032 20936
rect 47084 20924 47090 20936
rect 47213 20927 47271 20933
rect 47213 20924 47225 20927
rect 47084 20896 47225 20924
rect 47084 20884 47090 20896
rect 47213 20893 47225 20896
rect 47259 20893 47271 20927
rect 47213 20887 47271 20893
rect 47670 20884 47676 20936
rect 47728 20924 47734 20936
rect 47949 20927 48007 20933
rect 47949 20924 47961 20927
rect 47728 20896 47961 20924
rect 47728 20884 47734 20896
rect 47949 20893 47961 20896
rect 47995 20893 48007 20927
rect 47949 20887 48007 20893
rect 48222 20884 48228 20936
rect 48280 20924 48286 20936
rect 48593 20927 48651 20933
rect 48593 20924 48605 20927
rect 48280 20896 48605 20924
rect 48280 20884 48286 20896
rect 48593 20893 48605 20896
rect 48639 20893 48651 20927
rect 48593 20887 48651 20893
rect 49050 20884 49056 20936
rect 49108 20884 49114 20936
rect 33100 20828 33258 20856
rect 34072 20828 35650 20856
rect 36556 20828 38332 20856
rect 33100 20816 33106 20828
rect 33778 20788 33784 20800
rect 32232 20760 33784 20788
rect 32125 20751 32183 20757
rect 33778 20748 33784 20760
rect 33836 20748 33842 20800
rect 34146 20748 34152 20800
rect 34204 20788 34210 20800
rect 34241 20791 34299 20797
rect 34241 20788 34253 20791
rect 34204 20760 34253 20788
rect 34204 20748 34210 20760
rect 34241 20757 34253 20760
rect 34287 20788 34299 20791
rect 36556 20788 36584 20828
rect 34287 20760 36584 20788
rect 34287 20757 34299 20760
rect 34241 20751 34299 20757
rect 36630 20748 36636 20800
rect 36688 20748 36694 20800
rect 37274 20748 37280 20800
rect 37332 20748 37338 20800
rect 38304 20788 38332 20828
rect 38562 20816 38568 20868
rect 38620 20816 38626 20868
rect 40405 20859 40463 20865
rect 40405 20825 40417 20859
rect 40451 20856 40463 20859
rect 40451 20828 41276 20856
rect 40451 20825 40463 20828
rect 40405 20819 40463 20825
rect 40770 20788 40776 20800
rect 38304 20760 40776 20788
rect 40770 20748 40776 20760
rect 40828 20748 40834 20800
rect 41248 20797 41276 20828
rect 41322 20816 41328 20868
rect 41380 20856 41386 20868
rect 41693 20859 41751 20865
rect 41693 20856 41705 20859
rect 41380 20828 41705 20856
rect 41380 20816 41386 20828
rect 41693 20825 41705 20828
rect 41739 20856 41751 20859
rect 42978 20856 42984 20868
rect 41739 20828 42984 20856
rect 41739 20825 41751 20828
rect 41693 20819 41751 20825
rect 42978 20816 42984 20828
rect 43036 20816 43042 20868
rect 41233 20791 41291 20797
rect 41233 20757 41245 20791
rect 41279 20757 41291 20791
rect 41233 20751 41291 20757
rect 42794 20748 42800 20800
rect 42852 20788 42858 20800
rect 43717 20791 43775 20797
rect 43717 20788 43729 20791
rect 42852 20760 43729 20788
rect 42852 20748 42858 20760
rect 43717 20757 43729 20760
rect 43763 20757 43775 20791
rect 43717 20751 43775 20757
rect 44266 20748 44272 20800
rect 44324 20788 44330 20800
rect 46385 20791 46443 20797
rect 46385 20788 46397 20791
rect 44324 20760 46397 20788
rect 44324 20748 44330 20760
rect 46385 20757 46397 20760
rect 46431 20757 46443 20791
rect 46385 20751 46443 20757
rect 49234 20748 49240 20800
rect 49292 20748 49298 20800
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 7282 20584 7288 20596
rect 5552 20556 7288 20584
rect 5552 20525 5580 20556
rect 7282 20544 7288 20556
rect 7340 20544 7346 20596
rect 8297 20587 8355 20593
rect 8297 20553 8309 20587
rect 8343 20584 8355 20587
rect 8389 20587 8447 20593
rect 8389 20584 8401 20587
rect 8343 20556 8401 20584
rect 8343 20553 8355 20556
rect 8297 20547 8355 20553
rect 8389 20553 8401 20556
rect 8435 20584 8447 20587
rect 13357 20587 13415 20593
rect 8435 20556 12434 20584
rect 8435 20553 8447 20556
rect 8389 20547 8447 20553
rect 5537 20519 5595 20525
rect 5537 20485 5549 20519
rect 5583 20485 5595 20519
rect 5537 20479 5595 20485
rect 6181 20519 6239 20525
rect 6181 20485 6193 20519
rect 6227 20516 6239 20519
rect 6227 20488 10640 20516
rect 6227 20485 6239 20488
rect 6181 20479 6239 20485
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20448 1823 20451
rect 1854 20448 1860 20460
rect 1811 20420 1860 20448
rect 1811 20417 1823 20420
rect 1765 20411 1823 20417
rect 1854 20408 1860 20420
rect 1912 20408 1918 20460
rect 3602 20408 3608 20460
rect 3660 20408 3666 20460
rect 5353 20451 5411 20457
rect 5353 20417 5365 20451
rect 5399 20417 5411 20451
rect 5353 20411 5411 20417
rect 2777 20383 2835 20389
rect 2777 20349 2789 20383
rect 2823 20380 2835 20383
rect 2866 20380 2872 20392
rect 2823 20352 2872 20380
rect 2823 20349 2835 20352
rect 2777 20343 2835 20349
rect 2866 20340 2872 20352
rect 2924 20340 2930 20392
rect 3878 20340 3884 20392
rect 3936 20340 3942 20392
rect 5368 20380 5396 20411
rect 5902 20408 5908 20460
rect 5960 20448 5966 20460
rect 6549 20451 6607 20457
rect 6549 20448 6561 20451
rect 5960 20420 6561 20448
rect 5960 20408 5966 20420
rect 6549 20417 6561 20420
rect 6595 20417 6607 20451
rect 8846 20448 8852 20460
rect 6549 20411 6607 20417
rect 6656 20420 8852 20448
rect 6656 20380 6684 20420
rect 8846 20408 8852 20420
rect 8904 20408 8910 20460
rect 9122 20408 9128 20460
rect 9180 20408 9186 20460
rect 9861 20451 9919 20457
rect 9861 20417 9873 20451
rect 9907 20448 9919 20451
rect 10226 20448 10232 20460
rect 9907 20420 10232 20448
rect 9907 20417 9919 20420
rect 9861 20411 9919 20417
rect 5368 20352 6684 20380
rect 7190 20340 7196 20392
rect 7248 20340 7254 20392
rect 8294 20340 8300 20392
rect 8352 20380 8358 20392
rect 9309 20383 9367 20389
rect 9309 20380 9321 20383
rect 8352 20352 9321 20380
rect 8352 20340 8358 20352
rect 9309 20349 9321 20352
rect 9355 20349 9367 20383
rect 9309 20343 9367 20349
rect 9398 20340 9404 20392
rect 9456 20380 9462 20392
rect 10045 20383 10103 20389
rect 10045 20380 10057 20383
rect 9456 20352 10057 20380
rect 9456 20340 9462 20352
rect 10045 20349 10057 20352
rect 10091 20349 10103 20383
rect 10045 20343 10103 20349
rect 5997 20315 6055 20321
rect 5997 20281 6009 20315
rect 6043 20312 6055 20315
rect 10152 20312 10180 20420
rect 10226 20408 10232 20420
rect 10284 20408 10290 20460
rect 10502 20408 10508 20460
rect 10560 20408 10566 20460
rect 10612 20448 10640 20488
rect 11698 20476 11704 20528
rect 11756 20476 11762 20528
rect 12250 20476 12256 20528
rect 12308 20476 12314 20528
rect 12406 20516 12434 20556
rect 13357 20553 13369 20587
rect 13403 20584 13415 20587
rect 13906 20584 13912 20596
rect 13403 20556 13912 20584
rect 13403 20553 13415 20556
rect 13357 20547 13415 20553
rect 13906 20544 13912 20556
rect 13964 20544 13970 20596
rect 15102 20584 15108 20596
rect 14016 20556 15108 20584
rect 14016 20516 14044 20556
rect 15102 20544 15108 20556
rect 15160 20544 15166 20596
rect 15378 20544 15384 20596
rect 15436 20584 15442 20596
rect 19058 20584 19064 20596
rect 15436 20556 19064 20584
rect 15436 20544 15442 20556
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 20438 20584 20444 20596
rect 19168 20556 20444 20584
rect 12406 20488 14044 20516
rect 15930 20476 15936 20528
rect 15988 20516 15994 20528
rect 19168 20516 19196 20556
rect 20438 20544 20444 20556
rect 20496 20544 20502 20596
rect 20714 20544 20720 20596
rect 20772 20544 20778 20596
rect 22002 20544 22008 20596
rect 22060 20544 22066 20596
rect 22738 20544 22744 20596
rect 22796 20544 22802 20596
rect 25958 20584 25964 20596
rect 23216 20556 25964 20584
rect 20070 20516 20076 20528
rect 15988 20488 19196 20516
rect 20010 20488 20076 20516
rect 15988 20476 15994 20488
rect 20070 20476 20076 20488
rect 20128 20476 20134 20528
rect 20346 20476 20352 20528
rect 20404 20516 20410 20528
rect 22462 20516 22468 20528
rect 20404 20488 22468 20516
rect 20404 20476 20410 20488
rect 22462 20476 22468 20488
rect 22520 20476 22526 20528
rect 12066 20448 12072 20460
rect 10612 20420 12072 20448
rect 12066 20408 12072 20420
rect 12124 20408 12130 20460
rect 12710 20408 12716 20460
rect 12768 20408 12774 20460
rect 15194 20408 15200 20460
rect 15252 20408 15258 20460
rect 16114 20408 16120 20460
rect 16172 20408 16178 20460
rect 16758 20408 16764 20460
rect 16816 20448 16822 20460
rect 17313 20451 17371 20457
rect 17313 20448 17325 20451
rect 16816 20420 17325 20448
rect 16816 20408 16822 20420
rect 17313 20417 17325 20420
rect 17359 20417 17371 20451
rect 17313 20411 17371 20417
rect 17402 20408 17408 20460
rect 17460 20408 17466 20460
rect 18049 20451 18107 20457
rect 18049 20417 18061 20451
rect 18095 20448 18107 20451
rect 18141 20451 18199 20457
rect 18141 20448 18153 20451
rect 18095 20420 18153 20448
rect 18095 20417 18107 20420
rect 18049 20411 18107 20417
rect 18141 20417 18153 20420
rect 18187 20448 18199 20451
rect 18414 20448 18420 20460
rect 18187 20420 18420 20448
rect 18187 20417 18199 20420
rect 18141 20411 18199 20417
rect 18414 20408 18420 20420
rect 18472 20408 18478 20460
rect 21082 20408 21088 20460
rect 21140 20408 21146 20460
rect 22649 20451 22707 20457
rect 22649 20417 22661 20451
rect 22695 20448 22707 20451
rect 22830 20448 22836 20460
rect 22695 20420 22836 20448
rect 22695 20417 22707 20420
rect 22649 20411 22707 20417
rect 22830 20408 22836 20420
rect 22888 20408 22894 20460
rect 11606 20340 11612 20392
rect 11664 20380 11670 20392
rect 12342 20380 12348 20392
rect 11664 20352 12348 20380
rect 11664 20340 11670 20352
rect 12342 20340 12348 20352
rect 12400 20340 12406 20392
rect 12618 20340 12624 20392
rect 12676 20380 12682 20392
rect 12676 20352 13400 20380
rect 12676 20340 12682 20352
rect 6043 20284 10180 20312
rect 6043 20281 6055 20284
rect 5997 20275 6055 20281
rect 11514 20272 11520 20324
rect 11572 20312 11578 20324
rect 13078 20312 13084 20324
rect 11572 20284 13084 20312
rect 11572 20272 11578 20284
rect 13078 20272 13084 20284
rect 13136 20272 13142 20324
rect 13372 20312 13400 20352
rect 13814 20340 13820 20392
rect 13872 20340 13878 20392
rect 14093 20383 14151 20389
rect 14093 20380 14105 20383
rect 13924 20352 14105 20380
rect 13924 20312 13952 20352
rect 14093 20349 14105 20352
rect 14139 20349 14151 20383
rect 14093 20343 14151 20349
rect 14182 20340 14188 20392
rect 14240 20380 14246 20392
rect 15565 20383 15623 20389
rect 15565 20380 15577 20383
rect 14240 20352 15577 20380
rect 14240 20340 14246 20352
rect 15565 20349 15577 20352
rect 15611 20349 15623 20383
rect 15565 20343 15623 20349
rect 17034 20340 17040 20392
rect 17092 20380 17098 20392
rect 17497 20383 17555 20389
rect 17497 20380 17509 20383
rect 17092 20352 17509 20380
rect 17092 20340 17098 20352
rect 17497 20349 17509 20352
rect 17543 20349 17555 20383
rect 17497 20343 17555 20349
rect 17770 20340 17776 20392
rect 17828 20380 17834 20392
rect 18509 20383 18567 20389
rect 18509 20380 18521 20383
rect 17828 20352 18521 20380
rect 17828 20340 17834 20352
rect 18509 20349 18521 20352
rect 18555 20349 18567 20383
rect 18785 20383 18843 20389
rect 18785 20380 18797 20383
rect 18509 20343 18567 20349
rect 18616 20352 18797 20380
rect 13372 20284 13952 20312
rect 15470 20272 15476 20324
rect 15528 20312 15534 20324
rect 18616 20312 18644 20352
rect 18785 20349 18797 20352
rect 18831 20349 18843 20383
rect 18785 20343 18843 20349
rect 19794 20340 19800 20392
rect 19852 20380 19858 20392
rect 21174 20380 21180 20392
rect 19852 20352 21180 20380
rect 19852 20340 19858 20352
rect 21174 20340 21180 20352
rect 21232 20340 21238 20392
rect 21361 20383 21419 20389
rect 21361 20349 21373 20383
rect 21407 20380 21419 20383
rect 22925 20383 22983 20389
rect 21407 20352 22508 20380
rect 21407 20349 21419 20352
rect 21361 20343 21419 20349
rect 22281 20315 22339 20321
rect 22281 20312 22293 20315
rect 15528 20284 18644 20312
rect 19812 20284 22293 20312
rect 15528 20272 15534 20284
rect 11146 20204 11152 20256
rect 11204 20204 11210 20256
rect 12434 20204 12440 20256
rect 12492 20244 12498 20256
rect 13630 20244 13636 20256
rect 12492 20216 13636 20244
rect 12492 20204 12498 20216
rect 13630 20204 13636 20216
rect 13688 20204 13694 20256
rect 16206 20204 16212 20256
rect 16264 20204 16270 20256
rect 16758 20204 16764 20256
rect 16816 20204 16822 20256
rect 16850 20204 16856 20256
rect 16908 20244 16914 20256
rect 16945 20247 17003 20253
rect 16945 20244 16957 20247
rect 16908 20216 16957 20244
rect 16908 20204 16914 20216
rect 16945 20213 16957 20216
rect 16991 20213 17003 20247
rect 16945 20207 17003 20213
rect 18322 20204 18328 20256
rect 18380 20244 18386 20256
rect 19812 20244 19840 20284
rect 22281 20281 22293 20284
rect 22327 20281 22339 20315
rect 22480 20312 22508 20352
rect 22925 20349 22937 20383
rect 22971 20380 22983 20383
rect 23216 20380 23244 20556
rect 25958 20544 25964 20556
rect 26016 20544 26022 20596
rect 26050 20544 26056 20596
rect 26108 20584 26114 20596
rect 26697 20587 26755 20593
rect 26697 20584 26709 20587
rect 26108 20556 26709 20584
rect 26108 20544 26114 20556
rect 26697 20553 26709 20556
rect 26743 20553 26755 20587
rect 26697 20547 26755 20553
rect 27338 20544 27344 20596
rect 27396 20584 27402 20596
rect 28997 20587 29055 20593
rect 27396 20556 28856 20584
rect 27396 20544 27402 20556
rect 24394 20516 24400 20528
rect 23860 20488 24400 20516
rect 23293 20451 23351 20457
rect 23293 20417 23305 20451
rect 23339 20448 23351 20451
rect 23474 20448 23480 20460
rect 23339 20420 23480 20448
rect 23339 20417 23351 20420
rect 23293 20411 23351 20417
rect 23474 20408 23480 20420
rect 23532 20448 23538 20460
rect 23860 20448 23888 20488
rect 24394 20476 24400 20488
rect 24452 20516 24458 20528
rect 24578 20516 24584 20528
rect 24452 20488 24584 20516
rect 24452 20476 24458 20488
rect 24578 20476 24584 20488
rect 24636 20476 24642 20528
rect 25498 20476 25504 20528
rect 25556 20516 25562 20528
rect 26605 20519 26663 20525
rect 26605 20516 26617 20519
rect 25556 20488 26617 20516
rect 25556 20476 25562 20488
rect 26605 20485 26617 20488
rect 26651 20516 26663 20519
rect 27614 20516 27620 20528
rect 26651 20488 27620 20516
rect 26651 20485 26663 20488
rect 26605 20479 26663 20485
rect 27614 20476 27620 20488
rect 27672 20476 27678 20528
rect 26050 20448 26056 20460
rect 23532 20420 23888 20448
rect 25424 20420 26056 20448
rect 23532 20408 23538 20420
rect 25424 20392 25452 20420
rect 26050 20408 26056 20420
rect 26108 20408 26114 20460
rect 26234 20408 26240 20460
rect 26292 20408 26298 20460
rect 27246 20408 27252 20460
rect 27304 20408 27310 20460
rect 28828 20448 28856 20556
rect 28997 20553 29009 20587
rect 29043 20584 29055 20587
rect 29638 20584 29644 20596
rect 29043 20556 29644 20584
rect 29043 20553 29055 20556
rect 28997 20547 29055 20553
rect 29638 20544 29644 20556
rect 29696 20544 29702 20596
rect 29822 20544 29828 20596
rect 29880 20584 29886 20596
rect 29917 20587 29975 20593
rect 29917 20584 29929 20587
rect 29880 20556 29929 20584
rect 29880 20544 29886 20556
rect 29917 20553 29929 20556
rect 29963 20553 29975 20587
rect 29917 20547 29975 20553
rect 30098 20544 30104 20596
rect 30156 20584 30162 20596
rect 30156 20556 33916 20584
rect 30156 20544 30162 20556
rect 29270 20476 29276 20528
rect 29328 20516 29334 20528
rect 30006 20516 30012 20528
rect 29328 20488 30012 20516
rect 29328 20476 29334 20488
rect 30006 20476 30012 20488
rect 30064 20476 30070 20528
rect 30374 20476 30380 20528
rect 30432 20516 30438 20528
rect 31113 20519 31171 20525
rect 31113 20516 31125 20519
rect 30432 20488 31125 20516
rect 30432 20476 30438 20488
rect 31113 20485 31125 20488
rect 31159 20485 31171 20519
rect 31113 20479 31171 20485
rect 31202 20476 31208 20528
rect 31260 20516 31266 20528
rect 31849 20519 31907 20525
rect 31849 20516 31861 20519
rect 31260 20488 31861 20516
rect 31260 20476 31266 20488
rect 31849 20485 31861 20488
rect 31895 20485 31907 20519
rect 31849 20479 31907 20485
rect 33042 20476 33048 20528
rect 33100 20476 33106 20528
rect 33888 20516 33916 20556
rect 33962 20544 33968 20596
rect 34020 20584 34026 20596
rect 34057 20587 34115 20593
rect 34057 20584 34069 20587
rect 34020 20556 34069 20584
rect 34020 20544 34026 20556
rect 34057 20553 34069 20556
rect 34103 20553 34115 20587
rect 34057 20547 34115 20553
rect 34609 20587 34667 20593
rect 34609 20553 34621 20587
rect 34655 20584 34667 20587
rect 35802 20584 35808 20596
rect 34655 20556 35808 20584
rect 34655 20553 34667 20556
rect 34609 20547 34667 20553
rect 35802 20544 35808 20556
rect 35860 20544 35866 20596
rect 36081 20587 36139 20593
rect 36081 20553 36093 20587
rect 36127 20584 36139 20587
rect 36170 20584 36176 20596
rect 36127 20556 36176 20584
rect 36127 20553 36139 20556
rect 36081 20547 36139 20553
rect 36170 20544 36176 20556
rect 36228 20544 36234 20596
rect 36541 20587 36599 20593
rect 36541 20584 36553 20587
rect 36372 20556 36553 20584
rect 34333 20519 34391 20525
rect 34333 20516 34345 20519
rect 33888 20488 34345 20516
rect 34333 20485 34345 20488
rect 34379 20516 34391 20519
rect 36262 20516 36268 20528
rect 34379 20488 36268 20516
rect 34379 20485 34391 20488
rect 34333 20479 34391 20485
rect 36262 20476 36268 20488
rect 36320 20476 36326 20528
rect 29825 20451 29883 20457
rect 29825 20448 29837 20451
rect 22971 20352 23244 20380
rect 22971 20349 22983 20352
rect 22925 20343 22983 20349
rect 23382 20340 23388 20392
rect 23440 20380 23446 20392
rect 23750 20380 23756 20392
rect 23440 20352 23756 20380
rect 23440 20340 23446 20352
rect 23750 20340 23756 20352
rect 23808 20380 23814 20392
rect 23845 20383 23903 20389
rect 23845 20380 23857 20383
rect 23808 20352 23857 20380
rect 23808 20340 23814 20352
rect 23845 20349 23857 20352
rect 23891 20349 23903 20383
rect 23845 20343 23903 20349
rect 24118 20340 24124 20392
rect 24176 20340 24182 20392
rect 24578 20340 24584 20392
rect 24636 20380 24642 20392
rect 25406 20380 25412 20392
rect 24636 20352 25412 20380
rect 24636 20340 24642 20352
rect 25406 20340 25412 20352
rect 25464 20340 25470 20392
rect 25590 20340 25596 20392
rect 25648 20340 25654 20392
rect 27525 20383 27583 20389
rect 27525 20349 27537 20383
rect 27571 20380 27583 20383
rect 28534 20380 28540 20392
rect 27571 20352 28540 20380
rect 27571 20349 27583 20352
rect 27525 20343 27583 20349
rect 28534 20340 28540 20352
rect 28592 20340 28598 20392
rect 28644 20380 28672 20434
rect 28828 20420 29837 20448
rect 29825 20417 29837 20420
rect 29871 20417 29883 20451
rect 29825 20411 29883 20417
rect 31021 20451 31079 20457
rect 31021 20417 31033 20451
rect 31067 20417 31079 20451
rect 31021 20411 31079 20417
rect 29270 20380 29276 20392
rect 28644 20352 29276 20380
rect 29270 20340 29276 20352
rect 29328 20340 29334 20392
rect 29730 20340 29736 20392
rect 29788 20380 29794 20392
rect 30101 20383 30159 20389
rect 30101 20380 30113 20383
rect 29788 20352 30113 20380
rect 29788 20340 29794 20352
rect 30101 20349 30113 20352
rect 30147 20380 30159 20383
rect 30190 20380 30196 20392
rect 30147 20352 30196 20380
rect 30147 20349 30159 20352
rect 30101 20343 30159 20349
rect 30190 20340 30196 20352
rect 30248 20340 30254 20392
rect 26053 20315 26111 20321
rect 22480 20284 23980 20312
rect 22281 20275 22339 20281
rect 18380 20216 19840 20244
rect 20257 20247 20315 20253
rect 18380 20204 18386 20216
rect 20257 20213 20269 20247
rect 20303 20244 20315 20247
rect 20346 20244 20352 20256
rect 20303 20216 20352 20244
rect 20303 20213 20315 20216
rect 20257 20207 20315 20213
rect 20346 20204 20352 20216
rect 20404 20204 20410 20256
rect 21082 20204 21088 20256
rect 21140 20244 21146 20256
rect 23842 20244 23848 20256
rect 21140 20216 23848 20244
rect 21140 20204 21146 20216
rect 23842 20204 23848 20216
rect 23900 20204 23906 20256
rect 23952 20244 23980 20284
rect 26053 20281 26065 20315
rect 26099 20312 26111 20315
rect 27246 20312 27252 20324
rect 26099 20284 27252 20312
rect 26099 20281 26111 20284
rect 26053 20275 26111 20281
rect 27246 20272 27252 20284
rect 27304 20272 27310 20324
rect 29457 20315 29515 20321
rect 29457 20281 29469 20315
rect 29503 20312 29515 20315
rect 30374 20312 30380 20324
rect 29503 20284 30380 20312
rect 29503 20281 29515 20284
rect 29457 20275 29515 20281
rect 30374 20272 30380 20284
rect 30432 20272 30438 20324
rect 31036 20312 31064 20411
rect 34698 20408 34704 20460
rect 34756 20448 34762 20460
rect 35250 20448 35256 20460
rect 34756 20420 35256 20448
rect 34756 20408 34762 20420
rect 35250 20408 35256 20420
rect 35308 20408 35314 20460
rect 35345 20451 35403 20457
rect 35345 20417 35357 20451
rect 35391 20448 35403 20451
rect 35618 20448 35624 20460
rect 35391 20420 35624 20448
rect 35391 20417 35403 20420
rect 35345 20411 35403 20417
rect 35618 20408 35624 20420
rect 35676 20408 35682 20460
rect 35802 20408 35808 20460
rect 35860 20448 35866 20460
rect 36372 20448 36400 20556
rect 36541 20553 36553 20556
rect 36587 20584 36599 20587
rect 37274 20584 37280 20596
rect 36587 20556 37280 20584
rect 36587 20553 36599 20556
rect 36541 20547 36599 20553
rect 37274 20544 37280 20556
rect 37332 20584 37338 20596
rect 37918 20584 37924 20596
rect 37332 20556 37924 20584
rect 37332 20544 37338 20556
rect 37918 20544 37924 20556
rect 37976 20544 37982 20596
rect 42058 20584 42064 20596
rect 38028 20556 42064 20584
rect 38028 20525 38056 20556
rect 42058 20544 42064 20556
rect 42116 20544 42122 20596
rect 42150 20544 42156 20596
rect 42208 20584 42214 20596
rect 42702 20584 42708 20596
rect 42208 20556 42708 20584
rect 42208 20544 42214 20556
rect 42702 20544 42708 20556
rect 42760 20584 42766 20596
rect 43073 20587 43131 20593
rect 43073 20584 43085 20587
rect 42760 20556 43085 20584
rect 42760 20544 42766 20556
rect 43073 20553 43085 20556
rect 43119 20553 43131 20587
rect 43073 20547 43131 20553
rect 43806 20544 43812 20596
rect 43864 20544 43870 20596
rect 44269 20587 44327 20593
rect 44269 20553 44281 20587
rect 44315 20584 44327 20587
rect 44450 20584 44456 20596
rect 44315 20556 44456 20584
rect 44315 20553 44327 20556
rect 44269 20547 44327 20553
rect 44450 20544 44456 20556
rect 44508 20544 44514 20596
rect 44637 20587 44695 20593
rect 44637 20553 44649 20587
rect 44683 20584 44695 20587
rect 44726 20584 44732 20596
rect 44683 20556 44732 20584
rect 44683 20553 44695 20556
rect 44637 20547 44695 20553
rect 44726 20544 44732 20556
rect 44784 20544 44790 20596
rect 44818 20544 44824 20596
rect 44876 20544 44882 20596
rect 46569 20587 46627 20593
rect 46569 20553 46581 20587
rect 46615 20584 46627 20587
rect 46750 20584 46756 20596
rect 46615 20556 46756 20584
rect 46615 20553 46627 20556
rect 46569 20547 46627 20553
rect 46750 20544 46756 20556
rect 46808 20544 46814 20596
rect 47029 20587 47087 20593
rect 47029 20553 47041 20587
rect 47075 20584 47087 20587
rect 47118 20584 47124 20596
rect 47075 20556 47124 20584
rect 47075 20553 47087 20556
rect 47029 20547 47087 20553
rect 47118 20544 47124 20556
rect 47176 20544 47182 20596
rect 47670 20544 47676 20596
rect 47728 20584 47734 20596
rect 48041 20587 48099 20593
rect 48041 20584 48053 20587
rect 47728 20556 48053 20584
rect 47728 20544 47734 20556
rect 48041 20553 48053 20556
rect 48087 20553 48099 20587
rect 48041 20547 48099 20553
rect 38013 20519 38071 20525
rect 38013 20485 38025 20519
rect 38059 20485 38071 20519
rect 38013 20479 38071 20485
rect 38746 20476 38752 20528
rect 38804 20476 38810 20528
rect 39758 20476 39764 20528
rect 39816 20516 39822 20528
rect 40310 20516 40316 20528
rect 39816 20488 40316 20516
rect 39816 20476 39822 20488
rect 40310 20476 40316 20488
rect 40368 20476 40374 20528
rect 42613 20519 42671 20525
rect 42613 20516 42625 20519
rect 40420 20488 42625 20516
rect 35860 20420 36400 20448
rect 36449 20451 36507 20457
rect 35860 20408 35866 20420
rect 36449 20417 36461 20451
rect 36495 20448 36507 20451
rect 36814 20448 36820 20460
rect 36495 20420 36820 20448
rect 36495 20417 36507 20420
rect 36449 20411 36507 20417
rect 31202 20340 31208 20392
rect 31260 20340 31266 20392
rect 32306 20340 32312 20392
rect 32364 20340 32370 20392
rect 32585 20383 32643 20389
rect 32585 20349 32597 20383
rect 32631 20380 32643 20383
rect 32674 20380 32680 20392
rect 32631 20352 32680 20380
rect 32631 20349 32643 20352
rect 32585 20343 32643 20349
rect 32674 20340 32680 20352
rect 32732 20340 32738 20392
rect 35529 20383 35587 20389
rect 35529 20349 35541 20383
rect 35575 20349 35587 20383
rect 35529 20343 35587 20349
rect 31110 20312 31116 20324
rect 31036 20284 31116 20312
rect 31110 20272 31116 20284
rect 31168 20312 31174 20324
rect 31168 20284 31800 20312
rect 31168 20272 31174 20284
rect 25774 20244 25780 20256
rect 23952 20216 25780 20244
rect 25774 20204 25780 20216
rect 25832 20204 25838 20256
rect 27062 20204 27068 20256
rect 27120 20244 27126 20256
rect 27706 20244 27712 20256
rect 27120 20216 27712 20244
rect 27120 20204 27126 20216
rect 27706 20204 27712 20216
rect 27764 20204 27770 20256
rect 29178 20204 29184 20256
rect 29236 20244 29242 20256
rect 30282 20244 30288 20256
rect 29236 20216 30288 20244
rect 29236 20204 29242 20216
rect 30282 20204 30288 20216
rect 30340 20204 30346 20256
rect 30650 20204 30656 20256
rect 30708 20204 30714 20256
rect 30926 20204 30932 20256
rect 30984 20244 30990 20256
rect 31665 20247 31723 20253
rect 31665 20244 31677 20247
rect 30984 20216 31677 20244
rect 30984 20204 30990 20216
rect 31665 20213 31677 20216
rect 31711 20213 31723 20247
rect 31772 20244 31800 20284
rect 33686 20272 33692 20324
rect 33744 20312 33750 20324
rect 35544 20312 35572 20343
rect 35710 20340 35716 20392
rect 35768 20380 35774 20392
rect 36464 20380 36492 20411
rect 36814 20408 36820 20420
rect 36872 20408 36878 20460
rect 37182 20408 37188 20460
rect 37240 20448 37246 20460
rect 37277 20451 37335 20457
rect 37277 20448 37289 20451
rect 37240 20420 37289 20448
rect 37240 20408 37246 20420
rect 37277 20417 37289 20420
rect 37323 20417 37335 20451
rect 40420 20448 40448 20488
rect 42613 20485 42625 20488
rect 42659 20485 42671 20519
rect 42613 20479 42671 20485
rect 43898 20476 43904 20528
rect 43956 20516 43962 20528
rect 44361 20519 44419 20525
rect 44361 20516 44373 20519
rect 43956 20488 44373 20516
rect 43956 20476 43962 20488
rect 44361 20485 44373 20488
rect 44407 20485 44419 20519
rect 44361 20479 44419 20485
rect 46382 20476 46388 20528
rect 46440 20516 46446 20528
rect 46661 20519 46719 20525
rect 46661 20516 46673 20519
rect 46440 20488 46673 20516
rect 46440 20476 46446 20488
rect 46661 20485 46673 20488
rect 46707 20485 46719 20519
rect 46661 20479 46719 20485
rect 47213 20519 47271 20525
rect 47213 20485 47225 20519
rect 47259 20516 47271 20519
rect 49326 20516 49332 20528
rect 47259 20488 49332 20516
rect 47259 20485 47271 20488
rect 47213 20479 47271 20485
rect 49326 20476 49332 20488
rect 49384 20476 49390 20528
rect 37277 20411 37335 20417
rect 40328 20420 40448 20448
rect 35768 20352 36492 20380
rect 35768 20340 35774 20352
rect 36722 20340 36728 20392
rect 36780 20340 36786 20392
rect 37734 20340 37740 20392
rect 37792 20340 37798 20392
rect 40328 20380 40356 20420
rect 40954 20408 40960 20460
rect 41012 20448 41018 20460
rect 41141 20451 41199 20457
rect 41141 20448 41153 20451
rect 41012 20420 41153 20448
rect 41012 20408 41018 20420
rect 41141 20417 41153 20420
rect 41187 20417 41199 20451
rect 43533 20451 43591 20457
rect 43533 20448 43545 20451
rect 41141 20411 41199 20417
rect 41386 20420 43545 20448
rect 37844 20352 40356 20380
rect 40405 20383 40463 20389
rect 33744 20284 35572 20312
rect 33744 20272 33750 20284
rect 36446 20272 36452 20324
rect 36504 20312 36510 20324
rect 37844 20312 37872 20352
rect 40405 20349 40417 20383
rect 40451 20349 40463 20383
rect 40405 20343 40463 20349
rect 40589 20383 40647 20389
rect 40589 20349 40601 20383
rect 40635 20380 40647 20383
rect 41046 20380 41052 20392
rect 40635 20352 41052 20380
rect 40635 20349 40647 20352
rect 40589 20343 40647 20349
rect 36504 20284 37872 20312
rect 36504 20272 36510 20284
rect 39022 20272 39028 20324
rect 39080 20312 39086 20324
rect 40420 20312 40448 20343
rect 41046 20340 41052 20352
rect 41104 20340 41110 20392
rect 41138 20312 41144 20324
rect 39080 20284 40080 20312
rect 40420 20284 41144 20312
rect 39080 20272 39086 20284
rect 34054 20244 34060 20256
rect 31772 20216 34060 20244
rect 31665 20207 31723 20213
rect 34054 20204 34060 20216
rect 34112 20204 34118 20256
rect 34885 20247 34943 20253
rect 34885 20213 34897 20247
rect 34931 20244 34943 20247
rect 35526 20244 35532 20256
rect 34931 20216 35532 20244
rect 34931 20213 34943 20216
rect 34885 20207 34943 20213
rect 35526 20204 35532 20216
rect 35584 20204 35590 20256
rect 36078 20204 36084 20256
rect 36136 20244 36142 20256
rect 39485 20247 39543 20253
rect 39485 20244 39497 20247
rect 36136 20216 39497 20244
rect 36136 20204 36142 20216
rect 39485 20213 39497 20216
rect 39531 20244 39543 20247
rect 39758 20244 39764 20256
rect 39531 20216 39764 20244
rect 39531 20213 39543 20216
rect 39485 20207 39543 20213
rect 39758 20204 39764 20216
rect 39816 20204 39822 20256
rect 39942 20204 39948 20256
rect 40000 20204 40006 20256
rect 40052 20244 40080 20284
rect 41138 20272 41144 20284
rect 41196 20312 41202 20324
rect 41386 20312 41414 20420
rect 43533 20417 43545 20420
rect 43579 20448 43591 20451
rect 44082 20448 44088 20460
rect 43579 20420 44088 20448
rect 43579 20417 43591 20420
rect 43533 20411 43591 20417
rect 44082 20408 44088 20420
rect 44140 20408 44146 20460
rect 47026 20408 47032 20460
rect 47084 20448 47090 20460
rect 47305 20451 47363 20457
rect 47305 20448 47317 20451
rect 47084 20420 47317 20448
rect 47084 20408 47090 20420
rect 47305 20417 47317 20420
rect 47351 20417 47363 20451
rect 47305 20411 47363 20417
rect 47949 20451 48007 20457
rect 47949 20417 47961 20451
rect 47995 20448 48007 20451
rect 48590 20448 48596 20460
rect 47995 20420 48596 20448
rect 47995 20417 48007 20420
rect 47949 20411 48007 20417
rect 48590 20408 48596 20420
rect 48648 20408 48654 20460
rect 49050 20408 49056 20460
rect 49108 20408 49114 20460
rect 41506 20340 41512 20392
rect 41564 20380 41570 20392
rect 42610 20380 42616 20392
rect 41564 20352 42616 20380
rect 41564 20340 41570 20352
rect 42610 20340 42616 20352
rect 42668 20340 42674 20392
rect 42978 20340 42984 20392
rect 43036 20380 43042 20392
rect 43717 20383 43775 20389
rect 43717 20380 43729 20383
rect 43036 20352 43729 20380
rect 43036 20340 43042 20352
rect 43717 20349 43729 20352
rect 43763 20380 43775 20383
rect 45554 20380 45560 20392
rect 43763 20352 45560 20380
rect 43763 20349 43775 20352
rect 43717 20343 43775 20349
rect 45554 20340 45560 20352
rect 45612 20340 45618 20392
rect 47765 20383 47823 20389
rect 47765 20349 47777 20383
rect 47811 20380 47823 20383
rect 49068 20380 49096 20408
rect 47811 20352 49096 20380
rect 47811 20349 47823 20352
rect 47765 20343 47823 20349
rect 41966 20312 41972 20324
rect 41196 20284 41414 20312
rect 41708 20284 41972 20312
rect 41196 20272 41202 20284
rect 41708 20244 41736 20284
rect 41966 20272 41972 20284
rect 42024 20272 42030 20324
rect 43254 20272 43260 20324
rect 43312 20312 43318 20324
rect 43349 20315 43407 20321
rect 43349 20312 43361 20315
rect 43312 20284 43361 20312
rect 43312 20272 43318 20284
rect 43349 20281 43361 20284
rect 43395 20312 43407 20315
rect 49237 20315 49295 20321
rect 49237 20312 49249 20315
rect 43395 20284 49249 20312
rect 43395 20281 43407 20284
rect 43349 20275 43407 20281
rect 49237 20281 49249 20284
rect 49283 20281 49295 20315
rect 49237 20275 49295 20281
rect 40052 20216 41736 20244
rect 41782 20204 41788 20256
rect 41840 20204 41846 20256
rect 48314 20204 48320 20256
rect 48372 20244 48378 20256
rect 48409 20247 48467 20253
rect 48409 20244 48421 20247
rect 48372 20216 48421 20244
rect 48372 20204 48378 20216
rect 48409 20213 48421 20216
rect 48455 20213 48467 20247
rect 48409 20207 48467 20213
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 3602 20000 3608 20052
rect 3660 20040 3666 20052
rect 10321 20043 10379 20049
rect 10321 20040 10333 20043
rect 3660 20012 10333 20040
rect 3660 20000 3666 20012
rect 10321 20009 10333 20012
rect 10367 20009 10379 20043
rect 10321 20003 10379 20009
rect 11146 20000 11152 20052
rect 11204 20040 11210 20052
rect 12234 20043 12292 20049
rect 12234 20040 12246 20043
rect 11204 20012 12246 20040
rect 11204 20000 11210 20012
rect 12234 20009 12246 20012
rect 12280 20009 12292 20043
rect 12234 20003 12292 20009
rect 12342 20000 12348 20052
rect 12400 20040 12406 20052
rect 12434 20040 12440 20052
rect 12400 20012 12440 20040
rect 12400 20000 12406 20012
rect 12434 20000 12440 20012
rect 12492 20000 12498 20052
rect 12618 20000 12624 20052
rect 12676 20040 12682 20052
rect 15378 20040 15384 20052
rect 12676 20012 15384 20040
rect 12676 20000 12682 20012
rect 15378 20000 15384 20012
rect 15436 20000 15442 20052
rect 15470 20000 15476 20052
rect 15528 20000 15534 20052
rect 16942 20000 16948 20052
rect 17000 20040 17006 20052
rect 18785 20043 18843 20049
rect 18785 20040 18797 20043
rect 17000 20012 18797 20040
rect 17000 20000 17006 20012
rect 18785 20009 18797 20012
rect 18831 20009 18843 20043
rect 18785 20003 18843 20009
rect 19518 20000 19524 20052
rect 19576 20040 19582 20052
rect 19889 20043 19947 20049
rect 19889 20040 19901 20043
rect 19576 20012 19901 20040
rect 19576 20000 19582 20012
rect 19889 20009 19901 20012
rect 19935 20009 19947 20043
rect 19889 20003 19947 20009
rect 21266 20000 21272 20052
rect 21324 20040 21330 20052
rect 26694 20040 26700 20052
rect 21324 20012 26700 20040
rect 21324 20000 21330 20012
rect 26694 20000 26700 20012
rect 26752 20000 26758 20052
rect 26786 20000 26792 20052
rect 26844 20000 26850 20052
rect 27706 20000 27712 20052
rect 27764 20040 27770 20052
rect 28810 20040 28816 20052
rect 27764 20012 28816 20040
rect 27764 20000 27770 20012
rect 28810 20000 28816 20012
rect 28868 20000 28874 20052
rect 29270 20000 29276 20052
rect 29328 20000 29334 20052
rect 29362 20000 29368 20052
rect 29420 20040 29426 20052
rect 30929 20043 30987 20049
rect 29420 20012 30880 20040
rect 29420 20000 29426 20012
rect 5258 19932 5264 19984
rect 5316 19972 5322 19984
rect 10410 19972 10416 19984
rect 5316 19944 10416 19972
rect 5316 19932 5322 19944
rect 10410 19932 10416 19944
rect 10468 19932 10474 19984
rect 14185 19975 14243 19981
rect 14185 19972 14197 19975
rect 13372 19944 14197 19972
rect 4522 19864 4528 19916
rect 4580 19864 4586 19916
rect 6178 19864 6184 19916
rect 6236 19904 6242 19916
rect 6273 19907 6331 19913
rect 6273 19904 6285 19907
rect 6236 19876 6285 19904
rect 6236 19864 6242 19876
rect 6273 19873 6285 19876
rect 6319 19873 6331 19907
rect 6273 19867 6331 19873
rect 6362 19864 6368 19916
rect 6420 19904 6426 19916
rect 9950 19904 9956 19916
rect 6420 19876 9956 19904
rect 6420 19864 6426 19876
rect 9950 19864 9956 19876
rect 10008 19864 10014 19916
rect 11977 19907 12035 19913
rect 11977 19873 11989 19907
rect 12023 19904 12035 19907
rect 12342 19904 12348 19916
rect 12023 19876 12348 19904
rect 12023 19873 12035 19876
rect 11977 19867 12035 19873
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 1762 19796 1768 19848
rect 1820 19796 1826 19848
rect 4065 19839 4123 19845
rect 4065 19805 4077 19839
rect 4111 19836 4123 19839
rect 5718 19836 5724 19848
rect 4111 19808 5724 19836
rect 4111 19805 4123 19808
rect 4065 19799 4123 19805
rect 5718 19796 5724 19808
rect 5776 19796 5782 19848
rect 5994 19796 6000 19848
rect 6052 19796 6058 19848
rect 7834 19796 7840 19848
rect 7892 19796 7898 19848
rect 7926 19796 7932 19848
rect 7984 19836 7990 19848
rect 8389 19839 8447 19845
rect 8389 19836 8401 19839
rect 7984 19808 8401 19836
rect 7984 19796 7990 19808
rect 8389 19805 8401 19808
rect 8435 19836 8447 19839
rect 10873 19839 10931 19845
rect 8435 19808 10364 19836
rect 8435 19805 8447 19808
rect 8389 19799 8447 19805
rect 2774 19728 2780 19780
rect 2832 19728 2838 19780
rect 4246 19728 4252 19780
rect 4304 19768 4310 19780
rect 9861 19771 9919 19777
rect 4304 19740 7788 19768
rect 4304 19728 4310 19740
rect 7650 19660 7656 19712
rect 7708 19660 7714 19712
rect 7760 19700 7788 19740
rect 9861 19737 9873 19771
rect 9907 19768 9919 19771
rect 10134 19768 10140 19780
rect 9907 19740 10140 19768
rect 9907 19737 9919 19740
rect 9861 19731 9919 19737
rect 10134 19728 10140 19740
rect 10192 19728 10198 19780
rect 10229 19771 10287 19777
rect 10229 19737 10241 19771
rect 10275 19737 10287 19771
rect 10336 19768 10364 19808
rect 10873 19805 10885 19839
rect 10919 19836 10931 19839
rect 11698 19836 11704 19848
rect 10919 19808 11704 19836
rect 10919 19805 10931 19808
rect 10873 19799 10931 19805
rect 11698 19796 11704 19808
rect 11756 19796 11762 19848
rect 13372 19822 13400 19944
rect 14185 19941 14197 19944
rect 14231 19972 14243 19975
rect 14366 19972 14372 19984
rect 14231 19944 14372 19972
rect 14231 19941 14243 19944
rect 14185 19935 14243 19941
rect 14366 19932 14372 19944
rect 14424 19972 14430 19984
rect 15194 19972 15200 19984
rect 14424 19944 15200 19972
rect 14424 19932 14430 19944
rect 15194 19932 15200 19944
rect 15252 19972 15258 19984
rect 15838 19972 15844 19984
rect 15252 19944 15844 19972
rect 15252 19932 15258 19944
rect 15838 19932 15844 19944
rect 15896 19932 15902 19984
rect 19429 19975 19487 19981
rect 19429 19941 19441 19975
rect 19475 19972 19487 19975
rect 19794 19972 19800 19984
rect 19475 19944 19800 19972
rect 19475 19941 19487 19944
rect 19429 19935 19487 19941
rect 19794 19932 19800 19944
rect 19852 19932 19858 19984
rect 21818 19932 21824 19984
rect 21876 19972 21882 19984
rect 23201 19975 23259 19981
rect 23201 19972 23213 19975
rect 21876 19944 23213 19972
rect 21876 19932 21882 19944
rect 23201 19941 23213 19944
rect 23247 19941 23259 19975
rect 23934 19972 23940 19984
rect 23201 19935 23259 19941
rect 23676 19944 23940 19972
rect 13814 19864 13820 19916
rect 13872 19904 13878 19916
rect 17037 19907 17095 19913
rect 17037 19904 17049 19907
rect 13872 19876 17049 19904
rect 13872 19864 13878 19876
rect 17037 19873 17049 19876
rect 17083 19904 17095 19907
rect 17770 19904 17776 19916
rect 17083 19876 17776 19904
rect 17083 19873 17095 19876
rect 17037 19867 17095 19873
rect 17770 19864 17776 19876
rect 17828 19864 17834 19916
rect 17862 19864 17868 19916
rect 17920 19904 17926 19916
rect 20717 19907 20775 19913
rect 17920 19876 20392 19904
rect 17920 19864 17926 19876
rect 13630 19796 13636 19848
rect 13688 19836 13694 19848
rect 14090 19836 14096 19848
rect 13688 19808 14096 19836
rect 13688 19796 13694 19808
rect 14090 19796 14096 19808
rect 14148 19796 14154 19848
rect 14829 19839 14887 19845
rect 14829 19805 14841 19839
rect 14875 19805 14887 19839
rect 14829 19799 14887 19805
rect 14844 19768 14872 19799
rect 15930 19796 15936 19848
rect 15988 19796 15994 19848
rect 16942 19836 16948 19848
rect 16224 19808 16948 19836
rect 16224 19768 16252 19808
rect 16942 19796 16948 19808
rect 17000 19796 17006 19848
rect 18414 19796 18420 19848
rect 18472 19796 18478 19848
rect 10336 19740 12434 19768
rect 14844 19740 16252 19768
rect 10229 19731 10287 19737
rect 8481 19703 8539 19709
rect 8481 19700 8493 19703
rect 7760 19672 8493 19700
rect 8481 19669 8493 19672
rect 8527 19669 8539 19703
rect 8481 19663 8539 19669
rect 9125 19703 9183 19709
rect 9125 19669 9137 19703
rect 9171 19700 9183 19703
rect 9214 19700 9220 19712
rect 9171 19672 9220 19700
rect 9171 19669 9183 19672
rect 9125 19663 9183 19669
rect 9214 19660 9220 19672
rect 9272 19660 9278 19712
rect 10244 19700 10272 19731
rect 12406 19712 12434 19740
rect 16298 19728 16304 19780
rect 16356 19768 16362 19780
rect 17313 19771 17371 19777
rect 17313 19768 17325 19771
rect 16356 19740 17325 19768
rect 16356 19728 16362 19740
rect 17313 19737 17325 19740
rect 17359 19737 17371 19771
rect 17313 19731 17371 19737
rect 18598 19728 18604 19780
rect 18656 19768 18662 19780
rect 19797 19771 19855 19777
rect 18656 19740 19748 19768
rect 18656 19728 18662 19740
rect 10594 19700 10600 19712
rect 10244 19672 10600 19700
rect 10594 19660 10600 19672
rect 10652 19660 10658 19712
rect 10778 19660 10784 19712
rect 10836 19700 10842 19712
rect 11517 19703 11575 19709
rect 11517 19700 11529 19703
rect 10836 19672 11529 19700
rect 10836 19660 10842 19672
rect 11517 19669 11529 19672
rect 11563 19669 11575 19703
rect 12406 19672 12440 19712
rect 11517 19663 11575 19669
rect 12434 19660 12440 19672
rect 12492 19660 12498 19712
rect 12526 19660 12532 19712
rect 12584 19700 12590 19712
rect 13630 19700 13636 19712
rect 12584 19672 13636 19700
rect 12584 19660 12590 19672
rect 13630 19660 13636 19672
rect 13688 19700 13694 19712
rect 13725 19703 13783 19709
rect 13725 19700 13737 19703
rect 13688 19672 13737 19700
rect 13688 19660 13694 19672
rect 13725 19669 13737 19672
rect 13771 19669 13783 19703
rect 13725 19663 13783 19669
rect 14553 19703 14611 19709
rect 14553 19669 14565 19703
rect 14599 19700 14611 19703
rect 15102 19700 15108 19712
rect 14599 19672 15108 19700
rect 14599 19669 14611 19672
rect 14553 19663 14611 19669
rect 15102 19660 15108 19672
rect 15160 19660 15166 19712
rect 16577 19703 16635 19709
rect 16577 19669 16589 19703
rect 16623 19700 16635 19703
rect 17586 19700 17592 19712
rect 16623 19672 17592 19700
rect 16623 19669 16635 19672
rect 16577 19663 16635 19669
rect 17586 19660 17592 19672
rect 17644 19660 17650 19712
rect 19720 19700 19748 19740
rect 19797 19737 19809 19771
rect 19843 19768 19855 19771
rect 19886 19768 19892 19780
rect 19843 19740 19892 19768
rect 19843 19737 19855 19740
rect 19797 19731 19855 19737
rect 19886 19728 19892 19740
rect 19944 19728 19950 19780
rect 20364 19768 20392 19876
rect 20717 19873 20729 19907
rect 20763 19904 20775 19907
rect 23676 19904 23704 19944
rect 23934 19932 23940 19944
rect 23992 19932 23998 19984
rect 24118 19932 24124 19984
rect 24176 19972 24182 19984
rect 24176 19944 28856 19972
rect 24176 19932 24182 19944
rect 20763 19876 23704 19904
rect 20763 19873 20775 19876
rect 20717 19867 20775 19873
rect 23750 19864 23756 19916
rect 23808 19864 23814 19916
rect 25222 19904 25228 19916
rect 24504 19876 25228 19904
rect 20438 19796 20444 19848
rect 20496 19796 20502 19848
rect 21726 19796 21732 19848
rect 21784 19836 21790 19848
rect 21784 19808 21850 19836
rect 21784 19796 21790 19808
rect 22462 19796 22468 19848
rect 22520 19836 22526 19848
rect 24504 19836 24532 19876
rect 25222 19864 25228 19876
rect 25280 19904 25286 19916
rect 27356 19913 27384 19944
rect 26145 19907 26203 19913
rect 26145 19904 26157 19907
rect 25280 19876 26157 19904
rect 25280 19864 25286 19876
rect 26145 19873 26157 19876
rect 26191 19873 26203 19907
rect 26145 19867 26203 19873
rect 27341 19907 27399 19913
rect 27341 19873 27353 19907
rect 27387 19873 27399 19907
rect 27341 19867 27399 19873
rect 28626 19864 28632 19916
rect 28684 19864 28690 19916
rect 28828 19904 28856 19944
rect 28902 19932 28908 19984
rect 28960 19972 28966 19984
rect 29733 19975 29791 19981
rect 29733 19972 29745 19975
rect 28960 19944 29745 19972
rect 28960 19932 28966 19944
rect 29733 19941 29745 19944
rect 29779 19941 29791 19975
rect 30852 19972 30880 20012
rect 30929 20009 30941 20043
rect 30975 20040 30987 20043
rect 33502 20040 33508 20052
rect 30975 20012 33508 20040
rect 30975 20009 30987 20012
rect 30929 20003 30987 20009
rect 33502 20000 33508 20012
rect 33560 20000 33566 20052
rect 33962 20000 33968 20052
rect 34020 20040 34026 20052
rect 34020 20012 34652 20040
rect 34020 20000 34026 20012
rect 33413 19975 33471 19981
rect 30852 19944 31754 19972
rect 29733 19935 29791 19941
rect 29454 19904 29460 19916
rect 28828 19876 29460 19904
rect 29454 19864 29460 19876
rect 29512 19864 29518 19916
rect 29638 19864 29644 19916
rect 29696 19904 29702 19916
rect 30285 19907 30343 19913
rect 30285 19904 30297 19907
rect 29696 19876 30297 19904
rect 29696 19864 29702 19876
rect 30285 19873 30297 19876
rect 30331 19873 30343 19907
rect 30285 19867 30343 19873
rect 31386 19864 31392 19916
rect 31444 19864 31450 19916
rect 31478 19864 31484 19916
rect 31536 19864 31542 19916
rect 22520 19808 24532 19836
rect 22520 19796 22526 19808
rect 24670 19796 24676 19848
rect 24728 19796 24734 19848
rect 25133 19839 25191 19845
rect 25133 19805 25145 19839
rect 25179 19836 25191 19839
rect 27522 19836 27528 19848
rect 25179 19808 27528 19836
rect 25179 19805 25191 19808
rect 25133 19799 25191 19805
rect 27522 19796 27528 19808
rect 27580 19796 27586 19848
rect 27893 19839 27951 19845
rect 27893 19805 27905 19839
rect 27939 19836 27951 19839
rect 28445 19839 28503 19845
rect 28445 19836 28457 19839
rect 27939 19808 28457 19836
rect 27939 19805 27951 19808
rect 27893 19799 27951 19805
rect 28445 19805 28457 19808
rect 28491 19836 28503 19839
rect 28810 19836 28816 19848
rect 28491 19808 28816 19836
rect 28491 19805 28503 19808
rect 28445 19799 28503 19805
rect 28810 19796 28816 19808
rect 28868 19796 28874 19848
rect 30190 19796 30196 19848
rect 30248 19796 30254 19848
rect 30374 19796 30380 19848
rect 30432 19836 30438 19848
rect 31018 19836 31024 19848
rect 30432 19808 31024 19836
rect 30432 19796 30438 19808
rect 31018 19796 31024 19808
rect 31076 19796 31082 19848
rect 31294 19796 31300 19848
rect 31352 19796 31358 19848
rect 20990 19768 20996 19780
rect 20364 19740 20996 19768
rect 20990 19728 20996 19740
rect 21048 19728 21054 19780
rect 22094 19728 22100 19780
rect 22152 19768 22158 19780
rect 22649 19771 22707 19777
rect 22649 19768 22661 19771
rect 22152 19740 22661 19768
rect 22152 19728 22158 19740
rect 22649 19737 22661 19740
rect 22695 19737 22707 19771
rect 22649 19731 22707 19737
rect 22925 19771 22983 19777
rect 22925 19737 22937 19771
rect 22971 19768 22983 19771
rect 23290 19768 23296 19780
rect 22971 19740 23296 19768
rect 22971 19737 22983 19740
rect 22925 19731 22983 19737
rect 23290 19728 23296 19740
rect 23348 19728 23354 19780
rect 23661 19771 23719 19777
rect 23661 19737 23673 19771
rect 23707 19768 23719 19771
rect 28353 19771 28411 19777
rect 23707 19740 28028 19768
rect 23707 19737 23719 19740
rect 23661 19731 23719 19737
rect 21726 19700 21732 19712
rect 19720 19672 21732 19700
rect 21726 19660 21732 19672
rect 21784 19660 21790 19712
rect 22002 19660 22008 19712
rect 22060 19700 22066 19712
rect 22189 19703 22247 19709
rect 22189 19700 22201 19703
rect 22060 19672 22201 19700
rect 22060 19660 22066 19672
rect 22189 19669 22201 19672
rect 22235 19669 22247 19703
rect 22189 19663 22247 19669
rect 22462 19660 22468 19712
rect 22520 19660 22526 19712
rect 23566 19660 23572 19712
rect 23624 19660 23630 19712
rect 24486 19660 24492 19712
rect 24544 19660 24550 19712
rect 24946 19660 24952 19712
rect 25004 19660 25010 19712
rect 25038 19660 25044 19712
rect 25096 19700 25102 19712
rect 25593 19703 25651 19709
rect 25593 19700 25605 19703
rect 25096 19672 25605 19700
rect 25096 19660 25102 19672
rect 25593 19669 25605 19672
rect 25639 19669 25651 19703
rect 25593 19663 25651 19669
rect 25774 19660 25780 19712
rect 25832 19700 25838 19712
rect 25961 19703 26019 19709
rect 25961 19700 25973 19703
rect 25832 19672 25973 19700
rect 25832 19660 25838 19672
rect 25961 19669 25973 19672
rect 26007 19669 26019 19703
rect 25961 19663 26019 19669
rect 26053 19703 26111 19709
rect 26053 19669 26065 19703
rect 26099 19700 26111 19703
rect 26234 19700 26240 19712
rect 26099 19672 26240 19700
rect 26099 19669 26111 19672
rect 26053 19663 26111 19669
rect 26234 19660 26240 19672
rect 26292 19660 26298 19712
rect 27062 19660 27068 19712
rect 27120 19700 27126 19712
rect 27157 19703 27215 19709
rect 27157 19700 27169 19703
rect 27120 19672 27169 19700
rect 27120 19660 27126 19672
rect 27157 19669 27169 19672
rect 27203 19669 27215 19703
rect 27157 19663 27215 19669
rect 27246 19660 27252 19712
rect 27304 19660 27310 19712
rect 28000 19709 28028 19740
rect 28353 19737 28365 19771
rect 28399 19768 28411 19771
rect 31202 19768 31208 19780
rect 28399 19740 31208 19768
rect 28399 19737 28411 19740
rect 28353 19731 28411 19737
rect 31202 19728 31208 19740
rect 31260 19728 31266 19780
rect 31726 19768 31754 19944
rect 33413 19941 33425 19975
rect 33459 19972 33471 19975
rect 34422 19972 34428 19984
rect 33459 19944 34428 19972
rect 33459 19941 33471 19944
rect 33413 19935 33471 19941
rect 34422 19932 34428 19944
rect 34480 19932 34486 19984
rect 34624 19972 34652 20012
rect 34698 20000 34704 20052
rect 34756 20040 34762 20052
rect 35342 20040 35348 20052
rect 34756 20012 35348 20040
rect 34756 20000 34762 20012
rect 35342 20000 35348 20012
rect 35400 20000 35406 20052
rect 37182 20040 37188 20052
rect 35452 20012 37188 20040
rect 35452 19972 35480 20012
rect 37182 20000 37188 20012
rect 37240 20000 37246 20052
rect 37274 20000 37280 20052
rect 37332 20000 37338 20052
rect 38626 20012 42564 20040
rect 34624 19944 35480 19972
rect 35618 19932 35624 19984
rect 35676 19972 35682 19984
rect 38626 19972 38654 20012
rect 35676 19944 38654 19972
rect 35676 19932 35682 19944
rect 38746 19932 38752 19984
rect 38804 19972 38810 19984
rect 39485 19975 39543 19981
rect 39485 19972 39497 19975
rect 38804 19944 39497 19972
rect 38804 19932 38810 19944
rect 39485 19941 39497 19944
rect 39531 19941 39543 19975
rect 39485 19935 39543 19941
rect 40770 19932 40776 19984
rect 40828 19972 40834 19984
rect 41506 19972 41512 19984
rect 40828 19944 41512 19972
rect 40828 19932 40834 19944
rect 41506 19932 41512 19944
rect 41564 19932 41570 19984
rect 41966 19932 41972 19984
rect 42024 19972 42030 19984
rect 42337 19975 42395 19981
rect 42337 19972 42349 19975
rect 42024 19944 42349 19972
rect 42024 19932 42030 19944
rect 42337 19941 42349 19944
rect 42383 19941 42395 19975
rect 42536 19972 42564 20012
rect 42610 20000 42616 20052
rect 42668 20000 42674 20052
rect 43346 20000 43352 20052
rect 43404 20000 43410 20052
rect 46198 20000 46204 20052
rect 46256 20040 46262 20052
rect 47213 20043 47271 20049
rect 47213 20040 47225 20043
rect 46256 20012 47225 20040
rect 46256 20000 46262 20012
rect 47213 20009 47225 20012
rect 47259 20009 47271 20043
rect 47213 20003 47271 20009
rect 47486 20000 47492 20052
rect 47544 20000 47550 20052
rect 47765 20043 47823 20049
rect 47765 20009 47777 20043
rect 47811 20040 47823 20043
rect 48958 20040 48964 20052
rect 47811 20012 48964 20040
rect 47811 20009 47823 20012
rect 47765 20003 47823 20009
rect 48958 20000 48964 20012
rect 49016 20000 49022 20052
rect 43714 19972 43720 19984
rect 42536 19944 43720 19972
rect 42337 19935 42395 19941
rect 43714 19932 43720 19944
rect 43772 19932 43778 19984
rect 48409 19975 48467 19981
rect 48409 19941 48421 19975
rect 48455 19972 48467 19975
rect 48774 19972 48780 19984
rect 48455 19944 48780 19972
rect 48455 19941 48467 19944
rect 48409 19935 48467 19941
rect 48774 19932 48780 19944
rect 48832 19932 48838 19984
rect 32214 19864 32220 19916
rect 32272 19904 32278 19916
rect 32585 19907 32643 19913
rect 32585 19904 32597 19907
rect 32272 19876 32597 19904
rect 32272 19864 32278 19876
rect 32585 19873 32597 19876
rect 32631 19873 32643 19907
rect 32585 19867 32643 19873
rect 32677 19907 32735 19913
rect 32677 19873 32689 19907
rect 32723 19904 32735 19907
rect 32858 19904 32864 19916
rect 32723 19876 32864 19904
rect 32723 19873 32735 19876
rect 32677 19867 32735 19873
rect 32858 19864 32864 19876
rect 32916 19864 32922 19916
rect 32950 19864 32956 19916
rect 33008 19904 33014 19916
rect 33870 19904 33876 19916
rect 33008 19876 33876 19904
rect 33008 19864 33014 19876
rect 33870 19864 33876 19876
rect 33928 19864 33934 19916
rect 34054 19864 34060 19916
rect 34112 19864 34118 19916
rect 35529 19907 35587 19913
rect 35529 19873 35541 19907
rect 35575 19904 35587 19907
rect 36078 19904 36084 19916
rect 35575 19876 36084 19904
rect 35575 19873 35587 19876
rect 35529 19867 35587 19873
rect 36078 19864 36084 19876
rect 36136 19864 36142 19916
rect 36725 19907 36783 19913
rect 36725 19873 36737 19907
rect 36771 19904 36783 19907
rect 37366 19904 37372 19916
rect 36771 19876 37372 19904
rect 36771 19873 36783 19876
rect 36725 19867 36783 19873
rect 37366 19864 37372 19876
rect 37424 19864 37430 19916
rect 37458 19864 37464 19916
rect 37516 19904 37522 19916
rect 37829 19907 37887 19913
rect 37829 19904 37841 19907
rect 37516 19876 37841 19904
rect 37516 19864 37522 19876
rect 37829 19873 37841 19876
rect 37875 19873 37887 19907
rect 37829 19867 37887 19873
rect 37918 19864 37924 19916
rect 37976 19904 37982 19916
rect 38933 19907 38991 19913
rect 38933 19904 38945 19907
rect 37976 19876 38945 19904
rect 37976 19864 37982 19876
rect 38933 19873 38945 19876
rect 38979 19904 38991 19907
rect 39022 19904 39028 19916
rect 38979 19876 39028 19904
rect 38979 19873 38991 19876
rect 38933 19867 38991 19873
rect 39022 19864 39028 19876
rect 39080 19864 39086 19916
rect 39117 19907 39175 19913
rect 39117 19873 39129 19907
rect 39163 19904 39175 19907
rect 39574 19904 39580 19916
rect 39163 19876 39580 19904
rect 39163 19873 39175 19876
rect 39117 19867 39175 19873
rect 39574 19864 39580 19876
rect 39632 19864 39638 19916
rect 40126 19864 40132 19916
rect 40184 19904 40190 19916
rect 40589 19907 40647 19913
rect 40589 19904 40601 19907
rect 40184 19876 40601 19904
rect 40184 19864 40190 19876
rect 40589 19873 40601 19876
rect 40635 19873 40647 19907
rect 40589 19867 40647 19873
rect 42245 19907 42303 19913
rect 42245 19873 42257 19907
rect 42291 19904 42303 19907
rect 49329 19907 49387 19913
rect 49329 19904 49341 19907
rect 42291 19876 49341 19904
rect 42291 19873 42303 19876
rect 42245 19867 42303 19873
rect 49329 19873 49341 19876
rect 49375 19873 49387 19907
rect 49329 19867 49387 19873
rect 32490 19796 32496 19848
rect 32548 19796 32554 19848
rect 32766 19796 32772 19848
rect 32824 19836 32830 19848
rect 33781 19839 33839 19845
rect 33781 19836 33793 19839
rect 32824 19808 33793 19836
rect 32824 19796 32830 19808
rect 33781 19805 33793 19808
rect 33827 19836 33839 19839
rect 35894 19836 35900 19848
rect 33827 19808 33916 19836
rect 33827 19805 33839 19808
rect 33781 19799 33839 19805
rect 33888 19768 33916 19808
rect 34440 19808 35900 19836
rect 34440 19768 34468 19808
rect 35894 19796 35900 19808
rect 35952 19796 35958 19848
rect 38838 19796 38844 19848
rect 38896 19836 38902 19848
rect 38896 19808 40264 19836
rect 38896 19796 38902 19808
rect 31726 19740 33824 19768
rect 33888 19740 34468 19768
rect 34517 19771 34575 19777
rect 27985 19703 28043 19709
rect 27985 19669 27997 19703
rect 28031 19669 28043 19703
rect 27985 19663 28043 19669
rect 29089 19703 29147 19709
rect 29089 19669 29101 19703
rect 29135 19700 29147 19703
rect 29270 19700 29276 19712
rect 29135 19672 29276 19700
rect 29135 19669 29147 19672
rect 29089 19663 29147 19669
rect 29270 19660 29276 19672
rect 29328 19660 29334 19712
rect 29454 19660 29460 19712
rect 29512 19700 29518 19712
rect 30098 19700 30104 19712
rect 29512 19672 30104 19700
rect 29512 19660 29518 19672
rect 30098 19660 30104 19672
rect 30156 19660 30162 19712
rect 32122 19660 32128 19712
rect 32180 19660 32186 19712
rect 32398 19660 32404 19712
rect 32456 19700 32462 19712
rect 33042 19700 33048 19712
rect 32456 19672 33048 19700
rect 32456 19660 32462 19672
rect 33042 19660 33048 19672
rect 33100 19660 33106 19712
rect 33796 19700 33824 19740
rect 34517 19737 34529 19771
rect 34563 19768 34575 19771
rect 34698 19768 34704 19780
rect 34563 19740 34704 19768
rect 34563 19737 34575 19740
rect 34517 19731 34575 19737
rect 34532 19700 34560 19731
rect 34698 19728 34704 19740
rect 34756 19728 34762 19780
rect 36541 19771 36599 19777
rect 36541 19768 36553 19771
rect 34900 19740 36553 19768
rect 34900 19709 34928 19740
rect 36541 19737 36553 19740
rect 36587 19737 36599 19771
rect 36541 19731 36599 19737
rect 37274 19728 37280 19780
rect 37332 19768 37338 19780
rect 40236 19768 40264 19808
rect 40310 19796 40316 19848
rect 40368 19836 40374 19848
rect 40405 19839 40463 19845
rect 40405 19836 40417 19839
rect 40368 19808 40417 19836
rect 40368 19796 40374 19808
rect 40405 19805 40417 19808
rect 40451 19805 40463 19839
rect 40405 19799 40463 19805
rect 40494 19796 40500 19848
rect 40552 19796 40558 19848
rect 40604 19836 40632 19867
rect 41233 19839 41291 19845
rect 41233 19836 41245 19839
rect 40604 19808 41245 19836
rect 41233 19805 41245 19808
rect 41279 19805 41291 19839
rect 41233 19799 41291 19805
rect 42260 19768 42288 19867
rect 43165 19839 43223 19845
rect 43165 19805 43177 19839
rect 43211 19836 43223 19839
rect 43438 19836 43444 19848
rect 43211 19808 43444 19836
rect 43211 19805 43223 19808
rect 43165 19799 43223 19805
rect 43438 19796 43444 19808
rect 43496 19796 43502 19848
rect 48133 19839 48191 19845
rect 48133 19805 48145 19839
rect 48179 19836 48191 19839
rect 48593 19839 48651 19845
rect 48593 19836 48605 19839
rect 48179 19808 48605 19836
rect 48179 19805 48191 19808
rect 48133 19799 48191 19805
rect 48593 19805 48605 19808
rect 48639 19836 48651 19839
rect 48682 19836 48688 19848
rect 48639 19808 48688 19836
rect 48639 19805 48651 19808
rect 48593 19799 48651 19805
rect 48682 19796 48688 19808
rect 48740 19796 48746 19848
rect 37332 19740 40172 19768
rect 40236 19740 42288 19768
rect 37332 19728 37338 19740
rect 33796 19672 34560 19700
rect 34885 19703 34943 19709
rect 34885 19669 34897 19703
rect 34931 19669 34943 19703
rect 34885 19663 34943 19669
rect 35066 19660 35072 19712
rect 35124 19700 35130 19712
rect 35253 19703 35311 19709
rect 35253 19700 35265 19703
rect 35124 19672 35265 19700
rect 35124 19660 35130 19672
rect 35253 19669 35265 19672
rect 35299 19669 35311 19703
rect 35253 19663 35311 19669
rect 35342 19660 35348 19712
rect 35400 19700 35406 19712
rect 35802 19700 35808 19712
rect 35400 19672 35808 19700
rect 35400 19660 35406 19672
rect 35802 19660 35808 19672
rect 35860 19660 35866 19712
rect 35894 19660 35900 19712
rect 35952 19700 35958 19712
rect 36081 19703 36139 19709
rect 36081 19700 36093 19703
rect 35952 19672 36093 19700
rect 35952 19660 35958 19672
rect 36081 19669 36093 19672
rect 36127 19669 36139 19703
rect 36081 19663 36139 19669
rect 36446 19660 36452 19712
rect 36504 19660 36510 19712
rect 37642 19660 37648 19712
rect 37700 19660 37706 19712
rect 37737 19703 37795 19709
rect 37737 19669 37749 19703
rect 37783 19700 37795 19703
rect 38378 19700 38384 19712
rect 37783 19672 38384 19700
rect 37783 19669 37795 19672
rect 37737 19663 37795 19669
rect 38378 19660 38384 19672
rect 38436 19660 38442 19712
rect 38473 19703 38531 19709
rect 38473 19669 38485 19703
rect 38519 19700 38531 19703
rect 38562 19700 38568 19712
rect 38519 19672 38568 19700
rect 38519 19669 38531 19672
rect 38473 19663 38531 19669
rect 38562 19660 38568 19672
rect 38620 19660 38626 19712
rect 38654 19660 38660 19712
rect 38712 19700 38718 19712
rect 39850 19700 39856 19712
rect 38712 19672 39856 19700
rect 38712 19660 38718 19672
rect 39850 19660 39856 19672
rect 39908 19660 39914 19712
rect 40034 19660 40040 19712
rect 40092 19660 40098 19712
rect 40144 19700 40172 19740
rect 42334 19728 42340 19780
rect 42392 19768 42398 19780
rect 42797 19771 42855 19777
rect 42797 19768 42809 19771
rect 42392 19740 42809 19768
rect 42392 19728 42398 19740
rect 42797 19737 42809 19740
rect 42843 19768 42855 19771
rect 42981 19771 43039 19777
rect 42981 19768 42993 19771
rect 42843 19740 42993 19768
rect 42843 19737 42855 19740
rect 42797 19731 42855 19737
rect 42981 19737 42993 19740
rect 43027 19768 43039 19771
rect 44634 19768 44640 19780
rect 43027 19740 44640 19768
rect 43027 19737 43039 19740
rect 42981 19731 43039 19737
rect 44634 19728 44640 19740
rect 44692 19728 44698 19780
rect 47949 19771 48007 19777
rect 47949 19737 47961 19771
rect 47995 19768 48007 19771
rect 49145 19771 49203 19777
rect 49145 19768 49157 19771
rect 47995 19740 49157 19768
rect 47995 19737 48007 19740
rect 47949 19731 48007 19737
rect 49145 19737 49157 19740
rect 49191 19768 49203 19771
rect 49326 19768 49332 19780
rect 49191 19740 49332 19768
rect 49191 19737 49203 19740
rect 49145 19731 49203 19737
rect 49326 19728 49332 19740
rect 49384 19728 49390 19780
rect 40678 19700 40684 19712
rect 40144 19672 40684 19700
rect 40678 19660 40684 19672
rect 40736 19660 40742 19712
rect 40954 19660 40960 19712
rect 41012 19700 41018 19712
rect 41877 19703 41935 19709
rect 41877 19700 41889 19703
rect 41012 19672 41889 19700
rect 41012 19660 41018 19672
rect 41877 19669 41889 19672
rect 41923 19669 41935 19703
rect 41877 19663 41935 19669
rect 45278 19660 45284 19712
rect 45336 19700 45342 19712
rect 47029 19703 47087 19709
rect 47029 19700 47041 19703
rect 45336 19672 47041 19700
rect 45336 19660 45342 19672
rect 47029 19669 47041 19672
rect 47075 19669 47087 19703
rect 47029 19663 47087 19669
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 6270 19496 6276 19508
rect 2746 19468 6276 19496
rect 2746 19428 2774 19468
rect 6270 19456 6276 19468
rect 6328 19456 6334 19508
rect 7101 19499 7159 19505
rect 7101 19465 7113 19499
rect 7147 19496 7159 19499
rect 7926 19496 7932 19508
rect 7147 19468 7932 19496
rect 7147 19465 7159 19468
rect 7101 19459 7159 19465
rect 7926 19456 7932 19468
rect 7984 19456 7990 19508
rect 8573 19499 8631 19505
rect 8573 19465 8585 19499
rect 8619 19496 8631 19499
rect 8619 19468 9674 19496
rect 8619 19465 8631 19468
rect 8573 19459 8631 19465
rect 1780 19400 2774 19428
rect 1780 19369 1808 19400
rect 4614 19388 4620 19440
rect 4672 19388 4678 19440
rect 6086 19388 6092 19440
rect 6144 19428 6150 19440
rect 9646 19428 9674 19468
rect 9858 19456 9864 19508
rect 9916 19456 9922 19508
rect 9950 19456 9956 19508
rect 10008 19496 10014 19508
rect 12805 19499 12863 19505
rect 12805 19496 12817 19499
rect 10008 19468 12817 19496
rect 10008 19456 10014 19468
rect 12805 19465 12817 19468
rect 12851 19465 12863 19499
rect 12805 19459 12863 19465
rect 13354 19456 13360 19508
rect 13412 19496 13418 19508
rect 15197 19499 15255 19505
rect 15197 19496 15209 19499
rect 13412 19468 15209 19496
rect 13412 19456 13418 19468
rect 15197 19465 15209 19468
rect 15243 19465 15255 19499
rect 15197 19459 15255 19465
rect 16298 19456 16304 19508
rect 16356 19456 16362 19508
rect 16666 19456 16672 19508
rect 16724 19496 16730 19508
rect 16853 19499 16911 19505
rect 16853 19496 16865 19499
rect 16724 19468 16865 19496
rect 16724 19456 16730 19468
rect 16853 19465 16865 19468
rect 16899 19465 16911 19499
rect 16853 19459 16911 19465
rect 17313 19499 17371 19505
rect 17313 19465 17325 19499
rect 17359 19496 17371 19499
rect 20717 19499 20775 19505
rect 20717 19496 20729 19499
rect 17359 19468 20729 19496
rect 17359 19465 17371 19468
rect 17313 19459 17371 19465
rect 20717 19465 20729 19468
rect 20763 19465 20775 19499
rect 20717 19459 20775 19465
rect 21177 19499 21235 19505
rect 21177 19465 21189 19499
rect 21223 19496 21235 19499
rect 21266 19496 21272 19508
rect 21223 19468 21272 19496
rect 21223 19465 21235 19468
rect 21177 19459 21235 19465
rect 21266 19456 21272 19468
rect 21324 19456 21330 19508
rect 21726 19456 21732 19508
rect 21784 19496 21790 19508
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 21784 19468 22017 19496
rect 21784 19456 21790 19468
rect 22005 19465 22017 19468
rect 22051 19465 22063 19499
rect 22005 19459 22063 19465
rect 23566 19456 23572 19508
rect 23624 19496 23630 19508
rect 25869 19499 25927 19505
rect 25869 19496 25881 19499
rect 23624 19468 25881 19496
rect 23624 19456 23630 19468
rect 25869 19465 25881 19468
rect 25915 19465 25927 19499
rect 25869 19459 25927 19465
rect 26142 19456 26148 19508
rect 26200 19496 26206 19508
rect 26237 19499 26295 19505
rect 26237 19496 26249 19499
rect 26200 19468 26249 19496
rect 26200 19456 26206 19468
rect 26237 19465 26249 19468
rect 26283 19465 26295 19499
rect 26237 19459 26295 19465
rect 27617 19499 27675 19505
rect 27617 19465 27629 19499
rect 27663 19496 27675 19499
rect 28350 19496 28356 19508
rect 27663 19468 28356 19496
rect 27663 19465 27675 19468
rect 27617 19459 27675 19465
rect 28350 19456 28356 19468
rect 28408 19456 28414 19508
rect 28445 19499 28503 19505
rect 28445 19465 28457 19499
rect 28491 19496 28503 19499
rect 28718 19496 28724 19508
rect 28491 19468 28724 19496
rect 28491 19465 28503 19468
rect 28445 19459 28503 19465
rect 28718 19456 28724 19468
rect 28776 19456 28782 19508
rect 28813 19499 28871 19505
rect 28813 19465 28825 19499
rect 28859 19496 28871 19499
rect 32030 19496 32036 19508
rect 28859 19468 32036 19496
rect 28859 19465 28871 19468
rect 28813 19459 28871 19465
rect 32030 19456 32036 19468
rect 32088 19456 32094 19508
rect 32214 19456 32220 19508
rect 32272 19496 32278 19508
rect 32309 19499 32367 19505
rect 32309 19496 32321 19499
rect 32272 19468 32321 19496
rect 32272 19456 32278 19468
rect 32309 19465 32321 19468
rect 32355 19465 32367 19499
rect 32309 19459 32367 19465
rect 32677 19499 32735 19505
rect 32677 19465 32689 19499
rect 32723 19496 32735 19499
rect 32766 19496 32772 19508
rect 32723 19468 32772 19496
rect 32723 19465 32735 19468
rect 32677 19459 32735 19465
rect 32766 19456 32772 19468
rect 32824 19456 32830 19508
rect 33505 19499 33563 19505
rect 33505 19465 33517 19499
rect 33551 19496 33563 19499
rect 34606 19496 34612 19508
rect 33551 19468 34612 19496
rect 33551 19465 33563 19468
rect 33505 19459 33563 19465
rect 34606 19456 34612 19468
rect 34664 19456 34670 19508
rect 34698 19456 34704 19508
rect 34756 19456 34762 19508
rect 35158 19456 35164 19508
rect 35216 19456 35222 19508
rect 36446 19456 36452 19508
rect 36504 19496 36510 19508
rect 40129 19499 40187 19505
rect 40129 19496 40141 19499
rect 36504 19468 40141 19496
rect 36504 19456 36510 19468
rect 40129 19465 40141 19468
rect 40175 19465 40187 19499
rect 40129 19459 40187 19465
rect 40494 19456 40500 19508
rect 40552 19456 40558 19508
rect 40678 19456 40684 19508
rect 40736 19496 40742 19508
rect 40736 19468 41384 19496
rect 40736 19456 40742 19468
rect 10318 19428 10324 19440
rect 6144 19400 9260 19428
rect 9646 19400 10324 19428
rect 6144 19388 6150 19400
rect 1765 19363 1823 19369
rect 1765 19329 1777 19363
rect 1811 19329 1823 19363
rect 1765 19323 1823 19329
rect 2777 19363 2835 19369
rect 2777 19329 2789 19363
rect 2823 19360 2835 19363
rect 2866 19360 2872 19372
rect 2823 19332 2872 19360
rect 2823 19329 2835 19332
rect 2777 19323 2835 19329
rect 2866 19320 2872 19332
rect 2924 19320 2930 19372
rect 3605 19363 3663 19369
rect 3605 19329 3617 19363
rect 3651 19360 3663 19363
rect 5258 19360 5264 19372
rect 3651 19332 5264 19360
rect 3651 19329 3663 19332
rect 3605 19323 3663 19329
rect 5258 19320 5264 19332
rect 5316 19320 5322 19372
rect 5353 19363 5411 19369
rect 5353 19329 5365 19363
rect 5399 19329 5411 19363
rect 5353 19323 5411 19329
rect 5997 19363 6055 19369
rect 5997 19329 6009 19363
rect 6043 19360 6055 19363
rect 7285 19363 7343 19369
rect 6043 19332 6960 19360
rect 6043 19329 6055 19332
rect 5997 19323 6055 19329
rect 5368 19292 5396 19323
rect 5276 19264 5396 19292
rect 5276 19236 5304 19264
rect 6822 19252 6828 19304
rect 6880 19252 6886 19304
rect 5258 19184 5264 19236
rect 5316 19224 5322 19236
rect 6932 19224 6960 19332
rect 7285 19329 7297 19363
rect 7331 19360 7343 19363
rect 7742 19360 7748 19372
rect 7331 19332 7748 19360
rect 7331 19329 7343 19332
rect 7285 19323 7343 19329
rect 7742 19320 7748 19332
rect 7800 19320 7806 19372
rect 7837 19363 7895 19369
rect 7837 19329 7849 19363
rect 7883 19360 7895 19363
rect 7926 19360 7932 19372
rect 7883 19332 7932 19360
rect 7883 19329 7895 19332
rect 7837 19323 7895 19329
rect 7926 19320 7932 19332
rect 7984 19320 7990 19372
rect 8754 19320 8760 19372
rect 8812 19320 8818 19372
rect 7006 19252 7012 19304
rect 7064 19292 7070 19304
rect 8021 19295 8079 19301
rect 8021 19292 8033 19295
rect 7064 19264 8033 19292
rect 7064 19252 7070 19264
rect 8021 19261 8033 19264
rect 8067 19261 8079 19295
rect 8021 19255 8079 19261
rect 7834 19224 7840 19236
rect 5316 19196 6868 19224
rect 6932 19196 7840 19224
rect 5316 19184 5322 19196
rect 2314 19116 2320 19168
rect 2372 19156 2378 19168
rect 5445 19159 5503 19165
rect 5445 19156 5457 19159
rect 2372 19128 5457 19156
rect 2372 19116 2378 19128
rect 5445 19125 5457 19128
rect 5491 19125 5503 19159
rect 5445 19119 5503 19125
rect 6178 19116 6184 19168
rect 6236 19116 6242 19168
rect 6457 19159 6515 19165
rect 6457 19125 6469 19159
rect 6503 19156 6515 19159
rect 6546 19156 6552 19168
rect 6503 19128 6552 19156
rect 6503 19125 6515 19128
rect 6457 19119 6515 19125
rect 6546 19116 6552 19128
rect 6604 19116 6610 19168
rect 6638 19116 6644 19168
rect 6696 19116 6702 19168
rect 6840 19156 6868 19196
rect 7834 19184 7840 19196
rect 7892 19184 7898 19236
rect 7926 19184 7932 19236
rect 7984 19224 7990 19236
rect 8938 19224 8944 19236
rect 7984 19196 8944 19224
rect 7984 19184 7990 19196
rect 8938 19184 8944 19196
rect 8996 19184 9002 19236
rect 9232 19233 9260 19400
rect 10318 19388 10324 19400
rect 10376 19388 10382 19440
rect 11149 19431 11207 19437
rect 11149 19397 11161 19431
rect 11195 19428 11207 19431
rect 11330 19428 11336 19440
rect 11195 19400 11336 19428
rect 11195 19397 11207 19400
rect 11149 19391 11207 19397
rect 11330 19388 11336 19400
rect 11388 19388 11394 19440
rect 12066 19388 12072 19440
rect 12124 19428 12130 19440
rect 13725 19431 13783 19437
rect 13725 19428 13737 19431
rect 12124 19400 13737 19428
rect 12124 19388 12130 19400
rect 13725 19397 13737 19400
rect 13771 19397 13783 19431
rect 15562 19428 15568 19440
rect 13725 19391 13783 19397
rect 14476 19400 15568 19428
rect 9306 19320 9312 19372
rect 9364 19360 9370 19372
rect 9401 19363 9459 19369
rect 9401 19360 9413 19363
rect 9364 19332 9413 19360
rect 9364 19320 9370 19332
rect 9401 19329 9413 19332
rect 9447 19329 9459 19363
rect 9401 19323 9459 19329
rect 10045 19363 10103 19369
rect 10045 19329 10057 19363
rect 10091 19360 10103 19363
rect 10134 19360 10140 19372
rect 10091 19332 10140 19360
rect 10091 19329 10103 19332
rect 10045 19323 10103 19329
rect 10134 19320 10140 19332
rect 10192 19320 10198 19372
rect 10505 19363 10563 19369
rect 10505 19329 10517 19363
rect 10551 19360 10563 19363
rect 10551 19332 11468 19360
rect 10551 19329 10563 19332
rect 10505 19323 10563 19329
rect 9490 19252 9496 19304
rect 9548 19292 9554 19304
rect 11440 19292 11468 19332
rect 11790 19320 11796 19372
rect 11848 19320 11854 19372
rect 12897 19363 12955 19369
rect 12897 19329 12909 19363
rect 12943 19360 12955 19363
rect 14476 19360 14504 19400
rect 15562 19388 15568 19400
rect 15620 19388 15626 19440
rect 17862 19428 17868 19440
rect 15672 19400 17868 19428
rect 12943 19332 14504 19360
rect 12943 19329 12955 19332
rect 12897 19323 12955 19329
rect 14550 19320 14556 19372
rect 14608 19320 14614 19372
rect 15672 19369 15700 19400
rect 17862 19388 17868 19400
rect 17920 19388 17926 19440
rect 18598 19428 18604 19440
rect 18064 19400 18604 19428
rect 15657 19363 15715 19369
rect 15657 19329 15669 19363
rect 15703 19329 15715 19363
rect 15657 19323 15715 19329
rect 17218 19320 17224 19372
rect 17276 19320 17282 19372
rect 17770 19320 17776 19372
rect 17828 19360 17834 19372
rect 18064 19369 18092 19400
rect 18598 19388 18604 19400
rect 18656 19388 18662 19440
rect 20073 19431 20131 19437
rect 20073 19397 20085 19431
rect 20119 19428 20131 19431
rect 20530 19428 20536 19440
rect 20119 19400 20536 19428
rect 20119 19397 20131 19400
rect 20073 19391 20131 19397
rect 20530 19388 20536 19400
rect 20588 19388 20594 19440
rect 21085 19431 21143 19437
rect 21085 19397 21097 19431
rect 21131 19428 21143 19431
rect 24026 19428 24032 19440
rect 21131 19400 24032 19428
rect 21131 19397 21143 19400
rect 21085 19391 21143 19397
rect 24026 19388 24032 19400
rect 24084 19388 24090 19440
rect 24394 19388 24400 19440
rect 24452 19388 24458 19440
rect 25774 19388 25780 19440
rect 25832 19428 25838 19440
rect 29270 19428 29276 19440
rect 25832 19400 29276 19428
rect 25832 19388 25838 19400
rect 29270 19388 29276 19400
rect 29328 19388 29334 19440
rect 30745 19431 30803 19437
rect 29380 19400 30420 19428
rect 18049 19363 18107 19369
rect 18049 19360 18061 19363
rect 17828 19332 18061 19360
rect 17828 19320 17834 19332
rect 18049 19329 18061 19332
rect 18095 19329 18107 19363
rect 18049 19323 18107 19329
rect 19426 19320 19432 19372
rect 19484 19360 19490 19372
rect 19484 19332 20116 19360
rect 19484 19320 19490 19332
rect 20088 19304 20116 19332
rect 20714 19320 20720 19372
rect 20772 19360 20778 19372
rect 21818 19360 21824 19372
rect 20772 19332 21824 19360
rect 20772 19320 20778 19332
rect 21818 19320 21824 19332
rect 21876 19320 21882 19372
rect 22094 19320 22100 19372
rect 22152 19360 22158 19372
rect 22373 19363 22431 19369
rect 22373 19360 22385 19363
rect 22152 19332 22385 19360
rect 22152 19320 22158 19332
rect 22373 19329 22385 19332
rect 22419 19329 22431 19363
rect 22373 19323 22431 19329
rect 22462 19320 22468 19372
rect 22520 19320 22526 19372
rect 23382 19320 23388 19372
rect 23440 19360 23446 19372
rect 23477 19363 23535 19369
rect 23477 19360 23489 19363
rect 23440 19332 23489 19360
rect 23440 19320 23446 19332
rect 23477 19329 23489 19332
rect 23523 19329 23535 19363
rect 25958 19360 25964 19372
rect 23477 19323 23535 19329
rect 25424 19332 25964 19360
rect 13081 19295 13139 19301
rect 13081 19292 13093 19295
rect 9548 19264 11284 19292
rect 11440 19264 13093 19292
rect 9548 19252 9554 19264
rect 9217 19227 9275 19233
rect 9217 19193 9229 19227
rect 9263 19193 9275 19227
rect 11146 19224 11152 19236
rect 9217 19187 9275 19193
rect 10428 19196 11152 19224
rect 10428 19156 10456 19196
rect 11146 19184 11152 19196
rect 11204 19184 11210 19236
rect 11256 19224 11284 19264
rect 13081 19261 13093 19264
rect 13127 19292 13139 19295
rect 13446 19292 13452 19304
rect 13127 19264 13452 19292
rect 13127 19261 13139 19264
rect 13081 19255 13139 19261
rect 13446 19252 13452 19264
rect 13504 19252 13510 19304
rect 13909 19295 13967 19301
rect 13909 19261 13921 19295
rect 13955 19292 13967 19295
rect 13998 19292 14004 19304
rect 13955 19264 14004 19292
rect 13955 19261 13967 19264
rect 13909 19255 13967 19261
rect 13998 19252 14004 19264
rect 14056 19252 14062 19304
rect 16022 19252 16028 19304
rect 16080 19292 16086 19304
rect 16080 19264 16620 19292
rect 16080 19252 16086 19264
rect 11977 19227 12035 19233
rect 11977 19224 11989 19227
rect 11256 19196 11989 19224
rect 11977 19193 11989 19196
rect 12023 19193 12035 19227
rect 16592 19224 16620 19264
rect 16942 19252 16948 19304
rect 17000 19292 17006 19304
rect 17405 19295 17463 19301
rect 17405 19292 17417 19295
rect 17000 19264 17417 19292
rect 17000 19252 17006 19264
rect 17405 19261 17417 19264
rect 17451 19261 17463 19295
rect 17405 19255 17463 19261
rect 17586 19252 17592 19304
rect 17644 19292 17650 19304
rect 18325 19295 18383 19301
rect 18325 19292 18337 19295
rect 17644 19264 18337 19292
rect 17644 19252 17650 19264
rect 18325 19261 18337 19264
rect 18371 19261 18383 19295
rect 18325 19255 18383 19261
rect 20070 19252 20076 19304
rect 20128 19292 20134 19304
rect 20349 19295 20407 19301
rect 20349 19292 20361 19295
rect 20128 19264 20361 19292
rect 20128 19252 20134 19264
rect 20349 19261 20361 19264
rect 20395 19261 20407 19295
rect 20349 19255 20407 19261
rect 20990 19252 20996 19304
rect 21048 19292 21054 19304
rect 21269 19295 21327 19301
rect 21269 19292 21281 19295
rect 21048 19264 21281 19292
rect 21048 19252 21054 19264
rect 21269 19261 21281 19264
rect 21315 19292 21327 19295
rect 22002 19292 22008 19304
rect 21315 19264 22008 19292
rect 21315 19261 21327 19264
rect 21269 19255 21327 19261
rect 22002 19252 22008 19264
rect 22060 19252 22066 19304
rect 22646 19252 22652 19304
rect 22704 19252 22710 19304
rect 23753 19295 23811 19301
rect 23753 19261 23765 19295
rect 23799 19292 23811 19295
rect 25314 19292 25320 19304
rect 23799 19264 25320 19292
rect 23799 19261 23811 19264
rect 23753 19255 23811 19261
rect 25314 19252 25320 19264
rect 25372 19252 25378 19304
rect 16592 19196 17816 19224
rect 11977 19187 12035 19193
rect 6840 19128 10456 19156
rect 10502 19116 10508 19168
rect 10560 19156 10566 19168
rect 11790 19156 11796 19168
rect 10560 19128 11796 19156
rect 10560 19116 10566 19128
rect 11790 19116 11796 19128
rect 11848 19116 11854 19168
rect 12434 19116 12440 19168
rect 12492 19116 12498 19168
rect 14277 19159 14335 19165
rect 14277 19125 14289 19159
rect 14323 19156 14335 19159
rect 14366 19156 14372 19168
rect 14323 19128 14372 19156
rect 14323 19125 14335 19128
rect 14277 19119 14335 19125
rect 14366 19116 14372 19128
rect 14424 19116 14430 19168
rect 14918 19116 14924 19168
rect 14976 19156 14982 19168
rect 17678 19156 17684 19168
rect 14976 19128 17684 19156
rect 14976 19116 14982 19128
rect 17678 19116 17684 19128
rect 17736 19116 17742 19168
rect 17788 19156 17816 19196
rect 22370 19184 22376 19236
rect 22428 19224 22434 19236
rect 25225 19227 25283 19233
rect 22428 19196 23612 19224
rect 22428 19184 22434 19196
rect 23201 19159 23259 19165
rect 23201 19156 23213 19159
rect 17788 19128 23213 19156
rect 23201 19125 23213 19128
rect 23247 19156 23259 19159
rect 23474 19156 23480 19168
rect 23247 19128 23480 19156
rect 23247 19125 23259 19128
rect 23201 19119 23259 19125
rect 23474 19116 23480 19128
rect 23532 19116 23538 19168
rect 23584 19156 23612 19196
rect 25225 19193 25237 19227
rect 25271 19224 25283 19227
rect 25424 19224 25452 19332
rect 25958 19320 25964 19332
rect 26016 19320 26022 19372
rect 26694 19360 26700 19372
rect 26436 19332 26700 19360
rect 25682 19252 25688 19304
rect 25740 19292 25746 19304
rect 26329 19295 26387 19301
rect 25740 19264 26004 19292
rect 25740 19252 25746 19264
rect 25271 19196 25452 19224
rect 25271 19193 25283 19196
rect 25225 19187 25283 19193
rect 25498 19184 25504 19236
rect 25556 19224 25562 19236
rect 25866 19224 25872 19236
rect 25556 19196 25872 19224
rect 25556 19184 25562 19196
rect 25866 19184 25872 19196
rect 25924 19184 25930 19236
rect 25976 19224 26004 19264
rect 26329 19261 26341 19295
rect 26375 19292 26387 19295
rect 26436 19292 26464 19332
rect 26694 19320 26700 19332
rect 26752 19320 26758 19372
rect 28626 19360 28632 19372
rect 27540 19332 28632 19360
rect 26375 19264 26464 19292
rect 26513 19295 26571 19301
rect 26375 19261 26387 19264
rect 26329 19255 26387 19261
rect 26513 19261 26525 19295
rect 26559 19292 26571 19295
rect 27540 19292 27568 19332
rect 28626 19320 28632 19332
rect 28684 19320 28690 19372
rect 28718 19320 28724 19372
rect 28776 19360 28782 19372
rect 29380 19360 29408 19400
rect 28776 19332 29408 19360
rect 28776 19320 28782 19332
rect 26559 19264 27568 19292
rect 26559 19261 26571 19264
rect 26513 19255 26571 19261
rect 26528 19224 26556 19255
rect 27614 19252 27620 19304
rect 27672 19292 27678 19304
rect 27709 19295 27767 19301
rect 27709 19292 27721 19295
rect 27672 19264 27721 19292
rect 27672 19252 27678 19264
rect 27709 19261 27721 19264
rect 27755 19261 27767 19295
rect 27709 19255 27767 19261
rect 27801 19295 27859 19301
rect 27801 19261 27813 19295
rect 27847 19261 27859 19295
rect 27801 19255 27859 19261
rect 25976 19196 26556 19224
rect 27154 19156 27160 19168
rect 23584 19128 27160 19156
rect 27154 19116 27160 19128
rect 27212 19116 27218 19168
rect 27246 19116 27252 19168
rect 27304 19116 27310 19168
rect 27632 19156 27660 19252
rect 27816 19224 27844 19255
rect 27890 19252 27896 19304
rect 27948 19292 27954 19304
rect 28920 19301 28948 19332
rect 29638 19320 29644 19372
rect 29696 19320 29702 19372
rect 30282 19320 30288 19372
rect 30340 19320 30346 19372
rect 30392 19360 30420 19400
rect 30745 19397 30757 19431
rect 30791 19428 30803 19431
rect 30834 19428 30840 19440
rect 30791 19400 30840 19428
rect 30791 19397 30803 19400
rect 30745 19391 30803 19397
rect 30834 19388 30840 19400
rect 30892 19388 30898 19440
rect 31573 19431 31631 19437
rect 31573 19397 31585 19431
rect 31619 19428 31631 19431
rect 35618 19428 35624 19440
rect 31619 19400 35624 19428
rect 31619 19397 31631 19400
rect 31573 19391 31631 19397
rect 32324 19372 32352 19400
rect 35618 19388 35624 19400
rect 35676 19388 35682 19440
rect 36357 19431 36415 19437
rect 36357 19397 36369 19431
rect 36403 19428 36415 19431
rect 38470 19428 38476 19440
rect 36403 19400 38476 19428
rect 36403 19397 36415 19400
rect 36357 19391 36415 19397
rect 38470 19388 38476 19400
rect 38528 19388 38534 19440
rect 38746 19388 38752 19440
rect 38804 19388 38810 19440
rect 39850 19388 39856 19440
rect 39908 19428 39914 19440
rect 40589 19431 40647 19437
rect 40589 19428 40601 19431
rect 39908 19400 40601 19428
rect 39908 19388 39914 19400
rect 40589 19397 40601 19400
rect 40635 19397 40647 19431
rect 40589 19391 40647 19397
rect 30926 19360 30932 19372
rect 30392 19332 30932 19360
rect 30926 19320 30932 19332
rect 30984 19320 30990 19372
rect 31202 19320 31208 19372
rect 31260 19360 31266 19372
rect 31754 19360 31760 19372
rect 31260 19332 31760 19360
rect 31260 19320 31266 19332
rect 31754 19320 31760 19332
rect 31812 19320 31818 19372
rect 31846 19320 31852 19372
rect 31904 19360 31910 19372
rect 32214 19360 32220 19372
rect 31904 19332 32220 19360
rect 31904 19320 31910 19332
rect 32214 19320 32220 19332
rect 32272 19320 32278 19372
rect 32306 19320 32312 19372
rect 32364 19320 32370 19372
rect 32769 19363 32827 19369
rect 32769 19329 32781 19363
rect 32815 19360 32827 19363
rect 32950 19360 32956 19372
rect 32815 19332 32956 19360
rect 32815 19329 32827 19332
rect 32769 19323 32827 19329
rect 32950 19320 32956 19332
rect 33008 19320 33014 19372
rect 33042 19320 33048 19372
rect 33100 19360 33106 19372
rect 33100 19332 33824 19360
rect 33100 19320 33106 19332
rect 28905 19295 28963 19301
rect 27948 19264 28856 19292
rect 27948 19252 27954 19264
rect 28074 19224 28080 19236
rect 27816 19196 28080 19224
rect 28074 19184 28080 19196
rect 28132 19184 28138 19236
rect 28828 19224 28856 19264
rect 28905 19261 28917 19295
rect 28951 19261 28963 19295
rect 28905 19255 28963 19261
rect 28997 19295 29055 19301
rect 28997 19261 29009 19295
rect 29043 19261 29055 19295
rect 29656 19292 29684 19320
rect 32861 19295 32919 19301
rect 29656 19264 32352 19292
rect 28997 19255 29055 19261
rect 29012 19224 29040 19255
rect 28828 19196 29040 19224
rect 31570 19184 31576 19236
rect 31628 19224 31634 19236
rect 32324 19224 32352 19264
rect 32861 19261 32873 19295
rect 32907 19261 32919 19295
rect 32861 19255 32919 19261
rect 32876 19224 32904 19255
rect 33226 19252 33232 19304
rect 33284 19292 33290 19304
rect 33502 19292 33508 19304
rect 33284 19264 33508 19292
rect 33284 19252 33290 19264
rect 33502 19252 33508 19264
rect 33560 19252 33566 19304
rect 33796 19292 33824 19332
rect 33870 19320 33876 19372
rect 33928 19320 33934 19372
rect 33962 19320 33968 19372
rect 34020 19320 34026 19372
rect 34514 19320 34520 19372
rect 34572 19360 34578 19372
rect 35069 19363 35127 19369
rect 35069 19360 35081 19363
rect 34572 19332 35081 19360
rect 34572 19320 34578 19332
rect 35069 19329 35081 19332
rect 35115 19329 35127 19363
rect 35069 19323 35127 19329
rect 35158 19320 35164 19372
rect 35216 19360 35222 19372
rect 35710 19360 35716 19372
rect 35216 19332 35716 19360
rect 35216 19320 35222 19332
rect 35710 19320 35716 19332
rect 35768 19320 35774 19372
rect 35986 19320 35992 19372
rect 36044 19360 36050 19372
rect 36265 19363 36323 19369
rect 36265 19360 36277 19363
rect 36044 19332 36277 19360
rect 36044 19320 36050 19332
rect 36265 19329 36277 19332
rect 36311 19329 36323 19363
rect 36265 19323 36323 19329
rect 36464 19332 37136 19360
rect 33980 19292 34008 19320
rect 33796 19264 34008 19292
rect 34146 19252 34152 19304
rect 34204 19252 34210 19304
rect 34256 19264 34652 19292
rect 31628 19196 32168 19224
rect 32324 19196 32904 19224
rect 31628 19184 31634 19196
rect 32030 19156 32036 19168
rect 27632 19128 32036 19156
rect 32030 19116 32036 19128
rect 32088 19116 32094 19168
rect 32140 19156 32168 19196
rect 32950 19184 32956 19236
rect 33008 19224 33014 19236
rect 33962 19224 33968 19236
rect 33008 19196 33968 19224
rect 33008 19184 33014 19196
rect 33962 19184 33968 19196
rect 34020 19184 34026 19236
rect 34256 19156 34284 19264
rect 32140 19128 34284 19156
rect 34624 19156 34652 19264
rect 34974 19252 34980 19304
rect 35032 19292 35038 19304
rect 35253 19295 35311 19301
rect 35253 19292 35265 19295
rect 35032 19264 35265 19292
rect 35032 19252 35038 19264
rect 35253 19261 35265 19264
rect 35299 19261 35311 19295
rect 35253 19255 35311 19261
rect 35802 19252 35808 19304
rect 35860 19292 35866 19304
rect 36464 19292 36492 19332
rect 35860 19264 36492 19292
rect 36541 19295 36599 19301
rect 35860 19252 35866 19264
rect 36541 19261 36553 19295
rect 36587 19292 36599 19295
rect 36998 19292 37004 19304
rect 36587 19264 37004 19292
rect 36587 19261 36599 19264
rect 36541 19255 36599 19261
rect 36998 19252 37004 19264
rect 37056 19252 37062 19304
rect 37108 19292 37136 19332
rect 37182 19320 37188 19372
rect 37240 19360 37246 19372
rect 37240 19332 37504 19360
rect 37240 19320 37246 19332
rect 37476 19301 37504 19332
rect 37734 19320 37740 19372
rect 37792 19360 37798 19372
rect 37921 19363 37979 19369
rect 37921 19360 37933 19363
rect 37792 19332 37933 19360
rect 37792 19320 37798 19332
rect 37921 19329 37933 19332
rect 37967 19329 37979 19363
rect 40604 19360 40632 19391
rect 41356 19369 41384 19468
rect 42150 19456 42156 19508
rect 42208 19496 42214 19508
rect 42702 19496 42708 19508
rect 42208 19468 42708 19496
rect 42208 19456 42214 19468
rect 42702 19456 42708 19468
rect 42760 19456 42766 19508
rect 48866 19496 48872 19508
rect 42812 19468 48872 19496
rect 41325 19363 41384 19369
rect 40604 19332 41276 19360
rect 37921 19323 37979 19329
rect 37277 19295 37335 19301
rect 37277 19292 37289 19295
rect 37108 19264 37289 19292
rect 37277 19261 37289 19264
rect 37323 19261 37335 19295
rect 37277 19255 37335 19261
rect 37461 19295 37519 19301
rect 37461 19261 37473 19295
rect 37507 19292 37519 19295
rect 37826 19292 37832 19304
rect 37507 19264 37832 19292
rect 37507 19261 37519 19264
rect 37461 19255 37519 19261
rect 37826 19252 37832 19264
rect 37884 19252 37890 19304
rect 38197 19295 38255 19301
rect 38197 19261 38209 19295
rect 38243 19292 38255 19295
rect 40678 19292 40684 19304
rect 38243 19264 40684 19292
rect 38243 19261 38255 19264
rect 38197 19255 38255 19261
rect 40678 19252 40684 19264
rect 40736 19252 40742 19304
rect 40773 19295 40831 19301
rect 40773 19261 40785 19295
rect 40819 19261 40831 19295
rect 40773 19255 40831 19261
rect 35897 19227 35955 19233
rect 35897 19193 35909 19227
rect 35943 19224 35955 19227
rect 37182 19224 37188 19236
rect 35943 19196 37188 19224
rect 35943 19193 35955 19196
rect 35897 19187 35955 19193
rect 37182 19184 37188 19196
rect 37240 19184 37246 19236
rect 39758 19184 39764 19236
rect 39816 19224 39822 19236
rect 40788 19224 40816 19255
rect 39816 19196 40816 19224
rect 41248 19224 41276 19332
rect 41325 19329 41337 19363
rect 41371 19332 41384 19363
rect 41371 19329 41383 19332
rect 41325 19323 41383 19329
rect 41966 19320 41972 19372
rect 42024 19320 42030 19372
rect 42812 19233 42840 19468
rect 48866 19456 48872 19468
rect 48924 19456 48930 19508
rect 48593 19363 48651 19369
rect 48593 19329 48605 19363
rect 48639 19360 48651 19363
rect 49142 19360 49148 19372
rect 48639 19332 49148 19360
rect 48639 19329 48651 19332
rect 48593 19323 48651 19329
rect 49142 19320 49148 19332
rect 49200 19320 49206 19372
rect 47762 19252 47768 19304
rect 47820 19292 47826 19304
rect 48133 19295 48191 19301
rect 48133 19292 48145 19295
rect 47820 19264 48145 19292
rect 47820 19252 47826 19264
rect 48133 19261 48145 19264
rect 48179 19261 48191 19295
rect 48133 19255 48191 19261
rect 48406 19252 48412 19304
rect 48464 19252 48470 19304
rect 42797 19227 42855 19233
rect 42797 19224 42809 19227
rect 41248 19196 42809 19224
rect 39816 19184 39822 19196
rect 42797 19193 42809 19196
rect 42843 19193 42855 19227
rect 42797 19187 42855 19193
rect 47210 19184 47216 19236
rect 47268 19224 47274 19236
rect 47949 19227 48007 19233
rect 47949 19224 47961 19227
rect 47268 19196 47961 19224
rect 47268 19184 47274 19196
rect 47949 19193 47961 19196
rect 47995 19193 48007 19227
rect 47949 19187 48007 19193
rect 36630 19156 36636 19168
rect 34624 19128 36636 19156
rect 36630 19116 36636 19128
rect 36688 19116 36694 19168
rect 36906 19116 36912 19168
rect 36964 19116 36970 19168
rect 38746 19116 38752 19168
rect 38804 19156 38810 19168
rect 39666 19156 39672 19168
rect 38804 19128 39672 19156
rect 38804 19116 38810 19128
rect 39666 19116 39672 19128
rect 39724 19116 39730 19168
rect 42426 19116 42432 19168
rect 42484 19116 42490 19168
rect 47857 19159 47915 19165
rect 47857 19125 47869 19159
rect 47903 19156 47915 19159
rect 48498 19156 48504 19168
rect 47903 19128 48504 19156
rect 47903 19125 47915 19128
rect 47857 19119 47915 19125
rect 48498 19116 48504 19128
rect 48556 19116 48562 19168
rect 48777 19159 48835 19165
rect 48777 19125 48789 19159
rect 48823 19156 48835 19159
rect 49050 19156 49056 19168
rect 48823 19128 49056 19156
rect 48823 19125 48835 19128
rect 48777 19119 48835 19125
rect 49050 19116 49056 19128
rect 49108 19116 49114 19168
rect 49234 19116 49240 19168
rect 49292 19116 49298 19168
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 5994 18912 6000 18964
rect 6052 18952 6058 18964
rect 6181 18955 6239 18961
rect 6181 18952 6193 18955
rect 6052 18924 6193 18952
rect 6052 18912 6058 18924
rect 6181 18921 6193 18924
rect 6227 18921 6239 18955
rect 6181 18915 6239 18921
rect 7190 18912 7196 18964
rect 7248 18952 7254 18964
rect 12434 18952 12440 18964
rect 7248 18924 12440 18952
rect 7248 18912 7254 18924
rect 12434 18912 12440 18924
rect 12492 18912 12498 18964
rect 12526 18912 12532 18964
rect 12584 18952 12590 18964
rect 12713 18955 12771 18961
rect 12713 18952 12725 18955
rect 12584 18924 12725 18952
rect 12584 18912 12590 18924
rect 12713 18921 12725 18924
rect 12759 18921 12771 18955
rect 12713 18915 12771 18921
rect 14550 18912 14556 18964
rect 14608 18952 14614 18964
rect 16025 18955 16083 18961
rect 16025 18952 16037 18955
rect 14608 18924 16037 18952
rect 14608 18912 14614 18924
rect 16025 18921 16037 18924
rect 16071 18952 16083 18955
rect 16114 18952 16120 18964
rect 16071 18924 16120 18952
rect 16071 18921 16083 18924
rect 16025 18915 16083 18921
rect 16114 18912 16120 18924
rect 16172 18912 16178 18964
rect 16298 18912 16304 18964
rect 16356 18952 16362 18964
rect 16485 18955 16543 18961
rect 16485 18952 16497 18955
rect 16356 18924 16497 18952
rect 16356 18912 16362 18924
rect 16485 18921 16497 18924
rect 16531 18921 16543 18955
rect 16485 18915 16543 18921
rect 17310 18912 17316 18964
rect 17368 18952 17374 18964
rect 19797 18955 19855 18961
rect 19797 18952 19809 18955
rect 17368 18924 19809 18952
rect 17368 18912 17374 18924
rect 19797 18921 19809 18924
rect 19843 18921 19855 18955
rect 19797 18915 19855 18921
rect 19978 18912 19984 18964
rect 20036 18952 20042 18964
rect 22370 18952 22376 18964
rect 20036 18924 22376 18952
rect 20036 18912 20042 18924
rect 22370 18912 22376 18924
rect 22428 18912 22434 18964
rect 22544 18955 22602 18961
rect 22544 18921 22556 18955
rect 22590 18952 22602 18955
rect 22590 18924 23888 18952
rect 22590 18921 22602 18924
rect 22544 18915 22602 18921
rect 6638 18884 6644 18896
rect 2746 18856 6644 18884
rect 2746 18816 2774 18856
rect 6638 18844 6644 18856
rect 6696 18844 6702 18896
rect 7742 18844 7748 18896
rect 7800 18884 7806 18896
rect 9861 18887 9919 18893
rect 9861 18884 9873 18887
rect 7800 18856 9873 18884
rect 7800 18844 7806 18856
rect 9861 18853 9873 18856
rect 9907 18884 9919 18887
rect 10318 18884 10324 18896
rect 9907 18856 10324 18884
rect 9907 18853 9919 18856
rect 9861 18847 9919 18853
rect 10318 18844 10324 18856
rect 10376 18844 10382 18896
rect 11790 18844 11796 18896
rect 11848 18884 11854 18896
rect 12253 18887 12311 18893
rect 12253 18884 12265 18887
rect 11848 18856 12265 18884
rect 11848 18844 11854 18856
rect 12253 18853 12265 18856
rect 12299 18853 12311 18887
rect 12253 18847 12311 18853
rect 12621 18887 12679 18893
rect 12621 18853 12633 18887
rect 12667 18884 12679 18887
rect 13538 18884 13544 18896
rect 12667 18856 13544 18884
rect 12667 18853 12679 18856
rect 12621 18847 12679 18853
rect 13538 18844 13544 18856
rect 13596 18844 13602 18896
rect 16390 18844 16396 18896
rect 16448 18884 16454 18896
rect 16448 18856 17172 18884
rect 16448 18844 16454 18856
rect 1780 18788 2774 18816
rect 1780 18757 1808 18788
rect 3510 18776 3516 18828
rect 3568 18816 3574 18828
rect 4433 18819 4491 18825
rect 4433 18816 4445 18819
rect 3568 18788 4445 18816
rect 3568 18776 3574 18788
rect 4433 18785 4445 18788
rect 4479 18785 4491 18819
rect 4433 18779 4491 18785
rect 6178 18776 6184 18828
rect 6236 18816 6242 18828
rect 9030 18816 9036 18828
rect 6236 18788 9036 18816
rect 6236 18776 6242 18788
rect 9030 18776 9036 18788
rect 9088 18776 9094 18828
rect 9125 18819 9183 18825
rect 9125 18785 9137 18819
rect 9171 18816 9183 18819
rect 9217 18819 9275 18825
rect 9217 18816 9229 18819
rect 9171 18788 9229 18816
rect 9171 18785 9183 18788
rect 9125 18779 9183 18785
rect 9217 18785 9229 18788
rect 9263 18816 9275 18819
rect 9674 18816 9680 18828
rect 9263 18788 9680 18816
rect 9263 18785 9275 18788
rect 9217 18779 9275 18785
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 10505 18819 10563 18825
rect 10505 18785 10517 18819
rect 10551 18816 10563 18819
rect 13814 18816 13820 18828
rect 10551 18788 13820 18816
rect 10551 18785 10563 18788
rect 10505 18779 10563 18785
rect 13814 18776 13820 18788
rect 13872 18776 13878 18828
rect 15286 18816 15292 18828
rect 14292 18788 15292 18816
rect 14292 18760 14320 18788
rect 15286 18776 15292 18788
rect 15344 18776 15350 18828
rect 17034 18776 17040 18828
rect 17092 18776 17098 18828
rect 17144 18816 17172 18856
rect 17678 18844 17684 18896
rect 17736 18844 17742 18896
rect 18877 18887 18935 18893
rect 18877 18853 18889 18887
rect 18923 18884 18935 18887
rect 19886 18884 19892 18896
rect 18923 18856 19892 18884
rect 18923 18853 18935 18856
rect 18877 18847 18935 18853
rect 19886 18844 19892 18856
rect 19944 18844 19950 18896
rect 23860 18884 23888 18924
rect 24026 18912 24032 18964
rect 24084 18952 24090 18964
rect 24581 18955 24639 18961
rect 24581 18952 24593 18955
rect 24084 18924 24593 18952
rect 24084 18912 24090 18924
rect 24581 18921 24593 18924
rect 24627 18921 24639 18955
rect 24581 18915 24639 18921
rect 25130 18912 25136 18964
rect 25188 18912 25194 18964
rect 26510 18952 26516 18964
rect 25240 18924 26516 18952
rect 25148 18884 25176 18912
rect 23860 18856 25176 18884
rect 18233 18819 18291 18825
rect 18233 18816 18245 18819
rect 17144 18788 18245 18816
rect 18233 18785 18245 18788
rect 18279 18785 18291 18819
rect 20441 18819 20499 18825
rect 18233 18779 18291 18785
rect 19076 18788 20300 18816
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18717 1823 18751
rect 1765 18711 1823 18717
rect 4065 18751 4123 18757
rect 4065 18717 4077 18751
rect 4111 18748 4123 18751
rect 4246 18748 4252 18760
rect 4111 18720 4252 18748
rect 4111 18717 4123 18720
rect 4065 18711 4123 18717
rect 4246 18708 4252 18720
rect 4304 18708 4310 18760
rect 6365 18751 6423 18757
rect 6365 18717 6377 18751
rect 6411 18717 6423 18751
rect 6365 18711 6423 18717
rect 7009 18751 7067 18757
rect 7009 18717 7021 18751
rect 7055 18748 7067 18751
rect 7374 18748 7380 18760
rect 7055 18720 7380 18748
rect 7055 18717 7067 18720
rect 7009 18711 7067 18717
rect 2774 18640 2780 18692
rect 2832 18640 2838 18692
rect 6380 18680 6408 18711
rect 7374 18708 7380 18720
rect 7432 18708 7438 18760
rect 7469 18751 7527 18757
rect 7469 18717 7481 18751
rect 7515 18748 7527 18751
rect 7515 18720 9996 18748
rect 7515 18717 7527 18720
rect 7469 18711 7527 18717
rect 8205 18683 8263 18689
rect 6380 18652 8156 18680
rect 5258 18572 5264 18624
rect 5316 18612 5322 18624
rect 5629 18615 5687 18621
rect 5629 18612 5641 18615
rect 5316 18584 5641 18612
rect 5316 18572 5322 18584
rect 5629 18581 5641 18584
rect 5675 18581 5687 18615
rect 5629 18575 5687 18581
rect 6546 18572 6552 18624
rect 6604 18612 6610 18624
rect 6825 18615 6883 18621
rect 6825 18612 6837 18615
rect 6604 18584 6837 18612
rect 6604 18572 6610 18584
rect 6825 18581 6837 18584
rect 6871 18581 6883 18615
rect 8128 18612 8156 18652
rect 8205 18649 8217 18683
rect 8251 18680 8263 18683
rect 8294 18680 8300 18692
rect 8251 18652 8300 18680
rect 8251 18649 8263 18652
rect 8205 18643 8263 18649
rect 8294 18640 8300 18652
rect 8352 18640 8358 18692
rect 8389 18683 8447 18689
rect 8389 18649 8401 18683
rect 8435 18680 8447 18683
rect 8478 18680 8484 18692
rect 8435 18652 8484 18680
rect 8435 18649 8447 18652
rect 8389 18643 8447 18649
rect 8478 18640 8484 18652
rect 8536 18640 8542 18692
rect 9490 18680 9496 18692
rect 8588 18652 9496 18680
rect 8588 18612 8616 18652
rect 9490 18640 9496 18652
rect 9548 18640 9554 18692
rect 8128 18584 8616 18612
rect 6825 18575 6883 18581
rect 8662 18572 8668 18624
rect 8720 18612 8726 18624
rect 8757 18615 8815 18621
rect 8757 18612 8769 18615
rect 8720 18584 8769 18612
rect 8720 18572 8726 18584
rect 8757 18581 8769 18584
rect 8803 18612 8815 18615
rect 9858 18612 9864 18624
rect 8803 18584 9864 18612
rect 8803 18581 8815 18584
rect 8757 18575 8815 18581
rect 9858 18572 9864 18584
rect 9916 18572 9922 18624
rect 9968 18612 9996 18720
rect 10042 18708 10048 18760
rect 10100 18708 10106 18760
rect 12434 18748 12440 18760
rect 11914 18720 12440 18748
rect 12434 18708 12440 18720
rect 12492 18708 12498 18760
rect 13081 18751 13139 18757
rect 13081 18717 13093 18751
rect 13127 18748 13139 18751
rect 14182 18748 14188 18760
rect 13127 18720 14188 18748
rect 13127 18717 13139 18720
rect 13081 18711 13139 18717
rect 14182 18708 14188 18720
rect 14240 18708 14246 18760
rect 14274 18708 14280 18760
rect 14332 18708 14338 18760
rect 17126 18708 17132 18760
rect 17184 18748 17190 18760
rect 18141 18751 18199 18757
rect 18141 18748 18153 18751
rect 17184 18720 18153 18748
rect 17184 18708 17190 18720
rect 18141 18717 18153 18720
rect 18187 18748 18199 18751
rect 19076 18748 19104 18788
rect 18187 18720 19104 18748
rect 18187 18717 18199 18720
rect 18141 18711 18199 18717
rect 19242 18708 19248 18760
rect 19300 18748 19306 18760
rect 19426 18748 19432 18760
rect 19300 18720 19432 18748
rect 19300 18708 19306 18720
rect 19426 18708 19432 18720
rect 19484 18708 19490 18760
rect 19610 18708 19616 18760
rect 19668 18748 19674 18760
rect 20165 18751 20223 18757
rect 20165 18748 20177 18751
rect 19668 18720 20177 18748
rect 19668 18708 19674 18720
rect 20165 18717 20177 18720
rect 20211 18717 20223 18751
rect 20272 18748 20300 18788
rect 20441 18785 20453 18819
rect 20487 18816 20499 18819
rect 20622 18816 20628 18828
rect 20487 18788 20628 18816
rect 20487 18785 20499 18788
rect 20441 18779 20499 18785
rect 20622 18776 20628 18788
rect 20680 18776 20686 18828
rect 21729 18819 21787 18825
rect 21729 18785 21741 18819
rect 21775 18816 21787 18819
rect 21910 18816 21916 18828
rect 21775 18788 21916 18816
rect 21775 18785 21787 18788
rect 21729 18779 21787 18785
rect 21910 18776 21916 18788
rect 21968 18776 21974 18828
rect 25038 18816 25044 18828
rect 22066 18788 25044 18816
rect 21266 18748 21272 18760
rect 20272 18720 21272 18748
rect 20165 18711 20223 18717
rect 21266 18708 21272 18720
rect 21324 18708 21330 18760
rect 21545 18751 21603 18757
rect 21545 18717 21557 18751
rect 21591 18748 21603 18751
rect 22066 18748 22094 18788
rect 25038 18776 25044 18788
rect 25096 18776 25102 18828
rect 25240 18825 25268 18924
rect 26510 18912 26516 18924
rect 26568 18912 26574 18964
rect 28534 18912 28540 18964
rect 28592 18952 28598 18964
rect 28721 18955 28779 18961
rect 28721 18952 28733 18955
rect 28592 18924 28733 18952
rect 28592 18912 28598 18924
rect 28721 18921 28733 18924
rect 28767 18921 28779 18955
rect 28721 18915 28779 18921
rect 29546 18912 29552 18964
rect 29604 18952 29610 18964
rect 30098 18952 30104 18964
rect 29604 18924 30104 18952
rect 29604 18912 29610 18924
rect 30098 18912 30104 18924
rect 30156 18912 30162 18964
rect 30742 18912 30748 18964
rect 30800 18912 30806 18964
rect 32125 18955 32183 18961
rect 32125 18952 32137 18955
rect 31726 18924 32137 18952
rect 27522 18844 27528 18896
rect 27580 18884 27586 18896
rect 31726 18884 31754 18924
rect 32125 18921 32137 18924
rect 32171 18921 32183 18955
rect 33134 18952 33140 18964
rect 32125 18915 32183 18921
rect 32232 18924 33140 18952
rect 27580 18856 31754 18884
rect 27580 18844 27586 18856
rect 32030 18844 32036 18896
rect 32088 18884 32094 18896
rect 32232 18884 32260 18924
rect 33134 18912 33140 18924
rect 33192 18912 33198 18964
rect 33321 18955 33379 18961
rect 33321 18921 33333 18955
rect 33367 18952 33379 18955
rect 36538 18952 36544 18964
rect 33367 18924 36544 18952
rect 33367 18921 33379 18924
rect 33321 18915 33379 18921
rect 36538 18912 36544 18924
rect 36596 18912 36602 18964
rect 37369 18955 37427 18961
rect 37369 18921 37381 18955
rect 37415 18952 37427 18955
rect 40126 18952 40132 18964
rect 37415 18924 40132 18952
rect 37415 18921 37427 18924
rect 37369 18915 37427 18921
rect 40126 18912 40132 18924
rect 40184 18912 40190 18964
rect 41046 18912 41052 18964
rect 41104 18952 41110 18964
rect 41785 18955 41843 18961
rect 41785 18952 41797 18955
rect 41104 18924 41797 18952
rect 41104 18912 41110 18924
rect 41785 18921 41797 18924
rect 41831 18921 41843 18955
rect 41785 18915 41843 18921
rect 42150 18912 42156 18964
rect 42208 18952 42214 18964
rect 49234 18952 49240 18964
rect 42208 18924 49240 18952
rect 42208 18912 42214 18924
rect 49234 18912 49240 18924
rect 49292 18912 49298 18964
rect 35342 18884 35348 18896
rect 32088 18856 32260 18884
rect 32784 18856 35348 18884
rect 32088 18844 32094 18856
rect 25225 18819 25283 18825
rect 25225 18785 25237 18819
rect 25271 18785 25283 18819
rect 25225 18779 25283 18785
rect 26145 18819 26203 18825
rect 26145 18785 26157 18819
rect 26191 18816 26203 18819
rect 26602 18816 26608 18828
rect 26191 18788 26608 18816
rect 26191 18785 26203 18788
rect 26145 18779 26203 18785
rect 21591 18720 22094 18748
rect 21591 18717 21603 18720
rect 21545 18711 21603 18717
rect 22278 18708 22284 18760
rect 22336 18708 22342 18760
rect 23566 18708 23572 18760
rect 23624 18748 23630 18760
rect 23934 18748 23940 18760
rect 23624 18720 23940 18748
rect 23624 18708 23630 18720
rect 23934 18708 23940 18720
rect 23992 18708 23998 18760
rect 24026 18708 24032 18760
rect 24084 18748 24090 18760
rect 25240 18748 25268 18779
rect 26602 18776 26608 18788
rect 26660 18776 26666 18828
rect 27154 18776 27160 18828
rect 27212 18816 27218 18828
rect 27617 18819 27675 18825
rect 27212 18788 27476 18816
rect 27212 18776 27218 18788
rect 24084 18720 25268 18748
rect 25869 18751 25927 18757
rect 24084 18708 24090 18720
rect 25869 18717 25881 18751
rect 25915 18717 25927 18751
rect 25869 18711 25927 18717
rect 10778 18640 10784 18692
rect 10836 18640 10842 18692
rect 13725 18683 13783 18689
rect 12084 18652 13676 18680
rect 12084 18612 12112 18652
rect 9968 18584 12112 18612
rect 13648 18612 13676 18652
rect 13725 18649 13737 18683
rect 13771 18680 13783 18683
rect 14553 18683 14611 18689
rect 14553 18680 14565 18683
rect 13771 18652 14565 18680
rect 13771 18649 13783 18652
rect 13725 18643 13783 18649
rect 14553 18649 14565 18652
rect 14599 18649 14611 18683
rect 15838 18680 15844 18692
rect 15778 18652 15844 18680
rect 14553 18643 14611 18649
rect 15838 18640 15844 18652
rect 15896 18640 15902 18692
rect 16482 18640 16488 18692
rect 16540 18680 16546 18692
rect 16540 18652 17080 18680
rect 16540 18640 16546 18652
rect 15194 18612 15200 18624
rect 13648 18584 15200 18612
rect 15194 18572 15200 18584
rect 15252 18572 15258 18624
rect 15286 18572 15292 18624
rect 15344 18612 15350 18624
rect 16298 18612 16304 18624
rect 15344 18584 16304 18612
rect 15344 18572 15350 18584
rect 16298 18572 16304 18584
rect 16356 18612 16362 18624
rect 16853 18615 16911 18621
rect 16853 18612 16865 18615
rect 16356 18584 16865 18612
rect 16356 18572 16362 18584
rect 16853 18581 16865 18584
rect 16899 18581 16911 18615
rect 16853 18575 16911 18581
rect 16942 18572 16948 18624
rect 17000 18572 17006 18624
rect 17052 18612 17080 18652
rect 17862 18640 17868 18692
rect 17920 18680 17926 18692
rect 25884 18680 25912 18711
rect 17920 18652 21128 18680
rect 17920 18640 17926 18652
rect 18049 18615 18107 18621
rect 18049 18612 18061 18615
rect 17052 18584 18061 18612
rect 18049 18581 18061 18584
rect 18095 18581 18107 18615
rect 18049 18575 18107 18581
rect 19061 18615 19119 18621
rect 19061 18581 19073 18615
rect 19107 18612 19119 18615
rect 19242 18612 19248 18624
rect 19107 18584 19248 18612
rect 19107 18581 19119 18584
rect 19061 18575 19119 18581
rect 19242 18572 19248 18584
rect 19300 18572 19306 18624
rect 19334 18572 19340 18624
rect 19392 18572 19398 18624
rect 20257 18615 20315 18621
rect 20257 18581 20269 18615
rect 20303 18612 20315 18615
rect 20806 18612 20812 18624
rect 20303 18584 20812 18612
rect 20303 18581 20315 18584
rect 20257 18575 20315 18581
rect 20806 18572 20812 18584
rect 20864 18572 20870 18624
rect 21100 18621 21128 18652
rect 23860 18652 25912 18680
rect 21085 18615 21143 18621
rect 21085 18581 21097 18615
rect 21131 18581 21143 18615
rect 21085 18575 21143 18581
rect 21450 18572 21456 18624
rect 21508 18572 21514 18624
rect 21726 18572 21732 18624
rect 21784 18612 21790 18624
rect 22554 18612 22560 18624
rect 21784 18584 22560 18612
rect 21784 18572 21790 18584
rect 22554 18572 22560 18584
rect 22612 18572 22618 18624
rect 23382 18572 23388 18624
rect 23440 18612 23446 18624
rect 23860 18612 23888 18652
rect 26142 18640 26148 18692
rect 26200 18680 26206 18692
rect 26602 18680 26608 18692
rect 26200 18652 26608 18680
rect 26200 18640 26206 18652
rect 26602 18640 26608 18652
rect 26660 18640 26666 18692
rect 27448 18680 27476 18788
rect 27617 18785 27629 18819
rect 27663 18816 27675 18819
rect 29638 18816 29644 18828
rect 27663 18788 29644 18816
rect 27663 18785 27675 18788
rect 27617 18779 27675 18785
rect 29638 18776 29644 18788
rect 29696 18776 29702 18828
rect 29822 18776 29828 18828
rect 29880 18816 29886 18828
rect 30285 18819 30343 18825
rect 30285 18816 30297 18819
rect 29880 18788 30297 18816
rect 29880 18776 29886 18788
rect 30285 18785 30297 18788
rect 30331 18785 30343 18819
rect 30285 18779 30343 18785
rect 30742 18776 30748 18828
rect 30800 18816 30806 18828
rect 31389 18819 31447 18825
rect 31389 18816 31401 18819
rect 30800 18788 31401 18816
rect 30800 18776 30806 18788
rect 31389 18785 31401 18788
rect 31435 18785 31447 18819
rect 31389 18779 31447 18785
rect 31573 18819 31631 18825
rect 31573 18785 31585 18819
rect 31619 18816 31631 18819
rect 32214 18816 32220 18828
rect 31619 18788 32220 18816
rect 31619 18785 31631 18788
rect 31573 18779 31631 18785
rect 32214 18776 32220 18788
rect 32272 18776 32278 18828
rect 32784 18825 32812 18856
rect 35342 18844 35348 18856
rect 35400 18844 35406 18896
rect 37550 18844 37556 18896
rect 37608 18884 37614 18896
rect 38013 18887 38071 18893
rect 38013 18884 38025 18887
rect 37608 18856 38025 18884
rect 37608 18844 37614 18856
rect 38013 18853 38025 18856
rect 38059 18853 38071 18887
rect 38013 18847 38071 18853
rect 38194 18844 38200 18896
rect 38252 18884 38258 18896
rect 38252 18856 38608 18884
rect 38252 18844 38258 18856
rect 32769 18819 32827 18825
rect 32769 18785 32781 18819
rect 32815 18785 32827 18819
rect 32769 18779 32827 18785
rect 33502 18776 33508 18828
rect 33560 18816 33566 18828
rect 33870 18816 33876 18828
rect 33560 18788 33876 18816
rect 33560 18776 33566 18788
rect 33870 18776 33876 18788
rect 33928 18776 33934 18828
rect 33965 18819 34023 18825
rect 33965 18785 33977 18819
rect 34011 18816 34023 18819
rect 35250 18816 35256 18828
rect 34011 18788 35256 18816
rect 34011 18785 34023 18788
rect 33965 18779 34023 18785
rect 35250 18776 35256 18788
rect 35308 18776 35314 18828
rect 35618 18776 35624 18828
rect 35676 18776 35682 18828
rect 35897 18819 35955 18825
rect 35897 18785 35909 18819
rect 35943 18816 35955 18819
rect 38470 18816 38476 18828
rect 35943 18788 38476 18816
rect 35943 18785 35955 18788
rect 35897 18779 35955 18785
rect 38470 18776 38476 18788
rect 38528 18776 38534 18828
rect 38580 18825 38608 18856
rect 42242 18844 42248 18896
rect 42300 18884 42306 18896
rect 43165 18887 43223 18893
rect 43165 18884 43177 18887
rect 42300 18856 43177 18884
rect 42300 18844 42306 18856
rect 38565 18819 38623 18825
rect 38565 18785 38577 18819
rect 38611 18785 38623 18819
rect 38565 18779 38623 18785
rect 40313 18819 40371 18825
rect 40313 18785 40325 18819
rect 40359 18816 40371 18819
rect 42334 18816 42340 18828
rect 40359 18788 42340 18816
rect 40359 18785 40371 18788
rect 40313 18779 40371 18785
rect 42334 18776 42340 18788
rect 42392 18776 42398 18828
rect 27522 18708 27528 18760
rect 27580 18748 27586 18760
rect 28077 18751 28135 18757
rect 28077 18748 28089 18751
rect 27580 18720 28089 18748
rect 27580 18708 27586 18720
rect 28077 18717 28089 18720
rect 28123 18717 28135 18751
rect 28077 18711 28135 18717
rect 28626 18708 28632 18760
rect 28684 18748 28690 18760
rect 29178 18748 29184 18760
rect 28684 18720 29184 18748
rect 28684 18708 28690 18720
rect 29178 18708 29184 18720
rect 29236 18708 29242 18760
rect 29362 18708 29368 18760
rect 29420 18748 29426 18760
rect 30193 18751 30251 18757
rect 30193 18748 30205 18751
rect 29420 18720 30205 18748
rect 29420 18708 29426 18720
rect 30193 18717 30205 18720
rect 30239 18717 30251 18751
rect 30193 18711 30251 18717
rect 31202 18708 31208 18760
rect 31260 18748 31266 18760
rect 31297 18751 31355 18757
rect 31297 18748 31309 18751
rect 31260 18720 31309 18748
rect 31260 18708 31266 18720
rect 31297 18717 31309 18720
rect 31343 18717 31355 18751
rect 34333 18751 34391 18757
rect 34333 18748 34345 18751
rect 31297 18711 31355 18717
rect 31404 18720 34345 18748
rect 31404 18692 31432 18720
rect 34333 18717 34345 18720
rect 34379 18717 34391 18751
rect 34333 18711 34391 18717
rect 37182 18708 37188 18760
rect 37240 18748 37246 18760
rect 39393 18751 39451 18757
rect 39393 18748 39405 18751
rect 37240 18720 39405 18748
rect 37240 18708 37246 18720
rect 39393 18717 39405 18720
rect 39439 18717 39451 18751
rect 39393 18711 39451 18717
rect 40037 18751 40095 18757
rect 40037 18717 40049 18751
rect 40083 18717 40095 18751
rect 40037 18711 40095 18717
rect 29454 18680 29460 18692
rect 27448 18652 29460 18680
rect 29454 18640 29460 18652
rect 29512 18640 29518 18692
rect 31386 18640 31392 18692
rect 31444 18640 31450 18692
rect 32585 18683 32643 18689
rect 32585 18649 32597 18683
rect 32631 18680 32643 18683
rect 35894 18680 35900 18692
rect 32631 18652 35900 18680
rect 32631 18649 32643 18652
rect 32585 18643 32643 18649
rect 35894 18640 35900 18652
rect 35952 18640 35958 18692
rect 36630 18640 36636 18692
rect 36688 18640 36694 18692
rect 37826 18640 37832 18692
rect 37884 18680 37890 18692
rect 40052 18680 40080 18711
rect 41690 18708 41696 18760
rect 41748 18748 41754 18760
rect 42245 18751 42303 18757
rect 42245 18748 42257 18751
rect 41748 18720 42257 18748
rect 41748 18708 41754 18720
rect 42245 18717 42257 18720
rect 42291 18717 42303 18751
rect 42245 18711 42303 18717
rect 41598 18680 41604 18692
rect 37884 18652 40080 18680
rect 41538 18652 41604 18680
rect 37884 18640 37890 18652
rect 41598 18640 41604 18652
rect 41656 18680 41662 18692
rect 42444 18680 42472 18856
rect 43165 18853 43177 18856
rect 43211 18853 43223 18887
rect 43165 18847 43223 18853
rect 48593 18751 48651 18757
rect 48593 18717 48605 18751
rect 48639 18748 48651 18751
rect 48774 18748 48780 18760
rect 48639 18720 48780 18748
rect 48639 18717 48651 18720
rect 48593 18711 48651 18717
rect 48774 18708 48780 18720
rect 48832 18708 48838 18760
rect 49053 18751 49111 18757
rect 49053 18717 49065 18751
rect 49099 18748 49111 18751
rect 49142 18748 49148 18760
rect 49099 18720 49148 18748
rect 49099 18717 49111 18720
rect 49053 18711 49111 18717
rect 49142 18708 49148 18720
rect 49200 18708 49206 18760
rect 42610 18680 42616 18692
rect 41656 18652 42616 18680
rect 41656 18640 41662 18652
rect 42610 18640 42616 18652
rect 42668 18640 42674 18692
rect 23440 18584 23888 18612
rect 23440 18572 23446 18584
rect 24026 18572 24032 18624
rect 24084 18572 24090 18624
rect 24670 18572 24676 18624
rect 24728 18612 24734 18624
rect 24949 18615 25007 18621
rect 24949 18612 24961 18615
rect 24728 18584 24961 18612
rect 24728 18572 24734 18584
rect 24949 18581 24961 18584
rect 24995 18581 25007 18615
rect 24949 18575 25007 18581
rect 25041 18615 25099 18621
rect 25041 18581 25053 18615
rect 25087 18612 25099 18615
rect 25406 18612 25412 18624
rect 25087 18584 25412 18612
rect 25087 18581 25099 18584
rect 25041 18575 25099 18581
rect 25406 18572 25412 18584
rect 25464 18572 25470 18624
rect 26418 18572 26424 18624
rect 26476 18612 26482 18624
rect 28534 18612 28540 18624
rect 26476 18584 28540 18612
rect 26476 18572 26482 18584
rect 28534 18572 28540 18584
rect 28592 18572 28598 18624
rect 29086 18572 29092 18624
rect 29144 18572 29150 18624
rect 29733 18615 29791 18621
rect 29733 18581 29745 18615
rect 29779 18612 29791 18615
rect 30006 18612 30012 18624
rect 29779 18584 30012 18612
rect 29779 18581 29791 18584
rect 29733 18575 29791 18581
rect 30006 18572 30012 18584
rect 30064 18572 30070 18624
rect 30098 18572 30104 18624
rect 30156 18572 30162 18624
rect 30929 18615 30987 18621
rect 30929 18581 30941 18615
rect 30975 18612 30987 18615
rect 31294 18612 31300 18624
rect 30975 18584 31300 18612
rect 30975 18581 30987 18584
rect 30929 18575 30987 18581
rect 31294 18572 31300 18584
rect 31352 18572 31358 18624
rect 32030 18572 32036 18624
rect 32088 18612 32094 18624
rect 32493 18615 32551 18621
rect 32493 18612 32505 18615
rect 32088 18584 32505 18612
rect 32088 18572 32094 18584
rect 32493 18581 32505 18584
rect 32539 18581 32551 18615
rect 32493 18575 32551 18581
rect 33594 18572 33600 18624
rect 33652 18612 33658 18624
rect 33689 18615 33747 18621
rect 33689 18612 33701 18615
rect 33652 18584 33701 18612
rect 33652 18572 33658 18584
rect 33689 18581 33701 18584
rect 33735 18581 33747 18615
rect 33689 18575 33747 18581
rect 33781 18615 33839 18621
rect 33781 18581 33793 18615
rect 33827 18612 33839 18615
rect 33962 18612 33968 18624
rect 33827 18584 33968 18612
rect 33827 18581 33839 18584
rect 33781 18575 33839 18581
rect 33962 18572 33968 18584
rect 34020 18572 34026 18624
rect 34885 18615 34943 18621
rect 34885 18581 34897 18615
rect 34931 18612 34943 18615
rect 35802 18612 35808 18624
rect 34931 18584 35808 18612
rect 34931 18581 34943 18584
rect 34885 18575 34943 18581
rect 35802 18572 35808 18584
rect 35860 18572 35866 18624
rect 36906 18572 36912 18624
rect 36964 18612 36970 18624
rect 37645 18615 37703 18621
rect 37645 18612 37657 18615
rect 36964 18584 37657 18612
rect 36964 18572 36970 18584
rect 37645 18581 37657 18584
rect 37691 18581 37703 18615
rect 37645 18575 37703 18581
rect 37734 18572 37740 18624
rect 37792 18612 37798 18624
rect 38381 18615 38439 18621
rect 38381 18612 38393 18615
rect 37792 18584 38393 18612
rect 37792 18572 37798 18584
rect 38381 18581 38393 18584
rect 38427 18581 38439 18615
rect 38381 18575 38439 18581
rect 38470 18572 38476 18624
rect 38528 18572 38534 18624
rect 39206 18572 39212 18624
rect 39264 18572 39270 18624
rect 42794 18572 42800 18624
rect 42852 18612 42858 18624
rect 42889 18615 42947 18621
rect 42889 18612 42901 18615
rect 42852 18584 42901 18612
rect 42852 18572 42858 18584
rect 42889 18581 42901 18584
rect 42935 18581 42947 18615
rect 42889 18575 42947 18581
rect 48406 18572 48412 18624
rect 48464 18572 48470 18624
rect 48866 18572 48872 18624
rect 48924 18612 48930 18624
rect 49237 18615 49295 18621
rect 49237 18612 49249 18615
rect 48924 18584 49249 18612
rect 48924 18572 48930 18584
rect 49237 18581 49249 18584
rect 49283 18581 49295 18615
rect 49237 18575 49295 18581
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 7282 18368 7288 18420
rect 7340 18408 7346 18420
rect 7340 18380 10272 18408
rect 7340 18368 7346 18380
rect 3697 18343 3755 18349
rect 3697 18309 3709 18343
rect 3743 18340 3755 18343
rect 4062 18340 4068 18352
rect 3743 18312 4068 18340
rect 3743 18309 3755 18312
rect 3697 18303 3755 18309
rect 4062 18300 4068 18312
rect 4120 18300 4126 18352
rect 5813 18343 5871 18349
rect 5813 18309 5825 18343
rect 5859 18340 5871 18343
rect 6362 18340 6368 18352
rect 5859 18312 6368 18340
rect 5859 18309 5871 18312
rect 5813 18303 5871 18309
rect 6362 18300 6368 18312
rect 6420 18300 6426 18352
rect 6454 18300 6460 18352
rect 6512 18340 6518 18352
rect 6512 18312 7328 18340
rect 6512 18300 6518 18312
rect 1762 18232 1768 18284
rect 1820 18232 1826 18284
rect 3510 18232 3516 18284
rect 3568 18232 3574 18284
rect 4706 18232 4712 18284
rect 4764 18232 4770 18284
rect 5353 18275 5411 18281
rect 5353 18241 5365 18275
rect 5399 18241 5411 18275
rect 5353 18235 5411 18241
rect 2774 18164 2780 18216
rect 2832 18164 2838 18216
rect 5166 18096 5172 18148
rect 5224 18096 5230 18148
rect 5368 18136 5396 18235
rect 7190 18232 7196 18284
rect 7248 18232 7254 18284
rect 7300 18272 7328 18312
rect 7742 18300 7748 18352
rect 7800 18300 7806 18352
rect 8389 18343 8447 18349
rect 8389 18309 8401 18343
rect 8435 18340 8447 18343
rect 8662 18340 8668 18352
rect 8435 18312 8668 18340
rect 8435 18309 8447 18312
rect 8389 18303 8447 18309
rect 7929 18275 7987 18281
rect 7929 18272 7941 18275
rect 7300 18244 7941 18272
rect 7929 18241 7941 18244
rect 7975 18241 7987 18275
rect 7929 18235 7987 18241
rect 6086 18136 6092 18148
rect 5368 18108 6092 18136
rect 6086 18096 6092 18108
rect 6144 18096 6150 18148
rect 6733 18139 6791 18145
rect 6733 18105 6745 18139
rect 6779 18136 6791 18139
rect 8588 18136 8616 18312
rect 8662 18300 8668 18312
rect 8720 18300 8726 18352
rect 10244 18340 10272 18380
rect 10318 18368 10324 18420
rect 10376 18408 10382 18420
rect 12802 18408 12808 18420
rect 10376 18380 12808 18408
rect 10376 18368 10382 18380
rect 12802 18368 12808 18380
rect 12860 18368 12866 18420
rect 14829 18411 14887 18417
rect 14829 18408 14841 18411
rect 13280 18380 14841 18408
rect 13280 18340 13308 18380
rect 14829 18377 14841 18380
rect 14875 18377 14887 18411
rect 14829 18371 14887 18377
rect 15194 18368 15200 18420
rect 15252 18368 15258 18420
rect 16206 18368 16212 18420
rect 16264 18368 16270 18420
rect 17126 18368 17132 18420
rect 17184 18368 17190 18420
rect 17862 18368 17868 18420
rect 17920 18368 17926 18420
rect 18708 18380 21220 18408
rect 18708 18349 18736 18380
rect 18693 18343 18751 18349
rect 10244 18312 13308 18340
rect 17052 18312 18552 18340
rect 9950 18232 9956 18284
rect 10008 18272 10014 18284
rect 10008 18244 11100 18272
rect 10008 18232 10014 18244
rect 8665 18207 8723 18213
rect 8665 18173 8677 18207
rect 8711 18173 8723 18207
rect 8665 18167 8723 18173
rect 8941 18207 8999 18213
rect 8941 18173 8953 18207
rect 8987 18204 8999 18207
rect 9582 18204 9588 18216
rect 8987 18176 9588 18204
rect 8987 18173 8999 18176
rect 8941 18167 8999 18173
rect 6779 18108 8616 18136
rect 6779 18105 6791 18108
rect 6733 18099 6791 18105
rect 4525 18071 4583 18077
rect 4525 18037 4537 18071
rect 4571 18068 4583 18071
rect 6454 18068 6460 18080
rect 4571 18040 6460 18068
rect 4571 18037 4583 18040
rect 4525 18031 4583 18037
rect 6454 18028 6460 18040
rect 6512 18028 6518 18080
rect 7006 18028 7012 18080
rect 7064 18028 7070 18080
rect 8294 18028 8300 18080
rect 8352 18068 8358 18080
rect 8570 18068 8576 18080
rect 8352 18040 8576 18068
rect 8352 18028 8358 18040
rect 8570 18028 8576 18040
rect 8628 18028 8634 18080
rect 8680 18068 8708 18167
rect 9582 18164 9588 18176
rect 9640 18164 9646 18216
rect 10965 18207 11023 18213
rect 10965 18173 10977 18207
rect 11011 18173 11023 18207
rect 11072 18204 11100 18244
rect 11146 18232 11152 18284
rect 11204 18272 11210 18284
rect 11609 18275 11667 18281
rect 11609 18272 11621 18275
rect 11204 18244 11621 18272
rect 11204 18232 11210 18244
rect 11609 18241 11621 18244
rect 11655 18241 11667 18275
rect 11609 18235 11667 18241
rect 11624 18204 11652 18235
rect 11790 18232 11796 18284
rect 11848 18272 11854 18284
rect 12161 18275 12219 18281
rect 12161 18272 12173 18275
rect 11848 18244 12173 18272
rect 11848 18232 11854 18244
rect 12161 18241 12173 18244
rect 12207 18241 12219 18275
rect 12161 18235 12219 18241
rect 13998 18232 14004 18284
rect 14056 18232 14062 18284
rect 14182 18232 14188 18284
rect 14240 18272 14246 18284
rect 14240 18244 15424 18272
rect 14240 18232 14246 18244
rect 11072 18176 11376 18204
rect 11624 18176 12204 18204
rect 10965 18167 11023 18173
rect 10410 18096 10416 18148
rect 10468 18096 10474 18148
rect 10778 18068 10784 18080
rect 8680 18040 10784 18068
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 10873 18071 10931 18077
rect 10873 18037 10885 18071
rect 10919 18068 10931 18071
rect 10980 18068 11008 18167
rect 11054 18068 11060 18080
rect 10919 18040 11060 18068
rect 10919 18037 10931 18040
rect 10873 18031 10931 18037
rect 11054 18028 11060 18040
rect 11112 18028 11118 18080
rect 11238 18028 11244 18080
rect 11296 18068 11302 18080
rect 11348 18068 11376 18176
rect 11977 18139 12035 18145
rect 11977 18105 11989 18139
rect 12023 18136 12035 18139
rect 12066 18136 12072 18148
rect 12023 18108 12072 18136
rect 12023 18105 12035 18108
rect 11977 18099 12035 18105
rect 12066 18096 12072 18108
rect 12124 18096 12130 18148
rect 12176 18136 12204 18176
rect 12342 18164 12348 18216
rect 12400 18204 12406 18216
rect 12621 18207 12679 18213
rect 12621 18204 12633 18207
rect 12400 18176 12633 18204
rect 12400 18164 12406 18176
rect 12621 18173 12633 18176
rect 12667 18204 12679 18207
rect 12897 18207 12955 18213
rect 12667 18176 12756 18204
rect 12667 18173 12679 18176
rect 12621 18167 12679 18173
rect 12526 18136 12532 18148
rect 12176 18108 12532 18136
rect 12526 18096 12532 18108
rect 12584 18096 12590 18148
rect 12434 18068 12440 18080
rect 11296 18040 12440 18068
rect 11296 18028 11302 18040
rect 12434 18028 12440 18040
rect 12492 18028 12498 18080
rect 12728 18068 12756 18176
rect 12897 18173 12909 18207
rect 12943 18204 12955 18207
rect 13354 18204 13360 18216
rect 12943 18176 13360 18204
rect 12943 18173 12955 18176
rect 12897 18167 12955 18173
rect 13354 18164 13360 18176
rect 13412 18164 13418 18216
rect 13446 18164 13452 18216
rect 13504 18204 13510 18216
rect 15396 18213 15424 18244
rect 15470 18232 15476 18284
rect 15528 18272 15534 18284
rect 16117 18275 16175 18281
rect 16117 18272 16129 18275
rect 15528 18244 16129 18272
rect 15528 18232 15534 18244
rect 16117 18241 16129 18244
rect 16163 18272 16175 18275
rect 17052 18272 17080 18312
rect 16163 18244 17080 18272
rect 17773 18275 17831 18281
rect 16163 18241 16175 18244
rect 16117 18235 16175 18241
rect 17773 18241 17785 18275
rect 17819 18272 17831 18275
rect 18414 18272 18420 18284
rect 17819 18244 18420 18272
rect 17819 18241 17831 18244
rect 17773 18235 17831 18241
rect 18414 18232 18420 18244
rect 18472 18232 18478 18284
rect 18524 18272 18552 18312
rect 18693 18309 18705 18343
rect 18739 18309 18751 18343
rect 19978 18340 19984 18352
rect 18693 18303 18751 18309
rect 18800 18312 19984 18340
rect 18800 18272 18828 18312
rect 19978 18300 19984 18312
rect 20036 18300 20042 18352
rect 20162 18300 20168 18352
rect 20220 18340 20226 18352
rect 20220 18312 20378 18340
rect 20220 18300 20226 18312
rect 18524 18244 18828 18272
rect 19242 18232 19248 18284
rect 19300 18232 19306 18284
rect 14369 18207 14427 18213
rect 14369 18204 14381 18207
rect 13504 18176 14381 18204
rect 13504 18164 13510 18176
rect 14369 18173 14381 18176
rect 14415 18173 14427 18207
rect 14369 18167 14427 18173
rect 15289 18207 15347 18213
rect 15289 18173 15301 18207
rect 15335 18173 15347 18207
rect 15289 18167 15347 18173
rect 15381 18207 15439 18213
rect 15381 18173 15393 18207
rect 15427 18204 15439 18207
rect 16022 18204 16028 18216
rect 15427 18176 16028 18204
rect 15427 18173 15439 18176
rect 15381 18167 15439 18173
rect 13998 18096 14004 18148
rect 14056 18136 14062 18148
rect 15304 18136 15332 18167
rect 16022 18164 16028 18176
rect 16080 18164 16086 18216
rect 16758 18204 16764 18216
rect 16408 18176 16764 18204
rect 16408 18136 16436 18176
rect 16758 18164 16764 18176
rect 16816 18164 16822 18216
rect 17678 18164 17684 18216
rect 17736 18204 17742 18216
rect 17957 18207 18015 18213
rect 17957 18204 17969 18207
rect 17736 18176 17969 18204
rect 17736 18164 17742 18176
rect 17957 18173 17969 18176
rect 18003 18173 18015 18207
rect 17957 18167 18015 18173
rect 18598 18164 18604 18216
rect 18656 18204 18662 18216
rect 19613 18207 19671 18213
rect 19613 18204 19625 18207
rect 18656 18176 19625 18204
rect 18656 18164 18662 18176
rect 19613 18173 19625 18176
rect 19659 18173 19671 18207
rect 19613 18167 19671 18173
rect 19886 18164 19892 18216
rect 19944 18164 19950 18216
rect 14056 18108 14412 18136
rect 15304 18108 16436 18136
rect 14056 18096 14062 18108
rect 14274 18068 14280 18080
rect 12728 18040 14280 18068
rect 14274 18028 14280 18040
rect 14332 18028 14338 18080
rect 14384 18068 14412 18108
rect 16482 18096 16488 18148
rect 16540 18136 16546 18148
rect 16853 18139 16911 18145
rect 16853 18136 16865 18139
rect 16540 18108 16865 18136
rect 16540 18096 16546 18108
rect 16853 18105 16865 18108
rect 16899 18105 16911 18139
rect 16853 18099 16911 18105
rect 17034 18096 17040 18148
rect 17092 18136 17098 18148
rect 18877 18139 18935 18145
rect 18877 18136 18889 18139
rect 17092 18108 18889 18136
rect 17092 18096 17098 18108
rect 18877 18105 18889 18108
rect 18923 18105 18935 18139
rect 21192 18136 21220 18380
rect 21450 18368 21456 18420
rect 21508 18408 21514 18420
rect 24673 18411 24731 18417
rect 24673 18408 24685 18411
rect 21508 18380 24685 18408
rect 21508 18368 21514 18380
rect 24673 18377 24685 18380
rect 24719 18377 24731 18411
rect 24673 18371 24731 18377
rect 25130 18368 25136 18420
rect 25188 18408 25194 18420
rect 25498 18408 25504 18420
rect 25188 18380 25504 18408
rect 25188 18368 25194 18380
rect 25498 18368 25504 18380
rect 25556 18368 25562 18420
rect 26237 18411 26295 18417
rect 26237 18377 26249 18411
rect 26283 18408 26295 18411
rect 27246 18408 27252 18420
rect 26283 18380 27252 18408
rect 26283 18377 26295 18380
rect 26237 18371 26295 18377
rect 27246 18368 27252 18380
rect 27304 18368 27310 18420
rect 27706 18408 27712 18420
rect 27448 18380 27712 18408
rect 21266 18300 21272 18352
rect 21324 18340 21330 18352
rect 23198 18340 23204 18352
rect 21324 18312 23204 18340
rect 21324 18300 21330 18312
rect 23198 18300 23204 18312
rect 23256 18300 23262 18352
rect 23382 18300 23388 18352
rect 23440 18300 23446 18352
rect 23842 18300 23848 18352
rect 23900 18340 23906 18352
rect 24029 18343 24087 18349
rect 24029 18340 24041 18343
rect 23900 18312 24041 18340
rect 23900 18300 23906 18312
rect 24029 18309 24041 18312
rect 24075 18309 24087 18343
rect 27448 18340 27476 18380
rect 27706 18368 27712 18380
rect 27764 18368 27770 18420
rect 29457 18411 29515 18417
rect 29457 18408 29469 18411
rect 28736 18380 29469 18408
rect 24029 18303 24087 18309
rect 24964 18312 27476 18340
rect 27525 18343 27583 18349
rect 22189 18275 22247 18281
rect 22189 18241 22201 18275
rect 22235 18241 22247 18275
rect 22189 18235 22247 18241
rect 22649 18275 22707 18281
rect 22649 18241 22661 18275
rect 22695 18272 22707 18275
rect 23290 18272 23296 18284
rect 22695 18244 23296 18272
rect 22695 18241 22707 18244
rect 22649 18235 22707 18241
rect 22204 18204 22232 18235
rect 23290 18232 23296 18244
rect 23348 18232 23354 18284
rect 24854 18272 24860 18284
rect 23952 18244 24860 18272
rect 23952 18204 23980 18244
rect 24854 18232 24860 18244
rect 24912 18232 24918 18284
rect 22204 18176 23980 18204
rect 24578 18136 24584 18148
rect 21192 18108 24584 18136
rect 18877 18099 18935 18105
rect 24578 18096 24584 18108
rect 24636 18096 24642 18148
rect 15838 18068 15844 18080
rect 14384 18040 15844 18068
rect 15838 18028 15844 18040
rect 15896 18028 15902 18080
rect 16574 18028 16580 18080
rect 16632 18068 16638 18080
rect 16669 18071 16727 18077
rect 16669 18068 16681 18071
rect 16632 18040 16681 18068
rect 16632 18028 16638 18040
rect 16669 18037 16681 18040
rect 16715 18037 16727 18071
rect 16669 18031 16727 18037
rect 17402 18028 17408 18080
rect 17460 18028 17466 18080
rect 21361 18071 21419 18077
rect 21361 18037 21373 18071
rect 21407 18068 21419 18071
rect 21726 18068 21732 18080
rect 21407 18040 21732 18068
rect 21407 18037 21419 18040
rect 21361 18031 21419 18037
rect 21726 18028 21732 18040
rect 21784 18028 21790 18080
rect 22002 18028 22008 18080
rect 22060 18028 22066 18080
rect 23198 18028 23204 18080
rect 23256 18068 23262 18080
rect 24964 18068 24992 18312
rect 27525 18309 27537 18343
rect 27571 18340 27583 18343
rect 28736 18340 28764 18380
rect 29457 18377 29469 18380
rect 29503 18408 29515 18411
rect 30098 18408 30104 18420
rect 29503 18380 30104 18408
rect 29503 18377 29515 18380
rect 29457 18371 29515 18377
rect 30098 18368 30104 18380
rect 30156 18368 30162 18420
rect 30193 18411 30251 18417
rect 30193 18377 30205 18411
rect 30239 18408 30251 18411
rect 30374 18408 30380 18420
rect 30239 18380 30380 18408
rect 30239 18377 30251 18380
rect 30193 18371 30251 18377
rect 30374 18368 30380 18380
rect 30432 18368 30438 18420
rect 30929 18411 30987 18417
rect 30929 18377 30941 18411
rect 30975 18408 30987 18411
rect 31110 18408 31116 18420
rect 30975 18380 31116 18408
rect 30975 18377 30987 18380
rect 30929 18371 30987 18377
rect 31110 18368 31116 18380
rect 31168 18368 31174 18420
rect 31297 18411 31355 18417
rect 31297 18377 31309 18411
rect 31343 18408 31355 18411
rect 31343 18380 31892 18408
rect 31343 18377 31355 18380
rect 31297 18371 31355 18377
rect 27571 18312 28764 18340
rect 28813 18343 28871 18349
rect 27571 18309 27583 18312
rect 27525 18303 27583 18309
rect 28813 18309 28825 18343
rect 28859 18340 28871 18343
rect 31754 18340 31760 18352
rect 28859 18312 31760 18340
rect 28859 18309 28871 18312
rect 28813 18303 28871 18309
rect 31754 18300 31760 18312
rect 31812 18300 31818 18352
rect 25038 18232 25044 18284
rect 25096 18272 25102 18284
rect 26510 18272 26516 18284
rect 25096 18244 26516 18272
rect 25096 18232 25102 18244
rect 26510 18232 26516 18244
rect 26568 18232 26574 18284
rect 27617 18275 27675 18281
rect 27617 18241 27629 18275
rect 27663 18272 27675 18275
rect 28626 18272 28632 18284
rect 27663 18244 28632 18272
rect 27663 18241 27675 18244
rect 27617 18235 27675 18241
rect 28626 18232 28632 18244
rect 28684 18232 28690 18284
rect 28721 18275 28779 18281
rect 28721 18241 28733 18275
rect 28767 18241 28779 18275
rect 28721 18235 28779 18241
rect 25222 18164 25228 18216
rect 25280 18164 25286 18216
rect 26329 18207 26387 18213
rect 26329 18173 26341 18207
rect 26375 18173 26387 18207
rect 26329 18167 26387 18173
rect 26344 18136 26372 18167
rect 26418 18164 26424 18216
rect 26476 18164 26482 18216
rect 26786 18164 26792 18216
rect 26844 18204 26850 18216
rect 27709 18207 27767 18213
rect 27709 18204 27721 18207
rect 26844 18176 27721 18204
rect 26844 18164 26850 18176
rect 27709 18173 27721 18176
rect 27755 18173 27767 18207
rect 28736 18204 28764 18235
rect 30098 18232 30104 18284
rect 30156 18272 30162 18284
rect 31864 18272 31892 18380
rect 33410 18368 33416 18420
rect 33468 18408 33474 18420
rect 35897 18411 35955 18417
rect 35897 18408 35909 18411
rect 33468 18380 35909 18408
rect 33468 18368 33474 18380
rect 35897 18377 35909 18380
rect 35943 18377 35955 18411
rect 35897 18371 35955 18377
rect 36357 18411 36415 18417
rect 36357 18377 36369 18411
rect 36403 18408 36415 18411
rect 38470 18408 38476 18420
rect 36403 18380 38476 18408
rect 36403 18377 36415 18380
rect 36357 18371 36415 18377
rect 38470 18368 38476 18380
rect 38528 18368 38534 18420
rect 39758 18408 39764 18420
rect 38672 18380 39764 18408
rect 33594 18340 33600 18352
rect 32600 18312 33600 18340
rect 32600 18272 32628 18312
rect 33594 18300 33600 18312
rect 33652 18300 33658 18352
rect 34146 18300 34152 18352
rect 34204 18340 34210 18352
rect 37366 18340 37372 18352
rect 34204 18312 34362 18340
rect 36188 18312 37372 18340
rect 34204 18300 34210 18312
rect 30156 18244 31800 18272
rect 31864 18244 32628 18272
rect 32677 18275 32735 18281
rect 30156 18232 30162 18244
rect 28810 18204 28816 18216
rect 28736 18176 28816 18204
rect 27709 18167 27767 18173
rect 28810 18164 28816 18176
rect 28868 18164 28874 18216
rect 28902 18164 28908 18216
rect 28960 18164 28966 18216
rect 29546 18164 29552 18216
rect 29604 18204 29610 18216
rect 30285 18207 30343 18213
rect 30285 18204 30297 18207
rect 29604 18176 30297 18204
rect 29604 18164 29610 18176
rect 30285 18173 30297 18176
rect 30331 18204 30343 18207
rect 30558 18204 30564 18216
rect 30331 18176 30564 18204
rect 30331 18173 30343 18176
rect 30285 18167 30343 18173
rect 30558 18164 30564 18176
rect 30616 18164 30622 18216
rect 31386 18164 31392 18216
rect 31444 18164 31450 18216
rect 31570 18164 31576 18216
rect 31628 18164 31634 18216
rect 31772 18204 31800 18244
rect 32677 18241 32689 18275
rect 32723 18241 32735 18275
rect 32677 18235 32735 18241
rect 32769 18275 32827 18281
rect 32769 18241 32781 18275
rect 32815 18272 32827 18275
rect 33134 18272 33140 18284
rect 32815 18244 33140 18272
rect 32815 18241 32827 18244
rect 32769 18235 32827 18241
rect 32306 18204 32312 18216
rect 31772 18176 32312 18204
rect 32306 18164 32312 18176
rect 32364 18204 32370 18216
rect 32692 18204 32720 18235
rect 33134 18232 33140 18244
rect 33192 18232 33198 18284
rect 32364 18176 32720 18204
rect 32364 18164 32370 18176
rect 32858 18164 32864 18216
rect 32916 18164 32922 18216
rect 33597 18207 33655 18213
rect 33597 18173 33609 18207
rect 33643 18173 33655 18207
rect 33597 18167 33655 18173
rect 30466 18136 30472 18148
rect 26344 18108 30472 18136
rect 30466 18096 30472 18108
rect 30524 18096 30530 18148
rect 31404 18136 31432 18164
rect 31404 18108 31616 18136
rect 31588 18080 31616 18108
rect 32490 18096 32496 18148
rect 32548 18136 32554 18148
rect 33612 18136 33640 18167
rect 33870 18164 33876 18216
rect 33928 18204 33934 18216
rect 36188 18204 36216 18312
rect 37366 18300 37372 18312
rect 37424 18300 37430 18352
rect 37458 18300 37464 18352
rect 37516 18340 37522 18352
rect 38672 18340 38700 18380
rect 39758 18368 39764 18380
rect 39816 18368 39822 18420
rect 40034 18368 40040 18420
rect 40092 18408 40098 18420
rect 40865 18411 40923 18417
rect 40865 18408 40877 18411
rect 40092 18380 40877 18408
rect 40092 18368 40098 18380
rect 40865 18377 40877 18380
rect 40911 18377 40923 18411
rect 40865 18371 40923 18377
rect 42150 18368 42156 18420
rect 42208 18368 42214 18420
rect 48774 18368 48780 18420
rect 48832 18368 48838 18420
rect 37516 18312 38700 18340
rect 37516 18300 37522 18312
rect 38838 18300 38844 18352
rect 38896 18300 38902 18352
rect 40773 18343 40831 18349
rect 40773 18309 40785 18343
rect 40819 18340 40831 18343
rect 48406 18340 48412 18352
rect 40819 18312 48412 18340
rect 40819 18309 40831 18312
rect 40773 18303 40831 18309
rect 48406 18300 48412 18312
rect 48464 18300 48470 18352
rect 36265 18275 36323 18281
rect 36265 18241 36277 18275
rect 36311 18272 36323 18275
rect 37274 18272 37280 18284
rect 36311 18244 37280 18272
rect 36311 18241 36323 18244
rect 36265 18235 36323 18241
rect 37274 18232 37280 18244
rect 37332 18232 37338 18284
rect 37553 18275 37611 18281
rect 37553 18241 37565 18275
rect 37599 18272 37611 18275
rect 37918 18272 37924 18284
rect 37599 18244 37924 18272
rect 37599 18241 37611 18244
rect 37553 18235 37611 18241
rect 37918 18232 37924 18244
rect 37976 18232 37982 18284
rect 39666 18232 39672 18284
rect 39724 18272 39730 18284
rect 41690 18272 41696 18284
rect 39724 18244 41696 18272
rect 39724 18232 39730 18244
rect 33928 18176 36216 18204
rect 36541 18207 36599 18213
rect 33928 18164 33934 18176
rect 36541 18173 36553 18207
rect 36587 18204 36599 18207
rect 36814 18204 36820 18216
rect 36587 18176 36820 18204
rect 36587 18173 36599 18176
rect 36541 18167 36599 18173
rect 36814 18164 36820 18176
rect 36872 18164 36878 18216
rect 36906 18164 36912 18216
rect 36964 18164 36970 18216
rect 37369 18207 37427 18213
rect 37369 18173 37381 18207
rect 37415 18204 37427 18207
rect 37734 18204 37740 18216
rect 37415 18176 37740 18204
rect 37415 18173 37427 18176
rect 37369 18167 37427 18173
rect 37734 18164 37740 18176
rect 37792 18164 37798 18216
rect 38013 18207 38071 18213
rect 38013 18173 38025 18207
rect 38059 18173 38071 18207
rect 38013 18167 38071 18173
rect 32548 18108 33640 18136
rect 32548 18096 32554 18108
rect 35710 18096 35716 18148
rect 35768 18136 35774 18148
rect 37826 18136 37832 18148
rect 35768 18108 37832 18136
rect 35768 18096 35774 18108
rect 37826 18096 37832 18108
rect 37884 18136 37890 18148
rect 38028 18136 38056 18167
rect 38286 18164 38292 18216
rect 38344 18164 38350 18216
rect 38378 18164 38384 18216
rect 38436 18204 38442 18216
rect 40972 18213 41000 18244
rect 41690 18232 41696 18244
rect 41748 18232 41754 18284
rect 41785 18275 41843 18281
rect 41785 18241 41797 18275
rect 41831 18272 41843 18275
rect 41874 18272 41880 18284
rect 41831 18244 41880 18272
rect 41831 18241 41843 18244
rect 41785 18235 41843 18241
rect 41874 18232 41880 18244
rect 41932 18232 41938 18284
rect 42613 18275 42671 18281
rect 42613 18241 42625 18275
rect 42659 18241 42671 18275
rect 42613 18235 42671 18241
rect 48593 18275 48651 18281
rect 48593 18241 48605 18275
rect 48639 18272 48651 18275
rect 49050 18272 49056 18284
rect 48639 18244 49056 18272
rect 48639 18241 48651 18244
rect 48593 18235 48651 18241
rect 40957 18207 41015 18213
rect 38436 18176 40448 18204
rect 38436 18164 38442 18176
rect 40420 18145 40448 18176
rect 40957 18173 40969 18207
rect 41003 18173 41015 18207
rect 40957 18167 41015 18173
rect 41046 18164 41052 18216
rect 41104 18204 41110 18216
rect 42628 18204 42656 18235
rect 49050 18232 49056 18244
rect 49108 18232 49114 18284
rect 41104 18176 42656 18204
rect 41104 18164 41110 18176
rect 37884 18108 38056 18136
rect 40405 18139 40463 18145
rect 37884 18096 37890 18108
rect 40405 18105 40417 18139
rect 40451 18105 40463 18139
rect 40405 18099 40463 18105
rect 41598 18096 41604 18148
rect 41656 18096 41662 18148
rect 23256 18040 24992 18068
rect 23256 18028 23262 18040
rect 25038 18028 25044 18080
rect 25096 18068 25102 18080
rect 25869 18071 25927 18077
rect 25869 18068 25881 18071
rect 25096 18040 25881 18068
rect 25096 18028 25102 18040
rect 25869 18037 25881 18040
rect 25915 18037 25927 18071
rect 25869 18031 25927 18037
rect 27154 18028 27160 18080
rect 27212 18028 27218 18080
rect 27614 18028 27620 18080
rect 27672 18068 27678 18080
rect 28353 18071 28411 18077
rect 28353 18068 28365 18071
rect 27672 18040 28365 18068
rect 27672 18028 27678 18040
rect 28353 18037 28365 18040
rect 28399 18037 28411 18071
rect 28353 18031 28411 18037
rect 28626 18028 28632 18080
rect 28684 18068 28690 18080
rect 29086 18068 29092 18080
rect 28684 18040 29092 18068
rect 28684 18028 28690 18040
rect 29086 18028 29092 18040
rect 29144 18028 29150 18080
rect 29733 18071 29791 18077
rect 29733 18037 29745 18071
rect 29779 18068 29791 18071
rect 30926 18068 30932 18080
rect 29779 18040 30932 18068
rect 29779 18037 29791 18040
rect 29733 18031 29791 18037
rect 30926 18028 30932 18040
rect 30984 18028 30990 18080
rect 31570 18028 31576 18080
rect 31628 18028 31634 18080
rect 32309 18071 32367 18077
rect 32309 18037 32321 18071
rect 32355 18068 32367 18071
rect 34514 18068 34520 18080
rect 32355 18040 34520 18068
rect 32355 18037 32367 18040
rect 32309 18031 32367 18037
rect 34514 18028 34520 18040
rect 34572 18028 34578 18080
rect 35342 18028 35348 18080
rect 35400 18068 35406 18080
rect 37182 18068 37188 18080
rect 35400 18040 37188 18068
rect 35400 18028 35406 18040
rect 37182 18028 37188 18040
rect 37240 18028 37246 18080
rect 37458 18028 37464 18080
rect 37516 18068 37522 18080
rect 37737 18071 37795 18077
rect 37737 18068 37749 18071
rect 37516 18040 37749 18068
rect 37516 18028 37522 18040
rect 37737 18037 37749 18040
rect 37783 18068 37795 18071
rect 38838 18068 38844 18080
rect 37783 18040 38844 18068
rect 37783 18037 37795 18040
rect 37737 18031 37795 18037
rect 38838 18028 38844 18040
rect 38896 18068 38902 18080
rect 40037 18071 40095 18077
rect 40037 18068 40049 18071
rect 38896 18040 40049 18068
rect 38896 18028 38902 18040
rect 40037 18037 40049 18040
rect 40083 18068 40095 18071
rect 41506 18068 41512 18080
rect 40083 18040 41512 18068
rect 40083 18037 40095 18040
rect 40037 18031 40095 18037
rect 41506 18028 41512 18040
rect 41564 18028 41570 18080
rect 43257 18071 43315 18077
rect 43257 18037 43269 18071
rect 43303 18068 43315 18071
rect 43346 18068 43352 18080
rect 43303 18040 43352 18068
rect 43303 18037 43315 18040
rect 43257 18031 43315 18037
rect 43346 18028 43352 18040
rect 43404 18028 43410 18080
rect 48314 18028 48320 18080
rect 48372 18068 48378 18080
rect 49237 18071 49295 18077
rect 49237 18068 49249 18071
rect 48372 18040 49249 18068
rect 48372 18028 48378 18040
rect 49237 18037 49249 18040
rect 49283 18037 49295 18071
rect 49237 18031 49295 18037
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 8386 17824 8392 17876
rect 8444 17824 8450 17876
rect 9217 17867 9275 17873
rect 9217 17833 9229 17867
rect 9263 17864 9275 17867
rect 11146 17864 11152 17876
rect 9263 17836 11152 17864
rect 9263 17833 9275 17836
rect 9217 17827 9275 17833
rect 11146 17824 11152 17836
rect 11204 17824 11210 17876
rect 11422 17824 11428 17876
rect 11480 17864 11486 17876
rect 13633 17867 13691 17873
rect 13633 17864 13645 17867
rect 11480 17836 13645 17864
rect 11480 17824 11486 17836
rect 13633 17833 13645 17836
rect 13679 17833 13691 17867
rect 13633 17827 13691 17833
rect 14918 17824 14924 17876
rect 14976 17864 14982 17876
rect 14976 17836 15976 17864
rect 14976 17824 14982 17836
rect 1762 17756 1768 17808
rect 1820 17796 1826 17808
rect 8478 17796 8484 17808
rect 1820 17768 8484 17796
rect 1820 17756 1826 17768
rect 8478 17756 8484 17768
rect 8536 17756 8542 17808
rect 8846 17756 8852 17808
rect 8904 17796 8910 17808
rect 9950 17796 9956 17808
rect 8904 17768 9956 17796
rect 8904 17756 8910 17768
rect 9950 17756 9956 17768
rect 10008 17756 10014 17808
rect 13173 17799 13231 17805
rect 13173 17765 13185 17799
rect 13219 17796 13231 17799
rect 13354 17796 13360 17808
rect 13219 17768 13360 17796
rect 13219 17765 13231 17768
rect 13173 17759 13231 17765
rect 13354 17756 13360 17768
rect 13412 17756 13418 17808
rect 15948 17796 15976 17836
rect 16022 17824 16028 17876
rect 16080 17824 16086 17876
rect 17497 17867 17555 17873
rect 17497 17833 17509 17867
rect 17543 17864 17555 17867
rect 19886 17864 19892 17876
rect 17543 17836 19892 17864
rect 17543 17833 17555 17836
rect 17497 17827 17555 17833
rect 19886 17824 19892 17836
rect 19944 17824 19950 17876
rect 20254 17824 20260 17876
rect 20312 17864 20318 17876
rect 24486 17864 24492 17876
rect 20312 17836 24492 17864
rect 20312 17824 20318 17836
rect 24486 17824 24492 17836
rect 24544 17824 24550 17876
rect 24578 17824 24584 17876
rect 24636 17824 24642 17876
rect 25777 17867 25835 17873
rect 25777 17864 25789 17867
rect 24688 17836 25789 17864
rect 19429 17799 19487 17805
rect 19429 17796 19441 17799
rect 15948 17768 19441 17796
rect 19429 17765 19441 17768
rect 19475 17765 19487 17799
rect 19429 17759 19487 17765
rect 22830 17756 22836 17808
rect 22888 17796 22894 17808
rect 24688 17796 24716 17836
rect 25777 17833 25789 17836
rect 25823 17833 25835 17867
rect 25777 17827 25835 17833
rect 27328 17867 27386 17873
rect 27328 17833 27340 17867
rect 27374 17864 27386 17867
rect 30282 17864 30288 17876
rect 27374 17836 30288 17864
rect 27374 17833 27386 17836
rect 27328 17827 27386 17833
rect 30282 17824 30288 17836
rect 30340 17824 30346 17876
rect 30374 17824 30380 17876
rect 30432 17864 30438 17876
rect 30834 17864 30840 17876
rect 30432 17836 30840 17864
rect 30432 17824 30438 17836
rect 30834 17824 30840 17836
rect 30892 17864 30898 17876
rect 31938 17864 31944 17876
rect 30892 17836 31944 17864
rect 30892 17824 30898 17836
rect 31938 17824 31944 17836
rect 31996 17824 32002 17876
rect 32582 17824 32588 17876
rect 32640 17864 32646 17876
rect 32858 17864 32864 17876
rect 32640 17836 32864 17864
rect 32640 17824 32646 17836
rect 32858 17824 32864 17836
rect 32916 17824 32922 17876
rect 33778 17824 33784 17876
rect 33836 17824 33842 17876
rect 34698 17824 34704 17876
rect 34756 17864 34762 17876
rect 34756 17836 38148 17864
rect 34756 17824 34762 17836
rect 22888 17768 24716 17796
rect 22888 17756 22894 17768
rect 24762 17756 24768 17808
rect 24820 17796 24826 17808
rect 24820 17768 25176 17796
rect 24820 17756 24826 17768
rect 1210 17688 1216 17740
rect 1268 17728 1274 17740
rect 2041 17731 2099 17737
rect 2041 17728 2053 17731
rect 1268 17700 2053 17728
rect 1268 17688 1274 17700
rect 2041 17697 2053 17700
rect 2087 17697 2099 17731
rect 2041 17691 2099 17697
rect 3326 17688 3332 17740
rect 3384 17728 3390 17740
rect 4433 17731 4491 17737
rect 4433 17728 4445 17731
rect 3384 17700 4445 17728
rect 3384 17688 3390 17700
rect 4433 17697 4445 17700
rect 4479 17697 4491 17731
rect 4433 17691 4491 17697
rect 5813 17731 5871 17737
rect 5813 17697 5825 17731
rect 5859 17728 5871 17731
rect 7006 17728 7012 17740
rect 5859 17700 7012 17728
rect 5859 17697 5871 17700
rect 5813 17691 5871 17697
rect 7006 17688 7012 17700
rect 7064 17688 7070 17740
rect 7300 17700 10456 17728
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17629 1823 17663
rect 1765 17623 1823 17629
rect 4157 17663 4215 17669
rect 4157 17629 4169 17663
rect 4203 17660 4215 17663
rect 4338 17660 4344 17672
rect 4203 17632 4344 17660
rect 4203 17629 4215 17632
rect 4157 17623 4215 17629
rect 1780 17592 1808 17623
rect 4338 17620 4344 17632
rect 4396 17620 4402 17672
rect 4890 17620 4896 17672
rect 4948 17660 4954 17672
rect 7300 17669 7328 17700
rect 6089 17663 6147 17669
rect 6089 17660 6101 17663
rect 4948 17632 6101 17660
rect 4948 17620 4954 17632
rect 6089 17629 6101 17632
rect 6135 17629 6147 17663
rect 6089 17623 6147 17629
rect 7285 17663 7343 17669
rect 7285 17629 7297 17663
rect 7331 17629 7343 17663
rect 7285 17623 7343 17629
rect 8570 17620 8576 17672
rect 8628 17620 8634 17672
rect 9398 17620 9404 17672
rect 9456 17620 9462 17672
rect 7745 17595 7803 17601
rect 1780 17564 7236 17592
rect 4982 17484 4988 17536
rect 5040 17524 5046 17536
rect 7101 17527 7159 17533
rect 7101 17524 7113 17527
rect 5040 17496 7113 17524
rect 5040 17484 5046 17496
rect 7101 17493 7113 17496
rect 7147 17493 7159 17527
rect 7208 17524 7236 17564
rect 7745 17561 7757 17595
rect 7791 17592 7803 17595
rect 10229 17595 10287 17601
rect 10229 17592 10241 17595
rect 7791 17564 10241 17592
rect 7791 17561 7803 17564
rect 7745 17555 7803 17561
rect 10229 17561 10241 17564
rect 10275 17561 10287 17595
rect 10229 17555 10287 17561
rect 9674 17524 9680 17536
rect 7208 17496 9680 17524
rect 7101 17487 7159 17493
rect 9674 17484 9680 17496
rect 9732 17484 9738 17536
rect 9858 17484 9864 17536
rect 9916 17484 9922 17536
rect 10318 17484 10324 17536
rect 10376 17484 10382 17536
rect 10428 17524 10456 17700
rect 10502 17688 10508 17740
rect 10560 17688 10566 17740
rect 12342 17728 12348 17740
rect 11072 17700 12348 17728
rect 10778 17620 10784 17672
rect 10836 17660 10842 17672
rect 11072 17669 11100 17700
rect 12342 17688 12348 17700
rect 12400 17728 12406 17740
rect 12710 17728 12716 17740
rect 12400 17700 12716 17728
rect 12400 17688 12406 17700
rect 12710 17688 12716 17700
rect 12768 17688 12774 17740
rect 14274 17688 14280 17740
rect 14332 17728 14338 17740
rect 15102 17728 15108 17740
rect 14332 17700 15108 17728
rect 14332 17688 14338 17700
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 15194 17688 15200 17740
rect 15252 17728 15258 17740
rect 16666 17728 16672 17740
rect 15252 17700 16672 17728
rect 15252 17688 15258 17700
rect 16666 17688 16672 17700
rect 16724 17688 16730 17740
rect 16776 17700 18000 17728
rect 11057 17663 11115 17669
rect 11057 17660 11069 17663
rect 10836 17632 11069 17660
rect 10836 17620 10842 17632
rect 11057 17629 11069 17632
rect 11103 17629 11115 17663
rect 11057 17623 11115 17629
rect 12434 17620 12440 17672
rect 12492 17620 12498 17672
rect 13538 17620 13544 17672
rect 13596 17620 13602 17672
rect 15838 17660 15844 17672
rect 15686 17632 15844 17660
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 11330 17552 11336 17604
rect 11388 17552 11394 17604
rect 14550 17552 14556 17604
rect 14608 17552 14614 17604
rect 16776 17592 16804 17700
rect 16853 17663 16911 17669
rect 16853 17629 16865 17663
rect 16899 17660 16911 17663
rect 17862 17660 17868 17672
rect 16899 17632 17868 17660
rect 16899 17629 16911 17632
rect 16853 17623 16911 17629
rect 17862 17620 17868 17632
rect 17920 17620 17926 17672
rect 17972 17660 18000 17700
rect 18322 17688 18328 17740
rect 18380 17728 18386 17740
rect 18506 17728 18512 17740
rect 18380 17700 18512 17728
rect 18380 17688 18386 17700
rect 18506 17688 18512 17700
rect 18564 17688 18570 17740
rect 18598 17688 18604 17740
rect 18656 17728 18662 17740
rect 18693 17731 18751 17737
rect 18693 17728 18705 17731
rect 18656 17700 18705 17728
rect 18656 17688 18662 17700
rect 18693 17697 18705 17700
rect 18739 17697 18751 17731
rect 18693 17691 18751 17697
rect 19334 17688 19340 17740
rect 19392 17728 19398 17740
rect 20165 17731 20223 17737
rect 20165 17728 20177 17731
rect 19392 17700 20177 17728
rect 19392 17688 19398 17700
rect 20165 17697 20177 17700
rect 20211 17728 20223 17731
rect 20438 17728 20444 17740
rect 20211 17700 20444 17728
rect 20211 17697 20223 17700
rect 20165 17691 20223 17697
rect 20438 17688 20444 17700
rect 20496 17728 20502 17740
rect 21082 17728 21088 17740
rect 20496 17700 21088 17728
rect 20496 17688 20502 17700
rect 21082 17688 21088 17700
rect 21140 17728 21146 17740
rect 22278 17728 22284 17740
rect 21140 17700 22284 17728
rect 21140 17688 21146 17700
rect 22278 17688 22284 17700
rect 22336 17728 22342 17740
rect 23201 17731 23259 17737
rect 23201 17728 23213 17731
rect 22336 17700 23213 17728
rect 22336 17688 22342 17700
rect 23201 17697 23213 17700
rect 23247 17697 23259 17731
rect 23201 17691 23259 17697
rect 25038 17688 25044 17740
rect 25096 17688 25102 17740
rect 25148 17737 25176 17768
rect 28810 17756 28816 17808
rect 28868 17796 28874 17808
rect 28994 17796 29000 17808
rect 28868 17768 29000 17796
rect 28868 17756 28874 17768
rect 28994 17756 29000 17768
rect 29052 17756 29058 17808
rect 31297 17799 31355 17805
rect 31297 17765 31309 17799
rect 31343 17796 31355 17799
rect 33962 17796 33968 17808
rect 31343 17768 33968 17796
rect 31343 17765 31355 17768
rect 31297 17759 31355 17765
rect 33962 17756 33968 17768
rect 34020 17756 34026 17808
rect 37366 17756 37372 17808
rect 37424 17796 37430 17808
rect 37553 17799 37611 17805
rect 37553 17796 37565 17799
rect 37424 17768 37565 17796
rect 37424 17756 37430 17768
rect 37553 17765 37565 17768
rect 37599 17765 37611 17799
rect 37553 17759 37611 17765
rect 38013 17799 38071 17805
rect 38013 17765 38025 17799
rect 38059 17765 38071 17799
rect 38013 17759 38071 17765
rect 25133 17731 25191 17737
rect 25133 17697 25145 17731
rect 25179 17697 25191 17731
rect 25133 17691 25191 17697
rect 25590 17688 25596 17740
rect 25648 17728 25654 17740
rect 26329 17731 26387 17737
rect 26329 17728 26341 17731
rect 25648 17700 26341 17728
rect 25648 17688 25654 17700
rect 26329 17697 26341 17700
rect 26375 17697 26387 17731
rect 26329 17691 26387 17697
rect 26602 17688 26608 17740
rect 26660 17728 26666 17740
rect 27065 17731 27123 17737
rect 26660 17700 26924 17728
rect 26660 17688 26666 17700
rect 19518 17660 19524 17672
rect 17972 17632 19524 17660
rect 19518 17620 19524 17632
rect 19576 17620 19582 17672
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17629 19671 17663
rect 19613 17623 19671 17629
rect 15856 17564 16804 17592
rect 17957 17595 18015 17601
rect 11514 17524 11520 17536
rect 10428 17496 11520 17524
rect 11514 17484 11520 17496
rect 11572 17484 11578 17536
rect 11698 17484 11704 17536
rect 11756 17524 11762 17536
rect 12250 17524 12256 17536
rect 11756 17496 12256 17524
rect 11756 17484 11762 17496
rect 12250 17484 12256 17496
rect 12308 17524 12314 17536
rect 12805 17527 12863 17533
rect 12805 17524 12817 17527
rect 12308 17496 12817 17524
rect 12308 17484 12314 17496
rect 12805 17493 12817 17496
rect 12851 17493 12863 17527
rect 12805 17487 12863 17493
rect 13446 17484 13452 17536
rect 13504 17524 13510 17536
rect 14366 17524 14372 17536
rect 13504 17496 14372 17524
rect 13504 17484 13510 17496
rect 14366 17484 14372 17496
rect 14424 17524 14430 17536
rect 15856 17524 15884 17564
rect 17957 17561 17969 17595
rect 18003 17592 18015 17595
rect 18322 17592 18328 17604
rect 18003 17564 18328 17592
rect 18003 17561 18015 17564
rect 17957 17555 18015 17561
rect 18322 17552 18328 17564
rect 18380 17552 18386 17604
rect 14424 17496 15884 17524
rect 14424 17484 14430 17496
rect 15930 17484 15936 17536
rect 15988 17524 15994 17536
rect 16393 17527 16451 17533
rect 16393 17524 16405 17527
rect 15988 17496 16405 17524
rect 15988 17484 15994 17496
rect 16393 17493 16405 17496
rect 16439 17493 16451 17527
rect 16393 17487 16451 17493
rect 16574 17484 16580 17536
rect 16632 17524 16638 17536
rect 18966 17524 18972 17536
rect 16632 17496 18972 17524
rect 16632 17484 16638 17496
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 19628 17524 19656 17623
rect 22002 17620 22008 17672
rect 22060 17660 22066 17672
rect 24946 17660 24952 17672
rect 22060 17632 24952 17660
rect 22060 17620 22066 17632
rect 24946 17620 24952 17632
rect 25004 17660 25010 17672
rect 25222 17660 25228 17672
rect 25004 17632 25228 17660
rect 25004 17620 25010 17632
rect 25222 17620 25228 17632
rect 25280 17620 25286 17672
rect 25774 17620 25780 17672
rect 25832 17660 25838 17672
rect 25832 17632 26832 17660
rect 25832 17620 25838 17632
rect 20346 17552 20352 17604
rect 20404 17592 20410 17604
rect 20441 17595 20499 17601
rect 20441 17592 20453 17595
rect 20404 17564 20453 17592
rect 20404 17552 20410 17564
rect 20441 17561 20453 17564
rect 20487 17561 20499 17595
rect 20441 17555 20499 17561
rect 20898 17552 20904 17604
rect 20956 17552 20962 17604
rect 22465 17595 22523 17601
rect 22465 17561 22477 17595
rect 22511 17592 22523 17595
rect 23290 17592 23296 17604
rect 22511 17564 23296 17592
rect 22511 17561 22523 17564
rect 22465 17555 22523 17561
rect 23290 17552 23296 17564
rect 23348 17552 23354 17604
rect 23845 17595 23903 17601
rect 23845 17561 23857 17595
rect 23891 17592 23903 17595
rect 26145 17595 26203 17601
rect 26145 17592 26157 17595
rect 23891 17564 26157 17592
rect 23891 17561 23903 17564
rect 23845 17555 23903 17561
rect 26145 17561 26157 17564
rect 26191 17561 26203 17595
rect 26145 17555 26203 17561
rect 21358 17524 21364 17536
rect 19628 17496 21364 17524
rect 21358 17484 21364 17496
rect 21416 17484 21422 17536
rect 21910 17484 21916 17536
rect 21968 17484 21974 17536
rect 24949 17527 25007 17533
rect 24949 17493 24961 17527
rect 24995 17524 25007 17527
rect 25038 17524 25044 17536
rect 24995 17496 25044 17524
rect 24995 17493 25007 17496
rect 24949 17487 25007 17493
rect 25038 17484 25044 17496
rect 25096 17484 25102 17536
rect 26050 17484 26056 17536
rect 26108 17524 26114 17536
rect 26237 17527 26295 17533
rect 26237 17524 26249 17527
rect 26108 17496 26249 17524
rect 26108 17484 26114 17496
rect 26237 17493 26249 17496
rect 26283 17493 26295 17527
rect 26804 17524 26832 17632
rect 26896 17592 26924 17700
rect 27065 17697 27077 17731
rect 27111 17728 27123 17731
rect 28350 17728 28356 17740
rect 27111 17700 28356 17728
rect 27111 17697 27123 17700
rect 27065 17691 27123 17697
rect 28350 17688 28356 17700
rect 28408 17728 28414 17740
rect 28408 17700 30696 17728
rect 28408 17688 28414 17700
rect 28810 17620 28816 17672
rect 28868 17660 28874 17672
rect 29089 17663 29147 17669
rect 29089 17660 29101 17663
rect 28868 17632 29101 17660
rect 28868 17620 28874 17632
rect 29089 17629 29101 17632
rect 29135 17629 29147 17663
rect 29089 17623 29147 17629
rect 29825 17663 29883 17669
rect 29825 17629 29837 17663
rect 29871 17660 29883 17663
rect 30374 17660 30380 17672
rect 29871 17632 30380 17660
rect 29871 17629 29883 17632
rect 29825 17623 29883 17629
rect 30374 17620 30380 17632
rect 30432 17620 30438 17672
rect 30668 17601 30696 17700
rect 31662 17688 31668 17740
rect 31720 17728 31726 17740
rect 31849 17731 31907 17737
rect 31849 17728 31861 17731
rect 31720 17700 31861 17728
rect 31720 17688 31726 17700
rect 31849 17697 31861 17700
rect 31895 17697 31907 17731
rect 31849 17691 31907 17697
rect 33226 17688 33232 17740
rect 33284 17688 33290 17740
rect 33413 17731 33471 17737
rect 33413 17697 33425 17731
rect 33459 17728 33471 17731
rect 33686 17728 33692 17740
rect 33459 17700 33692 17728
rect 33459 17697 33471 17700
rect 33413 17691 33471 17697
rect 33686 17688 33692 17700
rect 33744 17728 33750 17740
rect 34054 17728 34060 17740
rect 33744 17700 34060 17728
rect 33744 17688 33750 17700
rect 34054 17688 34060 17700
rect 34112 17688 34118 17740
rect 34606 17728 34612 17740
rect 34164 17700 34612 17728
rect 31018 17620 31024 17672
rect 31076 17660 31082 17672
rect 31757 17663 31815 17669
rect 31757 17660 31769 17663
rect 31076 17632 31769 17660
rect 31076 17620 31082 17632
rect 31757 17629 31769 17632
rect 31803 17629 31815 17663
rect 31757 17623 31815 17629
rect 31938 17620 31944 17672
rect 31996 17660 32002 17672
rect 32401 17663 32459 17669
rect 32401 17660 32413 17663
rect 31996 17632 32413 17660
rect 31996 17620 32002 17632
rect 32401 17629 32413 17632
rect 32447 17660 32459 17663
rect 34164 17660 34192 17700
rect 34606 17688 34612 17700
rect 34664 17688 34670 17740
rect 34882 17688 34888 17740
rect 34940 17728 34946 17740
rect 35710 17728 35716 17740
rect 34940 17700 35716 17728
rect 34940 17688 34946 17700
rect 35710 17688 35716 17700
rect 35768 17728 35774 17740
rect 35805 17731 35863 17737
rect 35805 17728 35817 17731
rect 35768 17700 35817 17728
rect 35768 17688 35774 17700
rect 35805 17697 35817 17700
rect 35851 17697 35863 17731
rect 35805 17691 35863 17697
rect 36078 17688 36084 17740
rect 36136 17688 36142 17740
rect 36630 17688 36636 17740
rect 36688 17728 36694 17740
rect 36688 17700 37228 17728
rect 36688 17688 36694 17700
rect 37200 17672 37228 17700
rect 35618 17660 35624 17672
rect 32447 17632 34192 17660
rect 34348 17632 35624 17660
rect 32447 17629 32459 17632
rect 32401 17623 32459 17629
rect 30653 17595 30711 17601
rect 26896 17564 27830 17592
rect 30653 17561 30665 17595
rect 30699 17592 30711 17595
rect 32490 17592 32496 17604
rect 30699 17564 32496 17592
rect 30699 17561 30711 17564
rect 30653 17555 30711 17561
rect 32490 17552 32496 17564
rect 32548 17552 32554 17604
rect 34348 17592 34376 17632
rect 35618 17620 35624 17632
rect 35676 17620 35682 17672
rect 37182 17620 37188 17672
rect 37240 17660 37246 17672
rect 37458 17660 37464 17672
rect 37240 17632 37464 17660
rect 37240 17620 37246 17632
rect 37458 17620 37464 17632
rect 37516 17620 37522 17672
rect 38028 17660 38056 17759
rect 38120 17728 38148 17836
rect 38562 17824 38568 17876
rect 38620 17864 38626 17876
rect 40497 17867 40555 17873
rect 40497 17864 40509 17867
rect 38620 17836 40509 17864
rect 38620 17824 38626 17836
rect 40497 17833 40509 17836
rect 40543 17833 40555 17867
rect 40497 17827 40555 17833
rect 42334 17824 42340 17876
rect 42392 17824 42398 17876
rect 42610 17824 42616 17876
rect 42668 17824 42674 17876
rect 39758 17756 39764 17808
rect 39816 17796 39822 17808
rect 39816 17768 41414 17796
rect 39816 17756 39822 17768
rect 38473 17731 38531 17737
rect 38473 17728 38485 17731
rect 38120 17700 38485 17728
rect 38473 17697 38485 17700
rect 38519 17697 38531 17731
rect 38473 17691 38531 17697
rect 38562 17688 38568 17740
rect 38620 17688 38626 17740
rect 39206 17688 39212 17740
rect 39264 17688 39270 17740
rect 39942 17688 39948 17740
rect 40000 17728 40006 17740
rect 40957 17731 41015 17737
rect 40957 17728 40969 17731
rect 40000 17700 40969 17728
rect 40000 17688 40006 17700
rect 40957 17697 40969 17700
rect 41003 17697 41015 17731
rect 40957 17691 41015 17697
rect 41049 17731 41107 17737
rect 41049 17697 41061 17731
rect 41095 17697 41107 17731
rect 41049 17691 41107 17697
rect 38028 17632 40448 17660
rect 32692 17564 34376 17592
rect 28813 17527 28871 17533
rect 28813 17524 28825 17527
rect 26804 17496 28825 17524
rect 26237 17487 26295 17493
rect 28813 17493 28825 17496
rect 28859 17524 28871 17527
rect 28902 17524 28908 17536
rect 28859 17496 28908 17524
rect 28859 17493 28871 17496
rect 28813 17487 28871 17493
rect 28902 17484 28908 17496
rect 28960 17484 28966 17536
rect 29270 17484 29276 17536
rect 29328 17484 29334 17536
rect 31665 17527 31723 17533
rect 31665 17493 31677 17527
rect 31711 17524 31723 17527
rect 32692 17524 32720 17564
rect 34514 17552 34520 17604
rect 34572 17592 34578 17604
rect 34885 17595 34943 17601
rect 34885 17592 34897 17595
rect 34572 17564 34897 17592
rect 34572 17552 34578 17564
rect 34885 17561 34897 17564
rect 34931 17561 34943 17595
rect 34885 17555 34943 17561
rect 34974 17552 34980 17604
rect 35032 17592 35038 17604
rect 40310 17592 40316 17604
rect 35032 17564 35480 17592
rect 35032 17552 35038 17564
rect 31711 17496 32720 17524
rect 31711 17493 31723 17496
rect 31665 17487 31723 17493
rect 32766 17484 32772 17536
rect 32824 17484 32830 17536
rect 33137 17527 33195 17533
rect 33137 17493 33149 17527
rect 33183 17524 33195 17527
rect 33778 17524 33784 17536
rect 33183 17496 33784 17524
rect 33183 17493 33195 17496
rect 33137 17487 33195 17493
rect 33778 17484 33784 17496
rect 33836 17484 33842 17536
rect 34149 17527 34207 17533
rect 34149 17493 34161 17527
rect 34195 17524 34207 17527
rect 34698 17524 34704 17536
rect 34195 17496 34704 17524
rect 34195 17493 34207 17496
rect 34149 17487 34207 17493
rect 34698 17484 34704 17496
rect 34756 17484 34762 17536
rect 35342 17484 35348 17536
rect 35400 17484 35406 17536
rect 35452 17524 35480 17564
rect 37384 17564 40316 17592
rect 37384 17524 37412 17564
rect 40310 17552 40316 17564
rect 40368 17552 40374 17604
rect 35452 17496 37412 17524
rect 37826 17484 37832 17536
rect 37884 17524 37890 17536
rect 38381 17527 38439 17533
rect 38381 17524 38393 17527
rect 37884 17496 38393 17524
rect 37884 17484 37890 17496
rect 38381 17493 38393 17496
rect 38427 17493 38439 17527
rect 38381 17487 38439 17493
rect 38838 17484 38844 17536
rect 38896 17524 38902 17536
rect 39853 17527 39911 17533
rect 39853 17524 39865 17527
rect 38896 17496 39865 17524
rect 38896 17484 38902 17496
rect 39853 17493 39865 17496
rect 39899 17493 39911 17527
rect 39853 17487 39911 17493
rect 40129 17527 40187 17533
rect 40129 17493 40141 17527
rect 40175 17524 40187 17527
rect 40218 17524 40224 17536
rect 40175 17496 40224 17524
rect 40175 17493 40187 17496
rect 40129 17487 40187 17493
rect 40218 17484 40224 17496
rect 40276 17484 40282 17536
rect 40420 17524 40448 17632
rect 40586 17620 40592 17672
rect 40644 17660 40650 17672
rect 41064 17660 41092 17691
rect 40644 17632 41092 17660
rect 41386 17660 41414 17768
rect 41874 17756 41880 17808
rect 41932 17796 41938 17808
rect 42797 17799 42855 17805
rect 42797 17796 42809 17799
rect 41932 17768 42809 17796
rect 41932 17756 41938 17768
rect 42797 17765 42809 17768
rect 42843 17765 42855 17799
rect 42797 17759 42855 17765
rect 41693 17663 41751 17669
rect 41693 17660 41705 17663
rect 41386 17632 41705 17660
rect 40644 17620 40650 17632
rect 41693 17629 41705 17632
rect 41739 17629 41751 17663
rect 41693 17623 41751 17629
rect 48593 17663 48651 17669
rect 48593 17629 48605 17663
rect 48639 17660 48651 17663
rect 49050 17660 49056 17672
rect 48639 17632 49056 17660
rect 48639 17629 48651 17632
rect 48593 17623 48651 17629
rect 49050 17620 49056 17632
rect 49108 17620 49114 17672
rect 40865 17595 40923 17601
rect 40865 17561 40877 17595
rect 40911 17592 40923 17595
rect 48406 17592 48412 17604
rect 40911 17564 48412 17592
rect 40911 17561 40923 17564
rect 40865 17555 40923 17561
rect 48406 17552 48412 17564
rect 48464 17552 48470 17604
rect 42058 17524 42064 17536
rect 40420 17496 42064 17524
rect 42058 17484 42064 17496
rect 42116 17484 42122 17536
rect 48777 17527 48835 17533
rect 48777 17493 48789 17527
rect 48823 17524 48835 17527
rect 49142 17524 49148 17536
rect 48823 17496 49148 17524
rect 48823 17493 48835 17496
rect 48777 17487 48835 17493
rect 49142 17484 49148 17496
rect 49200 17484 49206 17536
rect 49234 17484 49240 17536
rect 49292 17484 49298 17536
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 3973 17323 4031 17329
rect 3973 17289 3985 17323
rect 4019 17320 4031 17323
rect 4430 17320 4436 17332
rect 4019 17292 4436 17320
rect 4019 17289 4031 17292
rect 3973 17283 4031 17289
rect 4430 17280 4436 17292
rect 4488 17280 4494 17332
rect 4798 17280 4804 17332
rect 4856 17280 4862 17332
rect 5074 17280 5080 17332
rect 5132 17320 5138 17332
rect 5445 17323 5503 17329
rect 5445 17320 5457 17323
rect 5132 17292 5457 17320
rect 5132 17280 5138 17292
rect 5445 17289 5457 17292
rect 5491 17289 5503 17323
rect 8294 17320 8300 17332
rect 5445 17283 5503 17289
rect 5552 17292 8300 17320
rect 5552 17252 5580 17292
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 8754 17280 8760 17332
rect 8812 17320 8818 17332
rect 9769 17323 9827 17329
rect 9769 17320 9781 17323
rect 8812 17292 9781 17320
rect 8812 17280 8818 17292
rect 9769 17289 9781 17292
rect 9815 17289 9827 17323
rect 9769 17283 9827 17289
rect 9950 17280 9956 17332
rect 10008 17320 10014 17332
rect 10781 17323 10839 17329
rect 10781 17320 10793 17323
rect 10008 17292 10793 17320
rect 10008 17280 10014 17292
rect 10781 17289 10793 17292
rect 10827 17289 10839 17323
rect 10781 17283 10839 17289
rect 12526 17280 12532 17332
rect 12584 17320 12590 17332
rect 13173 17323 13231 17329
rect 13173 17320 13185 17323
rect 12584 17292 13185 17320
rect 12584 17280 12590 17292
rect 13173 17289 13185 17292
rect 13219 17289 13231 17323
rect 13173 17283 13231 17289
rect 13998 17280 14004 17332
rect 14056 17280 14062 17332
rect 15378 17280 15384 17332
rect 15436 17320 15442 17332
rect 17678 17320 17684 17332
rect 15436 17292 17684 17320
rect 15436 17280 15442 17292
rect 17678 17280 17684 17292
rect 17736 17320 17742 17332
rect 18877 17323 18935 17329
rect 18877 17320 18889 17323
rect 17736 17292 18889 17320
rect 17736 17280 17742 17292
rect 18877 17289 18889 17292
rect 18923 17289 18935 17323
rect 18877 17283 18935 17289
rect 18966 17280 18972 17332
rect 19024 17320 19030 17332
rect 24210 17320 24216 17332
rect 19024 17292 24216 17320
rect 19024 17280 19030 17292
rect 24210 17280 24216 17292
rect 24268 17280 24274 17332
rect 24397 17323 24455 17329
rect 24397 17289 24409 17323
rect 24443 17320 24455 17323
rect 24762 17320 24768 17332
rect 24443 17292 24768 17320
rect 24443 17289 24455 17292
rect 24397 17283 24455 17289
rect 24762 17280 24768 17292
rect 24820 17280 24826 17332
rect 24854 17280 24860 17332
rect 24912 17280 24918 17332
rect 25317 17323 25375 17329
rect 25317 17289 25329 17323
rect 25363 17320 25375 17323
rect 27341 17323 27399 17329
rect 27341 17320 27353 17323
rect 25363 17292 27353 17320
rect 25363 17289 25375 17292
rect 25317 17283 25375 17289
rect 27341 17289 27353 17292
rect 27387 17289 27399 17323
rect 27341 17283 27399 17289
rect 27798 17280 27804 17332
rect 27856 17280 27862 17332
rect 29086 17280 29092 17332
rect 29144 17320 29150 17332
rect 29825 17323 29883 17329
rect 29825 17320 29837 17323
rect 29144 17292 29837 17320
rect 29144 17280 29150 17292
rect 29825 17289 29837 17292
rect 29871 17320 29883 17323
rect 29914 17320 29920 17332
rect 29871 17292 29920 17320
rect 29871 17289 29883 17292
rect 29825 17283 29883 17289
rect 29914 17280 29920 17292
rect 29972 17280 29978 17332
rect 30193 17323 30251 17329
rect 30193 17289 30205 17323
rect 30239 17320 30251 17323
rect 32030 17320 32036 17332
rect 30239 17292 32036 17320
rect 30239 17289 30251 17292
rect 30193 17283 30251 17289
rect 32030 17280 32036 17292
rect 32088 17280 32094 17332
rect 32766 17280 32772 17332
rect 32824 17320 32830 17332
rect 36262 17320 36268 17332
rect 32824 17292 36268 17320
rect 32824 17280 32830 17292
rect 36262 17280 36268 17292
rect 36320 17280 36326 17332
rect 37461 17323 37519 17329
rect 37461 17289 37473 17323
rect 37507 17320 37519 17323
rect 37642 17320 37648 17332
rect 37507 17292 37648 17320
rect 37507 17289 37519 17292
rect 37461 17283 37519 17289
rect 37642 17280 37648 17292
rect 37700 17280 37706 17332
rect 37921 17323 37979 17329
rect 37921 17289 37933 17323
rect 37967 17320 37979 17323
rect 38378 17320 38384 17332
rect 37967 17292 38384 17320
rect 37967 17289 37979 17292
rect 37921 17283 37979 17289
rect 38378 17280 38384 17292
rect 38436 17280 38442 17332
rect 41598 17320 41604 17332
rect 41386 17292 41604 17320
rect 9858 17252 9864 17264
rect 1780 17224 5580 17252
rect 8036 17224 9864 17252
rect 1780 17193 1808 17224
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17153 1823 17187
rect 1765 17147 1823 17153
rect 4157 17187 4215 17193
rect 4157 17153 4169 17187
rect 4203 17153 4215 17187
rect 4157 17147 4215 17153
rect 1302 17076 1308 17128
rect 1360 17116 1366 17128
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 1360 17088 2053 17116
rect 1360 17076 1366 17088
rect 2041 17085 2053 17088
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 4172 17048 4200 17147
rect 4982 17144 4988 17196
rect 5040 17144 5046 17196
rect 5626 17144 5632 17196
rect 5684 17144 5690 17196
rect 6546 17144 6552 17196
rect 6604 17144 6610 17196
rect 6825 17187 6883 17193
rect 6825 17153 6837 17187
rect 6871 17184 6883 17187
rect 7098 17184 7104 17196
rect 6871 17156 7104 17184
rect 6871 17153 6883 17156
rect 6825 17147 6883 17153
rect 7098 17144 7104 17156
rect 7156 17144 7162 17196
rect 8036 17193 8064 17224
rect 9858 17212 9864 17224
rect 9916 17212 9922 17264
rect 12434 17212 12440 17264
rect 12492 17252 12498 17264
rect 14016 17252 14044 17280
rect 12492 17224 14044 17252
rect 12492 17212 12498 17224
rect 20162 17212 20168 17264
rect 20220 17212 20226 17264
rect 20898 17212 20904 17264
rect 20956 17252 20962 17264
rect 21361 17255 21419 17261
rect 21361 17252 21373 17255
rect 20956 17224 21373 17252
rect 20956 17212 20962 17224
rect 21361 17221 21373 17224
rect 21407 17221 21419 17255
rect 21361 17215 21419 17221
rect 26510 17212 26516 17264
rect 26568 17212 26574 17264
rect 26789 17255 26847 17261
rect 26789 17221 26801 17255
rect 26835 17252 26847 17255
rect 27062 17252 27068 17264
rect 26835 17224 27068 17252
rect 26835 17221 26847 17224
rect 26789 17215 26847 17221
rect 27062 17212 27068 17224
rect 27120 17212 27126 17264
rect 27982 17212 27988 17264
rect 28040 17252 28046 17264
rect 30098 17252 30104 17264
rect 28040 17224 30104 17252
rect 28040 17212 28046 17224
rect 30098 17212 30104 17224
rect 30156 17212 30162 17264
rect 30742 17212 30748 17264
rect 30800 17252 30806 17264
rect 31849 17255 31907 17261
rect 31849 17252 31861 17255
rect 30800 17224 31861 17252
rect 30800 17212 30806 17224
rect 31849 17221 31861 17224
rect 31895 17221 31907 17255
rect 32490 17252 32496 17264
rect 31849 17215 31907 17221
rect 32324 17224 32496 17252
rect 8021 17187 8079 17193
rect 8021 17153 8033 17187
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 8665 17187 8723 17193
rect 8665 17153 8677 17187
rect 8711 17153 8723 17187
rect 8665 17147 8723 17153
rect 6638 17076 6644 17128
rect 6696 17116 6702 17128
rect 8680 17116 8708 17147
rect 9306 17144 9312 17196
rect 9364 17144 9370 17196
rect 9950 17144 9956 17196
rect 10008 17144 10014 17196
rect 11422 17144 11428 17196
rect 11480 17184 11486 17196
rect 11793 17187 11851 17193
rect 11793 17184 11805 17187
rect 11480 17156 11805 17184
rect 11480 17144 11486 17156
rect 11793 17153 11805 17156
rect 11839 17184 11851 17187
rect 12158 17184 12164 17196
rect 11839 17156 12164 17184
rect 11839 17153 11851 17156
rect 11793 17147 11851 17153
rect 12158 17144 12164 17156
rect 12216 17144 12222 17196
rect 12618 17144 12624 17196
rect 12676 17184 12682 17196
rect 13081 17187 13139 17193
rect 13081 17184 13093 17187
rect 12676 17156 13093 17184
rect 12676 17144 12682 17156
rect 13081 17153 13093 17156
rect 13127 17153 13139 17187
rect 13081 17147 13139 17153
rect 14461 17187 14519 17193
rect 14461 17153 14473 17187
rect 14507 17184 14519 17187
rect 15378 17184 15384 17196
rect 14507 17156 15384 17184
rect 14507 17153 14519 17156
rect 14461 17147 14519 17153
rect 15378 17144 15384 17156
rect 15436 17144 15442 17196
rect 15933 17187 15991 17193
rect 15933 17153 15945 17187
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 16025 17187 16083 17193
rect 16025 17153 16037 17187
rect 16071 17184 16083 17187
rect 16574 17184 16580 17196
rect 16071 17156 16580 17184
rect 16071 17153 16083 17156
rect 16025 17147 16083 17153
rect 10594 17116 10600 17128
rect 6696 17088 8616 17116
rect 8680 17088 10600 17116
rect 6696 17076 6702 17088
rect 7837 17051 7895 17057
rect 7837 17048 7849 17051
rect 4172 17020 7849 17048
rect 7837 17017 7849 17020
rect 7883 17017 7895 17051
rect 7837 17011 7895 17017
rect 4154 16940 4160 16992
rect 4212 16980 4218 16992
rect 8018 16980 8024 16992
rect 4212 16952 8024 16980
rect 4212 16940 4218 16952
rect 8018 16940 8024 16952
rect 8076 16980 8082 16992
rect 8481 16983 8539 16989
rect 8481 16980 8493 16983
rect 8076 16952 8493 16980
rect 8076 16940 8082 16952
rect 8481 16949 8493 16952
rect 8527 16949 8539 16983
rect 8588 16980 8616 17088
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 10870 17076 10876 17128
rect 10928 17076 10934 17128
rect 10965 17119 11023 17125
rect 10965 17085 10977 17119
rect 11011 17116 11023 17119
rect 13265 17119 13323 17125
rect 13265 17116 13277 17119
rect 11011 17088 13277 17116
rect 11011 17085 11023 17088
rect 10965 17079 11023 17085
rect 13265 17085 13277 17088
rect 13311 17085 13323 17119
rect 13265 17079 13323 17085
rect 13817 17119 13875 17125
rect 13817 17085 13829 17119
rect 13863 17116 13875 17119
rect 15470 17116 15476 17128
rect 13863 17088 15476 17116
rect 13863 17085 13875 17088
rect 13817 17079 13875 17085
rect 9122 17008 9128 17060
rect 9180 17008 9186 17060
rect 10413 17051 10471 17057
rect 10413 17017 10425 17051
rect 10459 17048 10471 17051
rect 12158 17048 12164 17060
rect 10459 17020 12164 17048
rect 10459 17017 10471 17020
rect 10413 17011 10471 17017
rect 12158 17008 12164 17020
rect 12216 17008 12222 17060
rect 12434 17008 12440 17060
rect 12492 17048 12498 17060
rect 13280 17048 13308 17079
rect 15470 17076 15476 17088
rect 15528 17116 15534 17128
rect 15948 17116 15976 17147
rect 16574 17144 16580 17156
rect 16632 17144 16638 17196
rect 18506 17144 18512 17196
rect 18564 17144 18570 17196
rect 19334 17144 19340 17196
rect 19392 17144 19398 17196
rect 21637 17187 21695 17193
rect 21637 17153 21649 17187
rect 21683 17184 21695 17187
rect 22186 17184 22192 17196
rect 21683 17156 22192 17184
rect 21683 17153 21695 17156
rect 21637 17147 21695 17153
rect 22186 17144 22192 17156
rect 22244 17144 22250 17196
rect 22278 17144 22284 17196
rect 22336 17184 22342 17196
rect 22649 17187 22707 17193
rect 22649 17184 22661 17187
rect 22336 17156 22661 17184
rect 22336 17144 22342 17156
rect 22649 17153 22661 17156
rect 22695 17153 22707 17187
rect 22649 17147 22707 17153
rect 24026 17144 24032 17196
rect 24084 17144 24090 17196
rect 24946 17144 24952 17196
rect 25004 17184 25010 17196
rect 25225 17187 25283 17193
rect 25225 17184 25237 17187
rect 25004 17156 25237 17184
rect 25004 17144 25010 17156
rect 25225 17153 25237 17156
rect 25271 17153 25283 17187
rect 25225 17147 25283 17153
rect 26237 17187 26295 17193
rect 26237 17153 26249 17187
rect 26283 17153 26295 17187
rect 26237 17147 26295 17153
rect 27709 17188 27767 17193
rect 27798 17188 27804 17196
rect 27709 17187 27804 17188
rect 27709 17153 27721 17187
rect 27755 17160 27804 17187
rect 27755 17153 27767 17160
rect 27709 17147 27767 17153
rect 15528 17088 15976 17116
rect 15528 17076 15534 17088
rect 16114 17076 16120 17128
rect 16172 17076 16178 17128
rect 17129 17119 17187 17125
rect 17129 17085 17141 17119
rect 17175 17085 17187 17119
rect 17129 17079 17187 17085
rect 14185 17051 14243 17057
rect 12492 17020 13216 17048
rect 13280 17020 14136 17048
rect 12492 17008 12498 17020
rect 11885 16983 11943 16989
rect 11885 16980 11897 16983
rect 8588 16952 11897 16980
rect 8481 16943 8539 16949
rect 11885 16949 11897 16952
rect 11931 16949 11943 16983
rect 11885 16943 11943 16949
rect 12526 16940 12532 16992
rect 12584 16980 12590 16992
rect 12713 16983 12771 16989
rect 12713 16980 12725 16983
rect 12584 16952 12725 16980
rect 12584 16940 12590 16952
rect 12713 16949 12725 16952
rect 12759 16949 12771 16983
rect 13188 16980 13216 17020
rect 13446 16980 13452 16992
rect 13188 16952 13452 16980
rect 12713 16943 12771 16949
rect 13446 16940 13452 16952
rect 13504 16940 13510 16992
rect 14108 16980 14136 17020
rect 14185 17017 14197 17051
rect 14231 17048 14243 17051
rect 14826 17048 14832 17060
rect 14231 17020 14832 17048
rect 14231 17017 14243 17020
rect 14185 17011 14243 17017
rect 14826 17008 14832 17020
rect 14884 17048 14890 17060
rect 14884 17020 15240 17048
rect 14884 17008 14890 17020
rect 14734 16980 14740 16992
rect 14108 16952 14740 16980
rect 14734 16940 14740 16952
rect 14792 16940 14798 16992
rect 15010 16940 15016 16992
rect 15068 16980 15074 16992
rect 15105 16983 15163 16989
rect 15105 16980 15117 16983
rect 15068 16952 15117 16980
rect 15068 16940 15074 16952
rect 15105 16949 15117 16952
rect 15151 16949 15163 16983
rect 15212 16980 15240 17020
rect 15562 17008 15568 17060
rect 15620 17008 15626 17060
rect 17034 17048 17040 17060
rect 15672 17020 17040 17048
rect 15672 16980 15700 17020
rect 17034 17008 17040 17020
rect 17092 17008 17098 17060
rect 15212 16952 15700 16980
rect 16761 16983 16819 16989
rect 15105 16943 15163 16949
rect 16761 16949 16773 16983
rect 16807 16980 16819 16983
rect 16942 16980 16948 16992
rect 16807 16952 16948 16980
rect 16807 16949 16819 16952
rect 16761 16943 16819 16949
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17144 16980 17172 17079
rect 17402 17076 17408 17128
rect 17460 17076 17466 17128
rect 17862 17076 17868 17128
rect 17920 17116 17926 17128
rect 19613 17119 19671 17125
rect 17920 17088 19472 17116
rect 17920 17076 17926 17088
rect 18598 16980 18604 16992
rect 17144 16952 18604 16980
rect 18598 16940 18604 16952
rect 18656 16940 18662 16992
rect 19444 16980 19472 17088
rect 19613 17085 19625 17119
rect 19659 17116 19671 17119
rect 20070 17116 20076 17128
rect 19659 17088 20076 17116
rect 19659 17085 19671 17088
rect 19613 17079 19671 17085
rect 20070 17076 20076 17088
rect 20128 17076 20134 17128
rect 22370 17076 22376 17128
rect 22428 17116 22434 17128
rect 22925 17119 22983 17125
rect 22925 17116 22937 17119
rect 22428 17088 22937 17116
rect 22428 17076 22434 17088
rect 22925 17085 22937 17088
rect 22971 17085 22983 17119
rect 22925 17079 22983 17085
rect 25498 17076 25504 17128
rect 25556 17076 25562 17128
rect 26252 17116 26280 17147
rect 27798 17144 27804 17160
rect 27856 17144 27862 17196
rect 28997 17187 29055 17193
rect 28997 17153 29009 17187
rect 29043 17184 29055 17187
rect 29362 17184 29368 17196
rect 29043 17156 29368 17184
rect 29043 17153 29055 17156
rect 28997 17147 29055 17153
rect 29362 17144 29368 17156
rect 29420 17144 29426 17196
rect 32324 17193 32352 17224
rect 32490 17212 32496 17224
rect 32548 17212 32554 17264
rect 32582 17212 32588 17264
rect 32640 17212 32646 17264
rect 34146 17252 34152 17264
rect 33810 17224 34152 17252
rect 34146 17212 34152 17224
rect 34204 17212 34210 17264
rect 35802 17212 35808 17264
rect 35860 17252 35866 17264
rect 41386 17252 41414 17292
rect 41598 17280 41604 17292
rect 41656 17320 41662 17332
rect 42061 17323 42119 17329
rect 42061 17320 42073 17323
rect 41656 17292 42073 17320
rect 41656 17280 41662 17292
rect 42061 17289 42073 17292
rect 42107 17320 42119 17323
rect 42610 17320 42616 17332
rect 42107 17292 42616 17320
rect 42107 17289 42119 17292
rect 42061 17283 42119 17289
rect 42610 17280 42616 17292
rect 42668 17280 42674 17332
rect 48406 17280 48412 17332
rect 48464 17280 48470 17332
rect 35860 17224 36492 17252
rect 40342 17224 41414 17252
rect 35860 17212 35866 17224
rect 30561 17187 30619 17193
rect 30561 17153 30573 17187
rect 30607 17184 30619 17187
rect 31389 17187 31447 17193
rect 31389 17184 31401 17187
rect 30607 17156 31401 17184
rect 30607 17153 30619 17156
rect 30561 17147 30619 17153
rect 31389 17153 31401 17156
rect 31435 17153 31447 17187
rect 31389 17147 31447 17153
rect 32309 17187 32367 17193
rect 32309 17153 32321 17187
rect 32355 17153 32367 17187
rect 32309 17147 32367 17153
rect 34606 17144 34612 17196
rect 34664 17144 34670 17196
rect 36354 17144 36360 17196
rect 36412 17144 36418 17196
rect 36464 17184 36492 17224
rect 37829 17187 37887 17193
rect 37829 17184 37841 17187
rect 36464 17156 37841 17184
rect 37829 17153 37841 17156
rect 37875 17153 37887 17187
rect 37829 17147 37887 17153
rect 38378 17144 38384 17196
rect 38436 17184 38442 17196
rect 38562 17184 38568 17196
rect 38436 17156 38568 17184
rect 38436 17144 38442 17156
rect 38562 17144 38568 17156
rect 38620 17144 38626 17196
rect 41046 17144 41052 17196
rect 41104 17144 41110 17196
rect 48593 17187 48651 17193
rect 48593 17153 48605 17187
rect 48639 17184 48651 17187
rect 48774 17184 48780 17196
rect 48639 17156 48780 17184
rect 48639 17153 48651 17156
rect 48593 17147 48651 17153
rect 48774 17144 48780 17156
rect 48832 17144 48838 17196
rect 49145 17187 49203 17193
rect 49145 17153 49157 17187
rect 49191 17184 49203 17187
rect 49234 17184 49240 17196
rect 49191 17156 49240 17184
rect 49191 17153 49203 17156
rect 49145 17147 49203 17153
rect 49234 17144 49240 17156
rect 49292 17144 49298 17196
rect 27985 17119 28043 17125
rect 26252 17088 27568 17116
rect 22002 17008 22008 17060
rect 22060 17008 22066 17060
rect 24486 17008 24492 17060
rect 24544 17048 24550 17060
rect 26053 17051 26111 17057
rect 26053 17048 26065 17051
rect 24544 17020 26065 17048
rect 24544 17008 24550 17020
rect 26053 17017 26065 17020
rect 26099 17017 26111 17051
rect 26053 17011 26111 17017
rect 20162 16980 20168 16992
rect 19444 16952 20168 16980
rect 20162 16940 20168 16952
rect 20220 16980 20226 16992
rect 21085 16983 21143 16989
rect 21085 16980 21097 16983
rect 20220 16952 21097 16980
rect 20220 16940 20226 16952
rect 21085 16949 21097 16952
rect 21131 16949 21143 16983
rect 21085 16943 21143 16949
rect 26602 16940 26608 16992
rect 26660 16980 26666 16992
rect 26973 16983 27031 16989
rect 26973 16980 26985 16983
rect 26660 16952 26985 16980
rect 26660 16940 26666 16952
rect 26973 16949 26985 16952
rect 27019 16949 27031 16983
rect 27540 16980 27568 17088
rect 27985 17085 27997 17119
rect 28031 17085 28043 17119
rect 27985 17079 28043 17085
rect 27890 17008 27896 17060
rect 27948 17048 27954 17060
rect 28000 17048 28028 17079
rect 28074 17076 28080 17128
rect 28132 17116 28138 17128
rect 29086 17116 29092 17128
rect 28132 17088 29092 17116
rect 28132 17076 28138 17088
rect 29086 17076 29092 17088
rect 29144 17076 29150 17128
rect 29273 17119 29331 17125
rect 29273 17085 29285 17119
rect 29319 17116 29331 17119
rect 29638 17116 29644 17128
rect 29319 17088 29644 17116
rect 29319 17085 29331 17088
rect 29273 17079 29331 17085
rect 29638 17076 29644 17088
rect 29696 17076 29702 17128
rect 30653 17119 30711 17125
rect 30653 17085 30665 17119
rect 30699 17116 30711 17119
rect 30742 17116 30748 17128
rect 30699 17088 30748 17116
rect 30699 17085 30711 17088
rect 30653 17079 30711 17085
rect 30742 17076 30748 17088
rect 30800 17076 30806 17128
rect 30837 17119 30895 17125
rect 30837 17085 30849 17119
rect 30883 17085 30895 17119
rect 30837 17079 30895 17085
rect 31726 17088 32444 17116
rect 27948 17020 28028 17048
rect 28629 17051 28687 17057
rect 27948 17008 27954 17020
rect 28629 17017 28641 17051
rect 28675 17048 28687 17051
rect 30852 17048 30880 17079
rect 31726 17048 31754 17088
rect 28675 17020 29132 17048
rect 28675 17017 28687 17020
rect 28629 17011 28687 17017
rect 28994 16980 29000 16992
rect 27540 16952 29000 16980
rect 26973 16943 27031 16949
rect 28994 16940 29000 16952
rect 29052 16940 29058 16992
rect 29104 16980 29132 17020
rect 29288 17020 30788 17048
rect 30852 17020 31754 17048
rect 29288 16980 29316 17020
rect 29104 16952 29316 16980
rect 29454 16940 29460 16992
rect 29512 16980 29518 16992
rect 29733 16983 29791 16989
rect 29733 16980 29745 16983
rect 29512 16952 29745 16980
rect 29512 16940 29518 16952
rect 29733 16949 29745 16952
rect 29779 16980 29791 16983
rect 30558 16980 30564 16992
rect 29779 16952 30564 16980
rect 29779 16949 29791 16952
rect 29733 16943 29791 16949
rect 30558 16940 30564 16952
rect 30616 16940 30622 16992
rect 30760 16980 30788 17020
rect 31202 16980 31208 16992
rect 30760 16952 31208 16980
rect 31202 16940 31208 16952
rect 31260 16940 31266 16992
rect 31386 16940 31392 16992
rect 31444 16980 31450 16992
rect 31754 16980 31760 16992
rect 31444 16952 31760 16980
rect 31444 16940 31450 16952
rect 31754 16940 31760 16952
rect 31812 16980 31818 16992
rect 31938 16980 31944 16992
rect 31812 16952 31944 16980
rect 31812 16940 31818 16952
rect 31938 16940 31944 16952
rect 31996 16940 32002 16992
rect 32416 16980 32444 17088
rect 33226 17076 33232 17128
rect 33284 17116 33290 17128
rect 34238 17116 34244 17128
rect 33284 17088 34244 17116
rect 33284 17076 33290 17088
rect 34238 17076 34244 17088
rect 34296 17076 34302 17128
rect 34882 17076 34888 17128
rect 34940 17116 34946 17128
rect 35345 17119 35403 17125
rect 35345 17116 35357 17119
rect 34940 17088 35357 17116
rect 34940 17076 34946 17088
rect 35345 17085 35357 17088
rect 35391 17085 35403 17119
rect 35345 17079 35403 17085
rect 35434 17076 35440 17128
rect 35492 17116 35498 17128
rect 36449 17119 36507 17125
rect 36449 17116 36461 17119
rect 35492 17088 36461 17116
rect 35492 17076 35498 17088
rect 36449 17085 36461 17088
rect 36495 17085 36507 17119
rect 36449 17079 36507 17085
rect 36538 17076 36544 17128
rect 36596 17076 36602 17128
rect 38105 17119 38163 17125
rect 38105 17085 38117 17119
rect 38151 17116 38163 17119
rect 38746 17116 38752 17128
rect 38151 17088 38752 17116
rect 38151 17085 38163 17088
rect 38105 17079 38163 17085
rect 38746 17076 38752 17088
rect 38804 17076 38810 17128
rect 38841 17119 38899 17125
rect 38841 17085 38853 17119
rect 38887 17085 38899 17119
rect 38841 17079 38899 17085
rect 39117 17119 39175 17125
rect 39117 17085 39129 17119
rect 39163 17116 39175 17119
rect 43346 17116 43352 17128
rect 39163 17088 43352 17116
rect 39163 17085 39175 17088
rect 39117 17079 39175 17085
rect 33686 17008 33692 17060
rect 33744 17048 33750 17060
rect 34057 17051 34115 17057
rect 34057 17048 34069 17051
rect 33744 17020 34069 17048
rect 33744 17008 33750 17020
rect 34057 17017 34069 17020
rect 34103 17048 34115 17051
rect 34974 17048 34980 17060
rect 34103 17020 34980 17048
rect 34103 17017 34115 17020
rect 34057 17011 34115 17017
rect 34974 17008 34980 17020
rect 35032 17008 35038 17060
rect 37001 17051 37059 17057
rect 37001 17048 37013 17051
rect 35084 17020 37013 17048
rect 33870 16980 33876 16992
rect 32416 16952 33876 16980
rect 33870 16940 33876 16952
rect 33928 16940 33934 16992
rect 34238 16940 34244 16992
rect 34296 16980 34302 16992
rect 35084 16980 35112 17020
rect 37001 17017 37013 17020
rect 37047 17017 37059 17051
rect 37001 17011 37059 17017
rect 37734 17008 37740 17060
rect 37792 17048 37798 17060
rect 38856 17048 38884 17079
rect 43346 17076 43352 17088
rect 43404 17076 43410 17128
rect 41693 17051 41751 17057
rect 41693 17048 41705 17051
rect 37792 17020 38884 17048
rect 40144 17020 41705 17048
rect 37792 17008 37798 17020
rect 34296 16952 35112 16980
rect 35989 16983 36047 16989
rect 34296 16940 34302 16952
rect 35989 16949 36001 16983
rect 36035 16980 36047 16983
rect 37090 16980 37096 16992
rect 36035 16952 37096 16980
rect 36035 16949 36047 16952
rect 35989 16943 36047 16949
rect 37090 16940 37096 16952
rect 37148 16940 37154 16992
rect 37366 16940 37372 16992
rect 37424 16980 37430 16992
rect 38473 16983 38531 16989
rect 38473 16980 38485 16983
rect 37424 16952 38485 16980
rect 37424 16940 37430 16952
rect 38473 16949 38485 16952
rect 38519 16949 38531 16983
rect 38473 16943 38531 16949
rect 38562 16940 38568 16992
rect 38620 16980 38626 16992
rect 40144 16980 40172 17020
rect 41693 17017 41705 17020
rect 41739 17017 41751 17051
rect 41693 17011 41751 17017
rect 38620 16952 40172 16980
rect 38620 16940 38626 16952
rect 40586 16940 40592 16992
rect 40644 16940 40650 16992
rect 48682 16940 48688 16992
rect 48740 16980 48746 16992
rect 49237 16983 49295 16989
rect 49237 16980 49249 16983
rect 48740 16952 49249 16980
rect 48740 16940 48746 16952
rect 49237 16949 49249 16952
rect 49283 16949 49295 16983
rect 49237 16943 49295 16949
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 4617 16779 4675 16785
rect 4617 16745 4629 16779
rect 4663 16776 4675 16779
rect 5810 16776 5816 16788
rect 4663 16748 5816 16776
rect 4663 16745 4675 16748
rect 4617 16739 4675 16745
rect 5810 16736 5816 16748
rect 5868 16736 5874 16788
rect 7469 16779 7527 16785
rect 7469 16745 7481 16779
rect 7515 16776 7527 16779
rect 8570 16776 8576 16788
rect 7515 16748 8576 16776
rect 7515 16745 7527 16748
rect 7469 16739 7527 16745
rect 8570 16736 8576 16748
rect 8628 16736 8634 16788
rect 8662 16736 8668 16788
rect 8720 16776 8726 16788
rect 8941 16779 8999 16785
rect 8941 16776 8953 16779
rect 8720 16748 8953 16776
rect 8720 16736 8726 16748
rect 8941 16745 8953 16748
rect 8987 16745 8999 16779
rect 8941 16739 8999 16745
rect 10226 16736 10232 16788
rect 10284 16776 10290 16788
rect 10870 16776 10876 16788
rect 10284 16748 10876 16776
rect 10284 16736 10290 16748
rect 10870 16736 10876 16748
rect 10928 16776 10934 16788
rect 14458 16776 14464 16788
rect 10928 16748 14464 16776
rect 10928 16736 10934 16748
rect 14458 16736 14464 16748
rect 14516 16736 14522 16788
rect 14734 16736 14740 16788
rect 14792 16776 14798 16788
rect 16206 16776 16212 16788
rect 14792 16748 16212 16776
rect 14792 16736 14798 16748
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 16393 16779 16451 16785
rect 16393 16745 16405 16779
rect 16439 16776 16451 16779
rect 16439 16748 16620 16776
rect 16439 16745 16451 16748
rect 16393 16739 16451 16745
rect 5626 16668 5632 16720
rect 5684 16708 5690 16720
rect 5684 16680 8248 16708
rect 5684 16668 5690 16680
rect 8220 16649 8248 16680
rect 8478 16668 8484 16720
rect 8536 16708 8542 16720
rect 9585 16711 9643 16717
rect 9585 16708 9597 16711
rect 8536 16680 9597 16708
rect 8536 16668 8542 16680
rect 9585 16677 9597 16680
rect 9631 16677 9643 16711
rect 16022 16708 16028 16720
rect 9585 16671 9643 16677
rect 14108 16680 16028 16708
rect 14108 16652 14136 16680
rect 16022 16668 16028 16680
rect 16080 16708 16086 16720
rect 16482 16708 16488 16720
rect 16080 16680 16488 16708
rect 16080 16668 16086 16680
rect 16482 16668 16488 16680
rect 16540 16668 16546 16720
rect 16592 16708 16620 16748
rect 16942 16736 16948 16788
rect 17000 16776 17006 16788
rect 17586 16776 17592 16788
rect 17000 16748 17592 16776
rect 17000 16736 17006 16748
rect 17586 16736 17592 16748
rect 17644 16736 17650 16788
rect 19242 16736 19248 16788
rect 19300 16776 19306 16788
rect 20441 16779 20499 16785
rect 20441 16776 20453 16779
rect 19300 16748 20453 16776
rect 19300 16736 19306 16748
rect 20441 16745 20453 16748
rect 20487 16776 20499 16779
rect 23290 16776 23296 16788
rect 20487 16748 23296 16776
rect 20487 16745 20499 16748
rect 20441 16739 20499 16745
rect 23290 16736 23296 16748
rect 23348 16776 23354 16788
rect 25317 16779 25375 16785
rect 25317 16776 25329 16779
rect 23348 16748 25329 16776
rect 23348 16736 23354 16748
rect 25317 16745 25329 16748
rect 25363 16776 25375 16779
rect 25363 16748 28994 16776
rect 25363 16745 25375 16748
rect 25317 16739 25375 16745
rect 28966 16720 28994 16748
rect 29362 16736 29368 16788
rect 29420 16776 29426 16788
rect 31113 16779 31171 16785
rect 31113 16776 31125 16779
rect 29420 16748 31125 16776
rect 29420 16736 29426 16748
rect 31113 16745 31125 16748
rect 31159 16745 31171 16779
rect 31113 16739 31171 16745
rect 32122 16736 32128 16788
rect 32180 16776 32186 16788
rect 33502 16776 33508 16788
rect 32180 16748 33508 16776
rect 32180 16736 32186 16748
rect 33502 16736 33508 16748
rect 33560 16736 33566 16788
rect 34146 16736 34152 16788
rect 34204 16776 34210 16788
rect 34517 16779 34575 16785
rect 34517 16776 34529 16779
rect 34204 16748 34529 16776
rect 34204 16736 34210 16748
rect 34517 16745 34529 16748
rect 34563 16745 34575 16779
rect 34517 16739 34575 16745
rect 34790 16736 34796 16788
rect 34848 16776 34854 16788
rect 35894 16776 35900 16788
rect 34848 16748 35900 16776
rect 34848 16736 34854 16748
rect 35894 16736 35900 16748
rect 35952 16736 35958 16788
rect 36265 16779 36323 16785
rect 36265 16745 36277 16779
rect 36311 16776 36323 16779
rect 36354 16776 36360 16788
rect 36311 16748 36360 16776
rect 36311 16745 36323 16748
rect 36265 16739 36323 16745
rect 36354 16736 36360 16748
rect 36412 16736 36418 16788
rect 36998 16736 37004 16788
rect 37056 16776 37062 16788
rect 39485 16779 39543 16785
rect 39485 16776 39497 16779
rect 37056 16748 39497 16776
rect 37056 16736 37062 16748
rect 39485 16745 39497 16748
rect 39531 16776 39543 16779
rect 41046 16776 41052 16788
rect 39531 16748 41052 16776
rect 39531 16745 39543 16748
rect 39485 16739 39543 16745
rect 41046 16736 41052 16748
rect 41104 16736 41110 16788
rect 48774 16736 48780 16788
rect 48832 16736 48838 16788
rect 17402 16708 17408 16720
rect 16592 16680 17408 16708
rect 17402 16668 17408 16680
rect 17460 16668 17466 16720
rect 20162 16708 20168 16720
rect 20088 16680 20168 16708
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16609 8263 16643
rect 8205 16603 8263 16609
rect 8294 16600 8300 16652
rect 8352 16600 8358 16652
rect 8938 16600 8944 16652
rect 8996 16640 9002 16652
rect 10134 16640 10140 16652
rect 8996 16612 10140 16640
rect 8996 16600 9002 16612
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 10410 16600 10416 16652
rect 10468 16640 10474 16652
rect 11701 16643 11759 16649
rect 11701 16640 11713 16643
rect 10468 16612 11713 16640
rect 10468 16600 10474 16612
rect 11701 16609 11713 16612
rect 11747 16609 11759 16643
rect 11701 16603 11759 16609
rect 13446 16600 13452 16652
rect 13504 16600 13510 16652
rect 13541 16643 13599 16649
rect 13541 16609 13553 16643
rect 13587 16640 13599 16643
rect 13998 16640 14004 16652
rect 13587 16612 14004 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 13998 16600 14004 16612
rect 14056 16600 14062 16652
rect 14090 16600 14096 16652
rect 14148 16600 14154 16652
rect 14366 16600 14372 16652
rect 14424 16640 14430 16652
rect 14921 16643 14979 16649
rect 14921 16640 14933 16643
rect 14424 16612 14933 16640
rect 14424 16600 14430 16612
rect 14921 16609 14933 16612
rect 14967 16609 14979 16643
rect 14921 16603 14979 16609
rect 15013 16643 15071 16649
rect 15013 16609 15025 16643
rect 15059 16609 15071 16643
rect 15013 16603 15071 16609
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16572 1823 16575
rect 4062 16572 4068 16584
rect 1811 16544 4068 16572
rect 1811 16541 1823 16544
rect 1765 16535 1823 16541
rect 4062 16532 4068 16544
rect 4120 16532 4126 16584
rect 4154 16532 4160 16584
rect 4212 16532 4218 16584
rect 4798 16532 4804 16584
rect 4856 16532 4862 16584
rect 5445 16575 5503 16581
rect 5445 16541 5457 16575
rect 5491 16572 5503 16575
rect 6362 16572 6368 16584
rect 5491 16544 6368 16572
rect 5491 16541 5503 16544
rect 5445 16535 5503 16541
rect 6362 16532 6368 16544
rect 6420 16532 6426 16584
rect 6454 16532 6460 16584
rect 6512 16572 6518 16584
rect 6733 16575 6791 16581
rect 6733 16572 6745 16575
rect 6512 16544 6745 16572
rect 6512 16532 6518 16544
rect 6733 16541 6745 16544
rect 6779 16541 6791 16575
rect 6733 16535 6791 16541
rect 8018 16532 8024 16584
rect 8076 16532 8082 16584
rect 10042 16532 10048 16584
rect 10100 16532 10106 16584
rect 11238 16572 11244 16584
rect 11072 16544 11244 16572
rect 1302 16464 1308 16516
rect 1360 16504 1366 16516
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1360 16476 2513 16504
rect 1360 16464 1366 16476
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 8036 16504 8064 16532
rect 8113 16507 8171 16513
rect 8113 16504 8125 16507
rect 8036 16476 8125 16504
rect 2501 16467 2559 16473
rect 8113 16473 8125 16476
rect 8159 16473 8171 16507
rect 8113 16467 8171 16473
rect 9398 16464 9404 16516
rect 9456 16464 9462 16516
rect 9582 16464 9588 16516
rect 9640 16504 9646 16516
rect 10689 16507 10747 16513
rect 10689 16504 10701 16507
rect 9640 16476 10701 16504
rect 9640 16464 9646 16476
rect 10689 16473 10701 16476
rect 10735 16473 10747 16507
rect 10689 16467 10747 16473
rect 3970 16396 3976 16448
rect 4028 16396 4034 16448
rect 5261 16439 5319 16445
rect 5261 16405 5273 16439
rect 5307 16436 5319 16439
rect 5350 16436 5356 16448
rect 5307 16408 5356 16436
rect 5307 16405 5319 16408
rect 5261 16399 5319 16405
rect 5350 16396 5356 16408
rect 5408 16396 5414 16448
rect 6549 16439 6607 16445
rect 6549 16405 6561 16439
rect 6595 16436 6607 16439
rect 6914 16436 6920 16448
rect 6595 16408 6920 16436
rect 6595 16405 6607 16408
rect 6549 16399 6607 16405
rect 6914 16396 6920 16408
rect 6972 16396 6978 16448
rect 7745 16439 7803 16445
rect 7745 16405 7757 16439
rect 7791 16436 7803 16439
rect 8846 16436 8852 16448
rect 7791 16408 8852 16436
rect 7791 16405 7803 16408
rect 7745 16399 7803 16405
rect 8846 16396 8852 16408
rect 8904 16396 8910 16448
rect 8938 16396 8944 16448
rect 8996 16436 9002 16448
rect 11072 16436 11100 16544
rect 11238 16532 11244 16544
rect 11296 16532 11302 16584
rect 11330 16532 11336 16584
rect 11388 16572 11394 16584
rect 12434 16572 12440 16584
rect 11388 16544 12440 16572
rect 11388 16532 11394 16544
rect 12434 16532 12440 16544
rect 12492 16532 12498 16584
rect 12529 16575 12587 16581
rect 12529 16541 12541 16575
rect 12575 16572 12587 16575
rect 13630 16572 13636 16584
rect 12575 16544 13636 16572
rect 12575 16541 12587 16544
rect 12529 16535 12587 16541
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 14826 16532 14832 16584
rect 14884 16532 14890 16584
rect 11882 16504 11888 16516
rect 11164 16476 11888 16504
rect 11164 16445 11192 16476
rect 11882 16464 11888 16476
rect 11940 16464 11946 16516
rect 12066 16464 12072 16516
rect 12124 16504 12130 16516
rect 13357 16507 13415 16513
rect 13357 16504 13369 16507
rect 12124 16476 13369 16504
rect 12124 16464 12130 16476
rect 13357 16473 13369 16476
rect 13403 16504 13415 16507
rect 14844 16504 14872 16532
rect 13403 16476 14872 16504
rect 15028 16504 15056 16603
rect 15102 16600 15108 16652
rect 15160 16640 15166 16652
rect 20088 16649 20116 16680
rect 20162 16668 20168 16680
rect 20220 16668 20226 16720
rect 20809 16711 20867 16717
rect 20809 16677 20821 16711
rect 20855 16708 20867 16711
rect 20898 16708 20904 16720
rect 20855 16680 20904 16708
rect 20855 16677 20867 16680
rect 20809 16671 20867 16677
rect 20898 16668 20904 16680
rect 20956 16668 20962 16720
rect 23934 16708 23940 16720
rect 23768 16680 23940 16708
rect 18693 16643 18751 16649
rect 18693 16640 18705 16643
rect 15160 16612 18705 16640
rect 15160 16600 15166 16612
rect 18693 16609 18705 16612
rect 18739 16609 18751 16643
rect 18693 16603 18751 16609
rect 20073 16643 20131 16649
rect 20073 16609 20085 16643
rect 20119 16609 20131 16643
rect 20073 16603 20131 16609
rect 21082 16600 21088 16652
rect 21140 16600 21146 16652
rect 21361 16643 21419 16649
rect 21361 16609 21373 16643
rect 21407 16640 21419 16643
rect 22738 16640 22744 16652
rect 21407 16612 22744 16640
rect 21407 16609 21419 16612
rect 21361 16603 21419 16609
rect 22738 16600 22744 16612
rect 22796 16600 22802 16652
rect 23768 16649 23796 16680
rect 23934 16668 23940 16680
rect 23992 16668 23998 16720
rect 24026 16668 24032 16720
rect 24084 16708 24090 16720
rect 25041 16711 25099 16717
rect 25041 16708 25053 16711
rect 24084 16680 25053 16708
rect 24084 16668 24090 16680
rect 25041 16677 25053 16680
rect 25087 16677 25099 16711
rect 28966 16680 29000 16720
rect 25041 16671 25099 16677
rect 28994 16668 29000 16680
rect 29052 16708 29058 16720
rect 30374 16708 30380 16720
rect 29052 16680 30380 16708
rect 29052 16668 29058 16680
rect 30374 16668 30380 16680
rect 30432 16668 30438 16720
rect 30466 16668 30472 16720
rect 30524 16708 30530 16720
rect 30929 16711 30987 16717
rect 30929 16708 30941 16711
rect 30524 16680 30941 16708
rect 30524 16668 30530 16680
rect 30929 16677 30941 16680
rect 30975 16708 30987 16711
rect 31018 16708 31024 16720
rect 30975 16680 31024 16708
rect 30975 16677 30987 16680
rect 30929 16671 30987 16677
rect 31018 16668 31024 16680
rect 31076 16668 31082 16720
rect 32858 16668 32864 16720
rect 32916 16708 32922 16720
rect 33229 16711 33287 16717
rect 33229 16708 33241 16711
rect 32916 16680 33241 16708
rect 32916 16668 32922 16680
rect 33229 16677 33241 16680
rect 33275 16677 33287 16711
rect 33229 16671 33287 16677
rect 34606 16668 34612 16720
rect 34664 16708 34670 16720
rect 37366 16708 37372 16720
rect 34664 16680 37372 16708
rect 34664 16668 34670 16680
rect 23753 16643 23811 16649
rect 23753 16609 23765 16643
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 23845 16643 23903 16649
rect 23845 16609 23857 16643
rect 23891 16640 23903 16643
rect 23891 16612 24808 16640
rect 23891 16609 23903 16612
rect 23845 16603 23903 16609
rect 15746 16532 15752 16584
rect 15804 16532 15810 16584
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16541 16911 16575
rect 16853 16535 16911 16541
rect 17497 16575 17555 16581
rect 17497 16541 17509 16575
rect 17543 16572 17555 16575
rect 17543 16544 20852 16572
rect 17543 16541 17555 16544
rect 17497 16535 17555 16541
rect 16666 16504 16672 16516
rect 15028 16476 16672 16504
rect 13403 16473 13415 16476
rect 13357 16467 13415 16473
rect 16666 16464 16672 16476
rect 16724 16464 16730 16516
rect 8996 16408 11100 16436
rect 11149 16439 11207 16445
rect 8996 16396 9002 16408
rect 11149 16405 11161 16439
rect 11195 16405 11207 16439
rect 11149 16399 11207 16405
rect 11514 16396 11520 16448
rect 11572 16396 11578 16448
rect 11606 16396 11612 16448
rect 11664 16396 11670 16448
rect 11974 16396 11980 16448
rect 12032 16436 12038 16448
rect 12345 16439 12403 16445
rect 12345 16436 12357 16439
rect 12032 16408 12357 16436
rect 12032 16396 12038 16408
rect 12345 16405 12357 16408
rect 12391 16405 12403 16439
rect 12345 16399 12403 16405
rect 12986 16396 12992 16448
rect 13044 16396 13050 16448
rect 14458 16396 14464 16448
rect 14516 16396 14522 16448
rect 16868 16436 16896 16535
rect 17957 16507 18015 16513
rect 17957 16473 17969 16507
rect 18003 16504 18015 16507
rect 18322 16504 18328 16516
rect 18003 16476 18328 16504
rect 18003 16473 18015 16476
rect 17957 16467 18015 16473
rect 18322 16464 18328 16476
rect 18380 16504 18386 16516
rect 19242 16504 19248 16516
rect 18380 16476 19248 16504
rect 18380 16464 18386 16476
rect 19242 16464 19248 16476
rect 19300 16464 19306 16516
rect 19889 16507 19947 16513
rect 19889 16473 19901 16507
rect 19935 16504 19947 16507
rect 20714 16504 20720 16516
rect 19935 16476 20720 16504
rect 19935 16473 19947 16476
rect 19889 16467 19947 16473
rect 20714 16464 20720 16476
rect 20772 16464 20778 16516
rect 19334 16436 19340 16448
rect 16868 16408 19340 16436
rect 19334 16396 19340 16408
rect 19392 16396 19398 16448
rect 19426 16396 19432 16448
rect 19484 16396 19490 16448
rect 19794 16396 19800 16448
rect 19852 16396 19858 16448
rect 20824 16436 20852 16544
rect 20898 16464 20904 16516
rect 20956 16504 20962 16516
rect 23750 16504 23756 16516
rect 20956 16476 21850 16504
rect 22848 16476 23756 16504
rect 20956 16464 20962 16476
rect 22848 16448 22876 16476
rect 23750 16464 23756 16476
rect 23808 16464 23814 16516
rect 24780 16504 24808 16612
rect 24854 16600 24860 16652
rect 24912 16640 24918 16652
rect 25593 16643 25651 16649
rect 25593 16640 25605 16643
rect 24912 16612 25605 16640
rect 24912 16600 24918 16612
rect 25593 16609 25605 16612
rect 25639 16640 25651 16643
rect 28350 16640 28356 16652
rect 25639 16612 28356 16640
rect 25639 16609 25651 16612
rect 25593 16603 25651 16609
rect 28350 16600 28356 16612
rect 28408 16600 28414 16652
rect 29178 16600 29184 16652
rect 29236 16640 29242 16652
rect 29236 16612 29868 16640
rect 29236 16600 29242 16612
rect 28077 16575 28135 16581
rect 28077 16541 28089 16575
rect 28123 16572 28135 16575
rect 28442 16572 28448 16584
rect 28123 16544 28448 16572
rect 28123 16541 28135 16544
rect 28077 16535 28135 16541
rect 28442 16532 28448 16544
rect 28500 16532 28506 16584
rect 28537 16575 28595 16581
rect 28537 16541 28549 16575
rect 28583 16541 28595 16575
rect 28537 16535 28595 16541
rect 24780 16476 25176 16504
rect 22370 16436 22376 16448
rect 20824 16408 22376 16436
rect 22370 16396 22376 16408
rect 22428 16396 22434 16448
rect 22830 16396 22836 16448
rect 22888 16396 22894 16448
rect 23290 16396 23296 16448
rect 23348 16396 23354 16448
rect 23474 16396 23480 16448
rect 23532 16436 23538 16448
rect 23661 16439 23719 16445
rect 23661 16436 23673 16439
rect 23532 16408 23673 16436
rect 23532 16396 23538 16408
rect 23661 16405 23673 16408
rect 23707 16405 23719 16439
rect 23661 16399 23719 16405
rect 24302 16396 24308 16448
rect 24360 16436 24366 16448
rect 24581 16439 24639 16445
rect 24581 16436 24593 16439
rect 24360 16408 24593 16436
rect 24360 16396 24366 16408
rect 24581 16405 24593 16408
rect 24627 16405 24639 16439
rect 25148 16436 25176 16476
rect 25774 16464 25780 16516
rect 25832 16504 25838 16516
rect 25869 16507 25927 16513
rect 25869 16504 25881 16507
rect 25832 16476 25881 16504
rect 25832 16464 25838 16476
rect 25869 16473 25881 16476
rect 25915 16473 25927 16507
rect 25869 16467 25927 16473
rect 26602 16464 26608 16516
rect 26660 16464 26666 16516
rect 27522 16504 27528 16516
rect 27356 16476 27528 16504
rect 27356 16445 27384 16476
rect 27522 16464 27528 16476
rect 27580 16464 27586 16516
rect 28552 16504 28580 16535
rect 28902 16532 28908 16584
rect 28960 16572 28966 16584
rect 29730 16572 29736 16584
rect 28960 16544 29736 16572
rect 28960 16532 28966 16544
rect 29730 16532 29736 16544
rect 29788 16532 29794 16584
rect 29840 16572 29868 16612
rect 29914 16600 29920 16652
rect 29972 16640 29978 16652
rect 30285 16643 30343 16649
rect 30285 16640 30297 16643
rect 29972 16612 30297 16640
rect 29972 16600 29978 16612
rect 30285 16609 30297 16612
rect 30331 16609 30343 16643
rect 31386 16640 31392 16652
rect 30285 16603 30343 16609
rect 30392 16612 31392 16640
rect 30193 16575 30251 16581
rect 30193 16572 30205 16575
rect 29840 16544 30205 16572
rect 30193 16541 30205 16544
rect 30239 16572 30251 16575
rect 30392 16572 30420 16612
rect 31386 16600 31392 16612
rect 31444 16600 31450 16652
rect 31481 16643 31539 16649
rect 31481 16609 31493 16643
rect 31527 16640 31539 16643
rect 32490 16640 32496 16652
rect 31527 16612 32496 16640
rect 31527 16609 31539 16612
rect 31481 16603 31539 16609
rect 32490 16600 32496 16612
rect 32548 16600 32554 16652
rect 32950 16600 32956 16652
rect 33008 16640 33014 16652
rect 34333 16643 34391 16649
rect 34333 16640 34345 16643
rect 33008 16612 34345 16640
rect 33008 16600 33014 16612
rect 34333 16609 34345 16612
rect 34379 16640 34391 16643
rect 34790 16640 34796 16652
rect 34379 16612 34796 16640
rect 34379 16609 34391 16612
rect 34333 16603 34391 16609
rect 34790 16600 34796 16612
rect 34848 16600 34854 16652
rect 30239 16544 30420 16572
rect 30239 16541 30251 16544
rect 30193 16535 30251 16541
rect 33594 16532 33600 16584
rect 33652 16572 33658 16584
rect 34900 16581 34928 16680
rect 37366 16668 37372 16680
rect 37424 16668 37430 16720
rect 35710 16600 35716 16652
rect 35768 16600 35774 16652
rect 36909 16643 36967 16649
rect 36909 16609 36921 16643
rect 36955 16609 36967 16643
rect 38013 16643 38071 16649
rect 38013 16640 38025 16643
rect 36909 16603 36967 16609
rect 37108 16612 38025 16640
rect 33781 16575 33839 16581
rect 33781 16572 33793 16575
rect 33652 16544 33793 16572
rect 33652 16532 33658 16544
rect 33781 16541 33793 16544
rect 33827 16541 33839 16575
rect 33781 16535 33839 16541
rect 34885 16575 34943 16581
rect 34885 16541 34897 16575
rect 34931 16541 34943 16575
rect 34885 16535 34943 16541
rect 36722 16532 36728 16584
rect 36780 16532 36786 16584
rect 36924 16572 36952 16603
rect 36998 16572 37004 16584
rect 36924 16544 37004 16572
rect 36998 16532 37004 16544
rect 37056 16532 37062 16584
rect 30374 16504 30380 16516
rect 28552 16476 30380 16504
rect 30374 16464 30380 16476
rect 30432 16504 30438 16516
rect 31662 16504 31668 16516
rect 30432 16476 31668 16504
rect 30432 16464 30438 16476
rect 31662 16464 31668 16476
rect 31720 16464 31726 16516
rect 31754 16464 31760 16516
rect 31812 16464 31818 16516
rect 32982 16476 33364 16504
rect 27341 16439 27399 16445
rect 27341 16436 27353 16439
rect 25148 16408 27353 16436
rect 24581 16399 24639 16405
rect 27341 16405 27353 16408
rect 27387 16405 27399 16439
rect 27341 16399 27399 16405
rect 27430 16396 27436 16448
rect 27488 16436 27494 16448
rect 27893 16439 27951 16445
rect 27893 16436 27905 16439
rect 27488 16408 27905 16436
rect 27488 16396 27494 16408
rect 27893 16405 27905 16408
rect 27939 16405 27951 16439
rect 27893 16399 27951 16405
rect 29178 16396 29184 16448
rect 29236 16396 29242 16448
rect 29730 16396 29736 16448
rect 29788 16396 29794 16448
rect 30101 16439 30159 16445
rect 30101 16405 30113 16439
rect 30147 16436 30159 16439
rect 30190 16436 30196 16448
rect 30147 16408 30196 16436
rect 30147 16405 30159 16408
rect 30101 16399 30159 16405
rect 30190 16396 30196 16408
rect 30248 16396 30254 16448
rect 30282 16396 30288 16448
rect 30340 16436 30346 16448
rect 30745 16439 30803 16445
rect 30745 16436 30757 16439
rect 30340 16408 30757 16436
rect 30340 16396 30346 16408
rect 30745 16405 30757 16408
rect 30791 16436 30803 16439
rect 33060 16436 33088 16476
rect 30791 16408 33088 16436
rect 33336 16436 33364 16476
rect 34146 16464 34152 16516
rect 34204 16504 34210 16516
rect 34204 16476 36768 16504
rect 34204 16464 34210 16476
rect 34238 16436 34244 16448
rect 33336 16408 34244 16436
rect 30791 16405 30803 16408
rect 30745 16399 30803 16405
rect 34238 16396 34244 16408
rect 34296 16396 34302 16448
rect 34974 16396 34980 16448
rect 35032 16436 35038 16448
rect 36630 16436 36636 16448
rect 35032 16408 36636 16436
rect 35032 16396 35038 16408
rect 36630 16396 36636 16408
rect 36688 16396 36694 16448
rect 36740 16436 36768 16476
rect 36906 16464 36912 16516
rect 36964 16504 36970 16516
rect 37108 16504 37136 16612
rect 38013 16609 38025 16612
rect 38059 16640 38071 16643
rect 40586 16640 40592 16652
rect 38059 16612 40592 16640
rect 38059 16609 38071 16612
rect 38013 16603 38071 16609
rect 40586 16600 40592 16612
rect 40644 16600 40650 16652
rect 37182 16532 37188 16584
rect 37240 16572 37246 16584
rect 37277 16575 37335 16581
rect 37277 16572 37289 16575
rect 37240 16544 37289 16572
rect 37240 16532 37246 16544
rect 37277 16541 37289 16544
rect 37323 16541 37335 16575
rect 37277 16535 37335 16541
rect 36964 16476 37136 16504
rect 37292 16504 37320 16535
rect 37458 16532 37464 16584
rect 37516 16572 37522 16584
rect 37734 16572 37740 16584
rect 37516 16544 37740 16572
rect 37516 16532 37522 16544
rect 37734 16532 37740 16544
rect 37792 16532 37798 16584
rect 40037 16575 40095 16581
rect 40037 16572 40049 16575
rect 39316 16544 40049 16572
rect 38470 16504 38476 16516
rect 37292 16476 38476 16504
rect 36964 16464 36970 16476
rect 38470 16464 38476 16476
rect 38528 16464 38534 16516
rect 39316 16436 39344 16544
rect 40037 16541 40049 16544
rect 40083 16541 40095 16575
rect 40037 16535 40095 16541
rect 40310 16532 40316 16584
rect 40368 16572 40374 16584
rect 41141 16575 41199 16581
rect 41141 16572 41153 16575
rect 40368 16544 41153 16572
rect 40368 16532 40374 16544
rect 41141 16541 41153 16544
rect 41187 16541 41199 16575
rect 41141 16535 41199 16541
rect 41322 16532 41328 16584
rect 41380 16572 41386 16584
rect 42245 16575 42303 16581
rect 42245 16572 42257 16575
rect 41380 16544 42257 16572
rect 41380 16532 41386 16544
rect 42245 16541 42257 16544
rect 42291 16541 42303 16575
rect 42245 16535 42303 16541
rect 48593 16575 48651 16581
rect 48593 16541 48605 16575
rect 48639 16572 48651 16575
rect 49053 16575 49111 16581
rect 49053 16572 49065 16575
rect 48639 16544 49065 16572
rect 48639 16541 48651 16544
rect 48593 16535 48651 16541
rect 49053 16541 49065 16544
rect 49099 16572 49111 16575
rect 49142 16572 49148 16584
rect 49099 16544 49148 16572
rect 49099 16541 49111 16544
rect 49053 16535 49111 16541
rect 49142 16532 49148 16544
rect 49200 16532 49206 16584
rect 40678 16464 40684 16516
rect 40736 16464 40742 16516
rect 36740 16408 39344 16436
rect 39666 16396 39672 16448
rect 39724 16436 39730 16448
rect 41785 16439 41843 16445
rect 41785 16436 41797 16439
rect 39724 16408 41797 16436
rect 39724 16396 39730 16408
rect 41785 16405 41797 16408
rect 41831 16405 41843 16439
rect 41785 16399 41843 16405
rect 42150 16396 42156 16448
rect 42208 16436 42214 16448
rect 42889 16439 42947 16445
rect 42889 16436 42901 16439
rect 42208 16408 42901 16436
rect 42208 16396 42214 16408
rect 42889 16405 42901 16408
rect 42935 16405 42947 16439
rect 42889 16399 42947 16405
rect 49234 16396 49240 16448
rect 49292 16396 49298 16448
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 3970 16192 3976 16244
rect 4028 16232 4034 16244
rect 5902 16232 5908 16244
rect 4028 16204 5908 16232
rect 4028 16192 4034 16204
rect 5902 16192 5908 16204
rect 5960 16192 5966 16244
rect 6362 16192 6368 16244
rect 6420 16232 6426 16244
rect 8389 16235 8447 16241
rect 8389 16232 8401 16235
rect 6420 16204 8401 16232
rect 6420 16192 6426 16204
rect 8389 16201 8401 16204
rect 8435 16232 8447 16235
rect 9122 16232 9128 16244
rect 8435 16204 9128 16232
rect 8435 16201 8447 16204
rect 8389 16195 8447 16201
rect 9122 16192 9128 16204
rect 9180 16192 9186 16244
rect 10134 16192 10140 16244
rect 10192 16192 10198 16244
rect 11422 16232 11428 16244
rect 10520 16204 11428 16232
rect 4062 16124 4068 16176
rect 4120 16164 4126 16176
rect 8938 16164 8944 16176
rect 4120 16136 8944 16164
rect 4120 16124 4126 16136
rect 8938 16124 8944 16136
rect 8996 16124 9002 16176
rect 9858 16124 9864 16176
rect 9916 16124 9922 16176
rect 10045 16167 10103 16173
rect 10045 16133 10057 16167
rect 10091 16164 10103 16167
rect 10520 16164 10548 16204
rect 11422 16192 11428 16204
rect 11480 16192 11486 16244
rect 11606 16192 11612 16244
rect 11664 16232 11670 16244
rect 11977 16235 12035 16241
rect 11977 16232 11989 16235
rect 11664 16204 11989 16232
rect 11664 16192 11670 16204
rect 11977 16201 11989 16204
rect 12023 16201 12035 16235
rect 11977 16195 12035 16201
rect 12437 16235 12495 16241
rect 12437 16201 12449 16235
rect 12483 16232 12495 16235
rect 13173 16235 13231 16241
rect 13173 16232 13185 16235
rect 12483 16204 13185 16232
rect 12483 16201 12495 16204
rect 12437 16195 12495 16201
rect 13173 16201 13185 16204
rect 13219 16201 13231 16235
rect 13173 16195 13231 16201
rect 13541 16235 13599 16241
rect 13541 16201 13553 16235
rect 13587 16232 13599 16235
rect 14369 16235 14427 16241
rect 14369 16232 14381 16235
rect 13587 16204 14381 16232
rect 13587 16201 13599 16204
rect 13541 16195 13599 16201
rect 14369 16201 14381 16204
rect 14415 16201 14427 16235
rect 14369 16195 14427 16201
rect 14458 16192 14464 16244
rect 14516 16232 14522 16244
rect 15654 16232 15660 16244
rect 14516 16204 15660 16232
rect 14516 16192 14522 16204
rect 15654 16192 15660 16204
rect 15712 16192 15718 16244
rect 16022 16192 16028 16244
rect 16080 16192 16086 16244
rect 17218 16192 17224 16244
rect 17276 16232 17282 16244
rect 17865 16235 17923 16241
rect 17865 16232 17877 16235
rect 17276 16204 17877 16232
rect 17276 16192 17282 16204
rect 17865 16201 17877 16204
rect 17911 16201 17923 16235
rect 17865 16195 17923 16201
rect 18325 16235 18383 16241
rect 18325 16201 18337 16235
rect 18371 16232 18383 16235
rect 19242 16232 19248 16244
rect 18371 16204 19248 16232
rect 18371 16201 18383 16204
rect 18325 16195 18383 16201
rect 19242 16192 19248 16204
rect 19300 16192 19306 16244
rect 20070 16192 20076 16244
rect 20128 16232 20134 16244
rect 22830 16232 22836 16244
rect 20128 16204 22836 16232
rect 20128 16192 20134 16204
rect 22830 16192 22836 16204
rect 22888 16192 22894 16244
rect 23109 16235 23167 16241
rect 23109 16201 23121 16235
rect 23155 16232 23167 16235
rect 25038 16232 25044 16244
rect 23155 16204 25044 16232
rect 23155 16201 23167 16204
rect 23109 16195 23167 16201
rect 25038 16192 25044 16204
rect 25096 16192 25102 16244
rect 25866 16232 25872 16244
rect 25148 16204 25872 16232
rect 10091 16136 10548 16164
rect 10091 16133 10103 16136
rect 10045 16127 10103 16133
rect 10594 16124 10600 16176
rect 10652 16124 10658 16176
rect 10962 16124 10968 16176
rect 11020 16164 11026 16176
rect 11241 16167 11299 16173
rect 11241 16164 11253 16167
rect 11020 16136 11253 16164
rect 11020 16124 11026 16136
rect 11241 16133 11253 16136
rect 11287 16164 11299 16167
rect 12066 16164 12072 16176
rect 11287 16136 12072 16164
rect 11287 16133 11299 16136
rect 11241 16127 11299 16133
rect 12066 16124 12072 16136
rect 12124 16124 12130 16176
rect 12986 16124 12992 16176
rect 13044 16164 13050 16176
rect 13633 16167 13691 16173
rect 13633 16164 13645 16167
rect 13044 16136 13645 16164
rect 13044 16124 13050 16136
rect 13633 16133 13645 16136
rect 13679 16133 13691 16167
rect 13633 16127 13691 16133
rect 15010 16124 15016 16176
rect 15068 16164 15074 16176
rect 19337 16167 19395 16173
rect 19337 16164 19349 16167
rect 15068 16136 19349 16164
rect 15068 16124 15074 16136
rect 19337 16133 19349 16136
rect 19383 16133 19395 16167
rect 20898 16164 20904 16176
rect 20562 16136 20904 16164
rect 19337 16127 19395 16133
rect 20898 16124 20904 16136
rect 20956 16164 20962 16176
rect 21177 16167 21235 16173
rect 21177 16164 21189 16167
rect 20956 16136 21189 16164
rect 20956 16124 20962 16136
rect 21177 16133 21189 16136
rect 21223 16133 21235 16167
rect 21177 16127 21235 16133
rect 21542 16124 21548 16176
rect 21600 16124 21606 16176
rect 23477 16167 23535 16173
rect 23477 16133 23489 16167
rect 23523 16164 23535 16167
rect 23658 16164 23664 16176
rect 23523 16136 23664 16164
rect 23523 16133 23535 16136
rect 23477 16127 23535 16133
rect 23658 16124 23664 16136
rect 23716 16124 23722 16176
rect 24762 16164 24768 16176
rect 24596 16136 24768 16164
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16096 1823 16099
rect 5442 16096 5448 16108
rect 1811 16068 5448 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 5442 16056 5448 16068
rect 5500 16056 5506 16108
rect 8294 16056 8300 16108
rect 8352 16096 8358 16108
rect 9309 16099 9367 16105
rect 8352 16068 8708 16096
rect 8352 16056 8358 16068
rect 8680 16040 8708 16068
rect 9309 16065 9321 16099
rect 9355 16096 9367 16099
rect 11974 16096 11980 16108
rect 9355 16068 11980 16096
rect 9355 16065 9367 16068
rect 9309 16059 9367 16065
rect 11974 16056 11980 16068
rect 12032 16056 12038 16108
rect 12342 16056 12348 16108
rect 12400 16056 12406 16108
rect 14737 16099 14795 16105
rect 14737 16096 14749 16099
rect 13924 16068 14749 16096
rect 1302 15988 1308 16040
rect 1360 16028 1366 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1360 16000 2053 16028
rect 1360 15988 1366 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 4338 15988 4344 16040
rect 4396 16028 4402 16040
rect 8481 16031 8539 16037
rect 8481 16028 8493 16031
rect 4396 16000 8493 16028
rect 4396 15988 4402 16000
rect 8481 15997 8493 16000
rect 8527 15997 8539 16031
rect 8481 15991 8539 15997
rect 8662 15988 8668 16040
rect 8720 15988 8726 16040
rect 9674 15988 9680 16040
rect 9732 16028 9738 16040
rect 9732 16000 9996 16028
rect 9732 15988 9738 16000
rect 8021 15963 8079 15969
rect 8021 15929 8033 15963
rect 8067 15960 8079 15963
rect 9858 15960 9864 15972
rect 8067 15932 9864 15960
rect 8067 15929 8079 15932
rect 8021 15923 8079 15929
rect 9858 15920 9864 15932
rect 9916 15920 9922 15972
rect 9968 15960 9996 16000
rect 10042 15988 10048 16040
rect 10100 16028 10106 16040
rect 12618 16028 12624 16040
rect 10100 16000 12624 16028
rect 10100 15988 10106 16000
rect 12618 15988 12624 16000
rect 12676 15988 12682 16040
rect 13722 15988 13728 16040
rect 13780 15988 13786 16040
rect 10781 15963 10839 15969
rect 10781 15960 10793 15963
rect 9968 15932 10793 15960
rect 10781 15929 10793 15932
rect 10827 15929 10839 15963
rect 13924 15960 13952 16068
rect 14737 16065 14749 16068
rect 14783 16065 14795 16099
rect 14737 16059 14795 16065
rect 14826 16056 14832 16108
rect 14884 16056 14890 16108
rect 15930 16056 15936 16108
rect 15988 16056 15994 16108
rect 16945 16099 17003 16105
rect 16945 16065 16957 16099
rect 16991 16065 17003 16099
rect 16945 16059 17003 16065
rect 13998 15988 14004 16040
rect 14056 16028 14062 16040
rect 15013 16031 15071 16037
rect 15013 16028 15025 16031
rect 14056 16000 15025 16028
rect 14056 15988 14062 16000
rect 15013 15997 15025 16000
rect 15059 16028 15071 16031
rect 16209 16031 16267 16037
rect 16209 16028 16221 16031
rect 15059 16000 16221 16028
rect 15059 15997 15071 16000
rect 15013 15991 15071 15997
rect 16209 15997 16221 16000
rect 16255 16028 16267 16031
rect 16298 16028 16304 16040
rect 16255 16000 16304 16028
rect 16255 15997 16267 16000
rect 16209 15991 16267 15997
rect 16298 15988 16304 16000
rect 16356 15988 16362 16040
rect 16960 15960 16988 16059
rect 17678 16056 17684 16108
rect 17736 16096 17742 16108
rect 18233 16099 18291 16105
rect 18233 16096 18245 16099
rect 17736 16068 18245 16096
rect 17736 16056 17742 16068
rect 18233 16065 18245 16068
rect 18279 16065 18291 16099
rect 18233 16059 18291 16065
rect 18598 16056 18604 16108
rect 18656 16096 18662 16108
rect 19061 16099 19119 16105
rect 19061 16096 19073 16099
rect 18656 16068 19073 16096
rect 18656 16056 18662 16068
rect 19061 16065 19073 16068
rect 19107 16065 19119 16099
rect 19061 16059 19119 16065
rect 22002 16056 22008 16108
rect 22060 16056 22066 16108
rect 24596 16105 24624 16136
rect 24762 16124 24768 16136
rect 24820 16124 24826 16176
rect 24857 16167 24915 16173
rect 24857 16133 24869 16167
rect 24903 16164 24915 16167
rect 25148 16164 25176 16204
rect 25866 16192 25872 16204
rect 25924 16192 25930 16244
rect 26329 16235 26387 16241
rect 26329 16201 26341 16235
rect 26375 16232 26387 16235
rect 26418 16232 26424 16244
rect 26375 16204 26424 16232
rect 26375 16201 26387 16204
rect 26329 16195 26387 16201
rect 26418 16192 26424 16204
rect 26476 16192 26482 16244
rect 26602 16192 26608 16244
rect 26660 16192 26666 16244
rect 27338 16192 27344 16244
rect 27396 16232 27402 16244
rect 27522 16232 27528 16244
rect 27396 16204 27528 16232
rect 27396 16192 27402 16204
rect 27522 16192 27528 16204
rect 27580 16232 27586 16244
rect 27617 16235 27675 16241
rect 27617 16232 27629 16235
rect 27580 16204 27629 16232
rect 27580 16192 27586 16204
rect 27617 16201 27629 16204
rect 27663 16201 27675 16235
rect 29270 16232 29276 16244
rect 27617 16195 27675 16201
rect 27724 16204 29276 16232
rect 26620 16164 26648 16192
rect 27154 16164 27160 16176
rect 24903 16136 25176 16164
rect 26082 16136 27160 16164
rect 24903 16133 24915 16136
rect 24857 16127 24915 16133
rect 27154 16124 27160 16136
rect 27212 16164 27218 16176
rect 27724 16164 27752 16204
rect 27212 16136 27752 16164
rect 28629 16167 28687 16173
rect 27212 16124 27218 16136
rect 28629 16133 28641 16167
rect 28675 16164 28687 16167
rect 28902 16164 28908 16176
rect 28675 16136 28908 16164
rect 28675 16133 28687 16136
rect 28629 16127 28687 16133
rect 28902 16124 28908 16136
rect 28960 16124 28966 16176
rect 29012 16164 29040 16204
rect 29270 16192 29276 16204
rect 29328 16232 29334 16244
rect 30101 16235 30159 16241
rect 29328 16204 30052 16232
rect 29328 16192 29334 16204
rect 30024 16164 30052 16204
rect 30101 16201 30113 16235
rect 30147 16232 30159 16235
rect 30374 16232 30380 16244
rect 30147 16204 30380 16232
rect 30147 16201 30159 16204
rect 30101 16195 30159 16201
rect 30374 16192 30380 16204
rect 30432 16192 30438 16244
rect 30650 16192 30656 16244
rect 30708 16232 30714 16244
rect 31021 16235 31079 16241
rect 31021 16232 31033 16235
rect 30708 16204 31033 16232
rect 30708 16192 30714 16204
rect 31021 16201 31033 16204
rect 31067 16201 31079 16235
rect 31021 16195 31079 16201
rect 31849 16235 31907 16241
rect 31849 16201 31861 16235
rect 31895 16232 31907 16235
rect 31938 16232 31944 16244
rect 31895 16204 31944 16232
rect 31895 16201 31907 16204
rect 31849 16195 31907 16201
rect 31938 16192 31944 16204
rect 31996 16192 32002 16244
rect 32674 16192 32680 16244
rect 32732 16232 32738 16244
rect 32769 16235 32827 16241
rect 32769 16232 32781 16235
rect 32732 16204 32781 16232
rect 32732 16192 32738 16204
rect 32769 16201 32781 16204
rect 32815 16201 32827 16235
rect 32769 16195 32827 16201
rect 33962 16192 33968 16244
rect 34020 16192 34026 16244
rect 34609 16235 34667 16241
rect 34609 16201 34621 16235
rect 34655 16232 34667 16235
rect 34974 16232 34980 16244
rect 34655 16204 34980 16232
rect 34655 16201 34667 16204
rect 34609 16195 34667 16201
rect 34974 16192 34980 16204
rect 35032 16192 35038 16244
rect 35342 16192 35348 16244
rect 35400 16232 35406 16244
rect 36906 16232 36912 16244
rect 35400 16204 36912 16232
rect 35400 16192 35406 16204
rect 36906 16192 36912 16204
rect 36964 16192 36970 16244
rect 37366 16192 37372 16244
rect 37424 16232 37430 16244
rect 37461 16235 37519 16241
rect 37461 16232 37473 16235
rect 37424 16204 37473 16232
rect 37424 16192 37430 16204
rect 37461 16201 37473 16204
rect 37507 16201 37519 16235
rect 37461 16195 37519 16201
rect 38654 16192 38660 16244
rect 38712 16232 38718 16244
rect 40957 16235 41015 16241
rect 40957 16232 40969 16235
rect 38712 16204 40969 16232
rect 38712 16192 38718 16204
rect 40957 16201 40969 16204
rect 41003 16201 41015 16235
rect 40957 16195 41015 16201
rect 41598 16192 41604 16244
rect 41656 16232 41662 16244
rect 41693 16235 41751 16241
rect 41693 16232 41705 16235
rect 41656 16204 41705 16232
rect 41656 16192 41662 16204
rect 41693 16201 41705 16204
rect 41739 16232 41751 16235
rect 41877 16235 41935 16241
rect 41877 16232 41889 16235
rect 41739 16204 41889 16232
rect 41739 16201 41751 16204
rect 41693 16195 41751 16201
rect 41877 16201 41889 16204
rect 41923 16201 41935 16235
rect 41877 16195 41935 16201
rect 30282 16164 30288 16176
rect 29012 16136 29118 16164
rect 30024 16136 30288 16164
rect 30282 16124 30288 16136
rect 30340 16124 30346 16176
rect 30926 16124 30932 16176
rect 30984 16124 30990 16176
rect 34790 16124 34796 16176
rect 34848 16124 34854 16176
rect 36722 16124 36728 16176
rect 36780 16164 36786 16176
rect 37645 16167 37703 16173
rect 37645 16164 37657 16167
rect 36780 16136 37657 16164
rect 36780 16124 36786 16136
rect 37645 16133 37657 16136
rect 37691 16133 37703 16167
rect 37645 16127 37703 16133
rect 38473 16167 38531 16173
rect 38473 16133 38485 16167
rect 38519 16164 38531 16167
rect 38562 16164 38568 16176
rect 38519 16136 38568 16164
rect 38519 16133 38531 16136
rect 38473 16127 38531 16133
rect 38562 16124 38568 16136
rect 38620 16124 38626 16176
rect 38746 16124 38752 16176
rect 38804 16164 38810 16176
rect 40865 16167 40923 16173
rect 38804 16136 38962 16164
rect 38804 16124 38810 16136
rect 40865 16133 40877 16167
rect 40911 16164 40923 16167
rect 48958 16164 48964 16176
rect 40911 16136 48964 16164
rect 40911 16133 40923 16136
rect 40865 16127 40923 16133
rect 48958 16124 48964 16136
rect 49016 16124 49022 16176
rect 24581 16099 24639 16105
rect 24581 16065 24593 16099
rect 24627 16065 24639 16099
rect 24581 16059 24639 16065
rect 27430 16056 27436 16108
rect 27488 16096 27494 16108
rect 27525 16099 27583 16105
rect 27525 16096 27537 16099
rect 27488 16068 27537 16096
rect 27488 16056 27494 16068
rect 27525 16065 27537 16068
rect 27571 16065 27583 16099
rect 27525 16059 27583 16065
rect 28350 16056 28356 16108
rect 28408 16056 28414 16108
rect 30190 16056 30196 16108
rect 30248 16096 30254 16108
rect 31573 16099 31631 16105
rect 31573 16096 31585 16099
rect 30248 16068 31585 16096
rect 30248 16056 30254 16068
rect 31573 16065 31585 16068
rect 31619 16065 31631 16099
rect 31573 16059 31631 16065
rect 32677 16099 32735 16105
rect 32677 16065 32689 16099
rect 32723 16065 32735 16099
rect 32677 16059 32735 16065
rect 18509 16031 18567 16037
rect 18509 15997 18521 16031
rect 18555 16028 18567 16031
rect 18555 16000 19196 16028
rect 18555 15997 18567 16000
rect 18509 15991 18567 15997
rect 18598 15960 18604 15972
rect 10781 15923 10839 15929
rect 10888 15932 15976 15960
rect 16960 15932 18604 15960
rect 6270 15852 6276 15904
rect 6328 15892 6334 15904
rect 9401 15895 9459 15901
rect 9401 15892 9413 15895
rect 6328 15864 9413 15892
rect 6328 15852 6334 15864
rect 9401 15861 9413 15864
rect 9447 15861 9459 15895
rect 9401 15855 9459 15861
rect 9490 15852 9496 15904
rect 9548 15892 9554 15904
rect 10888 15892 10916 15932
rect 9548 15864 10916 15892
rect 9548 15852 9554 15864
rect 11146 15852 11152 15904
rect 11204 15852 11210 15904
rect 11701 15895 11759 15901
rect 11701 15861 11713 15895
rect 11747 15892 11759 15895
rect 12066 15892 12072 15904
rect 11747 15864 12072 15892
rect 11747 15861 11759 15864
rect 11701 15855 11759 15861
rect 12066 15852 12072 15864
rect 12124 15892 12130 15904
rect 14826 15892 14832 15904
rect 12124 15864 14832 15892
rect 12124 15852 12130 15864
rect 14826 15852 14832 15864
rect 14884 15852 14890 15904
rect 15565 15895 15623 15901
rect 15565 15861 15577 15895
rect 15611 15892 15623 15895
rect 15838 15892 15844 15904
rect 15611 15864 15844 15892
rect 15611 15861 15623 15864
rect 15565 15855 15623 15861
rect 15838 15852 15844 15864
rect 15896 15852 15902 15904
rect 15948 15892 15976 15932
rect 18598 15920 18604 15932
rect 18656 15920 18662 15972
rect 17037 15895 17095 15901
rect 17037 15892 17049 15895
rect 15948 15864 17049 15892
rect 17037 15861 17049 15864
rect 17083 15892 17095 15895
rect 17218 15892 17224 15904
rect 17083 15864 17224 15892
rect 17083 15861 17095 15864
rect 17037 15855 17095 15861
rect 17218 15852 17224 15864
rect 17276 15852 17282 15904
rect 17589 15895 17647 15901
rect 17589 15861 17601 15895
rect 17635 15892 17647 15895
rect 17862 15892 17868 15904
rect 17635 15864 17868 15892
rect 17635 15861 17647 15864
rect 17589 15855 17647 15861
rect 17862 15852 17868 15864
rect 17920 15852 17926 15904
rect 17954 15852 17960 15904
rect 18012 15892 18018 15904
rect 18506 15892 18512 15904
rect 18012 15864 18512 15892
rect 18012 15852 18018 15864
rect 18506 15852 18512 15864
rect 18564 15852 18570 15904
rect 19168 15892 19196 16000
rect 19334 15988 19340 16040
rect 19392 16028 19398 16040
rect 19392 16000 22094 16028
rect 19392 15988 19398 16000
rect 20809 15963 20867 15969
rect 20809 15929 20821 15963
rect 20855 15960 20867 15963
rect 22066 15960 22094 16000
rect 23566 15988 23572 16040
rect 23624 15988 23630 16040
rect 23753 16031 23811 16037
rect 23753 15997 23765 16031
rect 23799 16028 23811 16031
rect 26418 16028 26424 16040
rect 23799 16000 26424 16028
rect 23799 15997 23811 16000
rect 23753 15991 23811 15997
rect 23768 15960 23796 15991
rect 26418 15988 26424 16000
rect 26476 15988 26482 16040
rect 27709 16031 27767 16037
rect 27709 15997 27721 16031
rect 27755 15997 27767 16031
rect 27709 15991 27767 15997
rect 27157 15963 27215 15969
rect 27157 15960 27169 15963
rect 20855 15932 21864 15960
rect 22066 15932 23796 15960
rect 25884 15932 27169 15960
rect 20855 15929 20867 15932
rect 20809 15923 20867 15929
rect 20990 15892 20996 15904
rect 19168 15864 20996 15892
rect 20990 15852 20996 15864
rect 21048 15852 21054 15904
rect 21836 15892 21864 15932
rect 22278 15892 22284 15904
rect 21836 15864 22284 15892
rect 22278 15852 22284 15864
rect 22336 15892 22342 15904
rect 22554 15892 22560 15904
rect 22336 15864 22560 15892
rect 22336 15852 22342 15864
rect 22554 15852 22560 15864
rect 22612 15852 22618 15904
rect 22646 15852 22652 15904
rect 22704 15852 22710 15904
rect 23934 15852 23940 15904
rect 23992 15892 23998 15904
rect 24121 15895 24179 15901
rect 24121 15892 24133 15895
rect 23992 15864 24133 15892
rect 23992 15852 23998 15864
rect 24121 15861 24133 15864
rect 24167 15861 24179 15895
rect 24121 15855 24179 15861
rect 24394 15852 24400 15904
rect 24452 15892 24458 15904
rect 25884 15892 25912 15932
rect 27157 15929 27169 15932
rect 27203 15929 27215 15963
rect 27157 15923 27215 15929
rect 27338 15920 27344 15972
rect 27396 15960 27402 15972
rect 27724 15960 27752 15991
rect 28718 15988 28724 16040
rect 28776 16028 28782 16040
rect 30834 16028 30840 16040
rect 28776 16000 30840 16028
rect 28776 15988 28782 16000
rect 30834 15988 30840 16000
rect 30892 15988 30898 16040
rect 31205 16031 31263 16037
rect 31205 15997 31217 16031
rect 31251 15997 31263 16031
rect 31205 15991 31263 15997
rect 27396 15932 27752 15960
rect 27396 15920 27402 15932
rect 30374 15920 30380 15972
rect 30432 15960 30438 15972
rect 30561 15963 30619 15969
rect 30561 15960 30573 15963
rect 30432 15932 30573 15960
rect 30432 15920 30438 15932
rect 30561 15929 30573 15932
rect 30607 15929 30619 15963
rect 30561 15923 30619 15929
rect 31110 15920 31116 15972
rect 31168 15960 31174 15972
rect 31220 15960 31248 15991
rect 31168 15932 31248 15960
rect 32692 15960 32720 16059
rect 33870 16056 33876 16108
rect 33928 16056 33934 16108
rect 36354 16056 36360 16108
rect 36412 16056 36418 16108
rect 37182 16096 37188 16108
rect 36478 16068 37188 16096
rect 37182 16056 37188 16068
rect 37240 16096 37246 16108
rect 37829 16099 37887 16105
rect 37829 16096 37841 16099
rect 37240 16068 37841 16096
rect 37240 16056 37246 16068
rect 37829 16065 37841 16068
rect 37875 16065 37887 16099
rect 37829 16059 37887 16065
rect 39758 16056 39764 16108
rect 39816 16096 39822 16108
rect 42242 16096 42248 16108
rect 39816 16068 42248 16096
rect 39816 16056 39822 16068
rect 42242 16056 42248 16068
rect 42300 16056 42306 16108
rect 42613 16099 42671 16105
rect 42613 16065 42625 16099
rect 42659 16065 42671 16099
rect 42613 16059 42671 16065
rect 48777 16099 48835 16105
rect 48777 16065 48789 16099
rect 48823 16096 48835 16099
rect 49050 16096 49056 16108
rect 48823 16068 49056 16096
rect 48823 16065 48835 16068
rect 48777 16059 48835 16065
rect 32950 15988 32956 16040
rect 33008 15988 33014 16040
rect 34146 15988 34152 16040
rect 34204 15988 34210 16040
rect 34882 15988 34888 16040
rect 34940 16028 34946 16040
rect 35069 16031 35127 16037
rect 35069 16028 35081 16031
rect 34940 16000 35081 16028
rect 34940 15988 34946 16000
rect 35069 15997 35081 16000
rect 35115 15997 35127 16031
rect 35069 15991 35127 15997
rect 35342 15988 35348 16040
rect 35400 15988 35406 16040
rect 35434 15988 35440 16040
rect 35492 16028 35498 16040
rect 36372 16028 36400 16056
rect 36817 16031 36875 16037
rect 36817 16028 36829 16031
rect 35492 16000 36829 16028
rect 35492 15988 35498 16000
rect 36817 15997 36829 16000
rect 36863 16028 36875 16031
rect 36998 16028 37004 16040
rect 36863 16000 37004 16028
rect 36863 15997 36875 16000
rect 36817 15991 36875 15997
rect 36998 15988 37004 16000
rect 37056 15988 37062 16040
rect 37458 15988 37464 16040
rect 37516 16028 37522 16040
rect 38197 16031 38255 16037
rect 38197 16028 38209 16031
rect 37516 16000 38209 16028
rect 37516 15988 37522 16000
rect 38197 15997 38209 16000
rect 38243 15997 38255 16031
rect 38197 15991 38255 15997
rect 41046 15988 41052 16040
rect 41104 15988 41110 16040
rect 33778 15960 33784 15972
rect 32692 15932 33784 15960
rect 31168 15920 31174 15932
rect 33778 15920 33784 15932
rect 33836 15960 33842 15972
rect 33836 15932 34652 15960
rect 33836 15920 33842 15932
rect 24452 15864 25912 15892
rect 32309 15895 32367 15901
rect 24452 15852 24458 15864
rect 32309 15861 32321 15895
rect 32355 15892 32367 15895
rect 33410 15892 33416 15904
rect 32355 15864 33416 15892
rect 32355 15861 32367 15864
rect 32309 15855 32367 15861
rect 33410 15852 33416 15864
rect 33468 15852 33474 15904
rect 33502 15852 33508 15904
rect 33560 15852 33566 15904
rect 34624 15892 34652 15932
rect 36354 15920 36360 15972
rect 36412 15960 36418 15972
rect 37277 15963 37335 15969
rect 37277 15960 37289 15963
rect 36412 15932 37289 15960
rect 36412 15920 36418 15932
rect 37277 15929 37289 15932
rect 37323 15960 37335 15963
rect 37642 15960 37648 15972
rect 37323 15932 37648 15960
rect 37323 15929 37335 15932
rect 37277 15923 37335 15929
rect 37642 15920 37648 15932
rect 37700 15960 37706 15972
rect 37700 15932 37964 15960
rect 37700 15920 37706 15932
rect 36372 15892 36400 15920
rect 34624 15864 36400 15892
rect 37936 15892 37964 15932
rect 39850 15920 39856 15972
rect 39908 15960 39914 15972
rect 40497 15963 40555 15969
rect 40497 15960 40509 15963
rect 39908 15932 40509 15960
rect 39908 15920 39914 15932
rect 40497 15929 40509 15932
rect 40543 15929 40555 15963
rect 42628 15960 42656 16059
rect 49050 16056 49056 16068
rect 49108 16056 49114 16108
rect 40497 15923 40555 15929
rect 41386 15932 42656 15960
rect 38562 15892 38568 15904
rect 37936 15864 38568 15892
rect 38562 15852 38568 15864
rect 38620 15852 38626 15904
rect 39574 15852 39580 15904
rect 39632 15892 39638 15904
rect 39945 15895 40003 15901
rect 39945 15892 39957 15895
rect 39632 15864 39957 15892
rect 39632 15852 39638 15864
rect 39945 15861 39957 15864
rect 39991 15892 40003 15895
rect 41386 15892 41414 15932
rect 39991 15864 41414 15892
rect 39991 15861 40003 15864
rect 39945 15855 40003 15861
rect 42334 15852 42340 15904
rect 42392 15892 42398 15904
rect 43257 15895 43315 15901
rect 43257 15892 43269 15895
rect 42392 15864 43269 15892
rect 42392 15852 42398 15864
rect 43257 15861 43269 15864
rect 43303 15861 43315 15895
rect 43257 15855 43315 15861
rect 48590 15852 48596 15904
rect 48648 15892 48654 15904
rect 49237 15895 49295 15901
rect 49237 15892 49249 15895
rect 48648 15864 49249 15892
rect 48648 15852 48654 15864
rect 49237 15861 49249 15864
rect 49283 15861 49295 15895
rect 49237 15855 49295 15861
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 3510 15648 3516 15700
rect 3568 15688 3574 15700
rect 9861 15691 9919 15697
rect 9861 15688 9873 15691
rect 3568 15660 9873 15688
rect 3568 15648 3574 15660
rect 9861 15657 9873 15660
rect 9907 15657 9919 15691
rect 11238 15688 11244 15700
rect 9861 15651 9919 15657
rect 10152 15660 11244 15688
rect 10152 15632 10180 15660
rect 11238 15648 11244 15660
rect 11296 15648 11302 15700
rect 11514 15648 11520 15700
rect 11572 15688 11578 15700
rect 12989 15691 13047 15697
rect 12989 15688 13001 15691
rect 11572 15660 13001 15688
rect 11572 15648 11578 15660
rect 12989 15657 13001 15660
rect 13035 15657 13047 15691
rect 12989 15651 13047 15657
rect 14550 15648 14556 15700
rect 14608 15688 14614 15700
rect 14921 15691 14979 15697
rect 14921 15688 14933 15691
rect 14608 15660 14933 15688
rect 14608 15648 14614 15660
rect 14921 15657 14933 15660
rect 14967 15657 14979 15691
rect 14921 15651 14979 15657
rect 15746 15648 15752 15700
rect 15804 15688 15810 15700
rect 18141 15691 18199 15697
rect 15804 15660 18092 15688
rect 15804 15648 15810 15660
rect 9766 15580 9772 15632
rect 9824 15620 9830 15632
rect 10134 15620 10140 15632
rect 9824 15592 10140 15620
rect 9824 15580 9830 15592
rect 10134 15580 10140 15592
rect 10192 15580 10198 15632
rect 12342 15580 12348 15632
rect 12400 15620 12406 15632
rect 15381 15623 15439 15629
rect 15381 15620 15393 15623
rect 12400 15592 15393 15620
rect 12400 15580 12406 15592
rect 15381 15589 15393 15592
rect 15427 15589 15439 15623
rect 16853 15623 16911 15629
rect 15381 15583 15439 15589
rect 15764 15592 15976 15620
rect 1302 15512 1308 15564
rect 1360 15552 1366 15564
rect 2041 15555 2099 15561
rect 2041 15552 2053 15555
rect 1360 15524 2053 15552
rect 1360 15512 1366 15524
rect 2041 15521 2053 15524
rect 2087 15521 2099 15555
rect 2041 15515 2099 15521
rect 10778 15512 10784 15564
rect 10836 15512 10842 15564
rect 11057 15555 11115 15561
rect 11057 15521 11069 15555
rect 11103 15552 11115 15555
rect 12529 15555 12587 15561
rect 11103 15524 12480 15552
rect 11103 15521 11115 15524
rect 11057 15515 11115 15521
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15484 1823 15487
rect 9674 15484 9680 15496
rect 1811 15456 9680 15484
rect 1811 15453 1823 15456
rect 1765 15447 1823 15453
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 10045 15487 10103 15493
rect 10045 15453 10057 15487
rect 10091 15484 10103 15487
rect 10686 15484 10692 15496
rect 10091 15456 10692 15484
rect 10091 15453 10103 15456
rect 10045 15447 10103 15453
rect 10686 15444 10692 15456
rect 10744 15444 10750 15496
rect 12452 15484 12480 15524
rect 12529 15521 12541 15555
rect 12575 15552 12587 15555
rect 12618 15552 12624 15564
rect 12575 15524 12624 15552
rect 12575 15521 12587 15524
rect 12529 15515 12587 15521
rect 12618 15512 12624 15524
rect 12676 15552 12682 15564
rect 13541 15555 13599 15561
rect 13541 15552 13553 15555
rect 12676 15524 13553 15552
rect 12676 15512 12682 15524
rect 13541 15521 13553 15524
rect 13587 15521 13599 15555
rect 15102 15552 15108 15564
rect 13541 15515 13599 15521
rect 13740 15524 15108 15552
rect 13740 15496 13768 15524
rect 15102 15512 15108 15524
rect 15160 15552 15166 15564
rect 15764 15552 15792 15592
rect 15160 15524 15792 15552
rect 15160 15512 15166 15524
rect 15838 15512 15844 15564
rect 15896 15512 15902 15564
rect 15948 15561 15976 15592
rect 16853 15589 16865 15623
rect 16899 15620 16911 15623
rect 17954 15620 17960 15632
rect 16899 15592 17960 15620
rect 16899 15589 16911 15592
rect 16853 15583 16911 15589
rect 17954 15580 17960 15592
rect 18012 15580 18018 15632
rect 15933 15555 15991 15561
rect 15933 15521 15945 15555
rect 15979 15521 15991 15555
rect 15933 15515 15991 15521
rect 17494 15512 17500 15564
rect 17552 15512 17558 15564
rect 18064 15552 18092 15660
rect 18141 15657 18153 15691
rect 18187 15688 18199 15691
rect 18414 15688 18420 15700
rect 18187 15660 18420 15688
rect 18187 15657 18199 15660
rect 18141 15651 18199 15657
rect 18414 15648 18420 15660
rect 18472 15648 18478 15700
rect 18598 15648 18604 15700
rect 18656 15688 18662 15700
rect 19797 15691 19855 15697
rect 19797 15688 19809 15691
rect 18656 15660 19809 15688
rect 18656 15648 18662 15660
rect 19797 15657 19809 15660
rect 19843 15657 19855 15691
rect 19797 15651 19855 15657
rect 20806 15648 20812 15700
rect 20864 15688 20870 15700
rect 21177 15691 21235 15697
rect 21177 15688 21189 15691
rect 20864 15660 21189 15688
rect 20864 15648 20870 15660
rect 21177 15657 21189 15660
rect 21223 15657 21235 15691
rect 21177 15651 21235 15657
rect 22646 15648 22652 15700
rect 22704 15688 22710 15700
rect 26142 15688 26148 15700
rect 22704 15660 26148 15688
rect 22704 15648 22710 15660
rect 26142 15648 26148 15660
rect 26200 15648 26206 15700
rect 26786 15688 26792 15700
rect 26252 15660 26792 15688
rect 21910 15620 21916 15632
rect 18708 15592 21916 15620
rect 18708 15561 18736 15592
rect 21910 15580 21916 15592
rect 21968 15580 21974 15632
rect 22002 15580 22008 15632
rect 22060 15620 22066 15632
rect 22060 15580 22094 15620
rect 22370 15580 22376 15632
rect 22428 15580 22434 15632
rect 22554 15580 22560 15632
rect 22612 15620 22618 15632
rect 24578 15620 24584 15632
rect 22612 15592 24584 15620
rect 22612 15580 22618 15592
rect 24578 15580 24584 15592
rect 24636 15580 24642 15632
rect 24673 15623 24731 15629
rect 24673 15589 24685 15623
rect 24719 15589 24731 15623
rect 24673 15583 24731 15589
rect 18693 15555 18751 15561
rect 18693 15552 18705 15555
rect 18064 15524 18705 15552
rect 18693 15521 18705 15524
rect 18739 15521 18751 15555
rect 18693 15515 18751 15521
rect 19334 15512 19340 15564
rect 19392 15512 19398 15564
rect 20346 15512 20352 15564
rect 20404 15512 20410 15564
rect 20898 15512 20904 15564
rect 20956 15512 20962 15564
rect 21726 15512 21732 15564
rect 21784 15512 21790 15564
rect 22066 15552 22094 15580
rect 22066 15524 23336 15552
rect 13722 15484 13728 15496
rect 12452 15456 13728 15484
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 14274 15444 14280 15496
rect 14332 15444 14338 15496
rect 17126 15444 17132 15496
rect 17184 15484 17190 15496
rect 17221 15487 17279 15493
rect 17221 15484 17233 15487
rect 17184 15456 17233 15484
rect 17184 15444 17190 15456
rect 17221 15453 17233 15456
rect 17267 15453 17279 15487
rect 17221 15447 17279 15453
rect 17678 15444 17684 15496
rect 17736 15484 17742 15496
rect 18509 15487 18567 15493
rect 18509 15484 18521 15487
rect 17736 15456 18521 15484
rect 17736 15444 17742 15456
rect 18509 15453 18521 15456
rect 18555 15453 18567 15487
rect 18509 15447 18567 15453
rect 18601 15487 18659 15493
rect 18601 15453 18613 15487
rect 18647 15484 18659 15487
rect 18966 15484 18972 15496
rect 18647 15456 18972 15484
rect 18647 15453 18659 15456
rect 18601 15447 18659 15453
rect 18966 15444 18972 15456
rect 19024 15484 19030 15496
rect 19352 15484 19380 15512
rect 19024 15456 19380 15484
rect 19024 15444 19030 15456
rect 22554 15444 22560 15496
rect 22612 15444 22618 15496
rect 6549 15419 6607 15425
rect 6549 15385 6561 15419
rect 6595 15416 6607 15419
rect 6914 15416 6920 15428
rect 6595 15388 6920 15416
rect 6595 15385 6607 15388
rect 6549 15379 6607 15385
rect 6914 15376 6920 15388
rect 6972 15416 6978 15428
rect 7650 15416 7656 15428
rect 6972 15388 7656 15416
rect 6972 15376 6978 15388
rect 7650 15376 7656 15388
rect 7708 15376 7714 15428
rect 9398 15376 9404 15428
rect 9456 15376 9462 15428
rect 11146 15376 11152 15428
rect 11204 15416 11210 15428
rect 11514 15416 11520 15428
rect 11204 15388 11520 15416
rect 11204 15376 11210 15388
rect 11514 15376 11520 15388
rect 11572 15376 11578 15428
rect 13357 15419 13415 15425
rect 13357 15385 13369 15419
rect 13403 15416 13415 15419
rect 15562 15416 15568 15428
rect 13403 15388 15568 15416
rect 13403 15385 13415 15388
rect 13357 15379 13415 15385
rect 15562 15376 15568 15388
rect 15620 15376 15626 15428
rect 15749 15419 15807 15425
rect 15749 15385 15761 15419
rect 15795 15416 15807 15419
rect 18414 15416 18420 15428
rect 15795 15388 18420 15416
rect 15795 15385 15807 15388
rect 15749 15379 15807 15385
rect 18414 15376 18420 15388
rect 18472 15376 18478 15428
rect 19242 15376 19248 15428
rect 19300 15416 19306 15428
rect 19429 15419 19487 15425
rect 19429 15416 19441 15419
rect 19300 15388 19441 15416
rect 19300 15376 19306 15388
rect 19429 15385 19441 15388
rect 19475 15385 19487 15419
rect 19429 15379 19487 15385
rect 20257 15419 20315 15425
rect 20257 15385 20269 15419
rect 20303 15416 20315 15419
rect 20303 15388 23060 15416
rect 20303 15385 20315 15388
rect 20257 15379 20315 15385
rect 6638 15308 6644 15360
rect 6696 15308 6702 15360
rect 8662 15308 8668 15360
rect 8720 15348 8726 15360
rect 9030 15348 9036 15360
rect 8720 15320 9036 15348
rect 8720 15308 8726 15320
rect 9030 15308 9036 15320
rect 9088 15308 9094 15360
rect 9490 15308 9496 15360
rect 9548 15348 9554 15360
rect 10226 15348 10232 15360
rect 9548 15320 10232 15348
rect 9548 15308 9554 15320
rect 10226 15308 10232 15320
rect 10284 15308 10290 15360
rect 10505 15351 10563 15357
rect 10505 15317 10517 15351
rect 10551 15348 10563 15351
rect 12066 15348 12072 15360
rect 10551 15320 12072 15348
rect 10551 15317 10563 15320
rect 10505 15311 10563 15317
rect 12066 15308 12072 15320
rect 12124 15308 12130 15360
rect 13449 15351 13507 15357
rect 13449 15317 13461 15351
rect 13495 15348 13507 15351
rect 14550 15348 14556 15360
rect 13495 15320 14556 15348
rect 13495 15317 13507 15320
rect 13449 15311 13507 15317
rect 14550 15308 14556 15320
rect 14608 15308 14614 15360
rect 16577 15351 16635 15357
rect 16577 15317 16589 15351
rect 16623 15348 16635 15351
rect 16850 15348 16856 15360
rect 16623 15320 16856 15348
rect 16623 15317 16635 15320
rect 16577 15311 16635 15317
rect 16850 15308 16856 15320
rect 16908 15308 16914 15360
rect 17313 15351 17371 15357
rect 17313 15317 17325 15351
rect 17359 15348 17371 15351
rect 17586 15348 17592 15360
rect 17359 15320 17592 15348
rect 17359 15317 17371 15320
rect 17313 15311 17371 15317
rect 17586 15308 17592 15320
rect 17644 15308 17650 15360
rect 19886 15308 19892 15360
rect 19944 15348 19950 15360
rect 20165 15351 20223 15357
rect 20165 15348 20177 15351
rect 19944 15320 20177 15348
rect 19944 15308 19950 15320
rect 20165 15317 20177 15320
rect 20211 15317 20223 15351
rect 20165 15311 20223 15317
rect 20530 15308 20536 15360
rect 20588 15348 20594 15360
rect 21266 15348 21272 15360
rect 20588 15320 21272 15348
rect 20588 15308 20594 15320
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 21542 15308 21548 15360
rect 21600 15308 21606 15360
rect 21634 15308 21640 15360
rect 21692 15308 21698 15360
rect 23032 15357 23060 15388
rect 23017 15351 23075 15357
rect 23017 15317 23029 15351
rect 23063 15317 23075 15351
rect 23308 15348 23336 15524
rect 23382 15512 23388 15564
rect 23440 15552 23446 15564
rect 23569 15555 23627 15561
rect 23569 15552 23581 15555
rect 23440 15524 23581 15552
rect 23440 15512 23446 15524
rect 23569 15521 23581 15524
rect 23615 15521 23627 15555
rect 24688 15552 24716 15583
rect 24762 15580 24768 15632
rect 24820 15620 24826 15632
rect 24820 15592 25360 15620
rect 24820 15580 24826 15592
rect 23569 15515 23627 15521
rect 23952 15524 24716 15552
rect 23477 15487 23535 15493
rect 23477 15453 23489 15487
rect 23523 15484 23535 15487
rect 23842 15484 23848 15496
rect 23523 15456 23848 15484
rect 23523 15453 23535 15456
rect 23477 15447 23535 15453
rect 23842 15444 23848 15456
rect 23900 15444 23906 15496
rect 23385 15419 23443 15425
rect 23385 15385 23397 15419
rect 23431 15416 23443 15419
rect 23952 15416 23980 15524
rect 25130 15512 25136 15564
rect 25188 15512 25194 15564
rect 25332 15561 25360 15592
rect 25317 15555 25375 15561
rect 25317 15521 25329 15555
rect 25363 15552 25375 15555
rect 26252 15552 26280 15660
rect 26786 15648 26792 15660
rect 26844 15648 26850 15700
rect 26970 15648 26976 15700
rect 27028 15648 27034 15700
rect 27522 15648 27528 15700
rect 27580 15688 27586 15700
rect 28813 15691 28871 15697
rect 28813 15688 28825 15691
rect 27580 15660 28825 15688
rect 27580 15648 27586 15660
rect 28813 15657 28825 15660
rect 28859 15688 28871 15691
rect 31846 15688 31852 15700
rect 28859 15660 31852 15688
rect 28859 15657 28871 15660
rect 28813 15651 28871 15657
rect 31846 15648 31852 15660
rect 31904 15648 31910 15700
rect 32217 15691 32275 15697
rect 32217 15657 32229 15691
rect 32263 15688 32275 15691
rect 34146 15688 34152 15700
rect 32263 15660 34152 15688
rect 32263 15657 32275 15660
rect 32217 15651 32275 15657
rect 34146 15648 34152 15660
rect 34204 15648 34210 15700
rect 34238 15648 34244 15700
rect 34296 15688 34302 15700
rect 34333 15691 34391 15697
rect 34333 15688 34345 15691
rect 34296 15660 34345 15688
rect 34296 15648 34302 15660
rect 34333 15657 34345 15660
rect 34379 15657 34391 15691
rect 37642 15688 37648 15700
rect 34333 15651 34391 15657
rect 34808 15660 37648 15688
rect 27062 15620 27068 15632
rect 26344 15592 27068 15620
rect 26344 15561 26372 15592
rect 27062 15580 27068 15592
rect 27120 15580 27126 15632
rect 27430 15580 27436 15632
rect 27488 15620 27494 15632
rect 28445 15623 28503 15629
rect 28445 15620 28457 15623
rect 27488 15592 28457 15620
rect 27488 15580 27494 15592
rect 28445 15589 28457 15592
rect 28491 15620 28503 15623
rect 28626 15620 28632 15632
rect 28491 15592 28632 15620
rect 28491 15589 28503 15592
rect 28445 15583 28503 15589
rect 28626 15580 28632 15592
rect 28684 15580 28690 15632
rect 28721 15623 28779 15629
rect 28721 15589 28733 15623
rect 28767 15620 28779 15623
rect 28902 15620 28908 15632
rect 28767 15592 28908 15620
rect 28767 15589 28779 15592
rect 28721 15583 28779 15589
rect 25363 15524 26280 15552
rect 26329 15555 26387 15561
rect 25363 15521 25375 15524
rect 25317 15515 25375 15521
rect 26329 15521 26341 15555
rect 26375 15521 26387 15555
rect 26329 15515 26387 15521
rect 26418 15512 26424 15564
rect 26476 15512 26482 15564
rect 26602 15512 26608 15564
rect 26660 15552 26666 15564
rect 27985 15555 28043 15561
rect 27985 15552 27997 15555
rect 26660 15524 27997 15552
rect 26660 15512 26666 15524
rect 27985 15521 27997 15524
rect 28031 15521 28043 15555
rect 27985 15515 28043 15521
rect 28534 15512 28540 15564
rect 28592 15552 28598 15564
rect 28736 15552 28764 15583
rect 28902 15580 28908 15592
rect 28960 15580 28966 15632
rect 32306 15580 32312 15632
rect 32364 15620 32370 15632
rect 33042 15620 33048 15632
rect 32364 15592 33048 15620
rect 32364 15580 32370 15592
rect 33042 15580 33048 15592
rect 33100 15580 33106 15632
rect 28592 15524 28764 15552
rect 28592 15512 28598 15524
rect 29178 15512 29184 15564
rect 29236 15552 29242 15564
rect 30745 15555 30803 15561
rect 30745 15552 30757 15555
rect 29236 15524 30757 15552
rect 29236 15512 29242 15524
rect 30745 15521 30757 15524
rect 30791 15521 30803 15555
rect 30745 15515 30803 15521
rect 32858 15512 32864 15564
rect 32916 15552 32922 15564
rect 33137 15555 33195 15561
rect 33137 15552 33149 15555
rect 32916 15524 33149 15552
rect 32916 15512 32922 15524
rect 33137 15521 33149 15524
rect 33183 15521 33195 15555
rect 33137 15515 33195 15521
rect 33321 15555 33379 15561
rect 33321 15521 33333 15555
rect 33367 15552 33379 15555
rect 34330 15552 34336 15564
rect 33367 15524 34336 15552
rect 33367 15521 33379 15524
rect 33321 15515 33379 15521
rect 34330 15512 34336 15524
rect 34388 15512 34394 15564
rect 27706 15444 27712 15496
rect 27764 15484 27770 15496
rect 27893 15487 27951 15493
rect 27893 15484 27905 15487
rect 27764 15456 27905 15484
rect 27764 15444 27770 15456
rect 27893 15453 27905 15456
rect 27939 15484 27951 15487
rect 28718 15484 28724 15496
rect 27939 15456 28724 15484
rect 27939 15453 27951 15456
rect 27893 15447 27951 15453
rect 28718 15444 28724 15456
rect 28776 15484 28782 15496
rect 29273 15487 29331 15493
rect 29273 15484 29285 15487
rect 28776 15456 29285 15484
rect 28776 15444 28782 15456
rect 29273 15453 29285 15456
rect 29319 15453 29331 15487
rect 29273 15447 29331 15453
rect 30282 15444 30288 15496
rect 30340 15484 30346 15496
rect 30469 15487 30527 15493
rect 30469 15484 30481 15487
rect 30340 15456 30481 15484
rect 30340 15444 30346 15456
rect 30469 15453 30481 15456
rect 30515 15453 30527 15487
rect 30469 15447 30527 15453
rect 32030 15444 32036 15496
rect 32088 15484 32094 15496
rect 32766 15484 32772 15496
rect 32088 15456 32772 15484
rect 32088 15444 32094 15456
rect 32766 15444 32772 15456
rect 32824 15444 32830 15496
rect 33873 15487 33931 15493
rect 33873 15453 33885 15487
rect 33919 15484 33931 15487
rect 34808 15484 34836 15660
rect 37642 15648 37648 15660
rect 37700 15648 37706 15700
rect 38000 15691 38058 15697
rect 38000 15657 38012 15691
rect 38046 15688 38058 15691
rect 42150 15688 42156 15700
rect 38046 15660 42156 15688
rect 38046 15657 38058 15660
rect 38000 15651 38058 15657
rect 42150 15648 42156 15660
rect 42208 15648 42214 15700
rect 48958 15648 48964 15700
rect 49016 15688 49022 15700
rect 49145 15691 49203 15697
rect 49145 15688 49157 15691
rect 49016 15660 49157 15688
rect 49016 15648 49022 15660
rect 49145 15657 49157 15660
rect 49191 15657 49203 15691
rect 49145 15651 49203 15657
rect 37182 15620 37188 15632
rect 36280 15592 37188 15620
rect 35158 15512 35164 15564
rect 35216 15512 35222 15564
rect 33919 15456 34836 15484
rect 33919 15453 33931 15456
rect 33873 15447 33931 15453
rect 34882 15444 34888 15496
rect 34940 15444 34946 15496
rect 36170 15444 36176 15496
rect 36228 15484 36234 15496
rect 36280 15484 36308 15592
rect 37182 15580 37188 15592
rect 37240 15580 37246 15632
rect 39482 15580 39488 15632
rect 39540 15580 39546 15632
rect 41322 15580 41328 15632
rect 41380 15620 41386 15632
rect 41785 15623 41843 15629
rect 41785 15620 41797 15623
rect 41380 15592 41797 15620
rect 41380 15580 41386 15592
rect 41785 15589 41797 15592
rect 41831 15589 41843 15623
rect 41785 15583 41843 15589
rect 40037 15555 40095 15561
rect 40037 15552 40049 15555
rect 37752 15524 40049 15552
rect 37277 15487 37335 15493
rect 37277 15484 37289 15487
rect 36228 15470 36308 15484
rect 36228 15456 36294 15470
rect 36464 15456 37289 15484
rect 36228 15444 36234 15456
rect 23431 15388 23980 15416
rect 24596 15388 26648 15416
rect 23431 15385 23443 15388
rect 23385 15379 23443 15385
rect 24596 15348 24624 15388
rect 23308 15320 24624 15348
rect 25041 15351 25099 15357
rect 23017 15311 23075 15317
rect 25041 15317 25053 15351
rect 25087 15348 25099 15351
rect 25406 15348 25412 15360
rect 25087 15320 25412 15348
rect 25087 15317 25099 15320
rect 25041 15311 25099 15317
rect 25406 15308 25412 15320
rect 25464 15308 25470 15360
rect 25866 15308 25872 15360
rect 25924 15308 25930 15360
rect 26234 15308 26240 15360
rect 26292 15308 26298 15360
rect 26620 15348 26648 15388
rect 26694 15376 26700 15428
rect 26752 15416 26758 15428
rect 27801 15419 27859 15425
rect 27801 15416 27813 15419
rect 26752 15388 27813 15416
rect 26752 15376 26758 15388
rect 27801 15385 27813 15388
rect 27847 15416 27859 15419
rect 28997 15419 29055 15425
rect 28997 15416 29009 15419
rect 27847 15388 29009 15416
rect 27847 15385 27859 15388
rect 27801 15379 27859 15385
rect 28997 15385 29009 15388
rect 29043 15416 29055 15419
rect 31018 15416 31024 15428
rect 29043 15388 31024 15416
rect 29043 15385 29055 15388
rect 28997 15379 29055 15385
rect 31018 15376 31024 15388
rect 31076 15376 31082 15428
rect 34238 15416 34244 15428
rect 31970 15388 34244 15416
rect 34238 15376 34244 15388
rect 34296 15376 34302 15428
rect 26786 15348 26792 15360
rect 26620 15320 26792 15348
rect 26786 15308 26792 15320
rect 26844 15308 26850 15360
rect 26970 15308 26976 15360
rect 27028 15348 27034 15360
rect 27065 15351 27123 15357
rect 27065 15348 27077 15351
rect 27028 15320 27077 15348
rect 27028 15308 27034 15320
rect 27065 15317 27077 15320
rect 27111 15317 27123 15351
rect 27065 15311 27123 15317
rect 27430 15308 27436 15360
rect 27488 15308 27494 15360
rect 29825 15351 29883 15357
rect 29825 15317 29837 15351
rect 29871 15348 29883 15351
rect 31110 15348 31116 15360
rect 29871 15320 31116 15348
rect 29871 15317 29883 15320
rect 29825 15311 29883 15317
rect 31110 15308 31116 15320
rect 31168 15308 31174 15360
rect 32677 15351 32735 15357
rect 32677 15317 32689 15351
rect 32723 15348 32735 15351
rect 32766 15348 32772 15360
rect 32723 15320 32772 15348
rect 32723 15317 32735 15320
rect 32677 15311 32735 15317
rect 32766 15308 32772 15320
rect 32824 15308 32830 15360
rect 33042 15308 33048 15360
rect 33100 15348 33106 15360
rect 35250 15348 35256 15360
rect 33100 15320 35256 15348
rect 33100 15308 33106 15320
rect 35250 15308 35256 15320
rect 35308 15308 35314 15360
rect 36078 15308 36084 15360
rect 36136 15348 36142 15360
rect 36464 15348 36492 15456
rect 37277 15453 37289 15456
rect 37323 15453 37335 15487
rect 37277 15447 37335 15453
rect 37458 15444 37464 15496
rect 37516 15484 37522 15496
rect 37752 15493 37780 15524
rect 40037 15521 40049 15524
rect 40083 15521 40095 15555
rect 40037 15515 40095 15521
rect 40313 15555 40371 15561
rect 40313 15521 40325 15555
rect 40359 15552 40371 15555
rect 42334 15552 42340 15564
rect 40359 15524 42340 15552
rect 40359 15521 40371 15524
rect 40313 15515 40371 15521
rect 42334 15512 42340 15524
rect 42392 15512 42398 15564
rect 37737 15487 37795 15493
rect 37737 15484 37749 15487
rect 37516 15456 37749 15484
rect 37516 15444 37522 15456
rect 37737 15453 37749 15456
rect 37783 15453 37795 15487
rect 37737 15447 37795 15453
rect 42242 15444 42248 15496
rect 42300 15444 42306 15496
rect 48869 15487 48927 15493
rect 48869 15453 48881 15487
rect 48915 15484 48927 15487
rect 49326 15484 49332 15496
rect 48915 15456 49332 15484
rect 48915 15453 48927 15456
rect 48869 15447 48927 15453
rect 49326 15444 49332 15456
rect 49384 15444 49390 15496
rect 36648 15388 38424 15416
rect 36648 15357 36676 15388
rect 38396 15360 38424 15388
rect 38470 15376 38476 15428
rect 38528 15376 38534 15428
rect 40310 15416 40316 15428
rect 39316 15388 40316 15416
rect 36136 15320 36492 15348
rect 36633 15351 36691 15357
rect 36136 15308 36142 15320
rect 36633 15317 36645 15351
rect 36679 15317 36691 15351
rect 36633 15311 36691 15317
rect 36906 15308 36912 15360
rect 36964 15308 36970 15360
rect 38378 15308 38384 15360
rect 38436 15348 38442 15360
rect 39316 15348 39344 15388
rect 40310 15376 40316 15388
rect 40368 15376 40374 15428
rect 41598 15416 41604 15428
rect 41538 15388 41604 15416
rect 41598 15376 41604 15388
rect 41656 15376 41662 15428
rect 42889 15419 42947 15425
rect 42889 15416 42901 15419
rect 41708 15388 42901 15416
rect 38436 15320 39344 15348
rect 38436 15308 38442 15320
rect 40034 15308 40040 15360
rect 40092 15348 40098 15360
rect 41708 15348 41736 15388
rect 42889 15385 42901 15388
rect 42935 15385 42947 15419
rect 42889 15379 42947 15385
rect 40092 15320 41736 15348
rect 40092 15308 40098 15320
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 9858 15104 9864 15156
rect 9916 15104 9922 15156
rect 10318 15104 10324 15156
rect 10376 15144 10382 15156
rect 11793 15147 11851 15153
rect 11793 15144 11805 15147
rect 10376 15116 11805 15144
rect 10376 15104 10382 15116
rect 11793 15113 11805 15116
rect 11839 15113 11851 15147
rect 11793 15107 11851 15113
rect 12066 15104 12072 15156
rect 12124 15144 12130 15156
rect 12253 15147 12311 15153
rect 12253 15144 12265 15147
rect 12124 15116 12265 15144
rect 12124 15104 12130 15116
rect 12253 15113 12265 15116
rect 12299 15113 12311 15147
rect 12253 15107 12311 15113
rect 12802 15104 12808 15156
rect 12860 15144 12866 15156
rect 14826 15144 14832 15156
rect 12860 15116 14832 15144
rect 12860 15104 12866 15116
rect 14826 15104 14832 15116
rect 14884 15104 14890 15156
rect 14918 15104 14924 15156
rect 14976 15144 14982 15156
rect 15105 15147 15163 15153
rect 15105 15144 15117 15147
rect 14976 15116 15117 15144
rect 14976 15104 14982 15116
rect 15105 15113 15117 15116
rect 15151 15113 15163 15147
rect 15105 15107 15163 15113
rect 8846 15036 8852 15088
rect 8904 15076 8910 15088
rect 9953 15079 10011 15085
rect 9953 15076 9965 15079
rect 8904 15048 9965 15076
rect 8904 15036 8910 15048
rect 9953 15045 9965 15048
rect 9999 15045 10011 15079
rect 9953 15039 10011 15045
rect 11974 15036 11980 15088
rect 12032 15076 12038 15088
rect 12526 15076 12532 15088
rect 12032 15048 12532 15076
rect 12032 15036 12038 15048
rect 12526 15036 12532 15048
rect 12584 15036 12590 15088
rect 13906 15036 13912 15088
rect 13964 15036 13970 15088
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 6638 15008 6644 15020
rect 1811 14980 6644 15008
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 6638 14968 6644 14980
rect 6696 14968 6702 15020
rect 9217 15011 9275 15017
rect 9217 14977 9229 15011
rect 9263 15008 9275 15011
rect 10962 15008 10968 15020
rect 9263 14980 10968 15008
rect 9263 14977 9275 14980
rect 9217 14971 9275 14977
rect 10962 14968 10968 14980
rect 11020 14968 11026 15020
rect 11146 14968 11152 15020
rect 11204 15008 11210 15020
rect 12161 15011 12219 15017
rect 12161 15008 12173 15011
rect 11204 14980 12173 15008
rect 11204 14968 11210 14980
rect 12161 14977 12173 14980
rect 12207 14977 12219 15011
rect 12161 14971 12219 14977
rect 12710 14968 12716 15020
rect 12768 15008 12774 15020
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12768 14980 13001 15008
rect 12768 14968 12774 14980
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 1302 14900 1308 14952
rect 1360 14940 1366 14952
rect 2041 14943 2099 14949
rect 2041 14940 2053 14943
rect 1360 14912 2053 14940
rect 1360 14900 1366 14912
rect 2041 14909 2053 14912
rect 2087 14909 2099 14943
rect 2041 14903 2099 14909
rect 10045 14943 10103 14949
rect 10045 14909 10057 14943
rect 10091 14909 10103 14943
rect 10045 14903 10103 14909
rect 10060 14872 10088 14903
rect 12250 14900 12256 14952
rect 12308 14940 12314 14952
rect 12345 14943 12403 14949
rect 12345 14940 12357 14943
rect 12308 14912 12357 14940
rect 12308 14900 12314 14912
rect 12345 14909 12357 14912
rect 12391 14909 12403 14943
rect 12345 14903 12403 14909
rect 12526 14900 12532 14952
rect 12584 14940 12590 14952
rect 13265 14943 13323 14949
rect 13265 14940 13277 14943
rect 12584 14912 13277 14940
rect 12584 14900 12590 14912
rect 13265 14909 13277 14912
rect 13311 14909 13323 14943
rect 15120 14940 15148 15107
rect 16758 15104 16764 15156
rect 16816 15144 16822 15156
rect 16853 15147 16911 15153
rect 16853 15144 16865 15147
rect 16816 15116 16865 15144
rect 16816 15104 16822 15116
rect 16853 15113 16865 15116
rect 16899 15113 16911 15147
rect 16853 15107 16911 15113
rect 17126 15104 17132 15156
rect 17184 15144 17190 15156
rect 18049 15147 18107 15153
rect 17184 15116 17448 15144
rect 17184 15104 17190 15116
rect 15286 15036 15292 15088
rect 15344 15076 15350 15088
rect 17221 15079 17279 15085
rect 17221 15076 17233 15079
rect 15344 15048 17233 15076
rect 15344 15036 15350 15048
rect 17221 15045 17233 15048
rect 17267 15045 17279 15079
rect 17221 15039 17279 15045
rect 17310 15036 17316 15088
rect 17368 15036 17374 15088
rect 17420 15076 17448 15116
rect 18049 15113 18061 15147
rect 18095 15144 18107 15147
rect 18690 15144 18696 15156
rect 18095 15116 18696 15144
rect 18095 15113 18107 15116
rect 18049 15107 18107 15113
rect 18690 15104 18696 15116
rect 18748 15104 18754 15156
rect 19521 15147 19579 15153
rect 19521 15113 19533 15147
rect 19567 15144 19579 15147
rect 19794 15144 19800 15156
rect 19567 15116 19800 15144
rect 19567 15113 19579 15116
rect 19521 15107 19579 15113
rect 19794 15104 19800 15116
rect 19852 15104 19858 15156
rect 20714 15104 20720 15156
rect 20772 15104 20778 15156
rect 21174 15104 21180 15156
rect 21232 15144 21238 15156
rect 21634 15144 21640 15156
rect 21232 15116 21640 15144
rect 21232 15104 21238 15116
rect 21634 15104 21640 15116
rect 21692 15144 21698 15156
rect 21913 15147 21971 15153
rect 21913 15144 21925 15147
rect 21692 15116 21925 15144
rect 21692 15104 21698 15116
rect 21913 15113 21925 15116
rect 21959 15113 21971 15147
rect 21913 15107 21971 15113
rect 22925 15147 22983 15153
rect 22925 15113 22937 15147
rect 22971 15144 22983 15147
rect 23474 15144 23480 15156
rect 22971 15116 23480 15144
rect 22971 15113 22983 15116
rect 22925 15107 22983 15113
rect 23474 15104 23480 15116
rect 23532 15104 23538 15156
rect 24121 15147 24179 15153
rect 24121 15113 24133 15147
rect 24167 15144 24179 15147
rect 26050 15144 26056 15156
rect 24167 15116 26056 15144
rect 24167 15113 24179 15116
rect 24121 15107 24179 15113
rect 26050 15104 26056 15116
rect 26108 15104 26114 15156
rect 27062 15104 27068 15156
rect 27120 15104 27126 15156
rect 27246 15104 27252 15156
rect 27304 15144 27310 15156
rect 27341 15147 27399 15153
rect 27341 15144 27353 15147
rect 27304 15116 27353 15144
rect 27304 15104 27310 15116
rect 27341 15113 27353 15116
rect 27387 15113 27399 15147
rect 27341 15107 27399 15113
rect 27617 15147 27675 15153
rect 27617 15113 27629 15147
rect 27663 15144 27675 15147
rect 28718 15144 28724 15156
rect 27663 15116 28724 15144
rect 27663 15113 27675 15116
rect 27617 15107 27675 15113
rect 21726 15076 21732 15088
rect 17420 15048 21732 15076
rect 21726 15036 21732 15048
rect 21784 15036 21790 15088
rect 25774 15076 25780 15088
rect 23584 15048 25780 15076
rect 15657 15011 15715 15017
rect 15657 14977 15669 15011
rect 15703 15008 15715 15011
rect 19794 15008 19800 15020
rect 15703 14980 19800 15008
rect 15703 14977 15715 14980
rect 15657 14971 15715 14977
rect 19794 14968 19800 14980
rect 19852 14968 19858 15020
rect 19889 15011 19947 15017
rect 19889 14977 19901 15011
rect 19935 15008 19947 15011
rect 20530 15008 20536 15020
rect 19935 14980 20536 15008
rect 19935 14977 19947 14980
rect 19889 14971 19947 14977
rect 20530 14968 20536 14980
rect 20588 14968 20594 15020
rect 21085 15011 21143 15017
rect 21085 14977 21097 15011
rect 21131 15008 21143 15011
rect 21450 15008 21456 15020
rect 21131 14980 21456 15008
rect 21131 14977 21143 14980
rect 21085 14971 21143 14977
rect 21450 14968 21456 14980
rect 21508 14968 21514 15020
rect 22281 15011 22339 15017
rect 22281 14977 22293 15011
rect 22327 15008 22339 15011
rect 23293 15011 23351 15017
rect 23293 15008 23305 15011
rect 22327 14980 23305 15008
rect 22327 14977 22339 14980
rect 22281 14971 22339 14977
rect 23293 14977 23305 14980
rect 23339 14977 23351 15011
rect 23293 14971 23351 14977
rect 17126 14940 17132 14952
rect 15120 14912 17132 14940
rect 13265 14903 13323 14909
rect 17126 14900 17132 14912
rect 17184 14900 17190 14952
rect 17405 14943 17463 14949
rect 17405 14909 17417 14943
rect 17451 14909 17463 14943
rect 17405 14903 17463 14909
rect 10060 14844 12434 14872
rect 9493 14807 9551 14813
rect 9493 14773 9505 14807
rect 9539 14804 9551 14807
rect 10410 14804 10416 14816
rect 9539 14776 10416 14804
rect 9539 14773 9551 14776
rect 9493 14767 9551 14773
rect 10410 14764 10416 14776
rect 10468 14764 10474 14816
rect 10597 14807 10655 14813
rect 10597 14773 10609 14807
rect 10643 14804 10655 14807
rect 10686 14804 10692 14816
rect 10643 14776 10692 14804
rect 10643 14773 10655 14776
rect 10597 14767 10655 14773
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 11054 14764 11060 14816
rect 11112 14764 11118 14816
rect 12406 14804 12434 14844
rect 14274 14832 14280 14884
rect 14332 14872 14338 14884
rect 14737 14875 14795 14881
rect 14737 14872 14749 14875
rect 14332 14844 14749 14872
rect 14332 14832 14338 14844
rect 14737 14841 14749 14844
rect 14783 14872 14795 14875
rect 17420 14872 17448 14903
rect 17862 14900 17868 14952
rect 17920 14940 17926 14952
rect 18782 14940 18788 14952
rect 17920 14912 18788 14940
rect 17920 14900 17926 14912
rect 18782 14900 18788 14912
rect 18840 14900 18846 14952
rect 18874 14900 18880 14952
rect 18932 14900 18938 14952
rect 19978 14900 19984 14952
rect 20036 14900 20042 14952
rect 20070 14900 20076 14952
rect 20128 14900 20134 14952
rect 20898 14900 20904 14952
rect 20956 14940 20962 14952
rect 21177 14943 21235 14949
rect 21177 14940 21189 14943
rect 20956 14912 21189 14940
rect 20956 14900 20962 14912
rect 21177 14909 21189 14912
rect 21223 14909 21235 14943
rect 21177 14903 21235 14909
rect 21266 14900 21272 14952
rect 21324 14900 21330 14952
rect 23584 14949 23612 15048
rect 25774 15036 25780 15048
rect 25832 15036 25838 15088
rect 26329 15079 26387 15085
rect 26329 15045 26341 15079
rect 26375 15076 26387 15079
rect 27264 15076 27292 15104
rect 26375 15048 27292 15076
rect 26375 15045 26387 15048
rect 26329 15039 26387 15045
rect 24486 14968 24492 15020
rect 24544 15008 24550 15020
rect 25133 15011 25191 15017
rect 25133 15008 25145 15011
rect 24544 14980 25145 15008
rect 24544 14968 24550 14980
rect 25133 14977 25145 14980
rect 25179 15008 25191 15011
rect 25682 15008 25688 15020
rect 25179 14980 25688 15008
rect 25179 14977 25191 14980
rect 25133 14971 25191 14977
rect 25682 14968 25688 14980
rect 25740 14968 25746 15020
rect 26237 15011 26295 15017
rect 26237 14977 26249 15011
rect 26283 15008 26295 15011
rect 27246 15008 27252 15020
rect 26283 14980 27252 15008
rect 26283 14977 26295 14980
rect 26237 14971 26295 14977
rect 23385 14943 23443 14949
rect 23385 14909 23397 14943
rect 23431 14909 23443 14943
rect 23385 14903 23443 14909
rect 23569 14943 23627 14949
rect 23569 14909 23581 14943
rect 23615 14909 23627 14943
rect 23569 14903 23627 14909
rect 14783 14844 17448 14872
rect 18325 14875 18383 14881
rect 14783 14841 14795 14844
rect 14737 14835 14795 14841
rect 18325 14841 18337 14875
rect 18371 14872 18383 14875
rect 18414 14872 18420 14884
rect 18371 14844 18420 14872
rect 18371 14841 18383 14844
rect 18325 14835 18383 14841
rect 18414 14832 18420 14844
rect 18472 14832 18478 14884
rect 13446 14804 13452 14816
rect 12406 14776 13452 14804
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 15286 14764 15292 14816
rect 15344 14764 15350 14816
rect 16301 14807 16359 14813
rect 16301 14773 16313 14807
rect 16347 14804 16359 14807
rect 16482 14804 16488 14816
rect 16347 14776 16488 14804
rect 16347 14773 16359 14776
rect 16301 14767 16359 14773
rect 16482 14764 16488 14776
rect 16540 14764 16546 14816
rect 16850 14764 16856 14816
rect 16908 14804 16914 14816
rect 17310 14804 17316 14816
rect 16908 14776 17316 14804
rect 16908 14764 16914 14776
rect 17310 14764 17316 14776
rect 17368 14764 17374 14816
rect 17494 14764 17500 14816
rect 17552 14804 17558 14816
rect 20438 14804 20444 14816
rect 17552 14776 20444 14804
rect 17552 14764 17558 14776
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 21450 14764 21456 14816
rect 21508 14804 21514 14816
rect 23400 14804 23428 14903
rect 24578 14900 24584 14952
rect 24636 14900 24642 14952
rect 24673 14943 24731 14949
rect 24673 14909 24685 14943
rect 24719 14909 24731 14943
rect 24673 14903 24731 14909
rect 24118 14832 24124 14884
rect 24176 14872 24182 14884
rect 24688 14872 24716 14903
rect 24762 14900 24768 14952
rect 24820 14940 24826 14952
rect 26252 14940 26280 14971
rect 27246 14968 27252 14980
rect 27304 14968 27310 15020
rect 24820 14912 26280 14940
rect 26421 14943 26479 14949
rect 24820 14900 24826 14912
rect 26421 14909 26433 14943
rect 26467 14909 26479 14943
rect 27632 14940 27660 15107
rect 28718 15104 28724 15116
rect 28776 15104 28782 15156
rect 29086 15104 29092 15156
rect 29144 15144 29150 15156
rect 32309 15147 32367 15153
rect 32309 15144 32321 15147
rect 29144 15116 32321 15144
rect 29144 15104 29150 15116
rect 32309 15113 32321 15116
rect 32355 15113 32367 15147
rect 33778 15144 33784 15156
rect 32309 15107 32367 15113
rect 32692 15116 33784 15144
rect 28350 15076 28356 15088
rect 28092 15048 28356 15076
rect 28092 15017 28120 15048
rect 28350 15036 28356 15048
rect 28408 15036 28414 15088
rect 28442 15036 28448 15088
rect 28500 15076 28506 15088
rect 28500 15048 28842 15076
rect 28500 15036 28506 15048
rect 29822 15036 29828 15088
rect 29880 15076 29886 15088
rect 31573 15079 31631 15085
rect 29880 15048 30880 15076
rect 29880 15036 29886 15048
rect 28077 15011 28135 15017
rect 28077 14977 28089 15011
rect 28123 14977 28135 15011
rect 28077 14971 28135 14977
rect 30653 15011 30711 15017
rect 30653 14977 30665 15011
rect 30699 14977 30711 15011
rect 30653 14971 30711 14977
rect 26421 14903 26479 14909
rect 26528 14912 27660 14940
rect 28353 14943 28411 14949
rect 26436 14872 26464 14903
rect 24176 14844 24716 14872
rect 24780 14844 26464 14872
rect 24176 14832 24182 14844
rect 23750 14804 23756 14816
rect 21508 14776 23756 14804
rect 21508 14764 21514 14776
rect 23750 14764 23756 14776
rect 23808 14764 23814 14816
rect 24486 14764 24492 14816
rect 24544 14804 24550 14816
rect 24780 14804 24808 14844
rect 24544 14776 24808 14804
rect 24544 14764 24550 14776
rect 25130 14764 25136 14816
rect 25188 14804 25194 14816
rect 25317 14807 25375 14813
rect 25317 14804 25329 14807
rect 25188 14776 25329 14804
rect 25188 14764 25194 14776
rect 25317 14773 25329 14776
rect 25363 14773 25375 14807
rect 25317 14767 25375 14773
rect 25406 14764 25412 14816
rect 25464 14804 25470 14816
rect 25501 14807 25559 14813
rect 25501 14804 25513 14807
rect 25464 14776 25513 14804
rect 25464 14764 25470 14776
rect 25501 14773 25513 14776
rect 25547 14773 25559 14807
rect 25501 14767 25559 14773
rect 25590 14764 25596 14816
rect 25648 14804 25654 14816
rect 25869 14807 25927 14813
rect 25869 14804 25881 14807
rect 25648 14776 25881 14804
rect 25648 14764 25654 14776
rect 25869 14773 25881 14776
rect 25915 14773 25927 14807
rect 25869 14767 25927 14773
rect 26234 14764 26240 14816
rect 26292 14804 26298 14816
rect 26528 14804 26556 14912
rect 28353 14909 28365 14943
rect 28399 14940 28411 14943
rect 28902 14940 28908 14952
rect 28399 14912 28908 14940
rect 28399 14909 28411 14912
rect 28353 14903 28411 14909
rect 28902 14900 28908 14912
rect 28960 14900 28966 14952
rect 29825 14943 29883 14949
rect 29825 14909 29837 14943
rect 29871 14940 29883 14943
rect 30098 14940 30104 14952
rect 29871 14912 30104 14940
rect 29871 14909 29883 14912
rect 29825 14903 29883 14909
rect 27154 14832 27160 14884
rect 27212 14872 27218 14884
rect 27709 14875 27767 14881
rect 27709 14872 27721 14875
rect 27212 14844 27721 14872
rect 27212 14832 27218 14844
rect 27709 14841 27721 14844
rect 27755 14872 27767 14875
rect 28074 14872 28080 14884
rect 27755 14844 28080 14872
rect 27755 14841 27767 14844
rect 27709 14835 27767 14841
rect 28074 14832 28080 14844
rect 28132 14832 28138 14884
rect 26292 14776 26556 14804
rect 26292 14764 26298 14776
rect 26786 14764 26792 14816
rect 26844 14804 26850 14816
rect 28810 14804 28816 14816
rect 26844 14776 28816 14804
rect 26844 14764 26850 14776
rect 28810 14764 28816 14776
rect 28868 14804 28874 14816
rect 29840 14804 29868 14903
rect 30098 14900 30104 14912
rect 30156 14900 30162 14952
rect 28868 14776 29868 14804
rect 28868 14764 28874 14776
rect 30098 14764 30104 14816
rect 30156 14804 30162 14816
rect 30285 14807 30343 14813
rect 30285 14804 30297 14807
rect 30156 14776 30297 14804
rect 30156 14764 30162 14776
rect 30285 14773 30297 14776
rect 30331 14773 30343 14807
rect 30668 14804 30696 14971
rect 30742 14900 30748 14952
rect 30800 14900 30806 14952
rect 30852 14949 30880 15048
rect 31573 15045 31585 15079
rect 31619 15076 31631 15079
rect 32692 15076 32720 15116
rect 33778 15104 33784 15116
rect 33836 15104 33842 15156
rect 33873 15147 33931 15153
rect 33873 15113 33885 15147
rect 33919 15144 33931 15147
rect 34514 15144 34520 15156
rect 33919 15116 34520 15144
rect 33919 15113 33931 15116
rect 33873 15107 33931 15113
rect 34514 15104 34520 15116
rect 34572 15104 34578 15156
rect 34698 15104 34704 15156
rect 34756 15144 34762 15156
rect 35069 15147 35127 15153
rect 35069 15144 35081 15147
rect 34756 15116 35081 15144
rect 34756 15104 34762 15116
rect 35069 15113 35081 15116
rect 35115 15113 35127 15147
rect 35069 15107 35127 15113
rect 36262 15104 36268 15156
rect 36320 15104 36326 15156
rect 39669 15147 39727 15153
rect 39669 15144 39681 15147
rect 36372 15116 39681 15144
rect 31619 15048 32720 15076
rect 32769 15079 32827 15085
rect 31619 15045 31631 15048
rect 31573 15039 31631 15045
rect 32769 15045 32781 15079
rect 32815 15076 32827 15079
rect 36372 15076 36400 15116
rect 39669 15113 39681 15116
rect 39715 15113 39727 15147
rect 39669 15107 39727 15113
rect 40126 15104 40132 15156
rect 40184 15144 40190 15156
rect 41509 15147 41567 15153
rect 41509 15144 41521 15147
rect 40184 15116 41521 15144
rect 40184 15104 40190 15116
rect 41509 15113 41521 15116
rect 41555 15113 41567 15147
rect 41509 15107 41567 15113
rect 41598 15104 41604 15156
rect 41656 15144 41662 15156
rect 41785 15147 41843 15153
rect 41785 15144 41797 15147
rect 41656 15116 41797 15144
rect 41656 15104 41662 15116
rect 41785 15113 41797 15116
rect 41831 15144 41843 15147
rect 41969 15147 42027 15153
rect 41969 15144 41981 15147
rect 41831 15116 41981 15144
rect 41831 15113 41843 15116
rect 41785 15107 41843 15113
rect 41969 15113 41981 15116
rect 42015 15113 42027 15147
rect 41969 15107 42027 15113
rect 32815 15048 36400 15076
rect 32815 15045 32827 15048
rect 32769 15039 32827 15045
rect 38470 15036 38476 15088
rect 38528 15036 38534 15088
rect 40037 15079 40095 15085
rect 40037 15045 40049 15079
rect 40083 15076 40095 15079
rect 48406 15076 48412 15088
rect 40083 15048 48412 15076
rect 40083 15045 40095 15048
rect 40037 15039 40095 15045
rect 48406 15036 48412 15048
rect 48464 15036 48470 15088
rect 32674 14968 32680 15020
rect 32732 14968 32738 15020
rect 35986 15008 35992 15020
rect 34716 14980 35992 15008
rect 30837 14943 30895 14949
rect 30837 14909 30849 14943
rect 30883 14909 30895 14943
rect 30837 14903 30895 14909
rect 31018 14900 31024 14952
rect 31076 14940 31082 14952
rect 32582 14940 32588 14952
rect 31076 14912 32588 14940
rect 31076 14900 31082 14912
rect 32582 14900 32588 14912
rect 32640 14900 32646 14952
rect 32953 14943 33011 14949
rect 32953 14909 32965 14943
rect 32999 14940 33011 14943
rect 33318 14940 33324 14952
rect 32999 14912 33324 14940
rect 32999 14909 33011 14912
rect 32953 14903 33011 14909
rect 33318 14900 33324 14912
rect 33376 14900 33382 14952
rect 33965 14943 34023 14949
rect 33965 14940 33977 14943
rect 33428 14912 33977 14940
rect 30926 14832 30932 14884
rect 30984 14872 30990 14884
rect 33428 14872 33456 14912
rect 33965 14909 33977 14912
rect 34011 14909 34023 14943
rect 33965 14903 34023 14909
rect 34146 14900 34152 14952
rect 34204 14900 34210 14952
rect 34716 14881 34744 14980
rect 35986 14968 35992 14980
rect 36044 14968 36050 15020
rect 39850 14968 39856 15020
rect 39908 15008 39914 15020
rect 40129 15011 40187 15017
rect 40129 15008 40141 15011
rect 39908 14980 40141 15008
rect 39908 14968 39914 14980
rect 40129 14977 40141 14980
rect 40175 14977 40187 15011
rect 40129 14971 40187 14977
rect 40310 14968 40316 15020
rect 40368 15008 40374 15020
rect 40865 15011 40923 15017
rect 40865 15008 40877 15011
rect 40368 14980 40877 15008
rect 40368 14968 40374 14980
rect 40865 14977 40877 14980
rect 40911 14977 40923 15011
rect 40865 14971 40923 14977
rect 42058 14968 42064 15020
rect 42116 15008 42122 15020
rect 42797 15011 42855 15017
rect 42797 15008 42809 15011
rect 42116 14980 42809 15008
rect 42116 14968 42122 14980
rect 42797 14977 42809 14980
rect 42843 14977 42855 15011
rect 42797 14971 42855 14977
rect 48777 15011 48835 15017
rect 48777 14977 48789 15011
rect 48823 15008 48835 15011
rect 49050 15008 49056 15020
rect 48823 14980 49056 15008
rect 48823 14977 48835 14980
rect 48777 14971 48835 14977
rect 49050 14968 49056 14980
rect 49108 14968 49114 15020
rect 35161 14943 35219 14949
rect 35161 14909 35173 14943
rect 35207 14909 35219 14943
rect 35161 14903 35219 14909
rect 35345 14943 35403 14949
rect 35345 14909 35357 14943
rect 35391 14909 35403 14943
rect 35345 14903 35403 14909
rect 30984 14844 33456 14872
rect 34701 14875 34759 14881
rect 30984 14832 30990 14844
rect 34701 14841 34713 14875
rect 34747 14841 34759 14875
rect 34701 14835 34759 14841
rect 33226 14804 33232 14816
rect 30668 14776 33232 14804
rect 30285 14767 30343 14773
rect 33226 14764 33232 14776
rect 33284 14764 33290 14816
rect 33505 14807 33563 14813
rect 33505 14773 33517 14807
rect 33551 14804 33563 14807
rect 35066 14804 35072 14816
rect 33551 14776 35072 14804
rect 33551 14773 33563 14776
rect 33505 14767 33563 14773
rect 35066 14764 35072 14776
rect 35124 14764 35130 14816
rect 35176 14804 35204 14903
rect 35360 14872 35388 14903
rect 35526 14900 35532 14952
rect 35584 14940 35590 14952
rect 36357 14943 36415 14949
rect 36357 14940 36369 14943
rect 35584 14912 36369 14940
rect 35584 14900 35590 14912
rect 36357 14909 36369 14912
rect 36403 14909 36415 14943
rect 36357 14903 36415 14909
rect 36541 14943 36599 14949
rect 36541 14909 36553 14943
rect 36587 14940 36599 14943
rect 36630 14940 36636 14952
rect 36587 14912 36636 14940
rect 36587 14909 36599 14912
rect 36541 14903 36599 14909
rect 36630 14900 36636 14912
rect 36688 14900 36694 14952
rect 37458 14900 37464 14952
rect 37516 14900 37522 14952
rect 37737 14943 37795 14949
rect 37737 14909 37749 14943
rect 37783 14940 37795 14943
rect 40034 14940 40040 14952
rect 37783 14912 40040 14940
rect 37783 14909 37795 14912
rect 37737 14903 37795 14909
rect 40034 14900 40040 14912
rect 40092 14900 40098 14952
rect 40221 14943 40279 14949
rect 40221 14909 40233 14943
rect 40267 14909 40279 14943
rect 40221 14903 40279 14909
rect 35802 14872 35808 14884
rect 35360 14844 35808 14872
rect 35802 14832 35808 14844
rect 35860 14832 35866 14884
rect 35897 14875 35955 14881
rect 35897 14841 35909 14875
rect 35943 14872 35955 14875
rect 37366 14872 37372 14884
rect 35943 14844 37372 14872
rect 35943 14841 35955 14844
rect 35897 14835 35955 14841
rect 37366 14832 37372 14844
rect 37424 14832 37430 14884
rect 39942 14832 39948 14884
rect 40000 14872 40006 14884
rect 40236 14872 40264 14903
rect 40000 14844 40264 14872
rect 40000 14832 40006 14844
rect 48314 14832 48320 14884
rect 48372 14872 48378 14884
rect 49237 14875 49295 14881
rect 49237 14872 49249 14875
rect 48372 14844 49249 14872
rect 48372 14832 48378 14844
rect 49237 14841 49249 14844
rect 49283 14841 49295 14875
rect 49237 14835 49295 14841
rect 36262 14804 36268 14816
rect 35176 14776 36268 14804
rect 36262 14764 36268 14776
rect 36320 14804 36326 14816
rect 36909 14807 36967 14813
rect 36909 14804 36921 14807
rect 36320 14776 36921 14804
rect 36320 14764 36326 14776
rect 36909 14773 36921 14776
rect 36955 14773 36967 14807
rect 36909 14767 36967 14773
rect 37090 14764 37096 14816
rect 37148 14804 37154 14816
rect 38194 14804 38200 14816
rect 37148 14776 38200 14804
rect 37148 14764 37154 14776
rect 38194 14764 38200 14776
rect 38252 14764 38258 14816
rect 38286 14764 38292 14816
rect 38344 14804 38350 14816
rect 39209 14807 39267 14813
rect 39209 14804 39221 14807
rect 38344 14776 39221 14804
rect 38344 14764 38350 14776
rect 39209 14773 39221 14776
rect 39255 14804 39267 14807
rect 41138 14804 41144 14816
rect 39255 14776 41144 14804
rect 39255 14773 39267 14776
rect 39209 14767 39267 14773
rect 41138 14764 41144 14776
rect 41196 14764 41202 14816
rect 42613 14807 42671 14813
rect 42613 14773 42625 14807
rect 42659 14804 42671 14807
rect 45830 14804 45836 14816
rect 42659 14776 45836 14804
rect 42659 14773 42671 14776
rect 42613 14767 42671 14773
rect 45830 14764 45836 14776
rect 45888 14764 45894 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 9674 14560 9680 14612
rect 9732 14600 9738 14612
rect 10413 14603 10471 14609
rect 10413 14600 10425 14603
rect 9732 14572 10425 14600
rect 9732 14560 9738 14572
rect 10413 14569 10425 14572
rect 10459 14569 10471 14603
rect 10413 14563 10471 14569
rect 10502 14560 10508 14612
rect 10560 14600 10566 14612
rect 14185 14603 14243 14609
rect 14185 14600 14197 14603
rect 10560 14572 14197 14600
rect 10560 14560 10566 14572
rect 14185 14569 14197 14572
rect 14231 14600 14243 14603
rect 16022 14600 16028 14612
rect 14231 14572 16028 14600
rect 14231 14569 14243 14572
rect 14185 14563 14243 14569
rect 16022 14560 16028 14572
rect 16080 14600 16086 14612
rect 16390 14600 16396 14612
rect 16080 14572 16396 14600
rect 16080 14560 16086 14572
rect 16390 14560 16396 14572
rect 16448 14560 16454 14612
rect 16942 14560 16948 14612
rect 17000 14600 17006 14612
rect 18690 14600 18696 14612
rect 17000 14572 18696 14600
rect 17000 14560 17006 14572
rect 18690 14560 18696 14572
rect 18748 14560 18754 14612
rect 21726 14560 21732 14612
rect 21784 14600 21790 14612
rect 23474 14600 23480 14612
rect 21784 14572 23480 14600
rect 21784 14560 21790 14572
rect 23474 14560 23480 14572
rect 23532 14560 23538 14612
rect 23750 14560 23756 14612
rect 23808 14560 23814 14612
rect 24213 14603 24271 14609
rect 24213 14569 24225 14603
rect 24259 14600 24271 14603
rect 24578 14600 24584 14612
rect 24259 14572 24584 14600
rect 24259 14569 24271 14572
rect 24213 14563 24271 14569
rect 24578 14560 24584 14572
rect 24636 14560 24642 14612
rect 25948 14603 26006 14609
rect 25948 14569 25960 14603
rect 25994 14600 26006 14603
rect 29086 14600 29092 14612
rect 25994 14572 29092 14600
rect 25994 14569 26006 14572
rect 25948 14563 26006 14569
rect 29086 14560 29092 14572
rect 29144 14560 29150 14612
rect 29733 14603 29791 14609
rect 29733 14569 29745 14603
rect 29779 14600 29791 14603
rect 30834 14600 30840 14612
rect 29779 14572 30840 14600
rect 29779 14569 29791 14572
rect 29733 14563 29791 14569
rect 30834 14560 30840 14572
rect 30892 14560 30898 14612
rect 30929 14603 30987 14609
rect 30929 14569 30941 14603
rect 30975 14600 30987 14603
rect 33870 14600 33876 14612
rect 30975 14572 33876 14600
rect 30975 14569 30987 14572
rect 30929 14563 30987 14569
rect 33870 14560 33876 14572
rect 33928 14560 33934 14612
rect 33962 14560 33968 14612
rect 34020 14600 34026 14612
rect 37734 14600 37740 14612
rect 34020 14572 37740 14600
rect 34020 14560 34026 14572
rect 37734 14560 37740 14572
rect 37792 14560 37798 14612
rect 41598 14560 41604 14612
rect 41656 14600 41662 14612
rect 42061 14603 42119 14609
rect 42061 14600 42073 14603
rect 41656 14572 42073 14600
rect 41656 14560 41662 14572
rect 42061 14569 42073 14572
rect 42107 14569 42119 14603
rect 42061 14563 42119 14569
rect 5442 14492 5448 14544
rect 5500 14532 5506 14544
rect 11054 14532 11060 14544
rect 5500 14504 11060 14532
rect 5500 14492 5506 14504
rect 11054 14492 11060 14504
rect 11112 14492 11118 14544
rect 11793 14535 11851 14541
rect 11793 14501 11805 14535
rect 11839 14532 11851 14535
rect 12342 14532 12348 14544
rect 11839 14504 12348 14532
rect 11839 14501 11851 14504
rect 11793 14495 11851 14501
rect 12342 14492 12348 14504
rect 12400 14492 12406 14544
rect 18141 14535 18199 14541
rect 18141 14532 18153 14535
rect 13464 14504 16436 14532
rect 1302 14424 1308 14476
rect 1360 14464 1366 14476
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1360 14436 2053 14464
rect 1360 14424 1366 14436
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 9033 14467 9091 14473
rect 9033 14433 9045 14467
rect 9079 14464 9091 14467
rect 12437 14467 12495 14473
rect 9079 14436 10364 14464
rect 9079 14433 9091 14436
rect 9033 14427 9091 14433
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 9769 14399 9827 14405
rect 9769 14396 9781 14399
rect 1811 14368 9781 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 9769 14365 9781 14368
rect 9815 14365 9827 14399
rect 9769 14359 9827 14365
rect 10336 14340 10364 14436
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 13354 14464 13360 14476
rect 12483 14436 13360 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 13464 14473 13492 14504
rect 13449 14467 13507 14473
rect 13449 14433 13461 14467
rect 13495 14433 13507 14467
rect 13449 14427 13507 14433
rect 13538 14424 13544 14476
rect 13596 14424 13602 14476
rect 13814 14424 13820 14476
rect 13872 14464 13878 14476
rect 15105 14467 15163 14473
rect 15105 14464 15117 14467
rect 13872 14436 15117 14464
rect 13872 14424 13878 14436
rect 15105 14433 15117 14436
rect 15151 14464 15163 14467
rect 15151 14436 16068 14464
rect 15151 14433 15163 14436
rect 15105 14427 15163 14433
rect 11422 14396 11428 14408
rect 11164 14368 11428 14396
rect 9582 14288 9588 14340
rect 9640 14288 9646 14340
rect 10318 14288 10324 14340
rect 10376 14288 10382 14340
rect 11164 14337 11192 14368
rect 11422 14356 11428 14368
rect 11480 14356 11486 14408
rect 11974 14356 11980 14408
rect 12032 14396 12038 14408
rect 12161 14399 12219 14405
rect 12161 14396 12173 14399
rect 12032 14368 12173 14396
rect 12032 14356 12038 14368
rect 12161 14365 12173 14368
rect 12207 14365 12219 14399
rect 16040 14396 16068 14436
rect 16206 14424 16212 14476
rect 16264 14424 16270 14476
rect 16408 14464 16436 14504
rect 16592 14504 18153 14532
rect 16592 14464 16620 14504
rect 18141 14501 18153 14504
rect 18187 14501 18199 14535
rect 18141 14495 18199 14501
rect 18414 14492 18420 14544
rect 18472 14532 18478 14544
rect 19613 14535 19671 14541
rect 19613 14532 19625 14535
rect 18472 14504 19625 14532
rect 18472 14492 18478 14504
rect 19613 14501 19625 14504
rect 19659 14501 19671 14535
rect 19613 14495 19671 14501
rect 19794 14492 19800 14544
rect 19852 14532 19858 14544
rect 19852 14504 21220 14532
rect 19852 14492 19858 14504
rect 16408 14436 16620 14464
rect 16666 14424 16672 14476
rect 16724 14464 16730 14476
rect 17034 14464 17040 14476
rect 16724 14436 17040 14464
rect 16724 14424 16730 14436
rect 17034 14424 17040 14436
rect 17092 14464 17098 14476
rect 17402 14464 17408 14476
rect 17092 14436 17408 14464
rect 17092 14424 17098 14436
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 18598 14464 18604 14476
rect 17512 14436 18604 14464
rect 16942 14396 16948 14408
rect 16040 14368 16948 14396
rect 12161 14359 12219 14365
rect 16942 14356 16948 14368
rect 17000 14356 17006 14408
rect 17218 14356 17224 14408
rect 17276 14356 17282 14408
rect 17310 14356 17316 14408
rect 17368 14396 17374 14408
rect 17512 14396 17540 14436
rect 18598 14424 18604 14436
rect 18656 14424 18662 14476
rect 18690 14424 18696 14476
rect 18748 14424 18754 14476
rect 19058 14424 19064 14476
rect 19116 14464 19122 14476
rect 20165 14467 20223 14473
rect 20165 14464 20177 14467
rect 19116 14436 20177 14464
rect 19116 14424 19122 14436
rect 20165 14433 20177 14436
rect 20211 14433 20223 14467
rect 20165 14427 20223 14433
rect 21082 14424 21088 14476
rect 21140 14424 21146 14476
rect 21192 14464 21220 14504
rect 22646 14492 22652 14544
rect 22704 14532 22710 14544
rect 25590 14532 25596 14544
rect 22704 14504 25596 14532
rect 22704 14492 22710 14504
rect 25590 14492 25596 14504
rect 25648 14492 25654 14544
rect 27893 14535 27951 14541
rect 27893 14501 27905 14535
rect 27939 14501 27951 14535
rect 28718 14532 28724 14544
rect 27893 14495 27951 14501
rect 28368 14504 28724 14532
rect 21726 14464 21732 14476
rect 21192 14436 21732 14464
rect 21726 14424 21732 14436
rect 21784 14424 21790 14476
rect 22738 14424 22744 14476
rect 22796 14464 22802 14476
rect 23109 14467 23167 14473
rect 23109 14464 23121 14467
rect 22796 14436 23121 14464
rect 22796 14424 22802 14436
rect 23109 14433 23121 14436
rect 23155 14433 23167 14467
rect 23109 14427 23167 14433
rect 24394 14424 24400 14476
rect 24452 14464 24458 14476
rect 24670 14464 24676 14476
rect 24452 14436 24676 14464
rect 24452 14424 24458 14436
rect 24670 14424 24676 14436
rect 24728 14424 24734 14476
rect 24854 14424 24860 14476
rect 24912 14464 24918 14476
rect 25685 14467 25743 14473
rect 25685 14464 25697 14467
rect 24912 14436 25697 14464
rect 24912 14424 24918 14436
rect 25685 14433 25697 14436
rect 25731 14464 25743 14467
rect 27154 14464 27160 14476
rect 25731 14436 27160 14464
rect 25731 14433 25743 14436
rect 25685 14427 25743 14433
rect 27154 14424 27160 14436
rect 27212 14424 27218 14476
rect 17368 14368 17540 14396
rect 17368 14356 17374 14368
rect 17678 14356 17684 14408
rect 17736 14396 17742 14408
rect 20346 14396 20352 14408
rect 17736 14368 20352 14396
rect 17736 14356 17742 14368
rect 20346 14356 20352 14368
rect 20404 14396 20410 14408
rect 20990 14396 20996 14408
rect 20404 14368 20996 14396
rect 20404 14356 20410 14368
rect 20990 14356 20996 14368
rect 21048 14356 21054 14408
rect 23934 14396 23940 14408
rect 23400 14368 23940 14396
rect 11149 14331 11207 14337
rect 11149 14297 11161 14331
rect 11195 14297 11207 14331
rect 11149 14291 11207 14297
rect 9217 14263 9275 14269
rect 9217 14229 9229 14263
rect 9263 14260 9275 14263
rect 11164 14260 11192 14291
rect 12250 14288 12256 14340
rect 12308 14288 12314 14340
rect 13357 14331 13415 14337
rect 13357 14297 13369 14331
rect 13403 14328 13415 14331
rect 13403 14300 14504 14328
rect 13403 14297 13415 14300
rect 13357 14291 13415 14297
rect 9263 14232 11192 14260
rect 9263 14229 9275 14232
rect 9217 14223 9275 14229
rect 11238 14220 11244 14272
rect 11296 14220 11302 14272
rect 11330 14220 11336 14272
rect 11388 14260 11394 14272
rect 12989 14263 13047 14269
rect 12989 14260 13001 14263
rect 11388 14232 13001 14260
rect 11388 14220 11394 14232
rect 12989 14229 13001 14232
rect 13035 14229 13047 14263
rect 12989 14223 13047 14229
rect 13906 14220 13912 14272
rect 13964 14260 13970 14272
rect 14182 14260 14188 14272
rect 13964 14232 14188 14260
rect 13964 14220 13970 14232
rect 14182 14220 14188 14232
rect 14240 14220 14246 14272
rect 14476 14269 14504 14300
rect 14826 14288 14832 14340
rect 14884 14288 14890 14340
rect 17862 14328 17868 14340
rect 15672 14300 17868 14328
rect 14461 14263 14519 14269
rect 14461 14229 14473 14263
rect 14507 14229 14519 14263
rect 14461 14223 14519 14229
rect 14918 14220 14924 14272
rect 14976 14220 14982 14272
rect 15672 14269 15700 14300
rect 17862 14288 17868 14300
rect 17920 14288 17926 14340
rect 21361 14331 21419 14337
rect 21361 14328 21373 14331
rect 17972 14300 21373 14328
rect 15657 14263 15715 14269
rect 15657 14229 15669 14263
rect 15703 14229 15715 14263
rect 15657 14223 15715 14229
rect 16022 14220 16028 14272
rect 16080 14220 16086 14272
rect 16114 14220 16120 14272
rect 16172 14220 16178 14272
rect 16206 14220 16212 14272
rect 16264 14260 16270 14272
rect 16853 14263 16911 14269
rect 16853 14260 16865 14263
rect 16264 14232 16865 14260
rect 16264 14220 16270 14232
rect 16853 14229 16865 14232
rect 16899 14229 16911 14263
rect 16853 14223 16911 14229
rect 17126 14220 17132 14272
rect 17184 14260 17190 14272
rect 17313 14263 17371 14269
rect 17313 14260 17325 14263
rect 17184 14232 17325 14260
rect 17184 14220 17190 14232
rect 17313 14229 17325 14232
rect 17359 14229 17371 14263
rect 17313 14223 17371 14229
rect 17402 14220 17408 14272
rect 17460 14260 17466 14272
rect 17972 14260 18000 14300
rect 21361 14297 21373 14300
rect 21407 14297 21419 14331
rect 21361 14291 21419 14297
rect 21910 14288 21916 14340
rect 21968 14288 21974 14340
rect 23014 14288 23020 14340
rect 23072 14328 23078 14340
rect 23400 14337 23428 14368
rect 23934 14356 23940 14368
rect 23992 14356 23998 14408
rect 24026 14356 24032 14408
rect 24084 14396 24090 14408
rect 24581 14399 24639 14405
rect 24581 14396 24593 14399
rect 24084 14368 24593 14396
rect 24084 14356 24090 14368
rect 24581 14365 24593 14368
rect 24627 14365 24639 14399
rect 24581 14359 24639 14365
rect 27062 14356 27068 14408
rect 27120 14356 27126 14408
rect 27908 14396 27936 14495
rect 28368 14473 28396 14504
rect 28718 14492 28724 14504
rect 28776 14492 28782 14544
rect 32030 14532 32036 14544
rect 30300 14504 32036 14532
rect 28353 14467 28411 14473
rect 28353 14433 28365 14467
rect 28399 14433 28411 14467
rect 28353 14427 28411 14433
rect 28534 14424 28540 14476
rect 28592 14464 28598 14476
rect 30300 14473 30328 14504
rect 32030 14492 32036 14504
rect 32088 14492 32094 14544
rect 32125 14535 32183 14541
rect 32125 14501 32137 14535
rect 32171 14532 32183 14535
rect 32858 14532 32864 14544
rect 32171 14504 32864 14532
rect 32171 14501 32183 14504
rect 32125 14495 32183 14501
rect 32858 14492 32864 14504
rect 32916 14492 32922 14544
rect 33321 14535 33379 14541
rect 33321 14501 33333 14535
rect 33367 14532 33379 14535
rect 34790 14532 34796 14544
rect 33367 14504 34796 14532
rect 33367 14501 33379 14504
rect 33321 14495 33379 14501
rect 34790 14492 34796 14504
rect 34848 14492 34854 14544
rect 36538 14492 36544 14544
rect 36596 14532 36602 14544
rect 36633 14535 36691 14541
rect 36633 14532 36645 14535
rect 36596 14504 36645 14532
rect 36596 14492 36602 14504
rect 36633 14501 36645 14504
rect 36679 14501 36691 14535
rect 39850 14532 39856 14544
rect 36633 14495 36691 14501
rect 38856 14504 39856 14532
rect 29089 14467 29147 14473
rect 29089 14464 29101 14467
rect 28592 14436 29101 14464
rect 28592 14424 28598 14436
rect 29089 14433 29101 14436
rect 29135 14464 29147 14467
rect 30285 14467 30343 14473
rect 29135 14436 30236 14464
rect 29135 14433 29147 14436
rect 29089 14427 29147 14433
rect 30208 14396 30236 14436
rect 30285 14433 30297 14467
rect 30331 14433 30343 14467
rect 30285 14427 30343 14433
rect 30374 14424 30380 14476
rect 30432 14464 30438 14476
rect 30742 14464 30748 14476
rect 30432 14436 30748 14464
rect 30432 14424 30438 14436
rect 30742 14424 30748 14436
rect 30800 14424 30806 14476
rect 31573 14467 31631 14473
rect 31573 14433 31585 14467
rect 31619 14464 31631 14467
rect 31662 14464 31668 14476
rect 31619 14436 31668 14464
rect 31619 14433 31631 14436
rect 31573 14427 31631 14433
rect 31662 14424 31668 14436
rect 31720 14424 31726 14476
rect 32769 14467 32827 14473
rect 32769 14433 32781 14467
rect 32815 14464 32827 14467
rect 32950 14464 32956 14476
rect 32815 14436 32956 14464
rect 32815 14433 32827 14436
rect 32769 14427 32827 14433
rect 32950 14424 32956 14436
rect 33008 14424 33014 14476
rect 33594 14424 33600 14476
rect 33652 14464 33658 14476
rect 33781 14467 33839 14473
rect 33781 14464 33793 14467
rect 33652 14436 33793 14464
rect 33652 14424 33658 14436
rect 33781 14433 33793 14436
rect 33827 14433 33839 14467
rect 33781 14427 33839 14433
rect 33965 14467 34023 14473
rect 33965 14433 33977 14467
rect 34011 14464 34023 14467
rect 34146 14464 34152 14476
rect 34011 14436 34152 14464
rect 34011 14433 34023 14436
rect 33965 14427 34023 14433
rect 34146 14424 34152 14436
rect 34204 14424 34210 14476
rect 34882 14424 34888 14476
rect 34940 14464 34946 14476
rect 37093 14467 37151 14473
rect 37093 14464 37105 14467
rect 34940 14436 37105 14464
rect 34940 14424 34946 14436
rect 37093 14433 37105 14436
rect 37139 14464 37151 14467
rect 37458 14464 37464 14476
rect 37139 14436 37464 14464
rect 37139 14433 37151 14436
rect 37093 14427 37151 14433
rect 37458 14424 37464 14436
rect 37516 14424 37522 14476
rect 37826 14424 37832 14476
rect 37884 14464 37890 14476
rect 38856 14464 38884 14504
rect 39850 14492 39856 14504
rect 39908 14492 39914 14544
rect 45554 14492 45560 14544
rect 45612 14532 45618 14544
rect 48590 14532 48596 14544
rect 45612 14504 48596 14532
rect 45612 14492 45618 14504
rect 48590 14492 48596 14504
rect 48648 14492 48654 14544
rect 37884 14436 38884 14464
rect 37884 14424 37890 14436
rect 38930 14424 38936 14476
rect 38988 14464 38994 14476
rect 39942 14464 39948 14476
rect 38988 14436 39948 14464
rect 38988 14424 38994 14436
rect 39942 14424 39948 14436
rect 40000 14464 40006 14476
rect 40000 14436 40080 14464
rect 40000 14424 40006 14436
rect 31018 14396 31024 14408
rect 27908 14368 29684 14396
rect 30208 14368 31024 14396
rect 23385 14331 23443 14337
rect 23385 14328 23397 14331
rect 23072 14300 23397 14328
rect 23072 14288 23078 14300
rect 23385 14297 23397 14300
rect 23431 14297 23443 14331
rect 23385 14291 23443 14297
rect 23474 14288 23480 14340
rect 23532 14328 23538 14340
rect 26234 14328 26240 14340
rect 23532 14300 26240 14328
rect 23532 14288 23538 14300
rect 26234 14288 26240 14300
rect 26292 14288 26298 14340
rect 28261 14331 28319 14337
rect 28261 14297 28273 14331
rect 28307 14328 28319 14331
rect 29656 14328 29684 14368
rect 31018 14356 31024 14368
rect 31076 14356 31082 14408
rect 31110 14356 31116 14408
rect 31168 14396 31174 14408
rect 31297 14399 31355 14405
rect 31297 14396 31309 14399
rect 31168 14368 31309 14396
rect 31168 14356 31174 14368
rect 31297 14365 31309 14368
rect 31343 14365 31355 14399
rect 31297 14359 31355 14365
rect 31478 14356 31484 14408
rect 31536 14396 31542 14408
rect 32585 14399 32643 14405
rect 32585 14396 32597 14399
rect 31536 14368 32597 14396
rect 31536 14356 31542 14368
rect 32585 14365 32597 14368
rect 32631 14396 32643 14399
rect 32631 14368 33272 14396
rect 32631 14365 32643 14368
rect 32585 14359 32643 14365
rect 31389 14331 31447 14337
rect 31389 14328 31401 14331
rect 28307 14300 28672 14328
rect 29656 14300 31401 14328
rect 28307 14297 28319 14300
rect 28261 14291 28319 14297
rect 28644 14272 28672 14300
rect 31389 14297 31401 14300
rect 31435 14297 31447 14331
rect 33134 14328 33140 14340
rect 31389 14291 31447 14297
rect 32508 14300 33140 14328
rect 17460 14232 18000 14260
rect 18509 14263 18567 14269
rect 17460 14220 17466 14232
rect 18509 14229 18521 14263
rect 18555 14260 18567 14263
rect 19150 14260 19156 14272
rect 18555 14232 19156 14260
rect 18555 14229 18567 14232
rect 18509 14223 18567 14229
rect 19150 14220 19156 14232
rect 19208 14220 19214 14272
rect 19337 14263 19395 14269
rect 19337 14229 19349 14263
rect 19383 14260 19395 14263
rect 19702 14260 19708 14272
rect 19383 14232 19708 14260
rect 19383 14229 19395 14232
rect 19337 14223 19395 14229
rect 19702 14220 19708 14232
rect 19760 14260 19766 14272
rect 19981 14263 20039 14269
rect 19981 14260 19993 14263
rect 19760 14232 19993 14260
rect 19760 14220 19766 14232
rect 19981 14229 19993 14232
rect 20027 14229 20039 14263
rect 19981 14223 20039 14229
rect 20070 14220 20076 14272
rect 20128 14220 20134 14272
rect 20717 14263 20775 14269
rect 20717 14229 20729 14263
rect 20763 14260 20775 14263
rect 20898 14260 20904 14272
rect 20763 14232 20904 14260
rect 20763 14229 20775 14232
rect 20717 14223 20775 14229
rect 20898 14220 20904 14232
rect 20956 14220 20962 14272
rect 21726 14220 21732 14272
rect 21784 14260 21790 14272
rect 23290 14260 23296 14272
rect 21784 14232 23296 14260
rect 21784 14220 21790 14232
rect 23290 14220 23296 14232
rect 23348 14220 23354 14272
rect 23661 14263 23719 14269
rect 23661 14229 23673 14263
rect 23707 14260 23719 14263
rect 23842 14260 23848 14272
rect 23707 14232 23848 14260
rect 23707 14229 23719 14232
rect 23661 14223 23719 14229
rect 23842 14220 23848 14232
rect 23900 14220 23906 14272
rect 24210 14220 24216 14272
rect 24268 14260 24274 14272
rect 25225 14263 25283 14269
rect 25225 14260 25237 14263
rect 24268 14232 25237 14260
rect 24268 14220 24274 14232
rect 25225 14229 25237 14232
rect 25271 14229 25283 14263
rect 25225 14223 25283 14229
rect 25498 14220 25504 14272
rect 25556 14260 25562 14272
rect 27433 14263 27491 14269
rect 27433 14260 27445 14263
rect 25556 14232 27445 14260
rect 25556 14220 25562 14232
rect 27433 14229 27445 14232
rect 27479 14229 27491 14263
rect 27433 14223 27491 14229
rect 28626 14220 28632 14272
rect 28684 14260 28690 14272
rect 28905 14263 28963 14269
rect 28905 14260 28917 14263
rect 28684 14232 28917 14260
rect 28684 14220 28690 14232
rect 28905 14229 28917 14232
rect 28951 14229 28963 14263
rect 28905 14223 28963 14229
rect 29270 14220 29276 14272
rect 29328 14220 29334 14272
rect 29454 14220 29460 14272
rect 29512 14260 29518 14272
rect 30101 14263 30159 14269
rect 30101 14260 30113 14263
rect 29512 14232 30113 14260
rect 29512 14220 29518 14232
rect 30101 14229 30113 14232
rect 30147 14229 30159 14263
rect 30101 14223 30159 14229
rect 30190 14220 30196 14272
rect 30248 14260 30254 14272
rect 30466 14260 30472 14272
rect 30248 14232 30472 14260
rect 30248 14220 30254 14232
rect 30466 14220 30472 14232
rect 30524 14260 30530 14272
rect 32030 14260 32036 14272
rect 30524 14232 32036 14260
rect 30524 14220 30530 14232
rect 32030 14220 32036 14232
rect 32088 14220 32094 14272
rect 32508 14269 32536 14300
rect 33134 14288 33140 14300
rect 33192 14288 33198 14340
rect 33244 14328 33272 14368
rect 33410 14356 33416 14408
rect 33468 14396 33474 14408
rect 33689 14399 33747 14405
rect 33689 14396 33701 14399
rect 33468 14368 33701 14396
rect 33468 14356 33474 14368
rect 33689 14365 33701 14368
rect 33735 14365 33747 14399
rect 33689 14359 33747 14365
rect 38470 14356 38476 14408
rect 38528 14356 38534 14408
rect 39482 14356 39488 14408
rect 39540 14356 39546 14408
rect 40052 14405 40080 14436
rect 40037 14399 40095 14405
rect 40037 14365 40049 14399
rect 40083 14365 40095 14399
rect 40037 14359 40095 14365
rect 41138 14356 41144 14408
rect 41196 14356 41202 14408
rect 48593 14399 48651 14405
rect 48593 14365 48605 14399
rect 48639 14396 48651 14399
rect 49050 14396 49056 14408
rect 48639 14368 49056 14396
rect 48639 14365 48651 14368
rect 48593 14359 48651 14365
rect 49050 14356 49056 14368
rect 49108 14356 49114 14408
rect 34333 14331 34391 14337
rect 34333 14328 34345 14331
rect 33244 14300 34345 14328
rect 34333 14297 34345 14300
rect 34379 14297 34391 14331
rect 34333 14291 34391 14297
rect 35158 14288 35164 14340
rect 35216 14328 35222 14340
rect 35434 14328 35440 14340
rect 35216 14300 35440 14328
rect 35216 14288 35222 14300
rect 35434 14288 35440 14300
rect 35492 14288 35498 14340
rect 36170 14288 36176 14340
rect 36228 14288 36234 14340
rect 37369 14331 37427 14337
rect 37369 14297 37381 14331
rect 37415 14297 37427 14331
rect 41785 14331 41843 14337
rect 41785 14328 41797 14331
rect 37369 14291 37427 14297
rect 38764 14300 41797 14328
rect 32493 14263 32551 14269
rect 32493 14229 32505 14263
rect 32539 14229 32551 14263
rect 32493 14223 32551 14229
rect 32582 14220 32588 14272
rect 32640 14260 32646 14272
rect 36078 14260 36084 14272
rect 32640 14232 36084 14260
rect 32640 14220 32646 14232
rect 36078 14220 36084 14232
rect 36136 14220 36142 14272
rect 37384 14260 37412 14291
rect 38764 14260 38792 14300
rect 41785 14297 41797 14300
rect 41831 14297 41843 14331
rect 41785 14291 41843 14297
rect 37384 14232 38792 14260
rect 38841 14263 38899 14269
rect 38841 14229 38853 14263
rect 38887 14260 38899 14263
rect 38930 14260 38936 14272
rect 38887 14232 38936 14260
rect 38887 14229 38899 14232
rect 38841 14223 38899 14229
rect 38930 14220 38936 14232
rect 38988 14220 38994 14272
rect 39298 14220 39304 14272
rect 39356 14220 39362 14272
rect 40678 14220 40684 14272
rect 40736 14220 40742 14272
rect 41414 14220 41420 14272
rect 41472 14260 41478 14272
rect 44174 14260 44180 14272
rect 41472 14232 44180 14260
rect 41472 14220 41478 14232
rect 44174 14220 44180 14232
rect 44232 14220 44238 14272
rect 48314 14220 48320 14272
rect 48372 14260 48378 14272
rect 48685 14263 48743 14269
rect 48685 14260 48697 14263
rect 48372 14232 48697 14260
rect 48372 14220 48378 14232
rect 48685 14229 48697 14232
rect 48731 14229 48743 14263
rect 48685 14223 48743 14229
rect 49234 14220 49240 14272
rect 49292 14220 49298 14272
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 3605 14059 3663 14065
rect 3605 14025 3617 14059
rect 3651 14056 3663 14059
rect 9766 14056 9772 14068
rect 3651 14028 9772 14056
rect 3651 14025 3663 14028
rect 3605 14019 3663 14025
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 9858 14016 9864 14068
rect 9916 14016 9922 14068
rect 11149 14059 11207 14065
rect 11149 14025 11161 14059
rect 11195 14056 11207 14059
rect 11195 14028 11468 14056
rect 11195 14025 11207 14028
rect 11149 14019 11207 14025
rect 11238 13988 11244 14000
rect 1780 13960 11244 13988
rect 1780 13929 1808 13960
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 11440 13988 11468 14028
rect 11514 14016 11520 14068
rect 11572 14056 11578 14068
rect 11609 14059 11667 14065
rect 11609 14056 11621 14059
rect 11572 14028 11621 14056
rect 11572 14016 11578 14028
rect 11609 14025 11621 14028
rect 11655 14025 11667 14059
rect 11609 14019 11667 14025
rect 15102 14016 15108 14068
rect 15160 14016 15166 14068
rect 16114 14056 16120 14068
rect 15580 14028 16120 14056
rect 12526 13988 12532 14000
rect 11440 13960 12532 13988
rect 12526 13948 12532 13960
rect 12584 13948 12590 14000
rect 13354 13948 13360 14000
rect 13412 13988 13418 14000
rect 13906 13988 13912 14000
rect 13412 13960 13912 13988
rect 13412 13948 13418 13960
rect 13906 13948 13912 13960
rect 13964 13948 13970 14000
rect 14182 13948 14188 14000
rect 14240 13948 14246 14000
rect 15580 13988 15608 14028
rect 16114 14016 16120 14028
rect 16172 14016 16178 14068
rect 16301 14059 16359 14065
rect 16301 14025 16313 14059
rect 16347 14056 16359 14059
rect 17402 14056 17408 14068
rect 16347 14028 17408 14056
rect 16347 14025 16359 14028
rect 16301 14019 16359 14025
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 17770 14016 17776 14068
rect 17828 14056 17834 14068
rect 17865 14059 17923 14065
rect 17865 14056 17877 14059
rect 17828 14028 17877 14056
rect 17828 14016 17834 14028
rect 17865 14025 17877 14028
rect 17911 14025 17923 14059
rect 17865 14019 17923 14025
rect 18233 14059 18291 14065
rect 18233 14025 18245 14059
rect 18279 14056 18291 14059
rect 20714 14056 20720 14068
rect 18279 14028 20720 14056
rect 18279 14025 18291 14028
rect 18233 14019 18291 14025
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 20990 14016 20996 14068
rect 21048 14056 21054 14068
rect 21453 14059 21511 14065
rect 21453 14056 21465 14059
rect 21048 14028 21465 14056
rect 21048 14016 21054 14028
rect 21453 14025 21465 14028
rect 21499 14025 21511 14059
rect 23290 14056 23296 14068
rect 21453 14019 21511 14025
rect 22020 14028 23296 14056
rect 17678 13988 17684 14000
rect 15028 13960 15608 13988
rect 15672 13960 17684 13988
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13889 1823 13923
rect 1765 13883 1823 13889
rect 3510 13880 3516 13932
rect 3568 13920 3574 13932
rect 3973 13923 4031 13929
rect 3973 13920 3985 13923
rect 3568 13892 3985 13920
rect 3568 13880 3574 13892
rect 3973 13889 3985 13892
rect 4019 13889 4031 13923
rect 3973 13883 4031 13889
rect 4062 13880 4068 13932
rect 4120 13920 4126 13932
rect 10226 13920 10232 13932
rect 4120 13892 10232 13920
rect 4120 13880 4126 13892
rect 10226 13880 10232 13892
rect 10284 13880 10290 13932
rect 10505 13923 10563 13929
rect 10505 13889 10517 13923
rect 10551 13889 10563 13923
rect 10505 13883 10563 13889
rect 12345 13923 12403 13929
rect 12345 13889 12357 13923
rect 12391 13920 12403 13923
rect 12710 13920 12716 13932
rect 12391 13892 12716 13920
rect 12391 13889 12403 13892
rect 12345 13883 12403 13889
rect 934 13812 940 13864
rect 992 13852 998 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 992 13824 2053 13852
rect 992 13812 998 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 7374 13812 7380 13864
rect 7432 13852 7438 13864
rect 7432 13824 9536 13852
rect 7432 13812 7438 13824
rect 9508 13716 9536 13824
rect 9582 13812 9588 13864
rect 9640 13852 9646 13864
rect 10318 13852 10324 13864
rect 9640 13824 10324 13852
rect 9640 13812 9646 13824
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 10520 13852 10548 13883
rect 12710 13880 12716 13892
rect 12768 13880 12774 13932
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 10520 13824 12112 13852
rect 11977 13719 12035 13725
rect 11977 13716 11989 13719
rect 9508 13688 11989 13716
rect 11977 13685 11989 13688
rect 12023 13685 12035 13719
rect 12084 13716 12112 13824
rect 12360 13824 12449 13852
rect 12360 13796 12388 13824
rect 12437 13821 12449 13824
rect 12483 13821 12495 13855
rect 12437 13815 12495 13821
rect 12529 13855 12587 13861
rect 12529 13821 12541 13855
rect 12575 13821 12587 13855
rect 12529 13815 12587 13821
rect 12342 13744 12348 13796
rect 12400 13744 12406 13796
rect 12250 13716 12256 13728
rect 12084 13688 12256 13716
rect 11977 13679 12035 13685
rect 12250 13676 12256 13688
rect 12308 13716 12314 13728
rect 12544 13716 12572 13815
rect 12618 13812 12624 13864
rect 12676 13852 12682 13864
rect 12989 13855 13047 13861
rect 12989 13852 13001 13855
rect 12676 13824 13001 13852
rect 12676 13812 12682 13824
rect 12989 13821 13001 13824
rect 13035 13852 13047 13855
rect 13035 13824 13308 13852
rect 13035 13821 13047 13824
rect 12989 13815 13047 13821
rect 13280 13784 13308 13824
rect 13354 13812 13360 13864
rect 13412 13812 13418 13864
rect 15028 13852 15056 13960
rect 15672 13929 15700 13960
rect 17678 13948 17684 13960
rect 17736 13948 17742 14000
rect 18325 13991 18383 13997
rect 18325 13957 18337 13991
rect 18371 13988 18383 13991
rect 18506 13988 18512 14000
rect 18371 13960 18512 13988
rect 18371 13957 18383 13960
rect 18325 13951 18383 13957
rect 18506 13948 18512 13960
rect 18564 13948 18570 14000
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13889 15715 13923
rect 15657 13883 15715 13889
rect 16761 13923 16819 13929
rect 16761 13889 16773 13923
rect 16807 13920 16819 13923
rect 17126 13920 17132 13932
rect 16807 13892 17132 13920
rect 16807 13889 16819 13892
rect 16761 13883 16819 13889
rect 17126 13880 17132 13892
rect 17184 13920 17190 13932
rect 17310 13920 17316 13932
rect 17184 13892 17316 13920
rect 17184 13880 17190 13892
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 17405 13923 17463 13929
rect 17405 13889 17417 13923
rect 17451 13920 17463 13923
rect 19518 13920 19524 13932
rect 17451 13892 19524 13920
rect 17451 13889 17463 13892
rect 17405 13883 17463 13889
rect 19518 13880 19524 13892
rect 19576 13880 19582 13932
rect 21082 13880 21088 13932
rect 21140 13880 21146 13932
rect 22020 13929 22048 14028
rect 23290 14016 23296 14028
rect 23348 14016 23354 14068
rect 24026 14016 24032 14068
rect 24084 14056 24090 14068
rect 26418 14056 26424 14068
rect 24084 14028 26424 14056
rect 24084 14016 24090 14028
rect 26418 14016 26424 14028
rect 26476 14056 26482 14068
rect 26605 14059 26663 14065
rect 26605 14056 26617 14059
rect 26476 14028 26617 14056
rect 26476 14016 26482 14028
rect 26605 14025 26617 14028
rect 26651 14025 26663 14059
rect 26605 14019 26663 14025
rect 28442 14016 28448 14068
rect 28500 14056 28506 14068
rect 28500 14028 29408 14056
rect 28500 14016 28506 14028
rect 22278 13948 22284 14000
rect 22336 13948 22342 14000
rect 24213 13991 24271 13997
rect 24213 13957 24225 13991
rect 24259 13988 24271 13991
rect 25222 13988 25228 14000
rect 24259 13960 25228 13988
rect 24259 13957 24271 13960
rect 24213 13951 24271 13957
rect 25222 13948 25228 13960
rect 25280 13948 25286 14000
rect 26786 13988 26792 14000
rect 26358 13960 26792 13988
rect 26786 13948 26792 13960
rect 26844 13988 26850 14000
rect 27062 13988 27068 14000
rect 26844 13960 27068 13988
rect 26844 13948 26850 13960
rect 27062 13948 27068 13960
rect 27120 13948 27126 14000
rect 27157 13991 27215 13997
rect 27157 13957 27169 13991
rect 27203 13988 27215 13991
rect 29270 13988 29276 14000
rect 27203 13960 29276 13988
rect 27203 13957 27215 13960
rect 27157 13951 27215 13957
rect 29270 13948 29276 13960
rect 29328 13948 29334 14000
rect 29380 13988 29408 14028
rect 30374 14016 30380 14068
rect 30432 14056 30438 14068
rect 31573 14059 31631 14065
rect 31573 14056 31585 14059
rect 30432 14028 31585 14056
rect 30432 14016 30438 14028
rect 31573 14025 31585 14028
rect 31619 14025 31631 14059
rect 31573 14019 31631 14025
rect 32766 14016 32772 14068
rect 32824 14056 32830 14068
rect 34885 14059 34943 14065
rect 34885 14056 34897 14059
rect 32824 14028 33916 14056
rect 32824 14016 32830 14028
rect 33888 13988 33916 14028
rect 34808 14028 34897 14056
rect 34808 13988 34836 14028
rect 34885 14025 34897 14028
rect 34931 14025 34943 14059
rect 34885 14019 34943 14025
rect 35066 14016 35072 14068
rect 35124 14056 35130 14068
rect 35618 14056 35624 14068
rect 35124 14028 35624 14056
rect 35124 14016 35130 14028
rect 35618 14016 35624 14028
rect 35676 14016 35682 14068
rect 35710 14016 35716 14068
rect 35768 14016 35774 14068
rect 36081 14059 36139 14065
rect 36081 14025 36093 14059
rect 36127 14056 36139 14059
rect 36817 14059 36875 14065
rect 36817 14056 36829 14059
rect 36127 14028 36829 14056
rect 36127 14025 36139 14028
rect 36081 14019 36139 14025
rect 36817 14025 36829 14028
rect 36863 14056 36875 14059
rect 37182 14056 37188 14068
rect 36863 14028 37188 14056
rect 36863 14025 36875 14028
rect 36817 14019 36875 14025
rect 34977 13991 35035 13997
rect 34977 13988 34989 13991
rect 29380 13960 30130 13988
rect 33888 13960 34836 13988
rect 34900 13960 34989 13988
rect 22005 13923 22063 13929
rect 22005 13889 22017 13923
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 13464 13824 15056 13852
rect 13464 13784 13492 13824
rect 15930 13812 15936 13864
rect 15988 13852 15994 13864
rect 15988 13824 17264 13852
rect 15988 13812 15994 13824
rect 13280 13756 13492 13784
rect 14642 13744 14648 13796
rect 14700 13784 14706 13796
rect 16390 13784 16396 13796
rect 14700 13756 16396 13784
rect 14700 13744 14706 13756
rect 16390 13744 16396 13756
rect 16448 13744 16454 13796
rect 16482 13744 16488 13796
rect 16540 13784 16546 13796
rect 17236 13793 17264 13824
rect 18138 13812 18144 13864
rect 18196 13852 18202 13864
rect 18417 13855 18475 13861
rect 18417 13852 18429 13855
rect 18196 13824 18429 13852
rect 18196 13812 18202 13824
rect 18417 13821 18429 13824
rect 18463 13821 18475 13855
rect 18417 13815 18475 13821
rect 19061 13855 19119 13861
rect 19061 13821 19073 13855
rect 19107 13852 19119 13855
rect 19610 13852 19616 13864
rect 19107 13824 19616 13852
rect 19107 13821 19119 13824
rect 19061 13815 19119 13821
rect 19610 13812 19616 13824
rect 19668 13812 19674 13864
rect 19702 13812 19708 13864
rect 19760 13812 19766 13864
rect 21100 13852 21128 13880
rect 21910 13852 21916 13864
rect 21100 13824 21916 13852
rect 21910 13812 21916 13824
rect 21968 13852 21974 13864
rect 23014 13852 23020 13864
rect 21968 13824 23020 13852
rect 21968 13812 21974 13824
rect 23014 13812 23020 13824
rect 23072 13852 23078 13864
rect 23400 13852 23428 13906
rect 24854 13880 24860 13932
rect 24912 13880 24918 13932
rect 28905 13923 28963 13929
rect 28905 13889 28917 13923
rect 28951 13920 28963 13923
rect 28994 13920 29000 13932
rect 28951 13892 29000 13920
rect 28951 13889 28963 13892
rect 28905 13883 28963 13889
rect 28994 13880 29000 13892
rect 29052 13880 29058 13932
rect 33686 13880 33692 13932
rect 33744 13880 33750 13932
rect 34422 13880 34428 13932
rect 34480 13920 34486 13932
rect 34900 13920 34928 13960
rect 34977 13957 34989 13960
rect 35023 13957 35035 13991
rect 36096 13988 36124 14019
rect 37182 14016 37188 14028
rect 37240 14016 37246 14068
rect 37274 14016 37280 14068
rect 37332 14056 37338 14068
rect 37461 14059 37519 14065
rect 37461 14056 37473 14059
rect 37332 14028 37473 14056
rect 37332 14016 37338 14028
rect 37461 14025 37473 14028
rect 37507 14025 37519 14059
rect 37461 14019 37519 14025
rect 37734 14016 37740 14068
rect 37792 14056 37798 14068
rect 37829 14059 37887 14065
rect 37829 14056 37841 14059
rect 37792 14028 37841 14056
rect 37792 14016 37798 14028
rect 37829 14025 37841 14028
rect 37875 14025 37887 14059
rect 37829 14019 37887 14025
rect 38657 14059 38715 14065
rect 38657 14025 38669 14059
rect 38703 14056 38715 14059
rect 39114 14056 39120 14068
rect 38703 14028 39120 14056
rect 38703 14025 38715 14028
rect 38657 14019 38715 14025
rect 39114 14016 39120 14028
rect 39172 14016 39178 14068
rect 40497 14059 40555 14065
rect 40497 14056 40509 14059
rect 39224 14028 40509 14056
rect 34977 13951 35035 13957
rect 35084 13960 36124 13988
rect 36173 13991 36231 13997
rect 35084 13920 35112 13960
rect 36173 13957 36185 13991
rect 36219 13988 36231 13991
rect 36354 13988 36360 14000
rect 36219 13960 36360 13988
rect 36219 13957 36231 13960
rect 36173 13951 36231 13957
rect 36354 13948 36360 13960
rect 36412 13948 36418 14000
rect 36722 13948 36728 14000
rect 36780 13988 36786 14000
rect 39224 13988 39252 14028
rect 40497 14025 40509 14028
rect 40543 14025 40555 14059
rect 40497 14019 40555 14025
rect 41325 14059 41383 14065
rect 41325 14025 41337 14059
rect 41371 14056 41383 14059
rect 41414 14056 41420 14068
rect 41371 14028 41420 14056
rect 41371 14025 41383 14028
rect 41325 14019 41383 14025
rect 41414 14016 41420 14028
rect 41472 14016 41478 14068
rect 41506 14016 41512 14068
rect 41564 14056 41570 14068
rect 41785 14059 41843 14065
rect 41785 14056 41797 14059
rect 41564 14028 41797 14056
rect 41564 14016 41570 14028
rect 41785 14025 41797 14028
rect 41831 14025 41843 14059
rect 41785 14019 41843 14025
rect 45649 14059 45707 14065
rect 45649 14025 45661 14059
rect 45695 14056 45707 14059
rect 47854 14056 47860 14068
rect 45695 14028 47860 14056
rect 45695 14025 45707 14028
rect 45649 14019 45707 14025
rect 47854 14016 47860 14028
rect 47912 14016 47918 14068
rect 48406 14016 48412 14068
rect 48464 14016 48470 14068
rect 48498 14016 48504 14068
rect 48556 14056 48562 14068
rect 49237 14059 49295 14065
rect 49237 14056 49249 14059
rect 48556 14028 49249 14056
rect 48556 14016 48562 14028
rect 49237 14025 49249 14028
rect 49283 14025 49295 14059
rect 49237 14019 49295 14025
rect 36780 13960 39252 13988
rect 36780 13948 36786 13960
rect 39298 13948 39304 14000
rect 39356 13988 39362 14000
rect 45005 13991 45063 13997
rect 45005 13988 45017 13991
rect 39356 13960 45017 13988
rect 39356 13948 39362 13960
rect 45005 13957 45017 13960
rect 45051 13957 45063 13991
rect 45005 13951 45063 13957
rect 48133 13991 48191 13997
rect 48133 13957 48145 13991
rect 48179 13988 48191 13991
rect 49142 13988 49148 14000
rect 48179 13960 49148 13988
rect 48179 13957 48191 13960
rect 48133 13951 48191 13957
rect 49142 13948 49148 13960
rect 49200 13948 49206 14000
rect 34480 13892 34928 13920
rect 34992 13892 35112 13920
rect 34480 13880 34486 13892
rect 23072 13824 23428 13852
rect 23072 13812 23078 13824
rect 23474 13812 23480 13864
rect 23532 13852 23538 13864
rect 23753 13855 23811 13861
rect 23753 13852 23765 13855
rect 23532 13824 23765 13852
rect 23532 13812 23538 13824
rect 23753 13821 23765 13824
rect 23799 13821 23811 13855
rect 23753 13815 23811 13821
rect 25130 13812 25136 13864
rect 25188 13812 25194 13864
rect 29365 13855 29423 13861
rect 29365 13821 29377 13855
rect 29411 13821 29423 13855
rect 29365 13815 29423 13821
rect 29641 13855 29699 13861
rect 29641 13821 29653 13855
rect 29687 13852 29699 13855
rect 29687 13824 30696 13852
rect 29687 13821 29699 13824
rect 29641 13815 29699 13821
rect 17221 13787 17279 13793
rect 16540 13756 17172 13784
rect 16540 13744 16546 13756
rect 12308 13688 12572 13716
rect 13620 13719 13678 13725
rect 12308 13676 12314 13688
rect 13620 13685 13632 13719
rect 13666 13716 13678 13719
rect 13998 13716 14004 13728
rect 13666 13688 14004 13716
rect 13666 13685 13678 13688
rect 13620 13679 13678 13685
rect 13998 13676 14004 13688
rect 14056 13676 14062 13728
rect 16298 13676 16304 13728
rect 16356 13716 16362 13728
rect 16942 13716 16948 13728
rect 16356 13688 16948 13716
rect 16356 13676 16362 13688
rect 16942 13676 16948 13688
rect 17000 13676 17006 13728
rect 17144 13716 17172 13756
rect 17221 13753 17233 13787
rect 17267 13753 17279 13787
rect 17221 13747 17279 13753
rect 29380 13728 29408 13815
rect 30668 13784 30696 13824
rect 30834 13812 30840 13864
rect 30892 13852 30898 13864
rect 31113 13855 31171 13861
rect 31113 13852 31125 13855
rect 30892 13824 31125 13852
rect 30892 13812 30898 13824
rect 31113 13821 31125 13824
rect 31159 13821 31171 13855
rect 31113 13815 31171 13821
rect 32214 13812 32220 13864
rect 32272 13852 32278 13864
rect 32309 13855 32367 13861
rect 32309 13852 32321 13855
rect 32272 13824 32321 13852
rect 32272 13812 32278 13824
rect 32309 13821 32321 13824
rect 32355 13821 32367 13855
rect 32309 13815 32367 13821
rect 32582 13812 32588 13864
rect 32640 13812 32646 13864
rect 33134 13812 33140 13864
rect 33192 13852 33198 13864
rect 33594 13852 33600 13864
rect 33192 13824 33600 13852
rect 33192 13812 33198 13824
rect 33594 13812 33600 13824
rect 33652 13852 33658 13864
rect 33652 13824 34008 13852
rect 33652 13812 33658 13824
rect 31846 13784 31852 13796
rect 30668 13756 31852 13784
rect 31846 13744 31852 13756
rect 31904 13744 31910 13796
rect 33980 13784 34008 13824
rect 34054 13812 34060 13864
rect 34112 13852 34118 13864
rect 34514 13852 34520 13864
rect 34112 13824 34520 13852
rect 34112 13812 34118 13824
rect 34514 13812 34520 13824
rect 34572 13812 34578 13864
rect 34992 13852 35020 13892
rect 36538 13880 36544 13932
rect 36596 13920 36602 13932
rect 37734 13920 37740 13932
rect 36596 13892 37740 13920
rect 36596 13880 36602 13892
rect 37734 13880 37740 13892
rect 37792 13880 37798 13932
rect 39025 13923 39083 13929
rect 39025 13920 39037 13923
rect 37844 13892 39037 13920
rect 34624 13824 35020 13852
rect 35069 13855 35127 13861
rect 34624 13784 34652 13824
rect 35069 13821 35081 13855
rect 35115 13821 35127 13855
rect 35069 13815 35127 13821
rect 36265 13855 36323 13861
rect 36265 13821 36277 13855
rect 36311 13821 36323 13855
rect 36265 13815 36323 13821
rect 33980 13756 34652 13784
rect 35084 13728 35112 13815
rect 36078 13744 36084 13796
rect 36136 13784 36142 13796
rect 36280 13784 36308 13815
rect 37090 13812 37096 13864
rect 37148 13852 37154 13864
rect 37844 13852 37872 13892
rect 39025 13889 39037 13892
rect 39071 13889 39083 13923
rect 39025 13883 39083 13889
rect 39206 13880 39212 13932
rect 39264 13920 39270 13932
rect 39264 13892 39804 13920
rect 39264 13880 39270 13892
rect 37148 13824 37872 13852
rect 37148 13812 37154 13824
rect 37918 13812 37924 13864
rect 37976 13812 37982 13864
rect 38105 13855 38163 13861
rect 38105 13821 38117 13855
rect 38151 13821 38163 13855
rect 38105 13815 38163 13821
rect 36136 13756 36308 13784
rect 36136 13744 36142 13756
rect 19962 13719 20020 13725
rect 19962 13716 19974 13719
rect 17144 13688 19974 13716
rect 19962 13685 19974 13688
rect 20008 13685 20020 13719
rect 19962 13679 20020 13685
rect 20070 13676 20076 13728
rect 20128 13716 20134 13728
rect 28534 13716 28540 13728
rect 20128 13688 28540 13716
rect 20128 13676 20134 13688
rect 28534 13676 28540 13688
rect 28592 13676 28598 13728
rect 29362 13676 29368 13728
rect 29420 13716 29426 13728
rect 30282 13716 30288 13728
rect 29420 13688 30288 13716
rect 29420 13676 29426 13688
rect 30282 13676 30288 13688
rect 30340 13676 30346 13728
rect 31294 13676 31300 13728
rect 31352 13716 31358 13728
rect 33962 13716 33968 13728
rect 31352 13688 33968 13716
rect 31352 13676 31358 13688
rect 33962 13676 33968 13688
rect 34020 13676 34026 13728
rect 34517 13719 34575 13725
rect 34517 13685 34529 13719
rect 34563 13716 34575 13719
rect 34974 13716 34980 13728
rect 34563 13688 34980 13716
rect 34563 13685 34575 13688
rect 34517 13679 34575 13685
rect 34974 13676 34980 13688
rect 35032 13676 35038 13728
rect 35066 13676 35072 13728
rect 35124 13676 35130 13728
rect 36170 13676 36176 13728
rect 36228 13716 36234 13728
rect 36909 13719 36967 13725
rect 36909 13716 36921 13719
rect 36228 13688 36921 13716
rect 36228 13676 36234 13688
rect 36909 13685 36921 13688
rect 36955 13716 36967 13719
rect 37182 13716 37188 13728
rect 36955 13688 37188 13716
rect 36955 13685 36967 13688
rect 36909 13679 36967 13685
rect 37182 13676 37188 13688
rect 37240 13676 37246 13728
rect 38120 13716 38148 13815
rect 38286 13812 38292 13864
rect 38344 13852 38350 13864
rect 39117 13855 39175 13861
rect 39117 13852 39129 13855
rect 38344 13824 39129 13852
rect 38344 13812 38350 13824
rect 39117 13821 39129 13824
rect 39163 13821 39175 13855
rect 39117 13815 39175 13821
rect 39301 13855 39359 13861
rect 39301 13821 39313 13855
rect 39347 13821 39359 13855
rect 39776 13852 39804 13892
rect 39850 13880 39856 13932
rect 39908 13880 39914 13932
rect 40862 13880 40868 13932
rect 40920 13880 40926 13932
rect 40954 13880 40960 13932
rect 41012 13880 41018 13932
rect 41509 13923 41567 13929
rect 41509 13889 41521 13923
rect 41555 13889 41567 13923
rect 41509 13883 41567 13889
rect 41524 13852 41552 13883
rect 45830 13880 45836 13932
rect 45888 13880 45894 13932
rect 48222 13880 48228 13932
rect 48280 13920 48286 13932
rect 48593 13923 48651 13929
rect 48593 13920 48605 13923
rect 48280 13892 48605 13920
rect 48280 13880 48286 13892
rect 48593 13889 48605 13892
rect 48639 13889 48651 13923
rect 48593 13883 48651 13889
rect 39776 13824 41552 13852
rect 45189 13855 45247 13861
rect 39301 13815 39359 13821
rect 45189 13821 45201 13855
rect 45235 13852 45247 13855
rect 46566 13852 46572 13864
rect 45235 13824 46572 13852
rect 45235 13821 45247 13824
rect 45189 13815 45247 13821
rect 38194 13744 38200 13796
rect 38252 13784 38258 13796
rect 39316 13784 39344 13815
rect 46566 13812 46572 13824
rect 46624 13812 46630 13864
rect 41138 13784 41144 13796
rect 38252 13756 41144 13784
rect 38252 13744 38258 13756
rect 41138 13744 41144 13756
rect 41196 13744 41202 13796
rect 41046 13716 41052 13728
rect 38120 13688 41052 13716
rect 41046 13676 41052 13688
rect 41104 13676 41110 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 9030 13472 9036 13524
rect 9088 13512 9094 13524
rect 9585 13515 9643 13521
rect 9585 13512 9597 13515
rect 9088 13484 9597 13512
rect 9088 13472 9094 13484
rect 9585 13481 9597 13484
rect 9631 13512 9643 13515
rect 11136 13515 11194 13521
rect 11136 13512 11148 13515
rect 9631 13484 11148 13512
rect 9631 13481 9643 13484
rect 9585 13475 9643 13481
rect 11136 13481 11148 13484
rect 11182 13512 11194 13515
rect 13081 13515 13139 13521
rect 13081 13512 13093 13515
rect 11182 13484 13093 13512
rect 11182 13481 11194 13484
rect 11136 13475 11194 13481
rect 13081 13481 13093 13484
rect 13127 13512 13139 13515
rect 13814 13512 13820 13524
rect 13127 13484 13820 13512
rect 13127 13481 13139 13484
rect 13081 13475 13139 13481
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 14458 13472 14464 13524
rect 14516 13472 14522 13524
rect 15194 13472 15200 13524
rect 15252 13472 15258 13524
rect 15562 13472 15568 13524
rect 15620 13512 15626 13524
rect 16393 13515 16451 13521
rect 16393 13512 16405 13515
rect 15620 13484 16405 13512
rect 15620 13472 15626 13484
rect 16393 13481 16405 13484
rect 16439 13481 16451 13515
rect 16393 13475 16451 13481
rect 18693 13515 18751 13521
rect 18693 13481 18705 13515
rect 18739 13512 18751 13515
rect 19242 13512 19248 13524
rect 18739 13484 19248 13512
rect 18739 13481 18751 13484
rect 18693 13475 18751 13481
rect 19242 13472 19248 13484
rect 19300 13472 19306 13524
rect 19521 13515 19579 13521
rect 19521 13481 19533 13515
rect 19567 13512 19579 13515
rect 19886 13512 19892 13524
rect 19567 13484 19892 13512
rect 19567 13481 19579 13484
rect 19521 13475 19579 13481
rect 19886 13472 19892 13484
rect 19944 13472 19950 13524
rect 19978 13472 19984 13524
rect 20036 13512 20042 13524
rect 20717 13515 20775 13521
rect 20717 13512 20729 13515
rect 20036 13484 20729 13512
rect 20036 13472 20042 13484
rect 20717 13481 20729 13484
rect 20763 13481 20775 13515
rect 20717 13475 20775 13481
rect 21358 13472 21364 13524
rect 21416 13512 21422 13524
rect 21913 13515 21971 13521
rect 21913 13512 21925 13515
rect 21416 13484 21925 13512
rect 21416 13472 21422 13484
rect 21913 13481 21925 13484
rect 21959 13481 21971 13515
rect 21913 13475 21971 13481
rect 22388 13484 23244 13512
rect 12434 13404 12440 13456
rect 12492 13444 12498 13456
rect 12802 13444 12808 13456
rect 12492 13416 12808 13444
rect 12492 13404 12498 13416
rect 12802 13404 12808 13416
rect 12860 13404 12866 13456
rect 13265 13447 13323 13453
rect 13265 13413 13277 13447
rect 13311 13444 13323 13447
rect 14182 13444 14188 13456
rect 13311 13416 14188 13444
rect 13311 13413 13323 13416
rect 13265 13407 13323 13413
rect 14182 13404 14188 13416
rect 14240 13404 14246 13456
rect 18138 13444 18144 13456
rect 16500 13416 18144 13444
rect 2774 13336 2780 13388
rect 2832 13336 2838 13388
rect 9769 13379 9827 13385
rect 9769 13345 9781 13379
rect 9815 13376 9827 13379
rect 9858 13376 9864 13388
rect 9815 13348 9864 13376
rect 9815 13345 9827 13348
rect 9769 13339 9827 13345
rect 9858 13336 9864 13348
rect 9916 13376 9922 13388
rect 11514 13376 11520 13388
rect 9916 13348 11520 13376
rect 9916 13336 9922 13348
rect 11514 13336 11520 13348
rect 11572 13336 11578 13388
rect 12526 13336 12532 13388
rect 12584 13376 12590 13388
rect 12621 13379 12679 13385
rect 12621 13376 12633 13379
rect 12584 13348 12633 13376
rect 12584 13336 12590 13348
rect 12621 13345 12633 13348
rect 12667 13376 12679 13379
rect 13538 13376 13544 13388
rect 12667 13348 13544 13376
rect 12667 13345 12679 13348
rect 12621 13339 12679 13345
rect 13538 13336 13544 13348
rect 13596 13336 13602 13388
rect 15654 13336 15660 13388
rect 15712 13336 15718 13388
rect 15841 13379 15899 13385
rect 15841 13345 15853 13379
rect 15887 13376 15899 13379
rect 16500 13376 16528 13416
rect 18138 13404 18144 13416
rect 18196 13444 18202 13456
rect 18598 13444 18604 13456
rect 18196 13416 18604 13444
rect 18196 13404 18202 13416
rect 18598 13404 18604 13416
rect 18656 13404 18662 13456
rect 18877 13447 18935 13453
rect 18877 13413 18889 13447
rect 18923 13444 18935 13447
rect 19058 13444 19064 13456
rect 18923 13416 19064 13444
rect 18923 13413 18935 13416
rect 18877 13407 18935 13413
rect 19058 13404 19064 13416
rect 19116 13404 19122 13456
rect 19260 13444 19288 13472
rect 19260 13416 20208 13444
rect 16853 13379 16911 13385
rect 16853 13376 16865 13379
rect 15887 13348 16528 13376
rect 16776 13348 16865 13376
rect 15887 13345 15899 13348
rect 15841 13339 15899 13345
rect 1762 13268 1768 13320
rect 1820 13268 1826 13320
rect 6914 13268 6920 13320
rect 6972 13308 6978 13320
rect 6972 13280 10088 13308
rect 6972 13268 6978 13280
rect 9950 13200 9956 13252
rect 10008 13200 10014 13252
rect 10060 13240 10088 13280
rect 10870 13268 10876 13320
rect 10928 13268 10934 13320
rect 13354 13268 13360 13320
rect 13412 13308 13418 13320
rect 13722 13308 13728 13320
rect 13412 13280 13728 13308
rect 13412 13268 13418 13280
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 15565 13311 15623 13317
rect 15565 13277 15577 13311
rect 15611 13308 15623 13311
rect 16206 13308 16212 13320
rect 15611 13280 16212 13308
rect 15611 13277 15623 13280
rect 15565 13271 15623 13277
rect 16206 13268 16212 13280
rect 16264 13268 16270 13320
rect 16482 13308 16488 13320
rect 16316 13280 16488 13308
rect 11054 13240 11060 13252
rect 10060 13212 11060 13240
rect 11054 13200 11060 13212
rect 11112 13200 11118 13252
rect 11606 13200 11612 13252
rect 11664 13200 11670 13252
rect 13541 13243 13599 13249
rect 13541 13209 13553 13243
rect 13587 13240 13599 13243
rect 14274 13240 14280 13252
rect 13587 13212 14280 13240
rect 13587 13209 13599 13212
rect 13541 13203 13599 13209
rect 14274 13200 14280 13212
rect 14332 13200 14338 13252
rect 14366 13200 14372 13252
rect 14424 13200 14430 13252
rect 15378 13200 15384 13252
rect 15436 13240 15442 13252
rect 16316 13240 16344 13280
rect 16482 13268 16488 13280
rect 16540 13308 16546 13320
rect 16776 13308 16804 13348
rect 16853 13345 16865 13348
rect 16899 13345 16911 13379
rect 16853 13339 16911 13345
rect 17037 13379 17095 13385
rect 17037 13345 17049 13379
rect 17083 13376 17095 13379
rect 17310 13376 17316 13388
rect 17083 13348 17316 13376
rect 17083 13345 17095 13348
rect 17037 13339 17095 13345
rect 17310 13336 17316 13348
rect 17368 13336 17374 13388
rect 17494 13336 17500 13388
rect 17552 13376 17558 13388
rect 18233 13379 18291 13385
rect 18233 13376 18245 13379
rect 17552 13348 18245 13376
rect 17552 13336 17558 13348
rect 18233 13345 18245 13348
rect 18279 13345 18291 13379
rect 18233 13339 18291 13345
rect 19794 13336 19800 13388
rect 19852 13376 19858 13388
rect 20073 13379 20131 13385
rect 20073 13376 20085 13379
rect 19852 13348 20085 13376
rect 19852 13336 19858 13348
rect 20073 13345 20085 13348
rect 20119 13345 20131 13379
rect 20073 13339 20131 13345
rect 16540 13280 16804 13308
rect 16540 13268 16546 13280
rect 17954 13268 17960 13320
rect 18012 13268 18018 13320
rect 18049 13311 18107 13317
rect 18049 13277 18061 13311
rect 18095 13308 18107 13311
rect 18414 13308 18420 13320
rect 18095 13280 18420 13308
rect 18095 13277 18107 13280
rect 18049 13271 18107 13277
rect 18414 13268 18420 13280
rect 18472 13268 18478 13320
rect 19610 13268 19616 13320
rect 19668 13308 19674 13320
rect 19889 13311 19947 13317
rect 19889 13308 19901 13311
rect 19668 13280 19901 13308
rect 19668 13268 19674 13280
rect 19889 13277 19901 13280
rect 19935 13277 19947 13311
rect 20180 13308 20208 13416
rect 21358 13336 21364 13388
rect 21416 13376 21422 13388
rect 22388 13385 22416 13484
rect 23106 13404 23112 13456
rect 23164 13404 23170 13456
rect 23216 13444 23244 13484
rect 23842 13472 23848 13524
rect 23900 13512 23906 13524
rect 24121 13515 24179 13521
rect 24121 13512 24133 13515
rect 23900 13484 24133 13512
rect 23900 13472 23906 13484
rect 24121 13481 24133 13484
rect 24167 13481 24179 13515
rect 24121 13475 24179 13481
rect 24857 13515 24915 13521
rect 24857 13481 24869 13515
rect 24903 13512 24915 13515
rect 24946 13512 24952 13524
rect 24903 13484 24952 13512
rect 24903 13481 24915 13484
rect 24857 13475 24915 13481
rect 24946 13472 24952 13484
rect 25004 13472 25010 13524
rect 25130 13472 25136 13524
rect 25188 13512 25194 13524
rect 26697 13515 26755 13521
rect 26697 13512 26709 13515
rect 25188 13484 26709 13512
rect 25188 13472 25194 13484
rect 26697 13481 26709 13484
rect 26743 13481 26755 13515
rect 26697 13475 26755 13481
rect 28997 13515 29055 13521
rect 28997 13481 29009 13515
rect 29043 13512 29055 13515
rect 29086 13512 29092 13524
rect 29043 13484 29092 13512
rect 29043 13481 29055 13484
rect 28997 13475 29055 13481
rect 29086 13472 29092 13484
rect 29144 13472 29150 13524
rect 29365 13515 29423 13521
rect 29365 13481 29377 13515
rect 29411 13512 29423 13515
rect 29454 13512 29460 13524
rect 29411 13484 29460 13512
rect 29411 13481 29423 13484
rect 29365 13475 29423 13481
rect 29454 13472 29460 13484
rect 29512 13472 29518 13524
rect 34422 13512 34428 13524
rect 29564 13484 34428 13512
rect 27430 13444 27436 13456
rect 23216 13416 27436 13444
rect 27430 13404 27436 13416
rect 27488 13404 27494 13456
rect 27614 13404 27620 13456
rect 27672 13444 27678 13456
rect 29564 13444 29592 13484
rect 34422 13472 34428 13484
rect 34480 13472 34486 13524
rect 34514 13472 34520 13524
rect 34572 13512 34578 13524
rect 34572 13484 38043 13512
rect 34572 13472 34578 13484
rect 30834 13444 30840 13456
rect 27672 13416 29592 13444
rect 30116 13416 30840 13444
rect 27672 13404 27678 13416
rect 22373 13379 22431 13385
rect 21416 13348 22324 13376
rect 21416 13336 21422 13348
rect 21085 13311 21143 13317
rect 21085 13308 21097 13311
rect 20180 13280 21097 13308
rect 19889 13271 19947 13277
rect 21085 13277 21097 13280
rect 21131 13308 21143 13311
rect 21266 13308 21272 13320
rect 21131 13280 21272 13308
rect 21131 13277 21143 13280
rect 21085 13271 21143 13277
rect 21266 13268 21272 13280
rect 21324 13308 21330 13320
rect 22094 13308 22100 13320
rect 21324 13280 22100 13308
rect 21324 13268 21330 13280
rect 22094 13268 22100 13280
rect 22152 13268 22158 13320
rect 15436 13212 16344 13240
rect 15436 13200 15442 13212
rect 16574 13200 16580 13252
rect 16632 13240 16638 13252
rect 16761 13243 16819 13249
rect 16761 13240 16773 13243
rect 16632 13212 16773 13240
rect 16632 13200 16638 13212
rect 16761 13209 16773 13212
rect 16807 13209 16819 13243
rect 18969 13243 19027 13249
rect 18969 13240 18981 13243
rect 16761 13203 16819 13209
rect 16868 13212 18981 13240
rect 10229 13175 10287 13181
rect 10229 13141 10241 13175
rect 10275 13172 10287 13175
rect 12066 13172 12072 13184
rect 10275 13144 12072 13172
rect 10275 13141 10287 13144
rect 10229 13135 10287 13141
rect 12066 13132 12072 13144
rect 12124 13132 12130 13184
rect 14826 13132 14832 13184
rect 14884 13132 14890 13184
rect 14918 13132 14924 13184
rect 14976 13172 14982 13184
rect 16868 13172 16896 13212
rect 18969 13209 18981 13212
rect 19015 13209 19027 13243
rect 18969 13203 19027 13209
rect 14976 13144 16896 13172
rect 14976 13132 14982 13144
rect 17586 13132 17592 13184
rect 17644 13132 17650 13184
rect 18984 13172 19012 13203
rect 19058 13200 19064 13252
rect 19116 13240 19122 13252
rect 19981 13243 20039 13249
rect 19981 13240 19993 13243
rect 19116 13212 19993 13240
rect 19116 13200 19122 13212
rect 19981 13209 19993 13212
rect 20027 13209 20039 13243
rect 22296 13240 22324 13348
rect 22373 13345 22385 13379
rect 22419 13345 22431 13379
rect 22373 13339 22431 13345
rect 22557 13379 22615 13385
rect 22557 13345 22569 13379
rect 22603 13345 22615 13379
rect 22557 13339 22615 13345
rect 22572 13308 22600 13339
rect 23750 13336 23756 13388
rect 23808 13336 23814 13388
rect 25409 13379 25467 13385
rect 25409 13345 25421 13379
rect 25455 13376 25467 13379
rect 27798 13376 27804 13388
rect 25455 13348 27804 13376
rect 25455 13345 25467 13348
rect 25409 13339 25467 13345
rect 27798 13336 27804 13348
rect 27856 13376 27862 13388
rect 30116 13376 30144 13416
rect 30834 13404 30840 13416
rect 30892 13404 30898 13456
rect 32950 13404 32956 13456
rect 33008 13444 33014 13456
rect 33008 13416 34100 13444
rect 33008 13404 33014 13416
rect 27856 13348 30144 13376
rect 27856 13336 27862 13348
rect 24946 13308 24952 13320
rect 22572 13280 24952 13308
rect 24946 13268 24952 13280
rect 25004 13268 25010 13320
rect 25222 13268 25228 13320
rect 25280 13268 25286 13320
rect 25498 13268 25504 13320
rect 25556 13308 25562 13320
rect 26053 13311 26111 13317
rect 26053 13308 26065 13311
rect 25556 13280 26065 13308
rect 25556 13268 25562 13280
rect 26053 13277 26065 13280
rect 26099 13277 26111 13311
rect 26053 13271 26111 13277
rect 27062 13268 27068 13320
rect 27120 13308 27126 13320
rect 28368 13317 28396 13348
rect 30190 13336 30196 13388
rect 30248 13376 30254 13388
rect 30285 13379 30343 13385
rect 30285 13376 30297 13379
rect 30248 13348 30297 13376
rect 30248 13336 30254 13348
rect 30285 13345 30297 13348
rect 30331 13345 30343 13379
rect 30285 13339 30343 13345
rect 31205 13379 31263 13385
rect 31205 13345 31217 13379
rect 31251 13376 31263 13379
rect 32214 13376 32220 13388
rect 31251 13348 32220 13376
rect 31251 13345 31263 13348
rect 31205 13339 31263 13345
rect 32214 13336 32220 13348
rect 32272 13336 32278 13388
rect 33962 13336 33968 13388
rect 34020 13336 34026 13388
rect 34072 13385 34100 13416
rect 35710 13404 35716 13456
rect 35768 13444 35774 13456
rect 35768 13416 36032 13444
rect 35768 13404 35774 13416
rect 34057 13379 34115 13385
rect 34057 13345 34069 13379
rect 34103 13345 34115 13379
rect 34057 13339 34115 13345
rect 34146 13336 34152 13388
rect 34204 13376 34210 13388
rect 34204 13348 35940 13376
rect 34204 13336 34210 13348
rect 27157 13311 27215 13317
rect 27157 13308 27169 13311
rect 27120 13280 27169 13308
rect 27120 13268 27126 13280
rect 27157 13277 27169 13280
rect 27203 13277 27215 13311
rect 27157 13271 27215 13277
rect 28353 13311 28411 13317
rect 28353 13277 28365 13311
rect 28399 13277 28411 13311
rect 28353 13271 28411 13277
rect 30098 13268 30104 13320
rect 30156 13268 30162 13320
rect 32858 13268 32864 13320
rect 32916 13308 32922 13320
rect 33873 13311 33931 13317
rect 33873 13308 33885 13311
rect 32916 13280 33885 13308
rect 32916 13268 32922 13280
rect 33873 13277 33885 13280
rect 33919 13277 33931 13311
rect 33873 13271 33931 13277
rect 34606 13268 34612 13320
rect 34664 13308 34670 13320
rect 34885 13311 34943 13317
rect 34885 13308 34897 13311
rect 34664 13280 34897 13308
rect 34664 13268 34670 13280
rect 34885 13277 34897 13280
rect 34931 13277 34943 13311
rect 34885 13271 34943 13277
rect 22738 13240 22744 13252
rect 22296 13212 22744 13240
rect 19981 13203 20039 13209
rect 22738 13200 22744 13212
rect 22796 13200 22802 13252
rect 23569 13243 23627 13249
rect 23569 13209 23581 13243
rect 23615 13240 23627 13243
rect 25866 13240 25872 13252
rect 23615 13212 25872 13240
rect 23615 13209 23627 13212
rect 23569 13203 23627 13209
rect 25866 13200 25872 13212
rect 25924 13200 25930 13252
rect 29748 13212 31432 13240
rect 20070 13172 20076 13184
rect 18984 13144 20076 13172
rect 20070 13132 20076 13144
rect 20128 13132 20134 13184
rect 20254 13132 20260 13184
rect 20312 13172 20318 13184
rect 21177 13175 21235 13181
rect 21177 13172 21189 13175
rect 20312 13144 21189 13172
rect 20312 13132 20318 13144
rect 21177 13141 21189 13144
rect 21223 13172 21235 13175
rect 21634 13172 21640 13184
rect 21223 13144 21640 13172
rect 21223 13141 21235 13144
rect 21177 13135 21235 13141
rect 21634 13132 21640 13144
rect 21692 13132 21698 13184
rect 22278 13132 22284 13184
rect 22336 13132 22342 13184
rect 23198 13132 23204 13184
rect 23256 13172 23262 13184
rect 23477 13175 23535 13181
rect 23477 13172 23489 13175
rect 23256 13144 23489 13172
rect 23256 13132 23262 13144
rect 23477 13141 23489 13144
rect 23523 13141 23535 13175
rect 23477 13135 23535 13141
rect 24486 13132 24492 13184
rect 24544 13172 24550 13184
rect 25317 13175 25375 13181
rect 25317 13172 25329 13175
rect 24544 13144 25329 13172
rect 24544 13132 24550 13144
rect 25317 13141 25329 13144
rect 25363 13172 25375 13175
rect 26050 13172 26056 13184
rect 25363 13144 26056 13172
rect 25363 13141 25375 13144
rect 25317 13135 25375 13141
rect 26050 13132 26056 13144
rect 26108 13132 26114 13184
rect 26970 13132 26976 13184
rect 27028 13172 27034 13184
rect 29748 13181 29776 13212
rect 27801 13175 27859 13181
rect 27801 13172 27813 13175
rect 27028 13144 27813 13172
rect 27028 13132 27034 13144
rect 27801 13141 27813 13144
rect 27847 13141 27859 13175
rect 27801 13135 27859 13141
rect 29733 13175 29791 13181
rect 29733 13141 29745 13175
rect 29779 13141 29791 13175
rect 29733 13135 29791 13141
rect 30006 13132 30012 13184
rect 30064 13172 30070 13184
rect 30193 13175 30251 13181
rect 30193 13172 30205 13175
rect 30064 13144 30205 13172
rect 30064 13132 30070 13144
rect 30193 13141 30205 13144
rect 30239 13141 30251 13175
rect 30193 13135 30251 13141
rect 30466 13132 30472 13184
rect 30524 13172 30530 13184
rect 30745 13175 30803 13181
rect 30745 13172 30757 13175
rect 30524 13144 30757 13172
rect 30524 13132 30530 13144
rect 30745 13141 30757 13144
rect 30791 13141 30803 13175
rect 31404 13172 31432 13212
rect 31478 13200 31484 13252
rect 31536 13200 31542 13252
rect 31938 13200 31944 13252
rect 31996 13200 32002 13252
rect 33318 13200 33324 13252
rect 33376 13240 33382 13252
rect 33594 13240 33600 13252
rect 33376 13212 33600 13240
rect 33376 13200 33382 13212
rect 33594 13200 33600 13212
rect 33652 13200 33658 13252
rect 34900 13240 34928 13271
rect 35710 13268 35716 13320
rect 35768 13268 35774 13320
rect 35802 13240 35808 13252
rect 34900 13212 35808 13240
rect 35802 13200 35808 13212
rect 35860 13200 35866 13252
rect 32122 13172 32128 13184
rect 31404 13144 32128 13172
rect 30745 13135 30803 13141
rect 32122 13132 32128 13144
rect 32180 13132 32186 13184
rect 32306 13132 32312 13184
rect 32364 13172 32370 13184
rect 32953 13175 33011 13181
rect 32953 13172 32965 13175
rect 32364 13144 32965 13172
rect 32364 13132 32370 13144
rect 32953 13141 32965 13144
rect 32999 13141 33011 13175
rect 32953 13135 33011 13141
rect 33505 13175 33563 13181
rect 33505 13141 33517 13175
rect 33551 13172 33563 13175
rect 35342 13172 35348 13184
rect 33551 13144 35348 13172
rect 33551 13141 33563 13144
rect 33505 13135 33563 13141
rect 35342 13132 35348 13144
rect 35400 13132 35406 13184
rect 35912 13172 35940 13348
rect 36004 13308 36032 13416
rect 36170 13404 36176 13456
rect 36228 13404 36234 13456
rect 36722 13336 36728 13388
rect 36780 13336 36786 13388
rect 36446 13308 36452 13320
rect 36004 13280 36452 13308
rect 36446 13268 36452 13280
rect 36504 13268 36510 13320
rect 38015 13308 38043 13484
rect 38194 13472 38200 13524
rect 38252 13472 38258 13524
rect 38562 13336 38568 13388
rect 38620 13376 38626 13388
rect 38620 13348 38792 13376
rect 38620 13336 38626 13348
rect 38657 13311 38715 13317
rect 38657 13308 38669 13311
rect 38015 13280 38669 13308
rect 38657 13277 38669 13280
rect 38703 13277 38715 13311
rect 38764 13308 38792 13348
rect 40037 13311 40095 13317
rect 40037 13308 40049 13311
rect 38764 13280 40049 13308
rect 38657 13271 38715 13277
rect 40037 13277 40049 13280
rect 40083 13277 40095 13311
rect 40037 13271 40095 13277
rect 41138 13268 41144 13320
rect 41196 13268 41202 13320
rect 46566 13268 46572 13320
rect 46624 13308 46630 13320
rect 47949 13311 48007 13317
rect 47949 13308 47961 13311
rect 46624 13280 47961 13308
rect 46624 13268 46630 13280
rect 47949 13277 47961 13280
rect 47995 13277 48007 13311
rect 47949 13271 48007 13277
rect 49142 13268 49148 13320
rect 49200 13268 49206 13320
rect 37182 13200 37188 13252
rect 37240 13200 37246 13252
rect 38746 13200 38752 13252
rect 38804 13240 38810 13252
rect 40681 13243 40739 13249
rect 40681 13240 40693 13243
rect 38804 13212 40693 13240
rect 38804 13200 38810 13212
rect 40681 13209 40693 13212
rect 40727 13209 40739 13243
rect 40681 13203 40739 13209
rect 39022 13172 39028 13184
rect 35912 13144 39028 13172
rect 39022 13132 39028 13144
rect 39080 13132 39086 13184
rect 39298 13132 39304 13184
rect 39356 13132 39362 13184
rect 39574 13132 39580 13184
rect 39632 13132 39638 13184
rect 41782 13132 41788 13184
rect 41840 13132 41846 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 2869 12971 2927 12977
rect 2869 12937 2881 12971
rect 2915 12968 2927 12971
rect 5626 12968 5632 12980
rect 2915 12940 5632 12968
rect 2915 12937 2927 12940
rect 2869 12931 2927 12937
rect 5626 12928 5632 12940
rect 5684 12928 5690 12980
rect 9858 12928 9864 12980
rect 9916 12928 9922 12980
rect 10410 12928 10416 12980
rect 10468 12968 10474 12980
rect 10873 12971 10931 12977
rect 10873 12968 10885 12971
rect 10468 12940 10885 12968
rect 10468 12928 10474 12940
rect 10873 12937 10885 12940
rect 10919 12937 10931 12971
rect 10873 12931 10931 12937
rect 11054 12928 11060 12980
rect 11112 12968 11118 12980
rect 11112 12940 11928 12968
rect 11112 12928 11118 12940
rect 1302 12792 1308 12844
rect 1360 12832 1366 12844
rect 3053 12835 3111 12841
rect 3053 12832 3065 12835
rect 1360 12804 3065 12832
rect 1360 12792 1366 12804
rect 3053 12801 3065 12804
rect 3099 12832 3111 12835
rect 3329 12835 3387 12841
rect 3329 12832 3341 12835
rect 3099 12804 3341 12832
rect 3099 12801 3111 12804
rect 3053 12795 3111 12801
rect 3329 12801 3341 12804
rect 3375 12801 3387 12835
rect 3329 12795 3387 12801
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12832 10839 12835
rect 11330 12832 11336 12844
rect 10827 12804 11336 12832
rect 10827 12801 10839 12804
rect 10781 12795 10839 12801
rect 11330 12792 11336 12804
rect 11388 12792 11394 12844
rect 11900 12832 11928 12940
rect 12066 12928 12072 12980
rect 12124 12928 12130 12980
rect 12250 12928 12256 12980
rect 12308 12968 12314 12980
rect 14829 12971 14887 12977
rect 14829 12968 14841 12971
rect 12308 12940 14841 12968
rect 12308 12928 12314 12940
rect 14829 12937 14841 12940
rect 14875 12937 14887 12971
rect 14829 12931 14887 12937
rect 15930 12928 15936 12980
rect 15988 12928 15994 12980
rect 16850 12928 16856 12980
rect 16908 12968 16914 12980
rect 19702 12968 19708 12980
rect 16908 12940 19708 12968
rect 16908 12928 16914 12940
rect 19702 12928 19708 12940
rect 19760 12928 19766 12980
rect 21085 12971 21143 12977
rect 21085 12937 21097 12971
rect 21131 12968 21143 12971
rect 22646 12968 22652 12980
rect 21131 12940 22652 12968
rect 21131 12937 21143 12940
rect 21085 12931 21143 12937
rect 22646 12928 22652 12940
rect 22704 12928 22710 12980
rect 22741 12971 22799 12977
rect 22741 12937 22753 12971
rect 22787 12968 22799 12971
rect 23566 12968 23572 12980
rect 22787 12940 23572 12968
rect 22787 12937 22799 12940
rect 22741 12931 22799 12937
rect 23566 12928 23572 12940
rect 23624 12928 23630 12980
rect 23750 12928 23756 12980
rect 23808 12968 23814 12980
rect 25685 12971 25743 12977
rect 25685 12968 25697 12971
rect 23808 12940 25697 12968
rect 23808 12928 23814 12940
rect 25685 12937 25697 12940
rect 25731 12968 25743 12971
rect 27062 12968 27068 12980
rect 25731 12940 27068 12968
rect 25731 12937 25743 12940
rect 25685 12931 25743 12937
rect 27062 12928 27068 12940
rect 27120 12928 27126 12980
rect 27154 12928 27160 12980
rect 27212 12968 27218 12980
rect 29362 12968 29368 12980
rect 27212 12940 29368 12968
rect 27212 12928 27218 12940
rect 29362 12928 29368 12940
rect 29420 12928 29426 12980
rect 32306 12968 32312 12980
rect 30576 12940 32312 12968
rect 13354 12900 13360 12912
rect 13096 12872 13360 12900
rect 12161 12835 12219 12841
rect 12161 12832 12173 12835
rect 11900 12804 12173 12832
rect 12161 12801 12173 12804
rect 12207 12801 12219 12835
rect 12161 12795 12219 12801
rect 12250 12792 12256 12844
rect 12308 12832 12314 12844
rect 12526 12832 12532 12844
rect 12308 12804 12532 12832
rect 12308 12792 12314 12804
rect 1210 12724 1216 12776
rect 1268 12764 1274 12776
rect 1581 12767 1639 12773
rect 1581 12764 1593 12767
rect 1268 12736 1593 12764
rect 1268 12724 1274 12736
rect 1581 12733 1593 12736
rect 1627 12733 1639 12767
rect 1581 12727 1639 12733
rect 1857 12767 1915 12773
rect 1857 12733 1869 12767
rect 1903 12764 1915 12767
rect 9490 12764 9496 12776
rect 1903 12736 9496 12764
rect 1903 12733 1915 12736
rect 1857 12727 1915 12733
rect 1596 12696 1624 12727
rect 9490 12724 9496 12736
rect 9548 12724 9554 12776
rect 10962 12724 10968 12776
rect 11020 12724 11026 12776
rect 12360 12773 12388 12804
rect 12526 12792 12532 12804
rect 12584 12792 12590 12844
rect 13096 12841 13124 12872
rect 13354 12860 13360 12872
rect 13412 12860 13418 12912
rect 14366 12860 14372 12912
rect 14424 12860 14430 12912
rect 16574 12860 16580 12912
rect 16632 12900 16638 12912
rect 17034 12900 17040 12912
rect 16632 12872 17040 12900
rect 16632 12860 16638 12872
rect 17034 12860 17040 12872
rect 17092 12900 17098 12912
rect 17129 12903 17187 12909
rect 17129 12900 17141 12903
rect 17092 12872 17141 12900
rect 17092 12860 17098 12872
rect 17129 12869 17141 12872
rect 17175 12869 17187 12903
rect 21174 12900 21180 12912
rect 17129 12863 17187 12869
rect 18432 12872 21180 12900
rect 13081 12835 13139 12841
rect 13081 12801 13093 12835
rect 13127 12801 13139 12835
rect 13081 12795 13139 12801
rect 12345 12767 12403 12773
rect 12345 12733 12357 12767
rect 12391 12764 12403 12767
rect 12391 12736 12425 12764
rect 12391 12733 12403 12736
rect 12345 12727 12403 12733
rect 12802 12724 12808 12776
rect 12860 12764 12866 12776
rect 13357 12767 13415 12773
rect 13357 12764 13369 12767
rect 12860 12736 13369 12764
rect 12860 12724 12866 12736
rect 13357 12733 13369 12736
rect 13403 12733 13415 12767
rect 14384 12764 14412 12860
rect 16022 12792 16028 12844
rect 16080 12792 16086 12844
rect 16850 12792 16856 12844
rect 16908 12792 16914 12844
rect 18230 12792 18236 12844
rect 18288 12792 18294 12844
rect 15197 12767 15255 12773
rect 15197 12764 15209 12767
rect 14384 12736 15209 12764
rect 13357 12727 13415 12733
rect 15197 12733 15209 12736
rect 15243 12764 15255 12767
rect 15286 12764 15292 12776
rect 15243 12736 15292 12764
rect 15243 12733 15255 12736
rect 15197 12727 15255 12733
rect 15286 12724 15292 12736
rect 15344 12724 15350 12776
rect 2774 12696 2780 12708
rect 1596 12668 2780 12696
rect 2774 12656 2780 12668
rect 2832 12656 2838 12708
rect 10042 12656 10048 12708
rect 10100 12696 10106 12708
rect 10137 12699 10195 12705
rect 10137 12696 10149 12699
rect 10100 12668 10149 12696
rect 10100 12656 10106 12668
rect 10137 12665 10149 12668
rect 10183 12696 10195 12699
rect 16040 12696 16068 12792
rect 16209 12767 16267 12773
rect 16209 12733 16221 12767
rect 16255 12733 16267 12767
rect 16209 12727 16267 12733
rect 10183 12668 13216 12696
rect 10183 12665 10195 12668
rect 10137 12659 10195 12665
rect 10410 12588 10416 12640
rect 10468 12588 10474 12640
rect 11422 12588 11428 12640
rect 11480 12628 11486 12640
rect 11701 12631 11759 12637
rect 11701 12628 11713 12631
rect 11480 12600 11713 12628
rect 11480 12588 11486 12600
rect 11701 12597 11713 12600
rect 11747 12597 11759 12631
rect 11701 12591 11759 12597
rect 12802 12588 12808 12640
rect 12860 12588 12866 12640
rect 13188 12628 13216 12668
rect 14384 12668 16068 12696
rect 16224 12696 16252 12727
rect 16482 12724 16488 12776
rect 16540 12764 16546 12776
rect 18432 12764 18460 12872
rect 21174 12860 21180 12872
rect 21232 12860 21238 12912
rect 21542 12860 21548 12912
rect 21600 12900 21606 12912
rect 23109 12903 23167 12909
rect 23109 12900 23121 12903
rect 21600 12872 23121 12900
rect 21600 12860 21606 12872
rect 23109 12869 23121 12872
rect 23155 12900 23167 12903
rect 23842 12900 23848 12912
rect 23155 12872 23848 12900
rect 23155 12869 23167 12872
rect 23109 12863 23167 12869
rect 23842 12860 23848 12872
rect 23900 12900 23906 12912
rect 24118 12900 24124 12912
rect 23900 12872 24124 12900
rect 23900 12860 23906 12872
rect 24118 12860 24124 12872
rect 24176 12860 24182 12912
rect 24210 12860 24216 12912
rect 24268 12860 24274 12912
rect 26786 12900 26792 12912
rect 25438 12872 26792 12900
rect 26786 12860 26792 12872
rect 26844 12860 26850 12912
rect 19518 12792 19524 12844
rect 19576 12792 19582 12844
rect 20993 12835 21051 12841
rect 20993 12801 21005 12835
rect 21039 12832 21051 12835
rect 21910 12832 21916 12844
rect 21039 12804 21916 12832
rect 21039 12801 21051 12804
rect 20993 12795 21051 12801
rect 21910 12792 21916 12804
rect 21968 12792 21974 12844
rect 22370 12792 22376 12844
rect 22428 12832 22434 12844
rect 22830 12832 22836 12844
rect 22428 12804 22836 12832
rect 22428 12792 22434 12804
rect 22830 12792 22836 12804
rect 22888 12832 22894 12844
rect 23201 12835 23259 12841
rect 23201 12832 23213 12835
rect 22888 12804 23213 12832
rect 22888 12792 22894 12804
rect 23201 12801 23213 12804
rect 23247 12801 23259 12835
rect 23201 12795 23259 12801
rect 23474 12792 23480 12844
rect 23532 12832 23538 12844
rect 27172 12841 27200 12928
rect 27433 12903 27491 12909
rect 27433 12869 27445 12903
rect 27479 12900 27491 12903
rect 27706 12900 27712 12912
rect 27479 12872 27712 12900
rect 27479 12869 27491 12872
rect 27433 12863 27491 12869
rect 27706 12860 27712 12872
rect 27764 12860 27770 12912
rect 28166 12860 28172 12912
rect 28224 12860 28230 12912
rect 28994 12860 29000 12912
rect 29052 12900 29058 12912
rect 29641 12903 29699 12909
rect 29641 12900 29653 12903
rect 29052 12872 29653 12900
rect 29052 12860 29058 12872
rect 29641 12869 29653 12872
rect 29687 12900 29699 12903
rect 29730 12900 29736 12912
rect 29687 12872 29736 12900
rect 29687 12869 29699 12872
rect 29641 12863 29699 12869
rect 29730 12860 29736 12872
rect 29788 12860 29794 12912
rect 30282 12860 30288 12912
rect 30340 12900 30346 12912
rect 30377 12903 30435 12909
rect 30377 12900 30389 12903
rect 30340 12872 30389 12900
rect 30340 12860 30346 12872
rect 30377 12869 30389 12872
rect 30423 12869 30435 12903
rect 30377 12863 30435 12869
rect 23937 12835 23995 12841
rect 23937 12832 23949 12835
rect 23532 12804 23949 12832
rect 23532 12792 23538 12804
rect 23937 12801 23949 12804
rect 23983 12801 23995 12835
rect 27157 12835 27215 12841
rect 23937 12795 23995 12801
rect 25976 12804 26280 12832
rect 25976 12776 26004 12804
rect 16540 12736 18460 12764
rect 16540 12724 16546 12736
rect 18598 12724 18604 12776
rect 18656 12764 18662 12776
rect 18874 12764 18880 12776
rect 18656 12736 18880 12764
rect 18656 12724 18662 12736
rect 18874 12724 18880 12736
rect 18932 12724 18938 12776
rect 19610 12724 19616 12776
rect 19668 12724 19674 12776
rect 19797 12767 19855 12773
rect 19797 12733 19809 12767
rect 19843 12764 19855 12767
rect 19843 12736 20760 12764
rect 19843 12733 19855 12736
rect 19797 12727 19855 12733
rect 16574 12696 16580 12708
rect 16224 12668 16580 12696
rect 14384 12628 14412 12668
rect 16574 12656 16580 12668
rect 16632 12656 16638 12708
rect 19150 12656 19156 12708
rect 19208 12656 19214 12708
rect 20622 12656 20628 12708
rect 20680 12656 20686 12708
rect 13188 12600 14412 12628
rect 15565 12631 15623 12637
rect 15565 12597 15577 12631
rect 15611 12628 15623 12631
rect 18414 12628 18420 12640
rect 15611 12600 18420 12628
rect 15611 12597 15623 12600
rect 15565 12591 15623 12597
rect 18414 12588 18420 12600
rect 18472 12588 18478 12640
rect 20254 12588 20260 12640
rect 20312 12588 20318 12640
rect 20732 12628 20760 12736
rect 21174 12724 21180 12776
rect 21232 12724 21238 12776
rect 22002 12724 22008 12776
rect 22060 12724 22066 12776
rect 22094 12724 22100 12776
rect 22152 12764 22158 12776
rect 23293 12767 23351 12773
rect 23293 12764 23305 12767
rect 22152 12736 23305 12764
rect 22152 12724 22158 12736
rect 23293 12733 23305 12736
rect 23339 12764 23351 12767
rect 25958 12764 25964 12776
rect 23339 12736 25964 12764
rect 23339 12733 23351 12736
rect 23293 12727 23351 12733
rect 25958 12724 25964 12736
rect 26016 12724 26022 12776
rect 26145 12767 26203 12773
rect 26145 12733 26157 12767
rect 26191 12733 26203 12767
rect 26252 12764 26280 12804
rect 27157 12801 27169 12835
rect 27203 12801 27215 12835
rect 27157 12795 27215 12801
rect 29270 12792 29276 12844
rect 29328 12832 29334 12844
rect 29546 12832 29552 12844
rect 29328 12804 29552 12832
rect 29328 12792 29334 12804
rect 29546 12792 29552 12804
rect 29604 12832 29610 12844
rect 30576 12832 30604 12940
rect 32306 12928 32312 12940
rect 32364 12928 32370 12980
rect 35710 12968 35716 12980
rect 32416 12940 35716 12968
rect 32416 12900 32444 12940
rect 35710 12928 35716 12940
rect 35768 12928 35774 12980
rect 35802 12928 35808 12980
rect 35860 12968 35866 12980
rect 36909 12971 36967 12977
rect 36909 12968 36921 12971
rect 35860 12940 36921 12968
rect 35860 12928 35866 12940
rect 36909 12937 36921 12940
rect 36955 12937 36967 12971
rect 41782 12968 41788 12980
rect 36909 12931 36967 12937
rect 37752 12940 41788 12968
rect 32324 12872 32444 12900
rect 29604 12804 30604 12832
rect 29604 12792 29610 12804
rect 31386 12792 31392 12844
rect 31444 12792 31450 12844
rect 32214 12792 32220 12844
rect 32272 12832 32278 12844
rect 32324 12841 32352 12872
rect 32490 12860 32496 12912
rect 32548 12900 32554 12912
rect 32585 12903 32643 12909
rect 32585 12900 32597 12903
rect 32548 12872 32597 12900
rect 32548 12860 32554 12872
rect 32585 12869 32597 12872
rect 32631 12869 32643 12903
rect 32585 12863 32643 12869
rect 34517 12903 34575 12909
rect 34517 12869 34529 12903
rect 34563 12900 34575 12903
rect 34606 12900 34612 12912
rect 34563 12872 34612 12900
rect 34563 12869 34575 12872
rect 34517 12863 34575 12869
rect 34606 12860 34612 12872
rect 34664 12860 34670 12912
rect 34790 12860 34796 12912
rect 34848 12900 34854 12912
rect 36357 12903 36415 12909
rect 36357 12900 36369 12903
rect 34848 12872 36369 12900
rect 34848 12860 34854 12872
rect 36357 12869 36369 12872
rect 36403 12869 36415 12903
rect 36357 12863 36415 12869
rect 36446 12860 36452 12912
rect 36504 12900 36510 12912
rect 37752 12909 37780 12940
rect 41782 12928 41788 12940
rect 41840 12928 41846 12980
rect 37737 12903 37795 12909
rect 36504 12872 37504 12900
rect 36504 12860 36510 12872
rect 32309 12835 32367 12841
rect 32309 12832 32321 12835
rect 32272 12804 32321 12832
rect 32272 12792 32278 12804
rect 32309 12801 32321 12804
rect 32355 12801 32367 12835
rect 32309 12795 32367 12801
rect 33686 12792 33692 12844
rect 33744 12792 33750 12844
rect 34422 12792 34428 12844
rect 34480 12832 34486 12844
rect 37476 12841 37504 12872
rect 37737 12869 37749 12903
rect 37783 12869 37795 12903
rect 37737 12863 37795 12869
rect 38470 12860 38476 12912
rect 38528 12860 38534 12912
rect 39850 12860 39856 12912
rect 39908 12900 39914 12912
rect 41141 12903 41199 12909
rect 41141 12900 41153 12903
rect 39908 12872 41153 12900
rect 39908 12860 39914 12872
rect 41141 12869 41153 12872
rect 41187 12900 41199 12903
rect 41877 12903 41935 12909
rect 41877 12900 41889 12903
rect 41187 12872 41889 12900
rect 41187 12869 41199 12872
rect 41141 12863 41199 12869
rect 41877 12869 41889 12872
rect 41923 12869 41935 12903
rect 41877 12863 41935 12869
rect 36265 12835 36323 12841
rect 36265 12832 36277 12835
rect 34480 12804 36277 12832
rect 34480 12792 34486 12804
rect 36265 12801 36277 12804
rect 36311 12801 36323 12835
rect 36265 12795 36323 12801
rect 37461 12835 37519 12841
rect 37461 12801 37473 12835
rect 37507 12801 37519 12835
rect 37461 12795 37519 12801
rect 39022 12792 39028 12844
rect 39080 12832 39086 12844
rect 39945 12835 40003 12841
rect 39945 12832 39957 12835
rect 39080 12804 39957 12832
rect 39080 12792 39086 12804
rect 39945 12801 39957 12804
rect 39991 12801 40003 12835
rect 39945 12795 40003 12801
rect 41598 12792 41604 12844
rect 41656 12792 41662 12844
rect 44174 12792 44180 12844
rect 44232 12832 44238 12844
rect 46201 12835 46259 12841
rect 46201 12832 46213 12835
rect 44232 12804 46213 12832
rect 44232 12792 44238 12804
rect 46201 12801 46213 12804
rect 46247 12801 46259 12835
rect 46201 12795 46259 12801
rect 47854 12792 47860 12844
rect 47912 12832 47918 12844
rect 47949 12835 48007 12841
rect 47949 12832 47961 12835
rect 47912 12804 47961 12832
rect 47912 12792 47918 12804
rect 47949 12801 47961 12804
rect 47995 12801 48007 12835
rect 47949 12795 48007 12801
rect 49142 12792 49148 12844
rect 49200 12792 49206 12844
rect 29181 12767 29239 12773
rect 29181 12764 29193 12767
rect 26252 12736 29193 12764
rect 26145 12727 26203 12733
rect 29181 12733 29193 12736
rect 29227 12733 29239 12767
rect 29181 12727 29239 12733
rect 31481 12767 31539 12773
rect 31481 12733 31493 12767
rect 31527 12764 31539 12767
rect 31570 12764 31576 12776
rect 31527 12736 31576 12764
rect 31527 12733 31539 12736
rect 31481 12727 31539 12733
rect 21266 12656 21272 12708
rect 21324 12696 21330 12708
rect 21324 12668 24072 12696
rect 21324 12656 21330 12668
rect 21818 12628 21824 12640
rect 20732 12600 21824 12628
rect 21818 12588 21824 12600
rect 21876 12588 21882 12640
rect 22462 12588 22468 12640
rect 22520 12628 22526 12640
rect 22830 12628 22836 12640
rect 22520 12600 22836 12628
rect 22520 12588 22526 12600
rect 22830 12588 22836 12600
rect 22888 12588 22894 12640
rect 24044 12628 24072 12668
rect 25222 12656 25228 12708
rect 25280 12696 25286 12708
rect 25406 12696 25412 12708
rect 25280 12668 25412 12696
rect 25280 12656 25286 12668
rect 25406 12656 25412 12668
rect 25464 12656 25470 12708
rect 26160 12628 26188 12727
rect 28534 12656 28540 12708
rect 28592 12696 28598 12708
rect 31496 12696 31524 12727
rect 31570 12724 31576 12736
rect 31628 12724 31634 12776
rect 31665 12767 31723 12773
rect 31665 12733 31677 12767
rect 31711 12733 31723 12767
rect 31665 12727 31723 12733
rect 28592 12668 31524 12696
rect 28592 12656 28598 12668
rect 24044 12600 26188 12628
rect 29454 12588 29460 12640
rect 29512 12628 29518 12640
rect 30098 12628 30104 12640
rect 29512 12600 30104 12628
rect 29512 12588 29518 12600
rect 30098 12588 30104 12600
rect 30156 12588 30162 12640
rect 31018 12588 31024 12640
rect 31076 12588 31082 12640
rect 31680 12628 31708 12727
rect 33318 12724 33324 12776
rect 33376 12764 33382 12776
rect 33704 12764 33732 12792
rect 33376 12736 33732 12764
rect 33376 12724 33382 12736
rect 34882 12724 34888 12776
rect 34940 12764 34946 12776
rect 35253 12767 35311 12773
rect 35253 12764 35265 12767
rect 34940 12736 35265 12764
rect 34940 12724 34946 12736
rect 35253 12733 35265 12736
rect 35299 12733 35311 12767
rect 35253 12727 35311 12733
rect 36446 12724 36452 12776
rect 36504 12724 36510 12776
rect 39485 12767 39543 12773
rect 39485 12764 39497 12767
rect 36556 12736 39497 12764
rect 33962 12656 33968 12708
rect 34020 12696 34026 12708
rect 34057 12699 34115 12705
rect 34057 12696 34069 12699
rect 34020 12668 34069 12696
rect 34020 12656 34026 12668
rect 34057 12665 34069 12668
rect 34103 12696 34115 12699
rect 34146 12696 34152 12708
rect 34103 12668 34152 12696
rect 34103 12665 34115 12668
rect 34057 12659 34115 12665
rect 34146 12656 34152 12668
rect 34204 12656 34210 12708
rect 35434 12656 35440 12708
rect 35492 12696 35498 12708
rect 36556 12696 36584 12736
rect 39485 12733 39497 12736
rect 39531 12733 39543 12767
rect 39485 12727 39543 12733
rect 35492 12668 36584 12696
rect 41325 12699 41383 12705
rect 35492 12656 35498 12668
rect 41325 12665 41337 12699
rect 41371 12696 41383 12699
rect 44174 12696 44180 12708
rect 41371 12668 44180 12696
rect 41371 12665 41383 12668
rect 41325 12659 41383 12665
rect 44174 12656 44180 12668
rect 44232 12656 44238 12708
rect 35158 12628 35164 12640
rect 31680 12600 35164 12628
rect 35158 12588 35164 12600
rect 35216 12588 35222 12640
rect 35897 12631 35955 12637
rect 35897 12597 35909 12631
rect 35943 12628 35955 12631
rect 38470 12628 38476 12640
rect 35943 12600 38476 12628
rect 35943 12597 35955 12600
rect 35897 12591 35955 12597
rect 38470 12588 38476 12600
rect 38528 12588 38534 12640
rect 38746 12588 38752 12640
rect 38804 12628 38810 12640
rect 40589 12631 40647 12637
rect 40589 12628 40601 12631
rect 38804 12600 40601 12628
rect 38804 12588 38810 12600
rect 40589 12597 40601 12600
rect 40635 12597 40647 12631
rect 40589 12591 40647 12597
rect 46017 12631 46075 12637
rect 46017 12597 46029 12631
rect 46063 12628 46075 12631
rect 47946 12628 47952 12640
rect 46063 12600 47952 12628
rect 46063 12597 46075 12600
rect 46017 12591 46075 12597
rect 47946 12588 47952 12600
rect 48004 12588 48010 12640
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 2774 12384 2780 12436
rect 2832 12384 2838 12436
rect 13078 12424 13084 12436
rect 9232 12396 13084 12424
rect 1857 12291 1915 12297
rect 1857 12257 1869 12291
rect 1903 12288 1915 12291
rect 5258 12288 5264 12300
rect 1903 12260 5264 12288
rect 1903 12257 1915 12260
rect 1857 12251 1915 12257
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 1302 12180 1308 12232
rect 1360 12220 1366 12232
rect 1581 12223 1639 12229
rect 1581 12220 1593 12223
rect 1360 12192 1593 12220
rect 1360 12180 1366 12192
rect 1581 12189 1593 12192
rect 1627 12189 1639 12223
rect 1581 12183 1639 12189
rect 1596 12152 1624 12183
rect 2869 12155 2927 12161
rect 2869 12152 2881 12155
rect 1596 12124 2881 12152
rect 2869 12121 2881 12124
rect 2915 12121 2927 12155
rect 2869 12115 2927 12121
rect 7558 12044 7564 12096
rect 7616 12084 7622 12096
rect 9232 12093 9260 12396
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 16761 12427 16819 12433
rect 16761 12424 16773 12427
rect 13464 12396 16773 12424
rect 10965 12291 11023 12297
rect 10965 12257 10977 12291
rect 11011 12288 11023 12291
rect 12250 12288 12256 12300
rect 11011 12260 12256 12288
rect 11011 12257 11023 12260
rect 10965 12251 11023 12257
rect 12250 12248 12256 12260
rect 12308 12248 12314 12300
rect 13464 12297 13492 12396
rect 16761 12393 16773 12396
rect 16807 12393 16819 12427
rect 16761 12387 16819 12393
rect 18598 12384 18604 12436
rect 18656 12424 18662 12436
rect 21634 12424 21640 12436
rect 18656 12396 21640 12424
rect 18656 12384 18662 12396
rect 21634 12384 21640 12396
rect 21692 12384 21698 12436
rect 22554 12384 22560 12436
rect 22612 12424 22618 12436
rect 23293 12427 23351 12433
rect 23293 12424 23305 12427
rect 22612 12396 23305 12424
rect 22612 12384 22618 12396
rect 23293 12393 23305 12396
rect 23339 12393 23351 12427
rect 25590 12424 25596 12436
rect 23293 12387 23351 12393
rect 23952 12396 25596 12424
rect 20901 12359 20959 12365
rect 20901 12325 20913 12359
rect 20947 12356 20959 12359
rect 23658 12356 23664 12368
rect 20947 12328 23664 12356
rect 20947 12325 20959 12328
rect 20901 12319 20959 12325
rect 23658 12316 23664 12328
rect 23716 12316 23722 12368
rect 13449 12291 13507 12297
rect 13449 12257 13461 12291
rect 13495 12257 13507 12291
rect 13449 12251 13507 12257
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 13906 12288 13912 12300
rect 13679 12260 13912 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 13906 12248 13912 12260
rect 13964 12248 13970 12300
rect 14645 12291 14703 12297
rect 14645 12257 14657 12291
rect 14691 12288 14703 12291
rect 16942 12288 16948 12300
rect 14691 12260 16948 12288
rect 14691 12257 14703 12260
rect 14645 12251 14703 12257
rect 16942 12248 16948 12260
rect 17000 12288 17006 12300
rect 17405 12291 17463 12297
rect 17405 12288 17417 12291
rect 17000 12260 17417 12288
rect 17000 12248 17006 12260
rect 17405 12257 17417 12260
rect 17451 12288 17463 12291
rect 17678 12288 17684 12300
rect 17451 12260 17684 12288
rect 17451 12257 17463 12260
rect 17405 12251 17463 12257
rect 17678 12248 17684 12260
rect 17736 12248 17742 12300
rect 19702 12248 19708 12300
rect 19760 12288 19766 12300
rect 20165 12291 20223 12297
rect 20165 12288 20177 12291
rect 19760 12260 20177 12288
rect 19760 12248 19766 12260
rect 20165 12257 20177 12260
rect 20211 12257 20223 12291
rect 20165 12251 20223 12257
rect 20806 12248 20812 12300
rect 20864 12288 20870 12300
rect 21453 12291 21511 12297
rect 21453 12288 21465 12291
rect 20864 12260 21465 12288
rect 20864 12248 20870 12260
rect 21453 12257 21465 12260
rect 21499 12257 21511 12291
rect 21453 12251 21511 12257
rect 22738 12248 22744 12300
rect 22796 12248 22802 12300
rect 23952 12297 23980 12396
rect 25590 12384 25596 12396
rect 25648 12384 25654 12436
rect 26050 12384 26056 12436
rect 26108 12424 26114 12436
rect 27614 12424 27620 12436
rect 26108 12396 27620 12424
rect 26108 12384 26114 12396
rect 27614 12384 27620 12396
rect 27672 12384 27678 12436
rect 29730 12384 29736 12436
rect 29788 12424 29794 12436
rect 31757 12427 31815 12433
rect 31757 12424 31769 12427
rect 29788 12396 31769 12424
rect 29788 12384 29794 12396
rect 31757 12393 31769 12396
rect 31803 12393 31815 12427
rect 33965 12427 34023 12433
rect 31757 12387 31815 12393
rect 32324 12396 33916 12424
rect 26326 12316 26332 12368
rect 26384 12356 26390 12368
rect 27338 12356 27344 12368
rect 26384 12328 27344 12356
rect 26384 12316 26390 12328
rect 27338 12316 27344 12328
rect 27396 12316 27402 12368
rect 31386 12316 31392 12368
rect 31444 12356 31450 12368
rect 32324 12356 32352 12396
rect 31444 12328 32352 12356
rect 33888 12356 33916 12396
rect 33965 12393 33977 12427
rect 34011 12424 34023 12427
rect 36446 12424 36452 12436
rect 34011 12396 36452 12424
rect 34011 12393 34023 12396
rect 33965 12387 34023 12393
rect 36446 12384 36452 12396
rect 36504 12384 36510 12436
rect 36630 12384 36636 12436
rect 36688 12384 36694 12436
rect 37090 12384 37096 12436
rect 37148 12384 37154 12436
rect 38194 12384 38200 12436
rect 38252 12424 38258 12436
rect 39209 12427 39267 12433
rect 39209 12424 39221 12427
rect 38252 12396 39221 12424
rect 38252 12384 38258 12396
rect 39209 12393 39221 12396
rect 39255 12424 39267 12427
rect 39393 12427 39451 12433
rect 39393 12424 39405 12427
rect 39255 12396 39405 12424
rect 39255 12393 39267 12396
rect 39209 12387 39267 12393
rect 39393 12393 39405 12396
rect 39439 12424 39451 12427
rect 39574 12424 39580 12436
rect 39439 12396 39580 12424
rect 39439 12393 39451 12396
rect 39393 12387 39451 12393
rect 39574 12384 39580 12396
rect 39632 12384 39638 12436
rect 34054 12356 34060 12368
rect 33888 12328 34060 12356
rect 31444 12316 31450 12328
rect 34054 12316 34060 12328
rect 34112 12356 34118 12368
rect 34241 12359 34299 12365
rect 34241 12356 34253 12359
rect 34112 12328 34253 12356
rect 34112 12316 34118 12328
rect 34241 12325 34253 12328
rect 34287 12325 34299 12359
rect 36648 12356 36676 12384
rect 37182 12356 37188 12368
rect 36648 12328 37188 12356
rect 34241 12319 34299 12325
rect 37182 12316 37188 12328
rect 37240 12316 37246 12368
rect 37274 12316 37280 12368
rect 37332 12356 37338 12368
rect 38930 12356 38936 12368
rect 37332 12328 38936 12356
rect 37332 12316 37338 12328
rect 38930 12316 38936 12328
rect 38988 12316 38994 12368
rect 41417 12359 41475 12365
rect 41417 12325 41429 12359
rect 41463 12356 41475 12359
rect 41463 12328 45554 12356
rect 41463 12325 41475 12328
rect 41417 12319 41475 12325
rect 23937 12291 23995 12297
rect 23308 12260 23704 12288
rect 9585 12223 9643 12229
rect 9585 12189 9597 12223
rect 9631 12220 9643 12223
rect 10689 12223 10747 12229
rect 9631 12192 10640 12220
rect 9631 12189 9643 12192
rect 9585 12183 9643 12189
rect 9217 12087 9275 12093
rect 9217 12084 9229 12087
rect 7616 12056 9229 12084
rect 7616 12044 7622 12056
rect 9217 12053 9229 12056
rect 9263 12053 9275 12087
rect 9217 12047 9275 12053
rect 10226 12044 10232 12096
rect 10284 12044 10290 12096
rect 10612 12084 10640 12192
rect 10689 12189 10701 12223
rect 10735 12189 10747 12223
rect 10689 12183 10747 12189
rect 10704 12152 10732 12183
rect 13722 12180 13728 12232
rect 13780 12220 13786 12232
rect 14274 12220 14280 12232
rect 13780 12192 14280 12220
rect 13780 12180 13786 12192
rect 14274 12180 14280 12192
rect 14332 12220 14338 12232
rect 14369 12223 14427 12229
rect 14369 12220 14381 12223
rect 14332 12192 14381 12220
rect 14332 12180 14338 12192
rect 14369 12189 14381 12192
rect 14415 12189 14427 12223
rect 14369 12183 14427 12189
rect 16482 12180 16488 12232
rect 16540 12220 16546 12232
rect 17957 12223 18015 12229
rect 17957 12220 17969 12223
rect 16540 12192 17969 12220
rect 16540 12180 16546 12192
rect 17957 12189 17969 12192
rect 18003 12220 18015 12223
rect 18322 12220 18328 12232
rect 18003 12192 18328 12220
rect 18003 12189 18015 12192
rect 17957 12183 18015 12189
rect 18322 12180 18328 12192
rect 18380 12220 18386 12232
rect 18380 12192 19472 12220
rect 18380 12180 18386 12192
rect 19444 12164 19472 12192
rect 21266 12180 21272 12232
rect 21324 12180 21330 12232
rect 23308 12220 23336 12260
rect 23676 12229 23704 12260
rect 23937 12257 23949 12291
rect 23983 12257 23995 12291
rect 23937 12251 23995 12257
rect 24857 12291 24915 12297
rect 24857 12257 24869 12291
rect 24903 12288 24915 12291
rect 26970 12288 26976 12300
rect 24903 12260 26976 12288
rect 24903 12257 24915 12260
rect 24857 12251 24915 12257
rect 26970 12248 26976 12260
rect 27028 12248 27034 12300
rect 27522 12248 27528 12300
rect 27580 12248 27586 12300
rect 28810 12248 28816 12300
rect 28868 12288 28874 12300
rect 28997 12291 29055 12297
rect 28997 12288 29009 12291
rect 28868 12260 29009 12288
rect 28868 12248 28874 12260
rect 28997 12257 29009 12260
rect 29043 12257 29055 12291
rect 28997 12251 29055 12257
rect 30006 12248 30012 12300
rect 30064 12248 30070 12300
rect 32214 12248 32220 12300
rect 32272 12248 32278 12300
rect 32493 12291 32551 12297
rect 32493 12257 32505 12291
rect 32539 12288 32551 12291
rect 34146 12288 34152 12300
rect 32539 12260 34152 12288
rect 32539 12257 32551 12260
rect 32493 12251 32551 12257
rect 34146 12248 34152 12260
rect 34204 12248 34210 12300
rect 34517 12291 34575 12297
rect 34517 12257 34529 12291
rect 34563 12288 34575 12291
rect 34698 12288 34704 12300
rect 34563 12260 34704 12288
rect 34563 12257 34575 12260
rect 34517 12251 34575 12257
rect 34698 12248 34704 12260
rect 34756 12248 34762 12300
rect 34885 12291 34943 12297
rect 34885 12257 34897 12291
rect 34931 12288 34943 12291
rect 35710 12288 35716 12300
rect 34931 12260 35716 12288
rect 34931 12257 34943 12260
rect 34885 12251 34943 12257
rect 35710 12248 35716 12260
rect 35768 12248 35774 12300
rect 36170 12248 36176 12300
rect 36228 12288 36234 12300
rect 36722 12288 36728 12300
rect 36228 12260 36728 12288
rect 36228 12248 36234 12260
rect 22112 12192 23336 12220
rect 23661 12223 23719 12229
rect 10870 12152 10876 12164
rect 10704 12124 10876 12152
rect 10870 12112 10876 12124
rect 10928 12112 10934 12164
rect 11606 12112 11612 12164
rect 11664 12112 11670 12164
rect 13078 12112 13084 12164
rect 13136 12152 13142 12164
rect 13357 12155 13415 12161
rect 13357 12152 13369 12155
rect 13136 12124 13369 12152
rect 13136 12112 13142 12124
rect 13357 12121 13369 12124
rect 13403 12152 13415 12155
rect 13446 12152 13452 12164
rect 13403 12124 13452 12152
rect 13403 12121 13415 12124
rect 13357 12115 13415 12121
rect 13446 12112 13452 12124
rect 13504 12112 13510 12164
rect 15286 12112 15292 12164
rect 15344 12112 15350 12164
rect 17494 12152 17500 12164
rect 16132 12124 17500 12152
rect 11054 12084 11060 12096
rect 10612 12056 11060 12084
rect 11054 12044 11060 12056
rect 11112 12084 11118 12096
rect 12250 12084 12256 12096
rect 11112 12056 12256 12084
rect 11112 12044 11118 12056
rect 12250 12044 12256 12056
rect 12308 12084 12314 12096
rect 12437 12087 12495 12093
rect 12437 12084 12449 12087
rect 12308 12056 12449 12084
rect 12308 12044 12314 12056
rect 12437 12053 12449 12056
rect 12483 12053 12495 12087
rect 12437 12047 12495 12053
rect 12989 12087 13047 12093
rect 12989 12053 13001 12087
rect 13035 12084 13047 12087
rect 15930 12084 15936 12096
rect 13035 12056 15936 12084
rect 13035 12053 13047 12056
rect 12989 12047 13047 12053
rect 15930 12044 15936 12056
rect 15988 12044 15994 12096
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 16132 12093 16160 12124
rect 17494 12112 17500 12124
rect 17552 12112 17558 12164
rect 17862 12112 17868 12164
rect 17920 12152 17926 12164
rect 18693 12155 18751 12161
rect 18693 12152 18705 12155
rect 17920 12124 18705 12152
rect 17920 12112 17926 12124
rect 18693 12121 18705 12124
rect 18739 12121 18751 12155
rect 18693 12115 18751 12121
rect 19426 12112 19432 12164
rect 19484 12112 19490 12164
rect 21174 12112 21180 12164
rect 21232 12152 21238 12164
rect 21634 12152 21640 12164
rect 21232 12124 21640 12152
rect 21232 12112 21238 12124
rect 21634 12112 21640 12124
rect 21692 12112 21698 12164
rect 16117 12087 16175 12093
rect 16117 12084 16129 12087
rect 16080 12056 16129 12084
rect 16080 12044 16086 12056
rect 16117 12053 16129 12056
rect 16163 12053 16175 12087
rect 16117 12047 16175 12053
rect 17126 12044 17132 12096
rect 17184 12044 17190 12096
rect 17218 12044 17224 12096
rect 17276 12044 17282 12096
rect 21266 12044 21272 12096
rect 21324 12084 21330 12096
rect 21361 12087 21419 12093
rect 21361 12084 21373 12087
rect 21324 12056 21373 12084
rect 21324 12044 21330 12056
rect 21361 12053 21373 12056
rect 21407 12084 21419 12087
rect 21450 12084 21456 12096
rect 21407 12056 21456 12084
rect 21407 12053 21419 12056
rect 21361 12047 21419 12053
rect 21450 12044 21456 12056
rect 21508 12044 21514 12096
rect 22112 12093 22140 12192
rect 23661 12189 23673 12223
rect 23707 12189 23719 12223
rect 23661 12183 23719 12189
rect 24486 12180 24492 12232
rect 24544 12220 24550 12232
rect 24581 12223 24639 12229
rect 24581 12220 24593 12223
rect 24544 12192 24593 12220
rect 24544 12180 24550 12192
rect 24581 12189 24593 12192
rect 24627 12189 24639 12223
rect 24581 12183 24639 12189
rect 25958 12180 25964 12232
rect 26016 12220 26022 12232
rect 26697 12223 26755 12229
rect 26697 12220 26709 12223
rect 26016 12192 26709 12220
rect 26016 12180 26022 12192
rect 26697 12189 26709 12192
rect 26743 12220 26755 12223
rect 26786 12220 26792 12232
rect 26743 12192 26792 12220
rect 26743 12189 26755 12192
rect 26697 12183 26755 12189
rect 26786 12180 26792 12192
rect 26844 12180 26850 12232
rect 27154 12180 27160 12232
rect 27212 12220 27218 12232
rect 28905 12223 28963 12229
rect 28905 12220 28917 12223
rect 27212 12192 28917 12220
rect 27212 12180 27218 12192
rect 28905 12189 28917 12192
rect 28951 12189 28963 12223
rect 28905 12183 28963 12189
rect 29086 12180 29092 12232
rect 29144 12220 29150 12232
rect 29362 12220 29368 12232
rect 29144 12192 29368 12220
rect 29144 12180 29150 12192
rect 29362 12180 29368 12192
rect 29420 12220 29426 12232
rect 29733 12223 29791 12229
rect 29733 12220 29745 12223
rect 29420 12192 29745 12220
rect 29420 12180 29426 12192
rect 29733 12189 29745 12192
rect 29779 12189 29791 12223
rect 29733 12183 29791 12189
rect 34238 12180 34244 12232
rect 34296 12220 34302 12232
rect 34296 12192 34652 12220
rect 36280 12206 36308 12260
rect 36722 12248 36728 12260
rect 36780 12248 36786 12300
rect 37550 12248 37556 12300
rect 37608 12248 37614 12300
rect 37734 12248 37740 12300
rect 37792 12248 37798 12300
rect 34296 12180 34302 12192
rect 30282 12152 30288 12164
rect 22572 12124 24808 12152
rect 22572 12096 22600 12124
rect 22097 12087 22155 12093
rect 22097 12053 22109 12087
rect 22143 12053 22155 12087
rect 22097 12047 22155 12053
rect 22462 12044 22468 12096
rect 22520 12044 22526 12096
rect 22554 12044 22560 12096
rect 22612 12044 22618 12096
rect 23753 12087 23811 12093
rect 23753 12053 23765 12087
rect 23799 12084 23811 12087
rect 24670 12084 24676 12096
rect 23799 12056 24676 12084
rect 23799 12053 23811 12056
rect 23753 12047 23811 12053
rect 24670 12044 24676 12056
rect 24728 12044 24734 12096
rect 24780 12084 24808 12124
rect 26988 12124 30288 12152
rect 26234 12084 26240 12096
rect 24780 12056 26240 12084
rect 26234 12044 26240 12056
rect 26292 12044 26298 12096
rect 26988 12093 27016 12124
rect 30282 12112 30288 12124
rect 30340 12112 30346 12164
rect 30466 12112 30472 12164
rect 30524 12112 30530 12164
rect 33226 12112 33232 12164
rect 33284 12112 33290 12164
rect 34624 12152 34652 12192
rect 37458 12180 37464 12232
rect 37516 12180 37522 12232
rect 38289 12223 38347 12229
rect 38289 12189 38301 12223
rect 38335 12189 38347 12223
rect 38289 12183 38347 12189
rect 35161 12155 35219 12161
rect 35161 12152 35173 12155
rect 34164 12124 34560 12152
rect 34624 12124 35173 12152
rect 26973 12087 27031 12093
rect 26973 12053 26985 12087
rect 27019 12053 27031 12087
rect 26973 12047 27031 12053
rect 27338 12044 27344 12096
rect 27396 12044 27402 12096
rect 27433 12087 27491 12093
rect 27433 12053 27445 12087
rect 27479 12084 27491 12087
rect 27614 12084 27620 12096
rect 27479 12056 27620 12084
rect 27479 12053 27491 12056
rect 27433 12047 27491 12053
rect 27614 12044 27620 12056
rect 27672 12084 27678 12096
rect 28077 12087 28135 12093
rect 28077 12084 28089 12087
rect 27672 12056 28089 12084
rect 27672 12044 27678 12056
rect 28077 12053 28089 12056
rect 28123 12084 28135 12087
rect 28350 12084 28356 12096
rect 28123 12056 28356 12084
rect 28123 12053 28135 12056
rect 28077 12047 28135 12053
rect 28350 12044 28356 12056
rect 28408 12044 28414 12096
rect 28442 12044 28448 12096
rect 28500 12044 28506 12096
rect 28813 12087 28871 12093
rect 28813 12053 28825 12087
rect 28859 12084 28871 12087
rect 30374 12084 30380 12096
rect 28859 12056 30380 12084
rect 28859 12053 28871 12056
rect 28813 12047 28871 12053
rect 30374 12044 30380 12056
rect 30432 12044 30438 12096
rect 31481 12087 31539 12093
rect 31481 12053 31493 12087
rect 31527 12084 31539 12087
rect 34164 12084 34192 12124
rect 34532 12096 34560 12124
rect 35161 12121 35173 12124
rect 35207 12152 35219 12155
rect 35434 12152 35440 12164
rect 35207 12124 35440 12152
rect 35207 12121 35219 12124
rect 35161 12115 35219 12121
rect 35434 12112 35440 12124
rect 35492 12112 35498 12164
rect 31527 12056 34192 12084
rect 31527 12053 31539 12056
rect 31481 12047 31539 12053
rect 34514 12044 34520 12096
rect 34572 12084 34578 12096
rect 38304 12084 38332 12183
rect 38470 12180 38476 12232
rect 38528 12220 38534 12232
rect 40957 12223 41015 12229
rect 40957 12220 40969 12223
rect 38528 12192 40969 12220
rect 38528 12180 38534 12192
rect 40957 12189 40969 12192
rect 41003 12189 41015 12223
rect 40957 12183 41015 12189
rect 41598 12180 41604 12232
rect 41656 12180 41662 12232
rect 45526 12220 45554 12328
rect 49142 12248 49148 12300
rect 49200 12248 49206 12300
rect 46109 12223 46167 12229
rect 46109 12220 46121 12223
rect 45526 12192 46121 12220
rect 46109 12189 46121 12192
rect 46155 12189 46167 12223
rect 46109 12183 46167 12189
rect 47946 12180 47952 12232
rect 48004 12180 48010 12232
rect 40126 12112 40132 12164
rect 40184 12112 40190 12164
rect 40313 12155 40371 12161
rect 40313 12121 40325 12155
rect 40359 12152 40371 12155
rect 47210 12152 47216 12164
rect 40359 12124 47216 12152
rect 40359 12121 40371 12124
rect 40313 12115 40371 12121
rect 47210 12112 47216 12124
rect 47268 12112 47274 12164
rect 34572 12056 38332 12084
rect 34572 12044 34578 12056
rect 38930 12044 38936 12096
rect 38988 12044 38994 12096
rect 40770 12044 40776 12096
rect 40828 12044 40834 12096
rect 45922 12044 45928 12096
rect 45980 12044 45986 12096
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 2317 11883 2375 11889
rect 2317 11849 2329 11883
rect 2363 11880 2375 11883
rect 4338 11880 4344 11892
rect 2363 11852 4344 11880
rect 2363 11849 2375 11852
rect 2317 11843 2375 11849
rect 4338 11840 4344 11852
rect 4396 11840 4402 11892
rect 9858 11840 9864 11892
rect 9916 11880 9922 11892
rect 9953 11883 10011 11889
rect 9953 11880 9965 11883
rect 9916 11852 9965 11880
rect 9916 11840 9922 11852
rect 9953 11849 9965 11852
rect 9999 11880 10011 11883
rect 10137 11883 10195 11889
rect 10137 11880 10149 11883
rect 9999 11852 10149 11880
rect 9999 11849 10011 11852
rect 9953 11843 10011 11849
rect 10137 11849 10149 11852
rect 10183 11849 10195 11883
rect 10137 11843 10195 11849
rect 10870 11840 10876 11892
rect 10928 11880 10934 11892
rect 13354 11880 13360 11892
rect 10928 11852 13360 11880
rect 10928 11840 10934 11852
rect 10594 11812 10600 11824
rect 6886 11784 10600 11812
rect 1210 11704 1216 11756
rect 1268 11744 1274 11756
rect 1581 11747 1639 11753
rect 1581 11744 1593 11747
rect 1268 11716 1593 11744
rect 1268 11704 1274 11716
rect 1581 11713 1593 11716
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11713 2559 11747
rect 2501 11707 2559 11713
rect 1302 11636 1308 11688
rect 1360 11676 1366 11688
rect 2516 11676 2544 11707
rect 2777 11679 2835 11685
rect 2777 11676 2789 11679
rect 1360 11648 2789 11676
rect 1360 11636 1366 11648
rect 2777 11645 2789 11648
rect 2823 11645 2835 11679
rect 2777 11639 2835 11645
rect 1765 11611 1823 11617
rect 1765 11577 1777 11611
rect 1811 11608 1823 11611
rect 6886 11608 6914 11784
rect 10594 11772 10600 11784
rect 10652 11772 10658 11824
rect 12360 11753 12388 11852
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 15470 11840 15476 11892
rect 15528 11880 15534 11892
rect 15565 11883 15623 11889
rect 15565 11880 15577 11883
rect 15528 11852 15577 11880
rect 15528 11840 15534 11852
rect 15565 11849 15577 11852
rect 15611 11849 15623 11883
rect 15565 11843 15623 11849
rect 16482 11840 16488 11892
rect 16540 11840 16546 11892
rect 16574 11840 16580 11892
rect 16632 11880 16638 11892
rect 19061 11883 19119 11889
rect 19061 11880 19073 11883
rect 16632 11852 19073 11880
rect 16632 11840 16638 11852
rect 19061 11849 19073 11852
rect 19107 11880 19119 11883
rect 19889 11883 19947 11889
rect 19889 11880 19901 11883
rect 19107 11852 19901 11880
rect 19107 11849 19119 11852
rect 19061 11843 19119 11849
rect 19889 11849 19901 11852
rect 19935 11880 19947 11883
rect 20070 11880 20076 11892
rect 19935 11852 20076 11880
rect 19935 11849 19947 11852
rect 19889 11843 19947 11849
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 20530 11840 20536 11892
rect 20588 11880 20594 11892
rect 20717 11883 20775 11889
rect 20717 11880 20729 11883
rect 20588 11852 20729 11880
rect 20588 11840 20594 11852
rect 20717 11849 20729 11852
rect 20763 11849 20775 11883
rect 20717 11843 20775 11849
rect 21085 11883 21143 11889
rect 21085 11849 21097 11883
rect 21131 11880 21143 11883
rect 22002 11880 22008 11892
rect 21131 11852 22008 11880
rect 21131 11849 21143 11852
rect 21085 11843 21143 11849
rect 22002 11840 22008 11852
rect 22060 11840 22066 11892
rect 22281 11883 22339 11889
rect 22281 11849 22293 11883
rect 22327 11880 22339 11883
rect 22370 11880 22376 11892
rect 22327 11852 22376 11880
rect 22327 11849 22339 11852
rect 22281 11843 22339 11849
rect 22370 11840 22376 11852
rect 22428 11840 22434 11892
rect 25590 11840 25596 11892
rect 25648 11880 25654 11892
rect 25685 11883 25743 11889
rect 25685 11880 25697 11883
rect 25648 11852 25697 11880
rect 25648 11840 25654 11852
rect 25685 11849 25697 11852
rect 25731 11849 25743 11883
rect 25685 11843 25743 11849
rect 25958 11840 25964 11892
rect 26016 11840 26022 11892
rect 26421 11883 26479 11889
rect 26421 11849 26433 11883
rect 26467 11880 26479 11883
rect 27338 11880 27344 11892
rect 26467 11852 27344 11880
rect 26467 11849 26479 11852
rect 26421 11843 26479 11849
rect 27338 11840 27344 11852
rect 27396 11840 27402 11892
rect 28442 11840 28448 11892
rect 28500 11880 28506 11892
rect 28500 11852 30144 11880
rect 28500 11840 28506 11852
rect 14182 11812 14188 11824
rect 13846 11784 14188 11812
rect 14182 11772 14188 11784
rect 14240 11772 14246 11824
rect 14274 11772 14280 11824
rect 14332 11812 14338 11824
rect 18969 11815 19027 11821
rect 14332 11784 16436 11812
rect 14332 11772 14338 11784
rect 10505 11747 10563 11753
rect 10505 11713 10517 11747
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 12345 11747 12403 11753
rect 12345 11713 12357 11747
rect 12391 11713 12403 11747
rect 12345 11707 12403 11713
rect 1811 11580 6914 11608
rect 10520 11608 10548 11707
rect 13998 11704 14004 11756
rect 14056 11744 14062 11756
rect 14369 11747 14427 11753
rect 14369 11744 14381 11747
rect 14056 11716 14381 11744
rect 14056 11704 14062 11716
rect 14369 11713 14381 11716
rect 14415 11744 14427 11747
rect 14734 11744 14740 11756
rect 14415 11716 14740 11744
rect 14415 11713 14427 11716
rect 14369 11707 14427 11713
rect 14734 11704 14740 11716
rect 14792 11704 14798 11756
rect 15470 11704 15476 11756
rect 15528 11704 15534 11756
rect 16408 11744 16436 11784
rect 18969 11781 18981 11815
rect 19015 11812 19027 11815
rect 20806 11812 20812 11824
rect 19015 11784 20812 11812
rect 19015 11781 19027 11784
rect 18969 11775 19027 11781
rect 20806 11772 20812 11784
rect 20864 11812 20870 11824
rect 22094 11812 22100 11824
rect 20864 11784 22100 11812
rect 20864 11772 20870 11784
rect 22094 11772 22100 11784
rect 22152 11772 22158 11824
rect 23382 11772 23388 11824
rect 23440 11812 23446 11824
rect 24486 11812 24492 11824
rect 23440 11784 24492 11812
rect 23440 11772 23446 11784
rect 16850 11744 16856 11756
rect 15580 11716 16344 11744
rect 16408 11716 16856 11744
rect 11701 11679 11759 11685
rect 11701 11645 11713 11679
rect 11747 11676 11759 11679
rect 12158 11676 12164 11688
rect 11747 11648 12164 11676
rect 11747 11645 11759 11648
rect 11701 11639 11759 11645
rect 12158 11636 12164 11648
rect 12216 11636 12222 11688
rect 12618 11636 12624 11688
rect 12676 11636 12682 11688
rect 15580 11676 15608 11716
rect 14660 11648 15608 11676
rect 15657 11679 15715 11685
rect 10520 11580 12434 11608
rect 1811 11577 1823 11580
rect 1765 11571 1823 11577
rect 11149 11543 11207 11549
rect 11149 11509 11161 11543
rect 11195 11540 11207 11543
rect 12066 11540 12072 11552
rect 11195 11512 12072 11540
rect 11195 11509 11207 11512
rect 11149 11503 11207 11509
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 12406 11540 12434 11580
rect 13630 11540 13636 11552
rect 12406 11512 13636 11540
rect 13630 11500 13636 11512
rect 13688 11540 13694 11552
rect 14660 11540 14688 11648
rect 15657 11645 15669 11679
rect 15703 11645 15715 11679
rect 15657 11639 15715 11645
rect 14734 11568 14740 11620
rect 14792 11608 14798 11620
rect 15672 11608 15700 11639
rect 14792 11580 15700 11608
rect 14792 11568 14798 11580
rect 13688 11512 14688 11540
rect 13688 11500 13694 11512
rect 14826 11500 14832 11552
rect 14884 11500 14890 11552
rect 15010 11500 15016 11552
rect 15068 11540 15074 11552
rect 15105 11543 15163 11549
rect 15105 11540 15117 11543
rect 15068 11512 15117 11540
rect 15068 11500 15074 11512
rect 15105 11509 15117 11512
rect 15151 11509 15163 11543
rect 15105 11503 15163 11509
rect 15470 11500 15476 11552
rect 15528 11540 15534 11552
rect 16206 11540 16212 11552
rect 15528 11512 16212 11540
rect 15528 11500 15534 11512
rect 16206 11500 16212 11512
rect 16264 11500 16270 11552
rect 16316 11540 16344 11716
rect 16850 11704 16856 11716
rect 16908 11704 16914 11756
rect 18230 11704 18236 11756
rect 18288 11704 18294 11756
rect 19797 11747 19855 11753
rect 19797 11713 19809 11747
rect 19843 11713 19855 11747
rect 19797 11707 19855 11713
rect 21913 11747 21971 11753
rect 21913 11713 21925 11747
rect 21959 11744 21971 11747
rect 22557 11747 22615 11753
rect 22557 11744 22569 11747
rect 21959 11716 22569 11744
rect 21959 11713 21971 11716
rect 21913 11707 21971 11713
rect 22557 11713 22569 11716
rect 22603 11744 22615 11747
rect 22646 11744 22652 11756
rect 22603 11716 22652 11744
rect 22603 11713 22615 11716
rect 22557 11707 22615 11713
rect 17129 11679 17187 11685
rect 17129 11645 17141 11679
rect 17175 11676 17187 11679
rect 19242 11676 19248 11688
rect 17175 11648 19248 11676
rect 17175 11645 17187 11648
rect 17129 11639 17187 11645
rect 19242 11636 19248 11648
rect 19300 11636 19306 11688
rect 19812 11676 19840 11707
rect 22646 11704 22652 11716
rect 22704 11704 22710 11756
rect 23952 11753 23980 11784
rect 24486 11772 24492 11784
rect 24544 11772 24550 11824
rect 25976 11812 26004 11840
rect 29086 11812 29092 11824
rect 25438 11784 26004 11812
rect 28552 11784 29092 11812
rect 23937 11747 23995 11753
rect 23937 11713 23949 11747
rect 23983 11713 23995 11747
rect 23937 11707 23995 11713
rect 27338 11704 27344 11756
rect 27396 11744 27402 11756
rect 27525 11747 27583 11753
rect 27525 11744 27537 11747
rect 27396 11716 27537 11744
rect 27396 11704 27402 11716
rect 27525 11713 27537 11716
rect 27571 11744 27583 11747
rect 28169 11747 28227 11753
rect 28169 11744 28181 11747
rect 27571 11716 28181 11744
rect 27571 11713 27583 11716
rect 27525 11707 27583 11713
rect 28169 11713 28181 11716
rect 28215 11744 28227 11747
rect 28442 11744 28448 11756
rect 28215 11716 28448 11744
rect 28215 11713 28227 11716
rect 28169 11707 28227 11713
rect 28442 11704 28448 11716
rect 28500 11704 28506 11756
rect 28552 11753 28580 11784
rect 29086 11772 29092 11784
rect 29144 11772 29150 11824
rect 29454 11772 29460 11824
rect 29512 11772 29518 11824
rect 30116 11812 30144 11852
rect 30282 11840 30288 11892
rect 30340 11880 30346 11892
rect 31205 11883 31263 11889
rect 31205 11880 31217 11883
rect 30340 11852 31217 11880
rect 30340 11840 30346 11852
rect 31205 11849 31217 11852
rect 31251 11849 31263 11883
rect 31205 11843 31263 11849
rect 31294 11840 31300 11892
rect 31352 11840 31358 11892
rect 32309 11883 32367 11889
rect 32309 11849 32321 11883
rect 32355 11880 32367 11883
rect 32674 11880 32680 11892
rect 32355 11852 32680 11880
rect 32355 11849 32367 11852
rect 32309 11843 32367 11849
rect 32674 11840 32680 11852
rect 32732 11840 32738 11892
rect 37274 11880 37280 11892
rect 33980 11852 37280 11880
rect 33873 11815 33931 11821
rect 33873 11812 33885 11815
rect 30116 11784 33885 11812
rect 33873 11781 33885 11784
rect 33919 11781 33931 11815
rect 33873 11775 33931 11781
rect 28537 11747 28595 11753
rect 28537 11713 28549 11747
rect 28583 11713 28595 11747
rect 28537 11707 28595 11713
rect 30098 11704 30104 11756
rect 30156 11744 30162 11756
rect 32677 11747 32735 11753
rect 32677 11744 32689 11747
rect 30156 11716 32689 11744
rect 30156 11704 30162 11716
rect 32677 11713 32689 11716
rect 32723 11713 32735 11747
rect 33980 11744 34008 11852
rect 37274 11840 37280 11852
rect 37332 11840 37338 11892
rect 37829 11883 37887 11889
rect 37829 11849 37841 11883
rect 37875 11880 37887 11883
rect 38657 11883 38715 11889
rect 38657 11880 38669 11883
rect 37875 11852 38669 11880
rect 37875 11849 37887 11852
rect 37829 11843 37887 11849
rect 38657 11849 38669 11852
rect 38703 11849 38715 11883
rect 38657 11843 38715 11849
rect 34609 11815 34667 11821
rect 34609 11781 34621 11815
rect 34655 11812 34667 11815
rect 34790 11812 34796 11824
rect 34655 11784 34796 11812
rect 34655 11781 34667 11784
rect 34609 11775 34667 11781
rect 34790 11772 34796 11784
rect 34848 11772 34854 11824
rect 36722 11812 36728 11824
rect 36662 11784 36728 11812
rect 36722 11772 36728 11784
rect 36780 11772 36786 11824
rect 37366 11772 37372 11824
rect 37424 11812 37430 11824
rect 37921 11815 37979 11821
rect 37921 11812 37933 11815
rect 37424 11784 37933 11812
rect 37424 11772 37430 11784
rect 37921 11781 37933 11784
rect 37967 11781 37979 11815
rect 37921 11775 37979 11781
rect 38120 11784 39896 11812
rect 32677 11707 32735 11713
rect 32876 11716 34008 11744
rect 19886 11676 19892 11688
rect 19812 11648 19892 11676
rect 19886 11636 19892 11648
rect 19944 11636 19950 11688
rect 19981 11679 20039 11685
rect 19981 11645 19993 11679
rect 20027 11645 20039 11679
rect 19981 11639 20039 11645
rect 18322 11568 18328 11620
rect 18380 11608 18386 11620
rect 19996 11608 20024 11639
rect 20162 11636 20168 11688
rect 20220 11676 20226 11688
rect 21177 11679 21235 11685
rect 21177 11676 21189 11679
rect 20220 11648 21189 11676
rect 20220 11636 20226 11648
rect 21177 11645 21189 11648
rect 21223 11676 21235 11679
rect 21266 11676 21272 11688
rect 21223 11648 21272 11676
rect 21223 11645 21235 11648
rect 21177 11639 21235 11645
rect 21266 11636 21272 11648
rect 21324 11636 21330 11688
rect 21358 11636 21364 11688
rect 21416 11636 21422 11688
rect 22066 11648 22600 11676
rect 18380 11580 20024 11608
rect 18380 11568 18386 11580
rect 20070 11568 20076 11620
rect 20128 11608 20134 11620
rect 22066 11608 22094 11648
rect 22572 11620 22600 11648
rect 22738 11636 22744 11688
rect 22796 11676 22802 11688
rect 24213 11679 24271 11685
rect 24213 11676 24225 11679
rect 22796 11648 24225 11676
rect 22796 11636 22802 11648
rect 24213 11645 24225 11648
rect 24259 11676 24271 11679
rect 26326 11676 26332 11688
rect 24259 11648 26332 11676
rect 24259 11645 24271 11648
rect 24213 11639 24271 11645
rect 26326 11636 26332 11648
rect 26384 11636 26390 11688
rect 27430 11636 27436 11688
rect 27488 11676 27494 11688
rect 27617 11679 27675 11685
rect 27617 11676 27629 11679
rect 27488 11648 27629 11676
rect 27488 11636 27494 11648
rect 27617 11645 27629 11648
rect 27663 11645 27675 11679
rect 27617 11639 27675 11645
rect 27801 11679 27859 11685
rect 27801 11645 27813 11679
rect 27847 11676 27859 11679
rect 27847 11648 28672 11676
rect 27847 11645 27859 11648
rect 27801 11639 27859 11645
rect 20128 11580 22094 11608
rect 20128 11568 20134 11580
rect 22554 11568 22560 11620
rect 22612 11568 22618 11620
rect 27154 11568 27160 11620
rect 27212 11568 27218 11620
rect 18601 11543 18659 11549
rect 18601 11540 18613 11543
rect 16316 11512 18613 11540
rect 18601 11509 18613 11512
rect 18647 11509 18659 11543
rect 18601 11503 18659 11509
rect 19334 11500 19340 11552
rect 19392 11540 19398 11552
rect 19429 11543 19487 11549
rect 19429 11540 19441 11543
rect 19392 11512 19441 11540
rect 19392 11500 19398 11512
rect 19429 11509 19441 11512
rect 19475 11509 19487 11543
rect 19429 11503 19487 11509
rect 19702 11500 19708 11552
rect 19760 11540 19766 11552
rect 22094 11540 22100 11552
rect 19760 11512 22100 11540
rect 19760 11500 19766 11512
rect 22094 11500 22100 11512
rect 22152 11500 22158 11552
rect 28644 11540 28672 11648
rect 28810 11636 28816 11688
rect 28868 11636 28874 11688
rect 29362 11636 29368 11688
rect 29420 11676 29426 11688
rect 31389 11679 31447 11685
rect 31389 11676 31401 11679
rect 29420 11648 31401 11676
rect 29420 11636 29426 11648
rect 31389 11645 31401 11648
rect 31435 11645 31447 11679
rect 31389 11639 31447 11645
rect 31938 11636 31944 11688
rect 31996 11676 32002 11688
rect 32306 11676 32312 11688
rect 31996 11648 32312 11676
rect 31996 11636 32002 11648
rect 32306 11636 32312 11648
rect 32364 11636 32370 11688
rect 32766 11636 32772 11688
rect 32824 11636 32830 11688
rect 32876 11685 32904 11716
rect 32861 11679 32919 11685
rect 32861 11645 32873 11679
rect 32907 11645 32919 11679
rect 33965 11679 34023 11685
rect 33965 11676 33977 11679
rect 32861 11639 32919 11645
rect 32968 11648 33977 11676
rect 29822 11568 29828 11620
rect 29880 11608 29886 11620
rect 30285 11611 30343 11617
rect 30285 11608 30297 11611
rect 29880 11580 30297 11608
rect 29880 11568 29886 11580
rect 30285 11577 30297 11580
rect 30331 11577 30343 11611
rect 30285 11571 30343 11577
rect 30742 11568 30748 11620
rect 30800 11608 30806 11620
rect 32968 11608 32996 11648
rect 33965 11645 33977 11648
rect 34011 11645 34023 11679
rect 33965 11639 34023 11645
rect 34149 11679 34207 11685
rect 34149 11645 34161 11679
rect 34195 11676 34207 11679
rect 34514 11676 34520 11688
rect 34195 11648 34520 11676
rect 34195 11645 34207 11648
rect 34149 11639 34207 11645
rect 34514 11636 34520 11648
rect 34572 11636 34578 11688
rect 34882 11636 34888 11688
rect 34940 11676 34946 11688
rect 38120 11685 38148 11784
rect 38378 11704 38384 11756
rect 38436 11744 38442 11756
rect 39868 11753 39896 11784
rect 40770 11772 40776 11824
rect 40828 11812 40834 11824
rect 45097 11815 45155 11821
rect 45097 11812 45109 11815
rect 40828 11784 45109 11812
rect 40828 11772 40834 11784
rect 45097 11781 45109 11784
rect 45143 11781 45155 11815
rect 45097 11775 45155 11781
rect 49142 11772 49148 11824
rect 49200 11772 49206 11824
rect 39025 11747 39083 11753
rect 39025 11744 39037 11747
rect 38436 11716 39037 11744
rect 38436 11704 38442 11716
rect 39025 11713 39037 11716
rect 39071 11713 39083 11747
rect 39025 11707 39083 11713
rect 39853 11747 39911 11753
rect 39853 11713 39865 11747
rect 39899 11713 39911 11747
rect 39853 11707 39911 11713
rect 45922 11704 45928 11756
rect 45980 11744 45986 11756
rect 47949 11747 48007 11753
rect 47949 11744 47961 11747
rect 45980 11716 47961 11744
rect 45980 11704 45986 11716
rect 47949 11713 47961 11716
rect 47995 11713 48007 11747
rect 47949 11707 48007 11713
rect 35161 11679 35219 11685
rect 35161 11676 35173 11679
rect 34940 11648 35173 11676
rect 34940 11636 34946 11648
rect 35161 11645 35173 11648
rect 35207 11676 35219 11679
rect 35437 11679 35495 11685
rect 35207 11648 35296 11676
rect 35207 11645 35219 11648
rect 35161 11639 35219 11645
rect 30800 11580 32996 11608
rect 33505 11611 33563 11617
rect 30800 11568 30806 11580
rect 33505 11577 33517 11611
rect 33551 11608 33563 11611
rect 35066 11608 35072 11620
rect 33551 11580 35072 11608
rect 33551 11577 33563 11580
rect 33505 11571 33563 11577
rect 35066 11568 35072 11580
rect 35124 11568 35130 11620
rect 29270 11540 29276 11552
rect 28644 11512 29276 11540
rect 29270 11500 29276 11512
rect 29328 11500 29334 11552
rect 29546 11500 29552 11552
rect 29604 11540 29610 11552
rect 29840 11540 29868 11568
rect 29604 11512 29868 11540
rect 30837 11543 30895 11549
rect 29604 11500 29610 11512
rect 30837 11509 30849 11543
rect 30883 11540 30895 11543
rect 31754 11540 31760 11552
rect 30883 11512 31760 11540
rect 30883 11509 30895 11512
rect 30837 11503 30895 11509
rect 31754 11500 31760 11512
rect 31812 11500 31818 11552
rect 31941 11543 31999 11549
rect 31941 11509 31953 11543
rect 31987 11540 31999 11543
rect 32306 11540 32312 11552
rect 31987 11512 32312 11540
rect 31987 11509 31999 11512
rect 31941 11503 31999 11509
rect 32306 11500 32312 11512
rect 32364 11500 32370 11552
rect 33594 11500 33600 11552
rect 33652 11540 33658 11552
rect 33870 11540 33876 11552
rect 33652 11512 33876 11540
rect 33652 11500 33658 11512
rect 33870 11500 33876 11512
rect 33928 11500 33934 11552
rect 34793 11543 34851 11549
rect 34793 11509 34805 11543
rect 34839 11540 34851 11543
rect 35158 11540 35164 11552
rect 34839 11512 35164 11540
rect 34839 11509 34851 11512
rect 34793 11503 34851 11509
rect 35158 11500 35164 11512
rect 35216 11500 35222 11552
rect 35268 11540 35296 11648
rect 35437 11645 35449 11679
rect 35483 11676 35495 11679
rect 36909 11679 36967 11685
rect 35483 11648 36860 11676
rect 35483 11645 35495 11648
rect 35437 11639 35495 11645
rect 36832 11608 36860 11648
rect 36909 11645 36921 11679
rect 36955 11676 36967 11679
rect 38105 11679 38163 11685
rect 38105 11676 38117 11679
rect 36955 11648 38117 11676
rect 36955 11645 36967 11648
rect 36909 11639 36967 11645
rect 38105 11645 38117 11648
rect 38151 11645 38163 11679
rect 38105 11639 38163 11645
rect 39114 11636 39120 11688
rect 39172 11636 39178 11688
rect 39206 11636 39212 11688
rect 39264 11636 39270 11688
rect 40126 11636 40132 11688
rect 40184 11676 40190 11688
rect 40773 11679 40831 11685
rect 40773 11676 40785 11679
rect 40184 11648 40785 11676
rect 40184 11636 40190 11648
rect 40773 11645 40785 11648
rect 40819 11645 40831 11679
rect 40773 11639 40831 11645
rect 37366 11608 37372 11620
rect 36832 11580 37372 11608
rect 37366 11568 37372 11580
rect 37424 11568 37430 11620
rect 37461 11611 37519 11617
rect 37461 11577 37473 11611
rect 37507 11608 37519 11611
rect 41598 11608 41604 11620
rect 37507 11580 41604 11608
rect 37507 11577 37519 11580
rect 37461 11571 37519 11577
rect 41598 11568 41604 11580
rect 41656 11568 41662 11620
rect 45281 11611 45339 11617
rect 45281 11577 45293 11611
rect 45327 11608 45339 11611
rect 46658 11608 46664 11620
rect 45327 11580 46664 11608
rect 45327 11577 45339 11580
rect 45281 11571 45339 11577
rect 46658 11568 46664 11580
rect 46716 11568 46722 11620
rect 35618 11540 35624 11552
rect 35268 11512 35624 11540
rect 35618 11500 35624 11512
rect 35676 11500 35682 11552
rect 35986 11500 35992 11552
rect 36044 11540 36050 11552
rect 40497 11543 40555 11549
rect 40497 11540 40509 11543
rect 36044 11512 40509 11540
rect 36044 11500 36050 11512
rect 40497 11509 40509 11512
rect 40543 11509 40555 11543
rect 40497 11503 40555 11509
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 1210 11296 1216 11348
rect 1268 11336 1274 11348
rect 2133 11339 2191 11345
rect 2133 11336 2145 11339
rect 1268 11308 2145 11336
rect 1268 11296 1274 11308
rect 2133 11305 2145 11308
rect 2179 11305 2191 11339
rect 2133 11299 2191 11305
rect 9858 11296 9864 11348
rect 9916 11336 9922 11348
rect 10413 11339 10471 11345
rect 10413 11336 10425 11339
rect 9916 11308 10425 11336
rect 9916 11296 9922 11308
rect 10413 11305 10425 11308
rect 10459 11305 10471 11339
rect 10413 11299 10471 11305
rect 10778 11296 10784 11348
rect 10836 11336 10842 11348
rect 10873 11339 10931 11345
rect 10873 11336 10885 11339
rect 10836 11308 10885 11336
rect 10836 11296 10842 11308
rect 10873 11305 10885 11308
rect 10919 11336 10931 11339
rect 10919 11308 14044 11336
rect 10919 11305 10931 11308
rect 10873 11299 10931 11305
rect 1762 11228 1768 11280
rect 1820 11228 1826 11280
rect 10226 11228 10232 11280
rect 10284 11268 10290 11280
rect 10284 11240 11284 11268
rect 10284 11228 10290 11240
rect 10870 11160 10876 11212
rect 10928 11200 10934 11212
rect 11149 11203 11207 11209
rect 11149 11200 11161 11203
rect 10928 11172 11161 11200
rect 10928 11160 10934 11172
rect 11149 11169 11161 11172
rect 11195 11169 11207 11203
rect 11256 11200 11284 11240
rect 13906 11228 13912 11280
rect 13964 11228 13970 11280
rect 14016 11268 14044 11308
rect 14550 11296 14556 11348
rect 14608 11296 14614 11348
rect 16206 11296 16212 11348
rect 16264 11336 16270 11348
rect 16482 11336 16488 11348
rect 16264 11308 16488 11336
rect 16264 11296 16270 11308
rect 16482 11296 16488 11308
rect 16540 11296 16546 11348
rect 16942 11296 16948 11348
rect 17000 11296 17006 11348
rect 18141 11339 18199 11345
rect 18141 11305 18153 11339
rect 18187 11336 18199 11339
rect 19058 11336 19064 11348
rect 18187 11308 19064 11336
rect 18187 11305 18199 11308
rect 18141 11299 18199 11305
rect 19058 11296 19064 11308
rect 19116 11296 19122 11348
rect 19429 11339 19487 11345
rect 19429 11305 19441 11339
rect 19475 11336 19487 11339
rect 20162 11336 20168 11348
rect 19475 11308 20168 11336
rect 19475 11305 19487 11308
rect 19429 11299 19487 11305
rect 20162 11296 20168 11308
rect 20220 11296 20226 11348
rect 20612 11339 20670 11345
rect 20612 11305 20624 11339
rect 20658 11336 20670 11339
rect 20658 11308 23244 11336
rect 20658 11305 20670 11308
rect 20612 11299 20670 11305
rect 15562 11268 15568 11280
rect 14016 11240 15568 11268
rect 15562 11228 15568 11240
rect 15620 11228 15626 11280
rect 16022 11228 16028 11280
rect 16080 11268 16086 11280
rect 20070 11268 20076 11280
rect 16080 11240 16344 11268
rect 16080 11228 16086 11240
rect 11425 11203 11483 11209
rect 11425 11200 11437 11203
rect 11256 11172 11437 11200
rect 11149 11163 11207 11169
rect 11425 11169 11437 11172
rect 11471 11169 11483 11203
rect 11425 11163 11483 11169
rect 12158 11160 12164 11212
rect 12216 11200 12222 11212
rect 12216 11172 12664 11200
rect 12216 11160 12222 11172
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 2317 11135 2375 11141
rect 2317 11132 2329 11135
rect 1636 11104 2329 11132
rect 1636 11092 1642 11104
rect 2317 11101 2329 11104
rect 2363 11101 2375 11135
rect 12636 11132 12664 11172
rect 12710 11160 12716 11212
rect 12768 11200 12774 11212
rect 13357 11203 13415 11209
rect 13357 11200 13369 11203
rect 12768 11172 13369 11200
rect 12768 11160 12774 11172
rect 13357 11169 13369 11172
rect 13403 11169 13415 11203
rect 13357 11163 13415 11169
rect 15010 11160 15016 11212
rect 15068 11160 15074 11212
rect 15102 11160 15108 11212
rect 15160 11160 15166 11212
rect 16114 11160 16120 11212
rect 16172 11200 16178 11212
rect 16316 11209 16344 11240
rect 17604 11240 20076 11268
rect 17604 11209 17632 11240
rect 20070 11228 20076 11240
rect 20128 11228 20134 11280
rect 23216 11268 23244 11308
rect 23290 11296 23296 11348
rect 23348 11296 23354 11348
rect 26329 11339 26387 11345
rect 26329 11305 26341 11339
rect 26375 11336 26387 11339
rect 26602 11336 26608 11348
rect 26375 11308 26608 11336
rect 26375 11305 26387 11308
rect 26329 11299 26387 11305
rect 26602 11296 26608 11308
rect 26660 11296 26666 11348
rect 27154 11296 27160 11348
rect 27212 11336 27218 11348
rect 27212 11308 28672 11336
rect 27212 11296 27218 11308
rect 23566 11268 23572 11280
rect 23216 11240 23572 11268
rect 23566 11228 23572 11240
rect 23624 11228 23630 11280
rect 28644 11277 28672 11308
rect 28994 11296 29000 11348
rect 29052 11296 29058 11348
rect 31386 11336 31392 11348
rect 31036 11308 31392 11336
rect 28629 11271 28687 11277
rect 28629 11237 28641 11271
rect 28675 11268 28687 11271
rect 29362 11268 29368 11280
rect 28675 11240 29368 11268
rect 28675 11237 28687 11240
rect 28629 11231 28687 11237
rect 29362 11228 29368 11240
rect 29420 11228 29426 11280
rect 16209 11203 16267 11209
rect 16209 11200 16221 11203
rect 16172 11172 16221 11200
rect 16172 11160 16178 11172
rect 16209 11169 16221 11172
rect 16255 11169 16267 11203
rect 16209 11163 16267 11169
rect 16301 11203 16359 11209
rect 16301 11169 16313 11203
rect 16347 11169 16359 11203
rect 16301 11163 16359 11169
rect 17589 11203 17647 11209
rect 17589 11169 17601 11203
rect 17635 11169 17647 11203
rect 17589 11163 17647 11169
rect 18598 11160 18604 11212
rect 18656 11160 18662 11212
rect 18785 11203 18843 11209
rect 18785 11169 18797 11203
rect 18831 11200 18843 11203
rect 19702 11200 19708 11212
rect 18831 11172 19708 11200
rect 18831 11169 18843 11172
rect 18785 11163 18843 11169
rect 19702 11160 19708 11172
rect 19760 11160 19766 11212
rect 20349 11203 20407 11209
rect 20349 11169 20361 11203
rect 20395 11200 20407 11203
rect 20622 11200 20628 11212
rect 20395 11172 20628 11200
rect 20395 11169 20407 11172
rect 20349 11163 20407 11169
rect 20622 11160 20628 11172
rect 20680 11160 20686 11212
rect 22462 11160 22468 11212
rect 22520 11200 22526 11212
rect 22557 11203 22615 11209
rect 22557 11200 22569 11203
rect 22520 11172 22569 11200
rect 22520 11160 22526 11172
rect 22557 11169 22569 11172
rect 22603 11169 22615 11203
rect 22557 11163 22615 11169
rect 23937 11203 23995 11209
rect 23937 11169 23949 11203
rect 23983 11200 23995 11203
rect 24026 11200 24032 11212
rect 23983 11172 24032 11200
rect 23983 11169 23995 11172
rect 23937 11163 23995 11169
rect 24026 11160 24032 11172
rect 24084 11160 24090 11212
rect 24486 11160 24492 11212
rect 24544 11200 24550 11212
rect 24581 11203 24639 11209
rect 24581 11200 24593 11203
rect 24544 11172 24593 11200
rect 24544 11160 24550 11172
rect 24581 11169 24593 11172
rect 24627 11169 24639 11203
rect 24581 11163 24639 11169
rect 27157 11203 27215 11209
rect 27157 11169 27169 11203
rect 27203 11200 27215 11203
rect 27522 11200 27528 11212
rect 27203 11172 27528 11200
rect 27203 11169 27215 11172
rect 27157 11163 27215 11169
rect 27522 11160 27528 11172
rect 27580 11200 27586 11212
rect 29178 11200 29184 11212
rect 27580 11172 29184 11200
rect 27580 11160 27586 11172
rect 29178 11160 29184 11172
rect 29236 11200 29242 11212
rect 29638 11200 29644 11212
rect 29236 11172 29644 11200
rect 29236 11160 29242 11172
rect 29638 11160 29644 11172
rect 29696 11160 29702 11212
rect 17313 11135 17371 11141
rect 17313 11132 17325 11135
rect 12636 11104 17325 11132
rect 2317 11095 2375 11101
rect 17313 11101 17325 11104
rect 17359 11101 17371 11135
rect 17313 11095 17371 11101
rect 18506 11092 18512 11144
rect 18564 11132 18570 11144
rect 18966 11132 18972 11144
rect 18564 11104 18972 11132
rect 18564 11092 18570 11104
rect 18966 11092 18972 11104
rect 19024 11092 19030 11144
rect 23661 11135 23719 11141
rect 23661 11101 23673 11135
rect 23707 11132 23719 11135
rect 24302 11132 24308 11144
rect 23707 11104 24308 11132
rect 23707 11101 23719 11104
rect 23661 11095 23719 11101
rect 24302 11092 24308 11104
rect 24360 11092 24366 11144
rect 25958 11092 25964 11144
rect 26016 11132 26022 11144
rect 26694 11132 26700 11144
rect 26016 11104 26700 11132
rect 26016 11092 26022 11104
rect 26694 11092 26700 11104
rect 26752 11132 26758 11144
rect 26752 11104 26832 11132
rect 26752 11092 26758 11104
rect 10594 11024 10600 11076
rect 10652 11064 10658 11076
rect 10652 11036 11836 11064
rect 10652 11024 10658 11036
rect 11422 10956 11428 11008
rect 11480 10996 11486 11008
rect 11698 10996 11704 11008
rect 11480 10968 11704 10996
rect 11480 10956 11486 10968
rect 11698 10956 11704 10968
rect 11756 10956 11762 11008
rect 11808 10996 11836 11036
rect 11882 11024 11888 11076
rect 11940 11024 11946 11076
rect 14277 11067 14335 11073
rect 12728 11036 14228 11064
rect 12728 10996 12756 11036
rect 11808 10968 12756 10996
rect 12897 10999 12955 11005
rect 12897 10965 12909 10999
rect 12943 10996 12955 10999
rect 13354 10996 13360 11008
rect 12943 10968 13360 10996
rect 12943 10965 12955 10968
rect 12897 10959 12955 10965
rect 13354 10956 13360 10968
rect 13412 10956 13418 11008
rect 14200 10996 14228 11036
rect 14277 11033 14289 11067
rect 14323 11064 14335 11067
rect 15102 11064 15108 11076
rect 14323 11036 15108 11064
rect 14323 11033 14335 11036
rect 14277 11027 14335 11033
rect 15102 11024 15108 11036
rect 15160 11024 15166 11076
rect 16114 11024 16120 11076
rect 16172 11024 16178 11076
rect 17405 11067 17463 11073
rect 17405 11033 17417 11067
rect 17451 11064 17463 11067
rect 19705 11067 19763 11073
rect 17451 11036 19656 11064
rect 17451 11033 17463 11036
rect 17405 11027 17463 11033
rect 14921 10999 14979 11005
rect 14921 10996 14933 10999
rect 14200 10968 14933 10996
rect 14921 10965 14933 10968
rect 14967 10996 14979 10999
rect 15010 10996 15016 11008
rect 14967 10968 15016 10996
rect 14967 10965 14979 10968
rect 14921 10959 14979 10965
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 15746 10956 15752 11008
rect 15804 10956 15810 11008
rect 17494 10956 17500 11008
rect 17552 10996 17558 11008
rect 18230 10996 18236 11008
rect 17552 10968 18236 10996
rect 17552 10956 17558 10968
rect 18230 10956 18236 10968
rect 18288 10956 18294 11008
rect 19628 10996 19656 11036
rect 19705 11033 19717 11067
rect 19751 11064 19763 11067
rect 20898 11064 20904 11076
rect 19751 11036 20904 11064
rect 19751 11033 19763 11036
rect 19705 11027 19763 11033
rect 20898 11024 20904 11036
rect 20956 11024 20962 11076
rect 21082 11024 21088 11076
rect 21140 11024 21146 11076
rect 23750 11024 23756 11076
rect 23808 11024 23814 11076
rect 24854 11024 24860 11076
rect 24912 11024 24918 11076
rect 26804 11064 26832 11104
rect 26878 11092 26884 11144
rect 26936 11092 26942 11144
rect 31036 11132 31064 11308
rect 31386 11296 31392 11308
rect 31444 11296 31450 11348
rect 34606 11296 34612 11348
rect 34664 11336 34670 11348
rect 34701 11339 34759 11345
rect 34701 11336 34713 11339
rect 34664 11308 34713 11336
rect 34664 11296 34670 11308
rect 34701 11305 34713 11308
rect 34747 11305 34759 11339
rect 34701 11299 34759 11305
rect 35066 11296 35072 11348
rect 35124 11336 35130 11348
rect 40221 11339 40279 11345
rect 35124 11308 39528 11336
rect 35124 11296 35130 11308
rect 33505 11271 33563 11277
rect 33505 11237 33517 11271
rect 33551 11268 33563 11271
rect 33551 11240 35848 11268
rect 33551 11237 33563 11240
rect 33505 11231 33563 11237
rect 31389 11203 31447 11209
rect 31389 11169 31401 11203
rect 31435 11200 31447 11203
rect 31754 11200 31760 11212
rect 31435 11172 31760 11200
rect 31435 11169 31447 11172
rect 31389 11163 31447 11169
rect 31754 11160 31760 11172
rect 31812 11160 31818 11212
rect 32674 11160 32680 11212
rect 32732 11200 32738 11212
rect 32858 11200 32864 11212
rect 32732 11172 32864 11200
rect 32732 11160 32738 11172
rect 32858 11160 32864 11172
rect 32916 11160 32922 11212
rect 33594 11160 33600 11212
rect 33652 11200 33658 11212
rect 34057 11203 34115 11209
rect 34057 11200 34069 11203
rect 33652 11172 34069 11200
rect 33652 11160 33658 11172
rect 34057 11169 34069 11172
rect 34103 11200 34115 11203
rect 34238 11200 34244 11212
rect 34103 11172 34244 11200
rect 34103 11169 34115 11172
rect 34057 11163 34115 11169
rect 34238 11160 34244 11172
rect 34296 11160 34302 11212
rect 35820 11200 35848 11240
rect 37366 11228 37372 11280
rect 37424 11268 37430 11280
rect 38841 11271 38899 11277
rect 38841 11268 38853 11271
rect 37424 11240 38853 11268
rect 37424 11228 37430 11240
rect 38841 11237 38853 11240
rect 38887 11237 38899 11271
rect 38841 11231 38899 11237
rect 39114 11200 39120 11212
rect 35820 11172 39120 11200
rect 39114 11160 39120 11172
rect 39172 11160 39178 11212
rect 28644 11104 31064 11132
rect 31113 11135 31171 11141
rect 26804 11036 27646 11064
rect 20806 10996 20812 11008
rect 19628 10968 20812 10996
rect 20806 10956 20812 10968
rect 20864 10956 20870 11008
rect 21634 10956 21640 11008
rect 21692 10996 21698 11008
rect 22097 10999 22155 11005
rect 22097 10996 22109 10999
rect 21692 10968 22109 10996
rect 21692 10956 21698 10968
rect 22097 10965 22109 10968
rect 22143 10965 22155 10999
rect 22097 10959 22155 10965
rect 24670 10956 24676 11008
rect 24728 10996 24734 11008
rect 28644 10996 28672 11104
rect 31113 11101 31125 11135
rect 31159 11101 31171 11135
rect 31113 11095 31171 11101
rect 29362 11024 29368 11076
rect 29420 11064 29426 11076
rect 29730 11064 29736 11076
rect 29420 11036 29736 11064
rect 29420 11024 29426 11036
rect 29730 11024 29736 11036
rect 29788 11024 29794 11076
rect 30374 11024 30380 11076
rect 30432 11064 30438 11076
rect 30469 11067 30527 11073
rect 30469 11064 30481 11067
rect 30432 11036 30481 11064
rect 30432 11024 30438 11036
rect 30469 11033 30481 11036
rect 30515 11064 30527 11067
rect 31128 11064 31156 11095
rect 33778 11092 33784 11144
rect 33836 11132 33842 11144
rect 33965 11135 34023 11141
rect 33965 11132 33977 11135
rect 33836 11104 33977 11132
rect 33836 11092 33842 11104
rect 33965 11101 33977 11104
rect 34011 11132 34023 11135
rect 34146 11132 34152 11144
rect 34011 11104 34152 11132
rect 34011 11101 34023 11104
rect 33965 11095 34023 11101
rect 34146 11092 34152 11104
rect 34204 11092 34210 11144
rect 35618 11092 35624 11144
rect 35676 11132 35682 11144
rect 35713 11135 35771 11141
rect 35713 11132 35725 11135
rect 35676 11104 35725 11132
rect 35676 11092 35682 11104
rect 35713 11101 35725 11104
rect 35759 11101 35771 11135
rect 35713 11095 35771 11101
rect 37274 11092 37280 11144
rect 37332 11132 37338 11144
rect 38197 11135 38255 11141
rect 38197 11132 38209 11135
rect 37332 11104 38209 11132
rect 37332 11092 37338 11104
rect 38197 11101 38209 11104
rect 38243 11132 38255 11135
rect 39206 11132 39212 11144
rect 38243 11104 39212 11132
rect 38243 11101 38255 11104
rect 38197 11095 38255 11101
rect 39206 11092 39212 11104
rect 39264 11092 39270 11144
rect 39500 11141 39528 11308
rect 40221 11305 40233 11339
rect 40267 11336 40279 11339
rect 47118 11336 47124 11348
rect 40267 11308 47124 11336
rect 40267 11305 40279 11308
rect 40221 11299 40279 11305
rect 47118 11296 47124 11308
rect 47176 11296 47182 11348
rect 41509 11271 41567 11277
rect 41509 11237 41521 11271
rect 41555 11237 41567 11271
rect 41509 11231 41567 11237
rect 41524 11200 41552 11231
rect 44174 11228 44180 11280
rect 44232 11268 44238 11280
rect 44232 11240 47992 11268
rect 44232 11228 44238 11240
rect 41524 11172 45554 11200
rect 39485 11135 39543 11141
rect 39485 11101 39497 11135
rect 39531 11101 39543 11135
rect 39485 11095 39543 11101
rect 40034 11092 40040 11144
rect 40092 11132 40098 11144
rect 41693 11135 41751 11141
rect 41693 11132 41705 11135
rect 40092 11104 41705 11132
rect 40092 11092 40098 11104
rect 41693 11101 41705 11104
rect 41739 11101 41751 11135
rect 45526 11132 45554 11172
rect 47964 11141 47992 11240
rect 49142 11160 49148 11212
rect 49200 11160 49206 11212
rect 45649 11135 45707 11141
rect 45649 11132 45661 11135
rect 45526 11104 45661 11132
rect 41693 11095 41751 11101
rect 45649 11101 45661 11104
rect 45695 11101 45707 11135
rect 45649 11095 45707 11101
rect 47949 11135 48007 11141
rect 47949 11101 47961 11135
rect 47995 11101 48007 11135
rect 47949 11095 48007 11101
rect 30515 11036 31156 11064
rect 31220 11036 31754 11064
rect 32614 11036 32720 11064
rect 30515 11033 30527 11036
rect 30469 11027 30527 11033
rect 24728 10968 28672 10996
rect 24728 10956 24734 10968
rect 28718 10956 28724 11008
rect 28776 10996 28782 11008
rect 29089 10999 29147 11005
rect 29089 10996 29101 10999
rect 28776 10968 29101 10996
rect 28776 10956 28782 10968
rect 29089 10965 29101 10968
rect 29135 10996 29147 10999
rect 29273 10999 29331 11005
rect 29273 10996 29285 10999
rect 29135 10968 29285 10996
rect 29135 10965 29147 10968
rect 29089 10959 29147 10965
rect 29273 10965 29285 10968
rect 29319 10996 29331 10999
rect 29454 10996 29460 11008
rect 29319 10968 29460 10996
rect 29319 10965 29331 10968
rect 29273 10959 29331 10965
rect 29454 10956 29460 10968
rect 29512 10996 29518 11008
rect 30282 10996 30288 11008
rect 29512 10968 30288 10996
rect 29512 10956 29518 10968
rect 30282 10956 30288 10968
rect 30340 10996 30346 11008
rect 31220 10996 31248 11036
rect 30340 10968 31248 10996
rect 31726 10996 31754 11036
rect 32306 10996 32312 11008
rect 31726 10968 32312 10996
rect 30340 10956 30346 10968
rect 32306 10956 32312 10968
rect 32364 10996 32370 11008
rect 32692 10996 32720 11036
rect 33870 11024 33876 11076
rect 33928 11064 33934 11076
rect 35250 11064 35256 11076
rect 33928 11036 35256 11064
rect 33928 11024 33934 11036
rect 35250 11024 35256 11036
rect 35308 11024 35314 11076
rect 35986 11024 35992 11076
rect 36044 11024 36050 11076
rect 36722 11024 36728 11076
rect 36780 11024 36786 11076
rect 37734 11024 37740 11076
rect 37792 11024 37798 11076
rect 40126 11024 40132 11076
rect 40184 11024 40190 11076
rect 40770 11024 40776 11076
rect 40828 11064 40834 11076
rect 40865 11067 40923 11073
rect 40865 11064 40877 11067
rect 40828 11036 40877 11064
rect 40828 11024 40834 11036
rect 40865 11033 40877 11036
rect 40911 11033 40923 11067
rect 40865 11027 40923 11033
rect 41049 11067 41107 11073
rect 41049 11033 41061 11067
rect 41095 11064 41107 11067
rect 44174 11064 44180 11076
rect 41095 11036 44180 11064
rect 41095 11033 41107 11036
rect 41049 11027 41107 11033
rect 44174 11024 44180 11036
rect 44232 11024 44238 11076
rect 45833 11067 45891 11073
rect 45833 11033 45845 11067
rect 45879 11064 45891 11067
rect 46934 11064 46940 11076
rect 45879 11036 46940 11064
rect 45879 11033 45891 11036
rect 45833 11027 45891 11033
rect 46934 11024 46940 11036
rect 46992 11024 46998 11076
rect 33229 10999 33287 11005
rect 33229 10996 33241 10999
rect 32364 10968 33241 10996
rect 32364 10956 32370 10968
rect 33229 10965 33241 10968
rect 33275 10996 33287 10999
rect 33318 10996 33324 11008
rect 33275 10968 33324 10996
rect 33275 10965 33287 10968
rect 33229 10959 33287 10965
rect 33318 10956 33324 10968
rect 33376 10996 33382 11008
rect 34977 10999 35035 11005
rect 34977 10996 34989 10999
rect 33376 10968 34989 10996
rect 33376 10956 33382 10968
rect 34977 10965 34989 10968
rect 35023 10996 35035 10999
rect 35158 10996 35164 11008
rect 35023 10968 35164 10996
rect 35023 10965 35035 10968
rect 34977 10959 35035 10965
rect 35158 10956 35164 10968
rect 35216 10956 35222 11008
rect 39298 10956 39304 11008
rect 39356 10956 39362 11008
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 1854 10752 1860 10804
rect 1912 10792 1918 10804
rect 11422 10792 11428 10804
rect 1912 10764 11428 10792
rect 1912 10752 1918 10764
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 11698 10752 11704 10804
rect 11756 10792 11762 10804
rect 12345 10795 12403 10801
rect 12345 10792 12357 10795
rect 11756 10764 12357 10792
rect 11756 10752 11762 10764
rect 12345 10761 12357 10764
rect 12391 10761 12403 10795
rect 12345 10755 12403 10761
rect 12526 10752 12532 10804
rect 12584 10792 12590 10804
rect 13633 10795 13691 10801
rect 13633 10792 13645 10795
rect 12584 10764 13645 10792
rect 12584 10752 12590 10764
rect 13633 10761 13645 10764
rect 13679 10761 13691 10795
rect 13633 10755 13691 10761
rect 14829 10795 14887 10801
rect 14829 10761 14841 10795
rect 14875 10792 14887 10795
rect 15194 10792 15200 10804
rect 14875 10764 15200 10792
rect 14875 10761 14887 10764
rect 14829 10755 14887 10761
rect 15194 10752 15200 10764
rect 15252 10752 15258 10804
rect 15565 10795 15623 10801
rect 15565 10761 15577 10795
rect 15611 10792 15623 10795
rect 17405 10795 17463 10801
rect 17405 10792 17417 10795
rect 15611 10764 17417 10792
rect 15611 10761 15623 10764
rect 15565 10755 15623 10761
rect 17405 10761 17417 10764
rect 17451 10761 17463 10795
rect 17405 10755 17463 10761
rect 18049 10795 18107 10801
rect 18049 10761 18061 10795
rect 18095 10792 18107 10795
rect 18322 10792 18328 10804
rect 18095 10764 18328 10792
rect 18095 10761 18107 10764
rect 18049 10755 18107 10761
rect 1210 10684 1216 10736
rect 1268 10724 1274 10736
rect 14918 10724 14924 10736
rect 1268 10696 2360 10724
rect 1268 10684 1274 10696
rect 1302 10616 1308 10668
rect 1360 10656 1366 10668
rect 2332 10665 2360 10696
rect 6886 10696 14924 10724
rect 1581 10659 1639 10665
rect 1581 10656 1593 10659
rect 1360 10628 1593 10656
rect 1360 10616 1366 10628
rect 1581 10625 1593 10628
rect 1627 10625 1639 10659
rect 1581 10619 1639 10625
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 2363 10628 2881 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 2869 10625 2881 10628
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 1596 10588 1624 10619
rect 3053 10591 3111 10597
rect 3053 10588 3065 10591
rect 1596 10560 3065 10588
rect 3053 10557 3065 10560
rect 3099 10557 3111 10591
rect 3053 10551 3111 10557
rect 1765 10523 1823 10529
rect 1765 10489 1777 10523
rect 1811 10520 1823 10523
rect 6886 10520 6914 10696
rect 14918 10684 14924 10696
rect 14976 10684 14982 10736
rect 17770 10724 17776 10736
rect 15856 10696 17776 10724
rect 10318 10616 10324 10668
rect 10376 10656 10382 10668
rect 11609 10659 11667 10665
rect 11609 10656 11621 10659
rect 10376 10628 11621 10656
rect 10376 10616 10382 10628
rect 11609 10625 11621 10628
rect 11655 10625 11667 10659
rect 11609 10619 11667 10625
rect 12250 10616 12256 10668
rect 12308 10656 12314 10668
rect 13541 10659 13599 10665
rect 12308 10628 12572 10656
rect 12308 10616 12314 10628
rect 12544 10597 12572 10628
rect 13541 10625 13553 10659
rect 13587 10656 13599 10659
rect 14737 10659 14795 10665
rect 13587 10628 14688 10656
rect 13587 10625 13599 10628
rect 13541 10619 13599 10625
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10557 12495 10591
rect 12437 10551 12495 10557
rect 12529 10591 12587 10597
rect 12529 10557 12541 10591
rect 12575 10557 12587 10591
rect 12529 10551 12587 10557
rect 1811 10492 6914 10520
rect 12452 10520 12480 10551
rect 13814 10548 13820 10600
rect 13872 10548 13878 10600
rect 14660 10588 14688 10628
rect 14737 10625 14749 10659
rect 14783 10656 14795 10659
rect 15856 10656 15884 10696
rect 17770 10684 17776 10696
rect 17828 10684 17834 10736
rect 14783 10628 15884 10656
rect 15933 10659 15991 10665
rect 14783 10625 14795 10628
rect 14737 10619 14795 10625
rect 15933 10625 15945 10659
rect 15979 10656 15991 10659
rect 16482 10656 16488 10668
rect 15979 10628 16488 10656
rect 15979 10625 15991 10628
rect 15933 10619 15991 10625
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 16574 10616 16580 10668
rect 16632 10656 16638 10668
rect 17313 10659 17371 10665
rect 17313 10656 17325 10659
rect 16632 10628 17325 10656
rect 16632 10616 16638 10628
rect 17313 10625 17325 10628
rect 17359 10625 17371 10659
rect 18064 10656 18092 10755
rect 18322 10752 18328 10764
rect 18380 10752 18386 10804
rect 18782 10752 18788 10804
rect 18840 10752 18846 10804
rect 19521 10795 19579 10801
rect 19521 10761 19533 10795
rect 19567 10792 19579 10795
rect 19610 10792 19616 10804
rect 19567 10764 19616 10792
rect 19567 10761 19579 10764
rect 19521 10755 19579 10761
rect 19610 10752 19616 10764
rect 19668 10752 19674 10804
rect 20714 10752 20720 10804
rect 20772 10752 20778 10804
rect 20898 10752 20904 10804
rect 20956 10792 20962 10804
rect 21085 10795 21143 10801
rect 21085 10792 21097 10795
rect 20956 10764 21097 10792
rect 20956 10752 20962 10764
rect 21085 10761 21097 10764
rect 21131 10761 21143 10795
rect 21085 10755 21143 10761
rect 21177 10795 21235 10801
rect 21177 10761 21189 10795
rect 21223 10792 21235 10795
rect 22646 10792 22652 10804
rect 21223 10764 22652 10792
rect 21223 10761 21235 10764
rect 21177 10755 21235 10761
rect 22646 10752 22652 10764
rect 22704 10752 22710 10804
rect 23566 10752 23572 10804
rect 23624 10792 23630 10804
rect 23753 10795 23811 10801
rect 23753 10792 23765 10795
rect 23624 10764 23765 10792
rect 23624 10752 23630 10764
rect 23753 10761 23765 10764
rect 23799 10792 23811 10795
rect 24394 10792 24400 10804
rect 23799 10764 24400 10792
rect 23799 10761 23811 10764
rect 23753 10755 23811 10761
rect 24394 10752 24400 10764
rect 24452 10752 24458 10804
rect 24486 10752 24492 10804
rect 24544 10792 24550 10804
rect 25314 10792 25320 10804
rect 24544 10764 25320 10792
rect 24544 10752 24550 10764
rect 25314 10752 25320 10764
rect 25372 10752 25378 10804
rect 25501 10795 25559 10801
rect 25501 10761 25513 10795
rect 25547 10792 25559 10795
rect 25685 10795 25743 10801
rect 25685 10792 25697 10795
rect 25547 10764 25697 10792
rect 25547 10761 25559 10764
rect 25501 10755 25559 10761
rect 25685 10761 25697 10764
rect 25731 10792 25743 10795
rect 25958 10792 25964 10804
rect 25731 10764 25964 10792
rect 25731 10761 25743 10764
rect 25685 10755 25743 10761
rect 25958 10752 25964 10764
rect 26016 10752 26022 10804
rect 27157 10795 27215 10801
rect 27157 10761 27169 10795
rect 27203 10792 27215 10795
rect 31389 10795 31447 10801
rect 31389 10792 31401 10795
rect 27203 10764 31401 10792
rect 27203 10761 27215 10764
rect 27157 10755 27215 10761
rect 31389 10761 31401 10764
rect 31435 10761 31447 10795
rect 31389 10755 31447 10761
rect 31478 10752 31484 10804
rect 31536 10792 31542 10804
rect 32769 10795 32827 10801
rect 32769 10792 32781 10795
rect 31536 10764 32781 10792
rect 31536 10752 31542 10764
rect 32769 10761 32781 10764
rect 32815 10761 32827 10795
rect 32769 10755 32827 10761
rect 33318 10752 33324 10804
rect 33376 10752 33382 10804
rect 39209 10795 39267 10801
rect 39209 10792 39221 10795
rect 34072 10764 39221 10792
rect 18598 10684 18604 10736
rect 18656 10724 18662 10736
rect 19981 10727 20039 10733
rect 19981 10724 19993 10727
rect 18656 10696 19993 10724
rect 18656 10684 18662 10696
rect 19981 10693 19993 10696
rect 20027 10724 20039 10727
rect 21450 10724 21456 10736
rect 20027 10696 21456 10724
rect 20027 10693 20039 10696
rect 19981 10687 20039 10693
rect 21450 10684 21456 10696
rect 21508 10684 21514 10736
rect 22020 10696 22770 10724
rect 17313 10619 17371 10625
rect 17420 10628 18092 10656
rect 15013 10591 15071 10597
rect 14660 10560 14964 10588
rect 12802 10520 12808 10532
rect 12452 10492 12808 10520
rect 1811 10489 1823 10492
rect 1765 10483 1823 10489
rect 12802 10480 12808 10492
rect 12860 10480 12866 10532
rect 13173 10523 13231 10529
rect 13173 10489 13185 10523
rect 13219 10520 13231 10523
rect 14826 10520 14832 10532
rect 13219 10492 14832 10520
rect 13219 10489 13231 10492
rect 13173 10483 13231 10489
rect 14826 10480 14832 10492
rect 14884 10480 14890 10532
rect 2498 10412 2504 10464
rect 2556 10412 2562 10464
rect 11238 10412 11244 10464
rect 11296 10412 11302 10464
rect 11977 10455 12035 10461
rect 11977 10421 11989 10455
rect 12023 10452 12035 10455
rect 12710 10452 12716 10464
rect 12023 10424 12716 10452
rect 12023 10421 12035 10424
rect 11977 10415 12035 10421
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 14366 10412 14372 10464
rect 14424 10412 14430 10464
rect 14936 10452 14964 10560
rect 15013 10557 15025 10591
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 15028 10520 15056 10551
rect 15378 10548 15384 10600
rect 15436 10588 15442 10600
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 15436 10560 16037 10588
rect 15436 10548 15442 10560
rect 16025 10557 16037 10560
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 16206 10548 16212 10600
rect 16264 10548 16270 10600
rect 16390 10548 16396 10600
rect 16448 10588 16454 10600
rect 17420 10588 17448 10628
rect 18690 10616 18696 10668
rect 18748 10616 18754 10668
rect 19886 10616 19892 10668
rect 19944 10616 19950 10668
rect 20530 10616 20536 10668
rect 20588 10656 20594 10668
rect 20990 10656 20996 10668
rect 20588 10628 20996 10656
rect 20588 10616 20594 10628
rect 20990 10616 20996 10628
rect 21048 10616 21054 10668
rect 21082 10616 21088 10668
rect 21140 10656 21146 10668
rect 22020 10656 22048 10696
rect 24026 10684 24032 10736
rect 24084 10724 24090 10736
rect 24670 10724 24676 10736
rect 24084 10696 24676 10724
rect 24084 10684 24090 10696
rect 24670 10684 24676 10696
rect 24728 10684 24734 10736
rect 27614 10684 27620 10736
rect 27672 10724 27678 10736
rect 28813 10727 28871 10733
rect 28813 10724 28825 10727
rect 27672 10696 28825 10724
rect 27672 10684 27678 10696
rect 28813 10693 28825 10696
rect 28859 10693 28871 10727
rect 28813 10687 28871 10693
rect 29270 10684 29276 10736
rect 29328 10724 29334 10736
rect 29328 10696 29868 10724
rect 29328 10684 29334 10696
rect 21140 10628 22048 10656
rect 21140 10616 21146 10628
rect 24578 10616 24584 10668
rect 24636 10616 24642 10668
rect 25961 10659 26019 10665
rect 25961 10656 25973 10659
rect 24872 10628 25973 10656
rect 16448 10560 17448 10588
rect 17589 10591 17647 10597
rect 16448 10548 16454 10560
rect 17589 10557 17601 10591
rect 17635 10588 17647 10591
rect 18782 10588 18788 10600
rect 17635 10560 18788 10588
rect 17635 10557 17647 10560
rect 17589 10551 17647 10557
rect 18782 10548 18788 10560
rect 18840 10548 18846 10600
rect 18874 10548 18880 10600
rect 18932 10548 18938 10600
rect 20165 10591 20223 10597
rect 20165 10557 20177 10591
rect 20211 10588 20223 10591
rect 21174 10588 21180 10600
rect 20211 10560 21180 10588
rect 20211 10557 20223 10560
rect 20165 10551 20223 10557
rect 21174 10548 21180 10560
rect 21232 10548 21238 10600
rect 21361 10591 21419 10597
rect 21361 10557 21373 10591
rect 21407 10557 21419 10591
rect 21361 10551 21419 10557
rect 16666 10520 16672 10532
rect 15028 10492 16672 10520
rect 16666 10480 16672 10492
rect 16724 10480 16730 10532
rect 16758 10480 16764 10532
rect 16816 10520 16822 10532
rect 16945 10523 17003 10529
rect 16945 10520 16957 10523
rect 16816 10492 16957 10520
rect 16816 10480 16822 10492
rect 16945 10489 16957 10492
rect 16991 10489 17003 10523
rect 21376 10520 21404 10551
rect 22002 10548 22008 10600
rect 22060 10548 22066 10600
rect 22278 10548 22284 10600
rect 22336 10548 22342 10600
rect 22370 10548 22376 10600
rect 22428 10588 22434 10600
rect 24872 10597 24900 10628
rect 25961 10625 25973 10628
rect 26007 10656 26019 10659
rect 26602 10656 26608 10668
rect 26007 10628 26608 10656
rect 26007 10625 26019 10628
rect 25961 10619 26019 10625
rect 26602 10616 26608 10628
rect 26660 10616 26666 10668
rect 27062 10616 27068 10668
rect 27120 10656 27126 10668
rect 27525 10659 27583 10665
rect 27525 10656 27537 10659
rect 27120 10628 27537 10656
rect 27120 10616 27126 10628
rect 27525 10625 27537 10628
rect 27571 10625 27583 10659
rect 27525 10619 27583 10625
rect 28721 10659 28779 10665
rect 28721 10625 28733 10659
rect 28767 10656 28779 10659
rect 29638 10656 29644 10668
rect 28767 10628 29644 10656
rect 28767 10625 28779 10628
rect 28721 10619 28779 10625
rect 29638 10616 29644 10628
rect 29696 10616 29702 10668
rect 29840 10665 29868 10696
rect 29914 10684 29920 10736
rect 29972 10724 29978 10736
rect 34072 10733 34100 10764
rect 39209 10761 39221 10764
rect 39255 10761 39267 10795
rect 39209 10755 39267 10761
rect 40126 10752 40132 10804
rect 40184 10792 40190 10804
rect 40221 10795 40279 10801
rect 40221 10792 40233 10795
rect 40184 10764 40233 10792
rect 40184 10752 40190 10764
rect 40221 10761 40233 10764
rect 40267 10761 40279 10795
rect 40221 10755 40279 10761
rect 40681 10795 40739 10801
rect 40681 10761 40693 10795
rect 40727 10792 40739 10795
rect 40770 10792 40776 10804
rect 40727 10764 40776 10792
rect 40727 10761 40739 10764
rect 40681 10755 40739 10761
rect 40770 10752 40776 10764
rect 40828 10752 40834 10804
rect 32677 10727 32735 10733
rect 32677 10724 32689 10727
rect 29972 10696 32689 10724
rect 29972 10684 29978 10696
rect 32677 10693 32689 10696
rect 32723 10693 32735 10727
rect 32677 10687 32735 10693
rect 34057 10727 34115 10733
rect 34057 10693 34069 10727
rect 34103 10693 34115 10727
rect 34057 10687 34115 10693
rect 35526 10684 35532 10736
rect 35584 10724 35590 10736
rect 36541 10727 36599 10733
rect 36541 10724 36553 10727
rect 35584 10696 36553 10724
rect 35584 10684 35590 10696
rect 36541 10693 36553 10696
rect 36587 10693 36599 10727
rect 36541 10687 36599 10693
rect 49145 10727 49203 10733
rect 49145 10693 49157 10727
rect 49191 10724 49203 10727
rect 49234 10724 49240 10736
rect 49191 10696 49240 10724
rect 49191 10693 49203 10696
rect 49145 10687 49203 10693
rect 49234 10684 49240 10696
rect 49292 10684 49298 10736
rect 29825 10659 29883 10665
rect 29825 10625 29837 10659
rect 29871 10625 29883 10659
rect 29825 10619 29883 10625
rect 31294 10616 31300 10668
rect 31352 10616 31358 10668
rect 35158 10616 35164 10668
rect 35216 10656 35222 10668
rect 35710 10656 35716 10668
rect 35216 10628 35716 10656
rect 35216 10616 35222 10628
rect 35710 10616 35716 10628
rect 35768 10616 35774 10668
rect 36446 10616 36452 10668
rect 36504 10616 36510 10668
rect 37274 10656 37280 10668
rect 36556 10628 37280 10656
rect 24857 10591 24915 10597
rect 22428 10560 24256 10588
rect 22428 10548 22434 10560
rect 24228 10529 24256 10560
rect 24857 10557 24869 10591
rect 24903 10557 24915 10591
rect 24857 10551 24915 10557
rect 27246 10548 27252 10600
rect 27304 10588 27310 10600
rect 27617 10591 27675 10597
rect 27617 10588 27629 10591
rect 27304 10560 27629 10588
rect 27304 10548 27310 10560
rect 27617 10557 27629 10560
rect 27663 10557 27675 10591
rect 27617 10551 27675 10557
rect 27801 10591 27859 10597
rect 27801 10557 27813 10591
rect 27847 10557 27859 10591
rect 27801 10551 27859 10557
rect 24213 10523 24271 10529
rect 21376 10492 22094 10520
rect 16945 10483 17003 10489
rect 17586 10452 17592 10464
rect 14936 10424 17592 10452
rect 17586 10412 17592 10424
rect 17644 10412 17650 10464
rect 18322 10412 18328 10464
rect 18380 10412 18386 10464
rect 22066 10452 22094 10492
rect 24213 10489 24225 10523
rect 24259 10489 24271 10523
rect 27816 10520 27844 10551
rect 28810 10548 28816 10600
rect 28868 10588 28874 10600
rect 28905 10591 28963 10597
rect 28905 10588 28917 10591
rect 28868 10560 28917 10588
rect 28868 10548 28874 10560
rect 28905 10557 28917 10560
rect 28951 10557 28963 10591
rect 28905 10551 28963 10557
rect 28994 10548 29000 10600
rect 29052 10588 29058 10600
rect 30469 10591 30527 10597
rect 30469 10588 30481 10591
rect 29052 10560 30481 10588
rect 29052 10548 29058 10560
rect 30469 10557 30481 10560
rect 30515 10557 30527 10591
rect 30469 10551 30527 10557
rect 31570 10548 31576 10600
rect 31628 10548 31634 10600
rect 32861 10591 32919 10597
rect 32861 10557 32873 10591
rect 32907 10557 32919 10591
rect 32861 10551 32919 10557
rect 27816 10492 29500 10520
rect 24213 10483 24271 10489
rect 22738 10452 22744 10464
rect 22066 10424 22744 10452
rect 22738 10412 22744 10424
rect 22796 10412 22802 10464
rect 26602 10412 26608 10464
rect 26660 10412 26666 10464
rect 28353 10455 28411 10461
rect 28353 10421 28365 10455
rect 28399 10452 28411 10455
rect 29270 10452 29276 10464
rect 28399 10424 29276 10452
rect 28399 10421 28411 10424
rect 28353 10415 28411 10421
rect 29270 10412 29276 10424
rect 29328 10412 29334 10464
rect 29472 10461 29500 10492
rect 30926 10480 30932 10532
rect 30984 10480 30990 10532
rect 32876 10520 32904 10551
rect 33778 10548 33784 10600
rect 33836 10548 33842 10600
rect 35802 10588 35808 10600
rect 33888 10560 35808 10588
rect 33888 10520 33916 10560
rect 35802 10548 35808 10560
rect 35860 10548 35866 10600
rect 36556 10588 36584 10628
rect 37274 10616 37280 10628
rect 37332 10656 37338 10668
rect 37461 10659 37519 10665
rect 37461 10656 37473 10659
rect 37332 10628 37473 10656
rect 37332 10616 37338 10628
rect 37461 10625 37473 10628
rect 37507 10625 37519 10659
rect 37461 10619 37519 10625
rect 38565 10659 38623 10665
rect 38565 10625 38577 10659
rect 38611 10625 38623 10659
rect 38565 10619 38623 10625
rect 35912 10560 36584 10588
rect 35912 10532 35940 10560
rect 36630 10548 36636 10600
rect 36688 10588 36694 10600
rect 36725 10591 36783 10597
rect 36725 10588 36737 10591
rect 36688 10560 36737 10588
rect 36688 10548 36694 10560
rect 36725 10557 36737 10560
rect 36771 10588 36783 10591
rect 38580 10588 38608 10619
rect 39482 10616 39488 10668
rect 39540 10656 39546 10668
rect 39761 10659 39819 10665
rect 39761 10656 39773 10659
rect 39540 10628 39773 10656
rect 39540 10616 39546 10628
rect 39761 10625 39773 10628
rect 39807 10625 39819 10659
rect 39761 10619 39819 10625
rect 46934 10616 46940 10668
rect 46992 10656 46998 10668
rect 47949 10659 48007 10665
rect 47949 10656 47961 10659
rect 46992 10628 47961 10656
rect 46992 10616 46998 10628
rect 47949 10625 47961 10628
rect 47995 10625 48007 10659
rect 47949 10619 48007 10625
rect 36771 10560 38608 10588
rect 39945 10591 40003 10597
rect 36771 10557 36783 10560
rect 36725 10551 36783 10557
rect 39945 10557 39957 10591
rect 39991 10588 40003 10591
rect 47026 10588 47032 10600
rect 39991 10560 47032 10588
rect 39991 10557 40003 10560
rect 39945 10551 40003 10557
rect 47026 10548 47032 10560
rect 47084 10548 47090 10600
rect 31726 10492 32904 10520
rect 33244 10492 33916 10520
rect 35529 10523 35587 10529
rect 29457 10455 29515 10461
rect 29457 10421 29469 10455
rect 29503 10452 29515 10455
rect 31386 10452 31392 10464
rect 29503 10424 31392 10452
rect 29503 10421 29515 10424
rect 29457 10415 29515 10421
rect 31386 10412 31392 10424
rect 31444 10412 31450 10464
rect 31478 10412 31484 10464
rect 31536 10452 31542 10464
rect 31726 10452 31754 10492
rect 31536 10424 31754 10452
rect 32309 10455 32367 10461
rect 31536 10412 31542 10424
rect 32309 10421 32321 10455
rect 32355 10452 32367 10455
rect 33244 10452 33272 10492
rect 35529 10489 35541 10523
rect 35575 10520 35587 10523
rect 35894 10520 35900 10532
rect 35575 10492 35900 10520
rect 35575 10489 35587 10492
rect 35529 10483 35587 10489
rect 32355 10424 33272 10452
rect 32355 10421 32367 10424
rect 32309 10415 32367 10421
rect 33410 10412 33416 10464
rect 33468 10452 33474 10464
rect 35544 10452 35572 10483
rect 35894 10480 35900 10492
rect 35952 10480 35958 10532
rect 36081 10523 36139 10529
rect 36081 10489 36093 10523
rect 36127 10520 36139 10523
rect 40034 10520 40040 10532
rect 36127 10492 40040 10520
rect 36127 10489 36139 10492
rect 36081 10483 36139 10489
rect 40034 10480 40040 10492
rect 40092 10480 40098 10532
rect 33468 10424 35572 10452
rect 33468 10412 33474 10424
rect 36538 10412 36544 10464
rect 36596 10452 36602 10464
rect 38105 10455 38163 10461
rect 38105 10452 38117 10455
rect 36596 10424 38117 10452
rect 36596 10412 36602 10424
rect 38105 10421 38117 10424
rect 38151 10421 38163 10455
rect 38105 10415 38163 10421
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 12529 10251 12587 10257
rect 12529 10217 12541 10251
rect 12575 10248 12587 10251
rect 12618 10248 12624 10260
rect 12575 10220 12624 10248
rect 12575 10217 12587 10220
rect 12529 10211 12587 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 12989 10251 13047 10257
rect 12989 10248 13001 10251
rect 12860 10220 13001 10248
rect 12860 10208 12866 10220
rect 12989 10217 13001 10220
rect 13035 10217 13047 10251
rect 12989 10211 13047 10217
rect 13262 10208 13268 10260
rect 13320 10248 13326 10260
rect 16482 10248 16488 10260
rect 13320 10220 16488 10248
rect 13320 10208 13326 10220
rect 16482 10208 16488 10220
rect 16540 10208 16546 10260
rect 16666 10208 16672 10260
rect 16724 10248 16730 10260
rect 17218 10248 17224 10260
rect 16724 10220 17224 10248
rect 16724 10208 16730 10220
rect 17218 10208 17224 10220
rect 17276 10248 17282 10260
rect 18509 10251 18567 10257
rect 18509 10248 18521 10251
rect 17276 10220 18521 10248
rect 17276 10208 17282 10220
rect 18509 10217 18521 10220
rect 18555 10248 18567 10251
rect 18966 10248 18972 10260
rect 18555 10220 18972 10248
rect 18555 10217 18567 10220
rect 18509 10211 18567 10217
rect 18966 10208 18972 10220
rect 19024 10208 19030 10260
rect 19337 10251 19395 10257
rect 19337 10217 19349 10251
rect 19383 10248 19395 10251
rect 19426 10248 19432 10260
rect 19383 10220 19432 10248
rect 19383 10217 19395 10220
rect 19337 10211 19395 10217
rect 19426 10208 19432 10220
rect 19484 10248 19490 10260
rect 22554 10248 22560 10260
rect 19484 10220 22560 10248
rect 19484 10208 19490 10220
rect 22554 10208 22560 10220
rect 22612 10208 22618 10260
rect 24844 10251 24902 10257
rect 24844 10217 24856 10251
rect 24890 10248 24902 10251
rect 26602 10248 26608 10260
rect 24890 10220 26608 10248
rect 24890 10217 24902 10220
rect 24844 10211 24902 10217
rect 26602 10208 26608 10220
rect 26660 10208 26666 10260
rect 26694 10208 26700 10260
rect 26752 10208 26758 10260
rect 27246 10208 27252 10260
rect 27304 10248 27310 10260
rect 27304 10220 28672 10248
rect 27304 10208 27310 10220
rect 19061 10183 19119 10189
rect 19061 10149 19073 10183
rect 19107 10180 19119 10183
rect 19794 10180 19800 10192
rect 19107 10152 19800 10180
rect 19107 10149 19119 10152
rect 19061 10143 19119 10149
rect 19794 10140 19800 10152
rect 19852 10140 19858 10192
rect 21726 10140 21732 10192
rect 21784 10180 21790 10192
rect 22097 10183 22155 10189
rect 22097 10180 22109 10183
rect 21784 10152 22109 10180
rect 21784 10140 21790 10152
rect 22097 10149 22109 10152
rect 22143 10149 22155 10183
rect 22097 10143 22155 10149
rect 1854 10072 1860 10124
rect 1912 10072 1918 10124
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 12526 10112 12532 10124
rect 10468 10084 12532 10112
rect 10468 10072 10474 10084
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 13538 10072 13544 10124
rect 13596 10072 13602 10124
rect 14274 10072 14280 10124
rect 14332 10072 14338 10124
rect 14553 10115 14611 10121
rect 14553 10081 14565 10115
rect 14599 10112 14611 10115
rect 16298 10112 16304 10124
rect 14599 10084 16304 10112
rect 14599 10081 14611 10084
rect 14553 10075 14611 10081
rect 16298 10072 16304 10084
rect 16356 10072 16362 10124
rect 17037 10115 17095 10121
rect 17037 10081 17049 10115
rect 17083 10112 17095 10115
rect 18506 10112 18512 10124
rect 17083 10084 18512 10112
rect 17083 10081 17095 10084
rect 17037 10075 17095 10081
rect 18506 10072 18512 10084
rect 18564 10112 18570 10124
rect 18874 10112 18880 10124
rect 18564 10084 18880 10112
rect 18564 10072 18570 10084
rect 18874 10072 18880 10084
rect 18932 10072 18938 10124
rect 19518 10072 19524 10124
rect 19576 10112 19582 10124
rect 19613 10115 19671 10121
rect 19613 10112 19625 10115
rect 19576 10084 19625 10112
rect 19576 10072 19582 10084
rect 19613 10081 19625 10084
rect 19659 10081 19671 10115
rect 19613 10075 19671 10081
rect 20349 10115 20407 10121
rect 20349 10081 20361 10115
rect 20395 10112 20407 10115
rect 20622 10112 20628 10124
rect 20395 10084 20628 10112
rect 20395 10081 20407 10084
rect 20349 10075 20407 10081
rect 20622 10072 20628 10084
rect 20680 10112 20686 10124
rect 22002 10112 22008 10124
rect 20680 10084 22008 10112
rect 20680 10072 20686 10084
rect 22002 10072 22008 10084
rect 22060 10112 22066 10124
rect 23290 10112 23296 10124
rect 22060 10084 23296 10112
rect 22060 10072 22066 10084
rect 23290 10072 23296 10084
rect 23348 10072 23354 10124
rect 24581 10115 24639 10121
rect 24581 10081 24593 10115
rect 24627 10112 24639 10115
rect 27249 10115 27307 10121
rect 24627 10084 27016 10112
rect 24627 10081 24639 10084
rect 24581 10075 24639 10081
rect 26988 10056 27016 10084
rect 27249 10081 27261 10115
rect 27295 10112 27307 10115
rect 27614 10112 27620 10124
rect 27295 10084 27620 10112
rect 27295 10081 27307 10084
rect 27249 10075 27307 10081
rect 27614 10072 27620 10084
rect 27672 10072 27678 10124
rect 28644 10112 28672 10220
rect 29362 10208 29368 10260
rect 29420 10208 29426 10260
rect 31754 10208 31760 10260
rect 31812 10248 31818 10260
rect 32125 10251 32183 10257
rect 32125 10248 32137 10251
rect 31812 10220 32137 10248
rect 31812 10208 31818 10220
rect 32125 10217 32137 10220
rect 32171 10217 32183 10251
rect 32125 10211 32183 10217
rect 32490 10208 32496 10260
rect 32548 10248 32554 10260
rect 36538 10248 36544 10260
rect 32548 10220 36544 10248
rect 32548 10208 32554 10220
rect 36538 10208 36544 10220
rect 36596 10208 36602 10260
rect 36630 10208 36636 10260
rect 36688 10208 36694 10260
rect 28721 10183 28779 10189
rect 28721 10149 28733 10183
rect 28767 10180 28779 10183
rect 28810 10180 28816 10192
rect 28767 10152 28816 10180
rect 28767 10149 28779 10152
rect 28721 10143 28779 10149
rect 28810 10140 28816 10152
rect 28868 10180 28874 10192
rect 29822 10180 29828 10192
rect 28868 10152 29828 10180
rect 28868 10140 28874 10152
rect 29822 10140 29828 10152
rect 29880 10180 29886 10192
rect 30190 10180 30196 10192
rect 29880 10152 30196 10180
rect 29880 10140 29886 10152
rect 30190 10140 30196 10152
rect 30248 10140 30254 10192
rect 33321 10183 33379 10189
rect 33321 10149 33333 10183
rect 33367 10180 33379 10183
rect 34790 10180 34796 10192
rect 33367 10152 34796 10180
rect 33367 10149 33379 10152
rect 33321 10143 33379 10149
rect 34790 10140 34796 10152
rect 34848 10140 34854 10192
rect 38473 10183 38531 10189
rect 38473 10149 38485 10183
rect 38519 10180 38531 10183
rect 46934 10180 46940 10192
rect 38519 10152 46940 10180
rect 38519 10149 38531 10152
rect 38473 10143 38531 10149
rect 46934 10140 46940 10152
rect 46992 10140 46998 10192
rect 29733 10115 29791 10121
rect 28644 10084 29684 10112
rect 1302 10004 1308 10056
rect 1360 10044 1366 10056
rect 1581 10047 1639 10053
rect 1581 10044 1593 10047
rect 1360 10016 1593 10044
rect 1360 10004 1366 10016
rect 1581 10013 1593 10016
rect 1627 10013 1639 10047
rect 1581 10007 1639 10013
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10044 11943 10047
rect 13354 10044 13360 10056
rect 11931 10016 13360 10044
rect 11931 10013 11943 10016
rect 11885 10007 11943 10013
rect 13354 10004 13360 10016
rect 13412 10004 13418 10056
rect 16758 10004 16764 10056
rect 16816 10004 16822 10056
rect 18598 10004 18604 10056
rect 18656 10044 18662 10056
rect 18785 10047 18843 10053
rect 18785 10044 18797 10047
rect 18656 10016 18797 10044
rect 18656 10004 18662 10016
rect 18785 10013 18797 10016
rect 18831 10013 18843 10047
rect 22830 10044 22836 10056
rect 18785 10007 18843 10013
rect 21928 10016 22836 10044
rect 11422 9936 11428 9988
rect 11480 9976 11486 9988
rect 14090 9976 14096 9988
rect 11480 9948 14096 9976
rect 11480 9936 11486 9948
rect 14090 9936 14096 9948
rect 14148 9936 14154 9988
rect 15286 9936 15292 9988
rect 15344 9936 15350 9988
rect 16301 9979 16359 9985
rect 16301 9945 16313 9979
rect 16347 9976 16359 9979
rect 16390 9976 16396 9988
rect 16347 9948 16396 9976
rect 16347 9945 16359 9948
rect 16301 9939 16359 9945
rect 16390 9936 16396 9948
rect 16448 9936 16454 9988
rect 16482 9936 16488 9988
rect 16540 9976 16546 9988
rect 17494 9976 17500 9988
rect 16540 9948 17500 9976
rect 16540 9936 16546 9948
rect 17494 9936 17500 9948
rect 17552 9936 17558 9988
rect 20612 9979 20670 9985
rect 20612 9945 20624 9979
rect 20658 9945 20670 9979
rect 20612 9939 20670 9945
rect 11238 9868 11244 9920
rect 11296 9908 11302 9920
rect 13262 9908 13268 9920
rect 11296 9880 13268 9908
rect 11296 9868 11302 9880
rect 13262 9868 13268 9880
rect 13320 9908 13326 9920
rect 13357 9911 13415 9917
rect 13357 9908 13369 9911
rect 13320 9880 13369 9908
rect 13320 9868 13326 9880
rect 13357 9877 13369 9880
rect 13403 9877 13415 9911
rect 13357 9871 13415 9877
rect 13449 9911 13507 9917
rect 13449 9877 13461 9911
rect 13495 9908 13507 9911
rect 19334 9908 19340 9920
rect 13495 9880 19340 9908
rect 13495 9877 13507 9880
rect 13449 9871 13507 9877
rect 19334 9868 19340 9880
rect 19392 9868 19398 9920
rect 20627 9908 20655 9939
rect 21082 9936 21088 9988
rect 21140 9936 21146 9988
rect 21358 9908 21364 9920
rect 20627 9880 21364 9908
rect 21358 9868 21364 9880
rect 21416 9868 21422 9920
rect 21450 9868 21456 9920
rect 21508 9908 21514 9920
rect 21928 9908 21956 10016
rect 22830 10004 22836 10016
rect 22888 10004 22894 10056
rect 25958 10004 25964 10056
rect 26016 10004 26022 10056
rect 26970 10004 26976 10056
rect 27028 10004 27034 10056
rect 28534 10044 28540 10056
rect 28382 10016 28540 10044
rect 28534 10004 28540 10016
rect 28592 10044 28598 10056
rect 29089 10047 29147 10053
rect 29089 10044 29101 10047
rect 28592 10016 29101 10044
rect 28592 10004 28598 10016
rect 29089 10013 29101 10016
rect 29135 10044 29147 10047
rect 29362 10044 29368 10056
rect 29135 10016 29368 10044
rect 29135 10013 29147 10016
rect 29089 10007 29147 10013
rect 29362 10004 29368 10016
rect 29420 10004 29426 10056
rect 22554 9936 22560 9988
rect 22612 9976 22618 9988
rect 24118 9976 24124 9988
rect 22612 9948 24124 9976
rect 22612 9936 22618 9948
rect 24118 9936 24124 9948
rect 24176 9936 24182 9988
rect 29656 9976 29684 10084
rect 29733 10081 29745 10115
rect 29779 10112 29791 10115
rect 31294 10112 31300 10124
rect 29779 10084 31300 10112
rect 29779 10081 29791 10084
rect 29733 10075 29791 10081
rect 31294 10072 31300 10084
rect 31352 10072 31358 10124
rect 31386 10072 31392 10124
rect 31444 10112 31450 10124
rect 33410 10112 33416 10124
rect 31444 10084 33416 10112
rect 31444 10072 31450 10084
rect 33410 10072 33416 10084
rect 33468 10072 33474 10124
rect 33965 10115 34023 10121
rect 33965 10081 33977 10115
rect 34011 10112 34023 10115
rect 34330 10112 34336 10124
rect 34011 10084 34336 10112
rect 34011 10081 34023 10084
rect 33965 10075 34023 10081
rect 34330 10072 34336 10084
rect 34388 10072 34394 10124
rect 34422 10072 34428 10124
rect 34480 10072 34486 10124
rect 35161 10115 35219 10121
rect 35161 10081 35173 10115
rect 35207 10112 35219 10115
rect 37737 10115 37795 10121
rect 37737 10112 37749 10115
rect 35207 10084 37749 10112
rect 35207 10081 35219 10084
rect 35161 10075 35219 10081
rect 37737 10081 37749 10084
rect 37783 10081 37795 10115
rect 37737 10075 37795 10081
rect 39482 10072 39488 10124
rect 39540 10072 39546 10124
rect 40313 10115 40371 10121
rect 40313 10081 40325 10115
rect 40359 10112 40371 10115
rect 45830 10112 45836 10124
rect 40359 10084 45836 10112
rect 40359 10081 40371 10084
rect 40313 10075 40371 10081
rect 45830 10072 45836 10084
rect 45888 10072 45894 10124
rect 49142 10072 49148 10124
rect 49200 10072 49206 10124
rect 30374 10004 30380 10056
rect 30432 10004 30438 10056
rect 32585 10047 32643 10053
rect 32585 10013 32597 10047
rect 32631 10044 32643 10047
rect 33318 10044 33324 10056
rect 32631 10016 33324 10044
rect 32631 10013 32643 10016
rect 32585 10007 32643 10013
rect 33318 10004 33324 10016
rect 33376 10004 33382 10056
rect 33686 10044 33692 10056
rect 33428 10016 33692 10044
rect 30558 9976 30564 9988
rect 28552 9948 29132 9976
rect 29656 9948 30564 9976
rect 21508 9880 21956 9908
rect 21508 9868 21514 9880
rect 22002 9868 22008 9920
rect 22060 9908 22066 9920
rect 23845 9911 23903 9917
rect 23845 9908 23857 9911
rect 22060 9880 23857 9908
rect 22060 9868 22066 9880
rect 23845 9877 23857 9880
rect 23891 9877 23903 9911
rect 23845 9871 23903 9877
rect 24026 9868 24032 9920
rect 24084 9868 24090 9920
rect 24946 9868 24952 9920
rect 25004 9908 25010 9920
rect 26329 9911 26387 9917
rect 26329 9908 26341 9911
rect 25004 9880 26341 9908
rect 25004 9868 25010 9880
rect 26329 9877 26341 9880
rect 26375 9877 26387 9911
rect 26329 9871 26387 9877
rect 26418 9868 26424 9920
rect 26476 9908 26482 9920
rect 28552 9908 28580 9948
rect 26476 9880 28580 9908
rect 29104 9908 29132 9948
rect 30558 9936 30564 9948
rect 30616 9936 30622 9988
rect 30650 9936 30656 9988
rect 30708 9936 30714 9988
rect 32306 9976 32312 9988
rect 31878 9948 32312 9976
rect 32306 9936 32312 9948
rect 32364 9936 32370 9988
rect 33428 9908 33456 10016
rect 33686 10004 33692 10016
rect 33744 10004 33750 10056
rect 33778 10004 33784 10056
rect 33836 10044 33842 10056
rect 34882 10044 34888 10056
rect 33836 10016 34888 10044
rect 33836 10004 33842 10016
rect 34882 10004 34888 10016
rect 34940 10004 34946 10056
rect 37093 10047 37151 10053
rect 37093 10013 37105 10047
rect 37139 10013 37151 10047
rect 37093 10007 37151 10013
rect 33502 9936 33508 9988
rect 33560 9976 33566 9988
rect 36538 9976 36544 9988
rect 33560 9948 33824 9976
rect 36386 9948 36544 9976
rect 33560 9936 33566 9948
rect 33796 9917 33824 9948
rect 36538 9936 36544 9948
rect 36596 9936 36602 9988
rect 29104 9880 33456 9908
rect 33781 9911 33839 9917
rect 26476 9868 26482 9880
rect 33781 9877 33793 9911
rect 33827 9908 33839 9911
rect 34238 9908 34244 9920
rect 33827 9880 34244 9908
rect 33827 9877 33839 9880
rect 33781 9871 33839 9877
rect 34238 9868 34244 9880
rect 34296 9868 34302 9920
rect 35434 9868 35440 9920
rect 35492 9908 35498 9920
rect 37108 9908 37136 10007
rect 39298 10004 39304 10056
rect 39356 10044 39362 10056
rect 39356 10016 42196 10044
rect 39356 10004 39362 10016
rect 38286 9936 38292 9988
rect 38344 9976 38350 9988
rect 38749 9979 38807 9985
rect 38749 9976 38761 9979
rect 38344 9948 38761 9976
rect 38344 9936 38350 9948
rect 38749 9945 38761 9948
rect 38795 9945 38807 9979
rect 38749 9939 38807 9945
rect 40129 9979 40187 9985
rect 40129 9945 40141 9979
rect 40175 9976 40187 9979
rect 40310 9976 40316 9988
rect 40175 9948 40316 9976
rect 40175 9945 40187 9948
rect 40129 9939 40187 9945
rect 40310 9936 40316 9948
rect 40368 9976 40374 9988
rect 40589 9979 40647 9985
rect 40589 9976 40601 9979
rect 40368 9948 40601 9976
rect 40368 9936 40374 9948
rect 40589 9945 40601 9948
rect 40635 9945 40647 9979
rect 42168 9976 42196 10016
rect 44174 10004 44180 10056
rect 44232 10044 44238 10056
rect 46109 10047 46167 10053
rect 46109 10044 46121 10047
rect 44232 10016 46121 10044
rect 44232 10004 44238 10016
rect 46109 10013 46121 10016
rect 46155 10013 46167 10047
rect 46109 10007 46167 10013
rect 46658 10004 46664 10056
rect 46716 10044 46722 10056
rect 47949 10047 48007 10053
rect 47949 10044 47961 10047
rect 46716 10016 47961 10044
rect 46716 10004 46722 10016
rect 47949 10013 47961 10016
rect 47995 10013 48007 10047
rect 47949 10007 48007 10013
rect 44361 9979 44419 9985
rect 44361 9976 44373 9979
rect 42168 9948 44373 9976
rect 40589 9939 40647 9945
rect 44361 9945 44373 9948
rect 44407 9945 44419 9979
rect 44361 9939 44419 9945
rect 44545 9979 44603 9985
rect 44545 9945 44557 9979
rect 44591 9976 44603 9979
rect 46750 9976 46756 9988
rect 44591 9948 46756 9976
rect 44591 9945 44603 9948
rect 44545 9939 44603 9945
rect 46750 9936 46756 9948
rect 46808 9936 46814 9988
rect 47302 9936 47308 9988
rect 47360 9936 47366 9988
rect 35492 9880 37136 9908
rect 35492 9868 35498 9880
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 1302 9664 1308 9716
rect 1360 9704 1366 9716
rect 2133 9707 2191 9713
rect 2133 9704 2145 9707
rect 1360 9676 2145 9704
rect 1360 9664 1366 9676
rect 2133 9673 2145 9676
rect 2179 9673 2191 9707
rect 2133 9667 2191 9673
rect 13814 9664 13820 9716
rect 13872 9704 13878 9716
rect 15381 9707 15439 9713
rect 15381 9704 15393 9707
rect 13872 9676 15393 9704
rect 13872 9664 13878 9676
rect 15381 9673 15393 9676
rect 15427 9673 15439 9707
rect 15381 9667 15439 9673
rect 16206 9664 16212 9716
rect 16264 9704 16270 9716
rect 19058 9704 19064 9716
rect 16264 9676 19064 9704
rect 16264 9664 16270 9676
rect 19058 9664 19064 9676
rect 19116 9664 19122 9716
rect 20438 9664 20444 9716
rect 20496 9704 20502 9716
rect 21082 9704 21088 9716
rect 20496 9676 21088 9704
rect 20496 9664 20502 9676
rect 21082 9664 21088 9676
rect 21140 9664 21146 9716
rect 22005 9707 22063 9713
rect 22005 9673 22017 9707
rect 22051 9673 22063 9707
rect 22005 9667 22063 9673
rect 12710 9596 12716 9648
rect 12768 9636 12774 9648
rect 12805 9639 12863 9645
rect 12805 9636 12817 9639
rect 12768 9608 12817 9636
rect 12768 9596 12774 9608
rect 12805 9605 12817 9608
rect 12851 9605 12863 9639
rect 13998 9636 14004 9648
rect 12805 9599 12863 9605
rect 13556 9608 14004 9636
rect 1302 9528 1308 9580
rect 1360 9568 1366 9580
rect 1673 9571 1731 9577
rect 1673 9568 1685 9571
rect 1360 9540 1685 9568
rect 1360 9528 1366 9540
rect 1673 9537 1685 9540
rect 1719 9568 1731 9571
rect 2317 9571 2375 9577
rect 2317 9568 2329 9571
rect 1719 9540 2329 9568
rect 1719 9537 1731 9540
rect 1673 9531 1731 9537
rect 2317 9537 2329 9540
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 12526 9528 12532 9580
rect 12584 9568 12590 9580
rect 12897 9571 12955 9577
rect 12897 9568 12909 9571
rect 12584 9540 12909 9568
rect 12584 9528 12590 9540
rect 12897 9537 12909 9540
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 1854 9460 1860 9512
rect 1912 9460 1918 9512
rect 13081 9503 13139 9509
rect 13081 9469 13093 9503
rect 13127 9500 13139 9503
rect 13354 9500 13360 9512
rect 13127 9472 13360 9500
rect 13127 9469 13139 9472
rect 13081 9463 13139 9469
rect 13354 9460 13360 9472
rect 13412 9460 13418 9512
rect 12437 9435 12495 9441
rect 12437 9401 12449 9435
rect 12483 9432 12495 9435
rect 13556 9432 13584 9608
rect 13998 9596 14004 9608
rect 14056 9596 14062 9648
rect 15194 9636 15200 9648
rect 15134 9608 15200 9636
rect 15194 9596 15200 9608
rect 15252 9596 15258 9648
rect 15838 9596 15844 9648
rect 15896 9596 15902 9648
rect 16117 9639 16175 9645
rect 16117 9605 16129 9639
rect 16163 9636 16175 9639
rect 16574 9636 16580 9648
rect 16163 9608 16580 9636
rect 16163 9605 16175 9608
rect 16117 9599 16175 9605
rect 16574 9596 16580 9608
rect 16632 9596 16638 9648
rect 17586 9596 17592 9648
rect 17644 9596 17650 9648
rect 20346 9596 20352 9648
rect 20404 9596 20410 9648
rect 21082 9528 21088 9580
rect 21140 9568 21146 9580
rect 21818 9568 21824 9580
rect 21140 9540 21824 9568
rect 21140 9528 21146 9540
rect 21818 9528 21824 9540
rect 21876 9528 21882 9580
rect 21910 9528 21916 9580
rect 21968 9568 21974 9580
rect 22020 9568 22048 9667
rect 23382 9664 23388 9716
rect 23440 9704 23446 9716
rect 26418 9704 26424 9716
rect 23440 9676 26424 9704
rect 23440 9664 23446 9676
rect 26418 9664 26424 9676
rect 26476 9664 26482 9716
rect 26970 9664 26976 9716
rect 27028 9704 27034 9716
rect 27028 9676 27568 9704
rect 27028 9664 27034 9676
rect 23106 9596 23112 9648
rect 23164 9596 23170 9648
rect 23750 9596 23756 9648
rect 23808 9636 23814 9648
rect 23808 9608 24334 9636
rect 23808 9596 23814 9608
rect 26050 9596 26056 9648
rect 26108 9636 26114 9648
rect 26237 9639 26295 9645
rect 26237 9636 26249 9639
rect 26108 9608 26249 9636
rect 26108 9596 26114 9608
rect 26237 9605 26249 9608
rect 26283 9605 26295 9639
rect 26237 9599 26295 9605
rect 21968 9540 22048 9568
rect 21968 9528 21974 9540
rect 22370 9528 22376 9580
rect 22428 9528 22434 9580
rect 23290 9528 23296 9580
rect 23348 9568 23354 9580
rect 23569 9571 23627 9577
rect 23569 9568 23581 9571
rect 23348 9540 23581 9568
rect 23348 9528 23354 9540
rect 23569 9537 23581 9540
rect 23615 9537 23627 9571
rect 23569 9531 23627 9537
rect 26142 9528 26148 9580
rect 26200 9528 26206 9580
rect 13633 9503 13691 9509
rect 13633 9469 13645 9503
rect 13679 9469 13691 9503
rect 13633 9463 13691 9469
rect 12483 9404 13584 9432
rect 12483 9401 12495 9404
rect 12437 9395 12495 9401
rect 11238 9324 11244 9376
rect 11296 9364 11302 9376
rect 12069 9367 12127 9373
rect 12069 9364 12081 9367
rect 11296 9336 12081 9364
rect 11296 9324 11302 9336
rect 12069 9333 12081 9336
rect 12115 9333 12127 9367
rect 13648 9364 13676 9463
rect 13906 9460 13912 9512
rect 13964 9460 13970 9512
rect 16850 9460 16856 9512
rect 16908 9460 16914 9512
rect 17126 9460 17132 9512
rect 17184 9460 17190 9512
rect 17678 9460 17684 9512
rect 17736 9500 17742 9512
rect 18877 9503 18935 9509
rect 18877 9500 18889 9503
rect 17736 9472 18889 9500
rect 17736 9460 17742 9472
rect 18877 9469 18889 9472
rect 18923 9469 18935 9503
rect 18877 9463 18935 9469
rect 19337 9503 19395 9509
rect 19337 9469 19349 9503
rect 19383 9469 19395 9503
rect 19337 9463 19395 9469
rect 14274 9364 14280 9376
rect 13648 9336 14280 9364
rect 12069 9327 12127 9333
rect 14274 9324 14280 9336
rect 14332 9324 14338 9376
rect 16850 9324 16856 9376
rect 16908 9364 16914 9376
rect 17862 9364 17868 9376
rect 16908 9336 17868 9364
rect 16908 9324 16914 9336
rect 17862 9324 17868 9336
rect 17920 9364 17926 9376
rect 19352 9364 19380 9463
rect 19610 9460 19616 9512
rect 19668 9460 19674 9512
rect 19702 9460 19708 9512
rect 19760 9500 19766 9512
rect 22186 9500 22192 9512
rect 19760 9472 22192 9500
rect 19760 9460 19766 9472
rect 22186 9460 22192 9472
rect 22244 9460 22250 9512
rect 22462 9460 22468 9512
rect 22520 9460 22526 9512
rect 22649 9503 22707 9509
rect 22649 9469 22661 9503
rect 22695 9500 22707 9503
rect 23474 9500 23480 9512
rect 22695 9472 23480 9500
rect 22695 9469 22707 9472
rect 22649 9463 22707 9469
rect 23474 9460 23480 9472
rect 23532 9460 23538 9512
rect 23845 9503 23903 9509
rect 23845 9469 23857 9503
rect 23891 9500 23903 9503
rect 25498 9500 25504 9512
rect 23891 9472 25504 9500
rect 23891 9469 23903 9472
rect 23845 9463 23903 9469
rect 25498 9460 25504 9472
rect 25556 9460 25562 9512
rect 26418 9460 26424 9512
rect 26476 9460 26482 9512
rect 27540 9509 27568 9676
rect 29270 9664 29276 9716
rect 29328 9704 29334 9716
rect 34330 9704 34336 9716
rect 29328 9676 31754 9704
rect 29328 9664 29334 9676
rect 30282 9636 30288 9648
rect 29748 9608 30288 9636
rect 29270 9568 29276 9580
rect 28934 9540 29276 9568
rect 29270 9528 29276 9540
rect 29328 9528 29334 9580
rect 27525 9503 27583 9509
rect 27525 9469 27537 9503
rect 27571 9469 27583 9503
rect 27525 9463 27583 9469
rect 27801 9503 27859 9509
rect 27801 9469 27813 9503
rect 27847 9500 27859 9503
rect 27847 9472 29040 9500
rect 27847 9469 27859 9472
rect 27801 9463 27859 9469
rect 21453 9435 21511 9441
rect 21453 9401 21465 9435
rect 21499 9432 21511 9435
rect 25777 9435 25835 9441
rect 21499 9404 21956 9432
rect 21499 9401 21511 9404
rect 21453 9395 21511 9401
rect 17920 9336 19380 9364
rect 21085 9367 21143 9373
rect 17920 9324 17926 9336
rect 21085 9333 21097 9367
rect 21131 9364 21143 9367
rect 21174 9364 21180 9376
rect 21131 9336 21180 9364
rect 21131 9333 21143 9336
rect 21085 9327 21143 9333
rect 21174 9324 21180 9336
rect 21232 9324 21238 9376
rect 21266 9324 21272 9376
rect 21324 9364 21330 9376
rect 21637 9367 21695 9373
rect 21637 9364 21649 9367
rect 21324 9336 21649 9364
rect 21324 9324 21330 9336
rect 21637 9333 21649 9336
rect 21683 9364 21695 9367
rect 21818 9364 21824 9376
rect 21683 9336 21824 9364
rect 21683 9333 21695 9336
rect 21637 9327 21695 9333
rect 21818 9324 21824 9336
rect 21876 9324 21882 9376
rect 21928 9364 21956 9404
rect 25777 9401 25789 9435
rect 25823 9432 25835 9435
rect 27430 9432 27436 9444
rect 25823 9404 27436 9432
rect 25823 9401 25835 9404
rect 25777 9395 25835 9401
rect 27430 9392 27436 9404
rect 27488 9392 27494 9444
rect 22554 9364 22560 9376
rect 21928 9336 22560 9364
rect 22554 9324 22560 9336
rect 22612 9324 22618 9376
rect 23842 9324 23848 9376
rect 23900 9364 23906 9376
rect 25317 9367 25375 9373
rect 25317 9364 25329 9367
rect 23900 9336 25329 9364
rect 23900 9324 23906 9336
rect 25317 9333 25329 9336
rect 25363 9333 25375 9367
rect 25317 9327 25375 9333
rect 27062 9324 27068 9376
rect 27120 9324 27126 9376
rect 27246 9324 27252 9376
rect 27304 9324 27310 9376
rect 27540 9364 27568 9463
rect 29012 9432 29040 9472
rect 29086 9460 29092 9512
rect 29144 9500 29150 9512
rect 29748 9509 29776 9608
rect 30282 9596 30288 9608
rect 30340 9596 30346 9648
rect 31726 9636 31754 9676
rect 34164 9676 34336 9704
rect 34164 9645 34192 9676
rect 34330 9664 34336 9676
rect 34388 9664 34394 9716
rect 34974 9664 34980 9716
rect 35032 9704 35038 9716
rect 35434 9704 35440 9716
rect 35032 9676 35440 9704
rect 35032 9664 35038 9676
rect 35434 9664 35440 9676
rect 35492 9704 35498 9716
rect 35621 9707 35679 9713
rect 35621 9704 35633 9707
rect 35492 9676 35633 9704
rect 35492 9664 35498 9676
rect 35621 9673 35633 9676
rect 35667 9673 35679 9707
rect 35621 9667 35679 9673
rect 37274 9664 37280 9716
rect 37332 9664 37338 9716
rect 32953 9639 33011 9645
rect 32953 9636 32965 9639
rect 31726 9608 32965 9636
rect 32953 9605 32965 9608
rect 32999 9605 33011 9639
rect 34149 9639 34207 9645
rect 34149 9636 34161 9639
rect 32953 9599 33011 9605
rect 33796 9608 34161 9636
rect 31849 9571 31907 9577
rect 31849 9568 31861 9571
rect 31142 9540 31861 9568
rect 31849 9537 31861 9540
rect 31895 9568 31907 9571
rect 32306 9568 32312 9580
rect 31895 9540 32312 9568
rect 31895 9537 31907 9540
rect 31849 9531 31907 9537
rect 32306 9528 32312 9540
rect 32364 9528 32370 9580
rect 32398 9528 32404 9580
rect 32456 9568 32462 9580
rect 33045 9571 33103 9577
rect 33045 9568 33057 9571
rect 32456 9540 33057 9568
rect 32456 9528 32462 9540
rect 33045 9537 33057 9540
rect 33091 9537 33103 9571
rect 33045 9531 33103 9537
rect 29733 9503 29791 9509
rect 29733 9500 29745 9503
rect 29144 9472 29745 9500
rect 29144 9460 29150 9472
rect 29733 9469 29745 9472
rect 29779 9469 29791 9503
rect 29733 9463 29791 9469
rect 30006 9460 30012 9512
rect 30064 9460 30070 9512
rect 32214 9460 32220 9512
rect 32272 9500 32278 9512
rect 33137 9503 33195 9509
rect 33137 9500 33149 9503
rect 32272 9472 33149 9500
rect 32272 9460 32278 9472
rect 33137 9469 33149 9472
rect 33183 9469 33195 9503
rect 33137 9463 33195 9469
rect 29546 9432 29552 9444
rect 29012 9404 29552 9432
rect 29546 9392 29552 9404
rect 29604 9392 29610 9444
rect 31662 9392 31668 9444
rect 31720 9432 31726 9444
rect 33796 9432 33824 9608
rect 34149 9605 34161 9608
rect 34195 9605 34207 9639
rect 35710 9636 35716 9648
rect 35374 9608 35716 9636
rect 34149 9599 34207 9605
rect 35710 9596 35716 9608
rect 35768 9636 35774 9648
rect 36538 9636 36544 9648
rect 35768 9608 36544 9636
rect 35768 9596 35774 9608
rect 36538 9596 36544 9608
rect 36596 9636 36602 9648
rect 37093 9639 37151 9645
rect 37093 9636 37105 9639
rect 36596 9608 37105 9636
rect 36596 9596 36602 9608
rect 37093 9605 37105 9608
rect 37139 9636 37151 9639
rect 37829 9639 37887 9645
rect 37829 9636 37841 9639
rect 37139 9608 37841 9636
rect 37139 9605 37151 9608
rect 37093 9599 37151 9605
rect 37829 9605 37841 9608
rect 37875 9605 37887 9639
rect 37829 9599 37887 9605
rect 49145 9639 49203 9645
rect 49145 9605 49157 9639
rect 49191 9636 49203 9639
rect 49326 9636 49332 9648
rect 49191 9608 49332 9636
rect 49191 9605 49203 9608
rect 49145 9599 49203 9605
rect 49326 9596 49332 9608
rect 49384 9596 49390 9648
rect 35526 9528 35532 9580
rect 35584 9568 35590 9580
rect 36081 9571 36139 9577
rect 36081 9568 36093 9571
rect 35584 9540 36093 9568
rect 35584 9528 35590 9540
rect 36081 9537 36093 9540
rect 36127 9537 36139 9571
rect 36081 9531 36139 9537
rect 47210 9528 47216 9580
rect 47268 9568 47274 9580
rect 47949 9571 48007 9577
rect 47949 9568 47961 9571
rect 47268 9540 47961 9568
rect 47268 9528 47274 9540
rect 47949 9537 47961 9540
rect 47995 9537 48007 9571
rect 47949 9531 48007 9537
rect 33870 9460 33876 9512
rect 33928 9460 33934 9512
rect 34514 9460 34520 9512
rect 34572 9500 34578 9512
rect 38378 9500 38384 9512
rect 34572 9472 38384 9500
rect 34572 9460 34578 9472
rect 38378 9460 38384 9472
rect 38436 9460 38442 9512
rect 31720 9404 33824 9432
rect 31720 9392 31726 9404
rect 29086 9364 29092 9376
rect 27540 9336 29092 9364
rect 29086 9324 29092 9336
rect 29144 9324 29150 9376
rect 29178 9324 29184 9376
rect 29236 9364 29242 9376
rect 29273 9367 29331 9373
rect 29273 9364 29285 9367
rect 29236 9336 29285 9364
rect 29236 9324 29242 9336
rect 29273 9333 29285 9336
rect 29319 9333 29331 9367
rect 29273 9327 29331 9333
rect 31478 9324 31484 9376
rect 31536 9324 31542 9376
rect 32585 9367 32643 9373
rect 32585 9333 32597 9367
rect 32631 9364 32643 9367
rect 35526 9364 35532 9376
rect 32631 9336 35532 9364
rect 32631 9333 32643 9336
rect 32585 9327 32643 9333
rect 35526 9324 35532 9336
rect 35584 9324 35590 9376
rect 36722 9324 36728 9376
rect 36780 9324 36786 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 12342 9120 12348 9172
rect 12400 9160 12406 9172
rect 12989 9163 13047 9169
rect 12989 9160 13001 9163
rect 12400 9132 13001 9160
rect 12400 9120 12406 9132
rect 12989 9129 13001 9132
rect 13035 9129 13047 9163
rect 13722 9160 13728 9172
rect 12989 9123 13047 9129
rect 13464 9132 13728 9160
rect 2406 8984 2412 9036
rect 2464 9024 2470 9036
rect 11146 9024 11152 9036
rect 2464 8996 11152 9024
rect 2464 8984 2470 8996
rect 11146 8984 11152 8996
rect 11204 8984 11210 9036
rect 13464 9033 13492 9132
rect 13722 9120 13728 9132
rect 13780 9160 13786 9172
rect 13780 9132 18460 9160
rect 13780 9120 13786 9132
rect 18432 9092 18460 9132
rect 18782 9120 18788 9172
rect 18840 9160 18846 9172
rect 18877 9163 18935 9169
rect 18877 9160 18889 9163
rect 18840 9132 18889 9160
rect 18840 9120 18846 9132
rect 18877 9129 18889 9132
rect 18923 9129 18935 9163
rect 19702 9160 19708 9172
rect 18877 9123 18935 9129
rect 18984 9132 19708 9160
rect 18984 9092 19012 9132
rect 19702 9120 19708 9132
rect 19760 9120 19766 9172
rect 19886 9120 19892 9172
rect 19944 9160 19950 9172
rect 19944 9132 20760 9160
rect 19944 9120 19950 9132
rect 18432 9064 19012 9092
rect 20732 9092 20760 9132
rect 20806 9120 20812 9172
rect 20864 9160 20870 9172
rect 21637 9163 21695 9169
rect 21637 9160 21649 9163
rect 20864 9132 21649 9160
rect 20864 9120 20870 9132
rect 21637 9129 21649 9132
rect 21683 9129 21695 9163
rect 21637 9123 21695 9129
rect 22646 9120 22652 9172
rect 22704 9160 22710 9172
rect 23109 9163 23167 9169
rect 23109 9160 23121 9163
rect 22704 9132 23121 9160
rect 22704 9120 22710 9132
rect 23109 9129 23121 9132
rect 23155 9129 23167 9163
rect 23109 9123 23167 9129
rect 23566 9120 23572 9172
rect 23624 9160 23630 9172
rect 24486 9160 24492 9172
rect 23624 9132 24492 9160
rect 23624 9120 23630 9132
rect 24486 9120 24492 9132
rect 24544 9120 24550 9172
rect 24854 9120 24860 9172
rect 24912 9160 24918 9172
rect 25961 9163 26019 9169
rect 25961 9160 25973 9163
rect 24912 9132 25973 9160
rect 24912 9120 24918 9132
rect 25961 9129 25973 9132
rect 26007 9129 26019 9163
rect 25961 9123 26019 9129
rect 27709 9163 27767 9169
rect 27709 9129 27721 9163
rect 27755 9160 27767 9163
rect 27798 9160 27804 9172
rect 27755 9132 27804 9160
rect 27755 9129 27767 9132
rect 27709 9123 27767 9129
rect 27798 9120 27804 9132
rect 27856 9120 27862 9172
rect 28169 9163 28227 9169
rect 28169 9129 28181 9163
rect 28215 9160 28227 9163
rect 29914 9160 29920 9172
rect 28215 9132 29920 9160
rect 28215 9129 28227 9132
rect 28169 9123 28227 9129
rect 29914 9120 29920 9132
rect 29972 9120 29978 9172
rect 30466 9160 30472 9172
rect 30208 9132 30472 9160
rect 21177 9095 21235 9101
rect 21177 9092 21189 9095
rect 20732 9064 21189 9092
rect 21177 9061 21189 9064
rect 21223 9061 21235 9095
rect 21177 9055 21235 9061
rect 21818 9052 21824 9104
rect 21876 9092 21882 9104
rect 21876 9064 22094 9092
rect 21876 9052 21882 9064
rect 13449 9027 13507 9033
rect 13449 8993 13461 9027
rect 13495 8993 13507 9027
rect 13449 8987 13507 8993
rect 13630 8984 13636 9036
rect 13688 8984 13694 9036
rect 14182 8984 14188 9036
rect 14240 9024 14246 9036
rect 22066 9024 22094 9064
rect 22370 9052 22376 9104
rect 22428 9092 22434 9104
rect 30208 9092 30236 9132
rect 30466 9120 30472 9132
rect 30524 9160 30530 9172
rect 32493 9163 32551 9169
rect 32493 9160 32505 9163
rect 30524 9132 32505 9160
rect 30524 9120 30530 9132
rect 32493 9129 32505 9132
rect 32539 9129 32551 9163
rect 32493 9123 32551 9129
rect 32953 9163 33011 9169
rect 32953 9129 32965 9163
rect 32999 9160 33011 9163
rect 34514 9160 34520 9172
rect 32999 9132 34520 9160
rect 32999 9129 33011 9132
rect 32953 9123 33011 9129
rect 34514 9120 34520 9132
rect 34572 9120 34578 9172
rect 34885 9163 34943 9169
rect 34885 9129 34897 9163
rect 34931 9160 34943 9163
rect 36446 9160 36452 9172
rect 34931 9132 36452 9160
rect 34931 9129 34943 9132
rect 34885 9123 34943 9129
rect 36446 9120 36452 9132
rect 36504 9120 36510 9172
rect 36814 9160 36820 9172
rect 36556 9132 36820 9160
rect 22428 9064 26464 9092
rect 22428 9052 22434 9064
rect 22189 9027 22247 9033
rect 22189 9024 22201 9027
rect 14240 8996 21036 9024
rect 22066 8996 22201 9024
rect 14240 8984 14246 8996
rect 1210 8916 1216 8968
rect 1268 8956 1274 8968
rect 2317 8959 2375 8965
rect 2317 8956 2329 8959
rect 1268 8928 2329 8956
rect 1268 8916 1274 8928
rect 2317 8925 2329 8928
rect 2363 8956 2375 8959
rect 2869 8959 2927 8965
rect 2869 8956 2881 8959
rect 2363 8928 2881 8956
rect 2363 8925 2375 8928
rect 2317 8919 2375 8925
rect 2869 8925 2881 8928
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 14274 8916 14280 8968
rect 14332 8916 14338 8968
rect 16669 8959 16727 8965
rect 16669 8956 16681 8959
rect 15856 8928 16681 8956
rect 1302 8848 1308 8900
rect 1360 8888 1366 8900
rect 1673 8891 1731 8897
rect 1673 8888 1685 8891
rect 1360 8860 1685 8888
rect 1360 8848 1366 8860
rect 1673 8857 1685 8860
rect 1719 8888 1731 8891
rect 3053 8891 3111 8897
rect 3053 8888 3065 8891
rect 1719 8860 3065 8888
rect 1719 8857 1731 8860
rect 1673 8851 1731 8857
rect 3053 8857 3065 8860
rect 3099 8857 3111 8891
rect 3053 8851 3111 8857
rect 12434 8848 12440 8900
rect 12492 8888 12498 8900
rect 13357 8891 13415 8897
rect 13357 8888 13369 8891
rect 12492 8860 13369 8888
rect 12492 8848 12498 8860
rect 13357 8857 13369 8860
rect 13403 8857 13415 8891
rect 13357 8851 13415 8857
rect 14550 8848 14556 8900
rect 14608 8848 14614 8900
rect 15194 8848 15200 8900
rect 15252 8848 15258 8900
rect 1762 8780 1768 8832
rect 1820 8780 1826 8832
rect 2498 8780 2504 8832
rect 2556 8780 2562 8832
rect 11974 8780 11980 8832
rect 12032 8820 12038 8832
rect 15856 8820 15884 8928
rect 16669 8925 16681 8928
rect 16715 8925 16727 8959
rect 16669 8919 16727 8925
rect 16850 8916 16856 8968
rect 16908 8956 16914 8968
rect 17129 8959 17187 8965
rect 17129 8956 17141 8959
rect 16908 8928 17141 8956
rect 16908 8916 16914 8928
rect 17129 8925 17141 8928
rect 17175 8925 17187 8959
rect 17129 8919 17187 8925
rect 19426 8916 19432 8968
rect 19484 8916 19490 8968
rect 17402 8848 17408 8900
rect 17460 8848 17466 8900
rect 17604 8860 17894 8888
rect 17604 8832 17632 8860
rect 19702 8848 19708 8900
rect 19760 8848 19766 8900
rect 20438 8848 20444 8900
rect 20496 8848 20502 8900
rect 21008 8888 21036 8996
rect 22189 8993 22201 8996
rect 22235 8993 22247 9027
rect 23753 9027 23811 9033
rect 22189 8987 22247 8993
rect 22296 8996 23704 9024
rect 21542 8916 21548 8968
rect 21600 8956 21606 8968
rect 22097 8959 22155 8965
rect 22097 8956 22109 8959
rect 21600 8928 22109 8956
rect 21600 8916 21606 8928
rect 22097 8925 22109 8928
rect 22143 8925 22155 8959
rect 22097 8919 22155 8925
rect 22296 8888 22324 8996
rect 22370 8916 22376 8968
rect 22428 8956 22434 8968
rect 23474 8956 23480 8968
rect 22428 8928 23480 8956
rect 22428 8916 22434 8928
rect 23474 8916 23480 8928
rect 23532 8916 23538 8968
rect 23566 8916 23572 8968
rect 23624 8916 23630 8968
rect 23676 8956 23704 8996
rect 23753 8993 23765 9027
rect 23799 9024 23811 9027
rect 23842 9024 23848 9036
rect 23799 8996 23848 9024
rect 23799 8993 23811 8996
rect 23753 8987 23811 8993
rect 23842 8984 23848 8996
rect 23900 8984 23906 9036
rect 24118 8984 24124 9036
rect 24176 8984 24182 9036
rect 24578 8984 24584 9036
rect 24636 9024 24642 9036
rect 26436 9033 26464 9064
rect 29012 9064 30236 9092
rect 29012 9036 29040 9064
rect 32030 9052 32036 9104
rect 32088 9092 32094 9104
rect 36556 9092 36584 9132
rect 36814 9120 36820 9132
rect 36872 9120 36878 9172
rect 32088 9064 36584 9092
rect 36633 9095 36691 9101
rect 32088 9052 32094 9064
rect 36633 9061 36645 9095
rect 36679 9092 36691 9095
rect 40034 9092 40040 9104
rect 36679 9064 40040 9092
rect 36679 9061 36691 9064
rect 36633 9055 36691 9061
rect 40034 9052 40040 9064
rect 40092 9052 40098 9104
rect 24673 9027 24731 9033
rect 24673 9024 24685 9027
rect 24636 8996 24685 9024
rect 24636 8984 24642 8996
rect 24673 8993 24685 8996
rect 24719 8993 24731 9027
rect 24673 8987 24731 8993
rect 26421 9027 26479 9033
rect 26421 8993 26433 9027
rect 26467 8993 26479 9027
rect 26421 8987 26479 8993
rect 28813 9027 28871 9033
rect 28813 8993 28825 9027
rect 28859 9024 28871 9027
rect 28994 9024 29000 9036
rect 28859 8996 29000 9024
rect 28859 8993 28871 8996
rect 28813 8987 28871 8993
rect 28994 8984 29000 8996
rect 29052 8984 29058 9036
rect 29733 9027 29791 9033
rect 29733 8993 29745 9027
rect 29779 9024 29791 9027
rect 30098 9024 30104 9036
rect 29779 8996 30104 9024
rect 29779 8993 29791 8996
rect 29733 8987 29791 8993
rect 30098 8984 30104 8996
rect 30156 8984 30162 9036
rect 31021 9027 31079 9033
rect 31021 8993 31033 9027
rect 31067 9024 31079 9027
rect 32858 9024 32864 9036
rect 31067 8996 32864 9024
rect 31067 8993 31079 8996
rect 31021 8987 31079 8993
rect 32858 8984 32864 8996
rect 32916 8984 32922 9036
rect 33594 8984 33600 9036
rect 33652 8984 33658 9036
rect 34057 9027 34115 9033
rect 34057 8993 34069 9027
rect 34103 9024 34115 9027
rect 34606 9024 34612 9036
rect 34103 8996 34612 9024
rect 34103 8993 34115 8996
rect 34057 8987 34115 8993
rect 34606 8984 34612 8996
rect 34664 8984 34670 9036
rect 34790 8984 34796 9036
rect 34848 9024 34854 9036
rect 35345 9027 35403 9033
rect 35345 9024 35357 9027
rect 34848 8996 35357 9024
rect 34848 8984 34854 8996
rect 35345 8993 35357 8996
rect 35391 8993 35403 9027
rect 35345 8987 35403 8993
rect 35434 8984 35440 9036
rect 35492 8984 35498 9036
rect 35526 8984 35532 9036
rect 35584 9024 35590 9036
rect 49145 9027 49203 9033
rect 35584 8996 37872 9024
rect 35584 8984 35590 8996
rect 25317 8959 25375 8965
rect 23676 8928 23796 8956
rect 21008 8860 22324 8888
rect 22554 8848 22560 8900
rect 22612 8888 22618 8900
rect 22741 8891 22799 8897
rect 22741 8888 22753 8891
rect 22612 8860 22753 8888
rect 22612 8848 22618 8860
rect 22741 8857 22753 8860
rect 22787 8888 22799 8891
rect 23658 8888 23664 8900
rect 22787 8860 23664 8888
rect 22787 8857 22799 8860
rect 22741 8851 22799 8857
rect 23658 8848 23664 8860
rect 23716 8848 23722 8900
rect 23768 8888 23796 8928
rect 25317 8925 25329 8959
rect 25363 8956 25375 8959
rect 25590 8956 25596 8968
rect 25363 8928 25596 8956
rect 25363 8925 25375 8928
rect 25317 8919 25375 8925
rect 25590 8916 25596 8928
rect 25648 8916 25654 8968
rect 27065 8959 27123 8965
rect 27065 8925 27077 8959
rect 27111 8956 27123 8959
rect 27154 8956 27160 8968
rect 27111 8928 27160 8956
rect 27111 8925 27123 8928
rect 27065 8919 27123 8925
rect 27154 8916 27160 8928
rect 27212 8916 27218 8968
rect 30377 8959 30435 8965
rect 30377 8956 30389 8959
rect 27724 8928 30389 8956
rect 27246 8888 27252 8900
rect 23768 8860 27252 8888
rect 27246 8848 27252 8860
rect 27304 8848 27310 8900
rect 12032 8792 15884 8820
rect 12032 8780 12038 8792
rect 16022 8780 16028 8832
rect 16080 8780 16086 8832
rect 16482 8780 16488 8832
rect 16540 8780 16546 8832
rect 17586 8780 17592 8832
rect 17644 8780 17650 8832
rect 19058 8780 19064 8832
rect 19116 8820 19122 8832
rect 19886 8820 19892 8832
rect 19116 8792 19892 8820
rect 19116 8780 19122 8792
rect 19886 8780 19892 8792
rect 19944 8780 19950 8832
rect 20070 8780 20076 8832
rect 20128 8820 20134 8832
rect 20990 8820 20996 8832
rect 20128 8792 20996 8820
rect 20128 8780 20134 8792
rect 20990 8780 20996 8792
rect 21048 8780 21054 8832
rect 21266 8780 21272 8832
rect 21324 8820 21330 8832
rect 22005 8823 22063 8829
rect 22005 8820 22017 8823
rect 21324 8792 22017 8820
rect 21324 8780 21330 8792
rect 22005 8789 22017 8792
rect 22051 8820 22063 8823
rect 27724 8820 27752 8928
rect 30377 8925 30389 8928
rect 30423 8925 30435 8959
rect 30377 8919 30435 8925
rect 28537 8891 28595 8897
rect 28537 8857 28549 8891
rect 28583 8888 28595 8891
rect 28994 8888 29000 8900
rect 28583 8860 29000 8888
rect 28583 8857 28595 8860
rect 28537 8851 28595 8857
rect 28994 8848 29000 8860
rect 29052 8848 29058 8900
rect 30392 8888 30420 8919
rect 30742 8916 30748 8968
rect 30800 8916 30806 8968
rect 33318 8916 33324 8968
rect 33376 8916 33382 8968
rect 33410 8916 33416 8968
rect 33468 8916 33474 8968
rect 33962 8916 33968 8968
rect 34020 8956 34026 8968
rect 34149 8959 34207 8965
rect 34149 8956 34161 8959
rect 34020 8928 34161 8956
rect 34020 8916 34026 8928
rect 34149 8925 34161 8928
rect 34195 8956 34207 8959
rect 34195 8928 36768 8956
rect 34195 8925 34207 8928
rect 34149 8919 34207 8925
rect 31294 8888 31300 8900
rect 30392 8860 31300 8888
rect 31294 8848 31300 8860
rect 31352 8848 31358 8900
rect 32306 8888 32312 8900
rect 32246 8860 32312 8888
rect 32306 8848 32312 8860
rect 32364 8848 32370 8900
rect 35253 8891 35311 8897
rect 35253 8888 35265 8891
rect 33520 8860 35265 8888
rect 22051 8792 27752 8820
rect 22051 8789 22063 8792
rect 22005 8783 22063 8789
rect 27798 8780 27804 8832
rect 27856 8820 27862 8832
rect 28629 8823 28687 8829
rect 28629 8820 28641 8823
rect 27856 8792 28641 8820
rect 27856 8780 27862 8792
rect 28629 8789 28641 8792
rect 28675 8789 28687 8823
rect 28629 8783 28687 8789
rect 29270 8780 29276 8832
rect 29328 8820 29334 8832
rect 30193 8823 30251 8829
rect 30193 8820 30205 8823
rect 29328 8792 30205 8820
rect 29328 8780 29334 8792
rect 30193 8789 30205 8792
rect 30239 8820 30251 8823
rect 30374 8820 30380 8832
rect 30239 8792 30380 8820
rect 30239 8789 30251 8792
rect 30193 8783 30251 8789
rect 30374 8780 30380 8792
rect 30432 8780 30438 8832
rect 31018 8780 31024 8832
rect 31076 8820 31082 8832
rect 33520 8820 33548 8860
rect 35253 8857 35265 8860
rect 35299 8857 35311 8891
rect 35253 8851 35311 8857
rect 35989 8891 36047 8897
rect 35989 8857 36001 8891
rect 36035 8888 36047 8891
rect 36173 8891 36231 8897
rect 36173 8888 36185 8891
rect 36035 8860 36185 8888
rect 36035 8857 36047 8860
rect 35989 8851 36047 8857
rect 36173 8857 36185 8860
rect 36219 8888 36231 8891
rect 36538 8888 36544 8900
rect 36219 8860 36544 8888
rect 36219 8857 36231 8860
rect 36173 8851 36231 8857
rect 31076 8792 33548 8820
rect 31076 8780 31082 8792
rect 34146 8780 34152 8832
rect 34204 8820 34210 8832
rect 34514 8820 34520 8832
rect 34204 8792 34520 8820
rect 34204 8780 34210 8792
rect 34514 8780 34520 8792
rect 34572 8780 34578 8832
rect 34606 8780 34612 8832
rect 34664 8820 34670 8832
rect 36004 8820 36032 8851
rect 36538 8848 36544 8860
rect 36596 8848 36602 8900
rect 36740 8888 36768 8928
rect 36814 8916 36820 8968
rect 36872 8916 36878 8968
rect 37844 8965 37872 8996
rect 49145 8993 49157 9027
rect 49191 9024 49203 9027
rect 49234 9024 49240 9036
rect 49191 8996 49240 9024
rect 49191 8993 49203 8996
rect 49145 8987 49203 8993
rect 49234 8984 49240 8996
rect 49292 8984 49298 9036
rect 37829 8959 37887 8965
rect 37829 8925 37841 8959
rect 37875 8925 37887 8959
rect 39853 8959 39911 8965
rect 39853 8956 39865 8959
rect 37829 8919 37887 8925
rect 39316 8928 39865 8956
rect 37274 8888 37280 8900
rect 36740 8860 37280 8888
rect 37274 8848 37280 8860
rect 37332 8848 37338 8900
rect 39316 8897 39344 8928
rect 39853 8925 39865 8928
rect 39899 8925 39911 8959
rect 39853 8919 39911 8925
rect 47118 8916 47124 8968
rect 47176 8956 47182 8968
rect 47949 8959 48007 8965
rect 47949 8956 47961 8959
rect 47176 8928 47961 8956
rect 47176 8916 47182 8928
rect 47949 8925 47961 8928
rect 47995 8925 48007 8959
rect 47949 8919 48007 8925
rect 39301 8891 39359 8897
rect 39301 8888 39313 8891
rect 37384 8860 39313 8888
rect 34664 8792 36032 8820
rect 34664 8780 34670 8792
rect 36262 8780 36268 8832
rect 36320 8820 36326 8832
rect 37384 8820 37412 8860
rect 39301 8857 39313 8860
rect 39347 8857 39359 8891
rect 39301 8851 39359 8857
rect 39485 8891 39543 8897
rect 39485 8857 39497 8891
rect 39531 8888 39543 8891
rect 42702 8888 42708 8900
rect 39531 8860 42708 8888
rect 39531 8857 39543 8860
rect 39485 8851 39543 8857
rect 42702 8848 42708 8860
rect 42760 8848 42766 8900
rect 36320 8792 37412 8820
rect 37645 8823 37703 8829
rect 36320 8780 36326 8792
rect 37645 8789 37657 8823
rect 37691 8820 37703 8823
rect 39574 8820 39580 8832
rect 37691 8792 39580 8820
rect 37691 8789 37703 8792
rect 37645 8783 37703 8789
rect 39574 8780 39580 8792
rect 39632 8780 39638 8832
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 13722 8576 13728 8628
rect 13780 8576 13786 8628
rect 14550 8576 14556 8628
rect 14608 8616 14614 8628
rect 14737 8619 14795 8625
rect 14737 8616 14749 8619
rect 14608 8588 14749 8616
rect 14608 8576 14614 8588
rect 14737 8585 14749 8588
rect 14783 8585 14795 8619
rect 14737 8579 14795 8585
rect 15102 8576 15108 8628
rect 15160 8576 15166 8628
rect 15746 8576 15752 8628
rect 15804 8576 15810 8628
rect 15841 8619 15899 8625
rect 15841 8585 15853 8619
rect 15887 8616 15899 8619
rect 15930 8616 15936 8628
rect 15887 8588 15936 8616
rect 15887 8585 15899 8588
rect 15841 8579 15899 8585
rect 15930 8576 15936 8588
rect 15988 8576 15994 8628
rect 16390 8576 16396 8628
rect 16448 8616 16454 8628
rect 16448 8588 17356 8616
rect 16448 8576 16454 8588
rect 1762 8508 1768 8560
rect 1820 8548 1826 8560
rect 14182 8548 14188 8560
rect 1820 8520 14188 8548
rect 1820 8508 1826 8520
rect 14182 8508 14188 8520
rect 14240 8508 14246 8560
rect 14274 8508 14280 8560
rect 14332 8548 14338 8560
rect 17129 8551 17187 8557
rect 14332 8520 16436 8548
rect 14332 8508 14338 8520
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 4062 8480 4068 8492
rect 1903 8452 4068 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 13814 8440 13820 8492
rect 13872 8480 13878 8492
rect 14093 8483 14151 8489
rect 14093 8480 14105 8483
rect 13872 8452 14105 8480
rect 13872 8440 13878 8452
rect 14093 8449 14105 8452
rect 14139 8480 14151 8483
rect 16408 8480 16436 8520
rect 17129 8517 17141 8551
rect 17175 8548 17187 8551
rect 17218 8548 17224 8560
rect 17175 8520 17224 8548
rect 17175 8517 17187 8520
rect 17129 8511 17187 8517
rect 17218 8508 17224 8520
rect 17276 8508 17282 8560
rect 17328 8548 17356 8588
rect 18690 8576 18696 8628
rect 18748 8616 18754 8628
rect 19061 8619 19119 8625
rect 19061 8616 19073 8619
rect 18748 8588 19073 8616
rect 18748 8576 18754 8588
rect 19061 8585 19073 8588
rect 19107 8585 19119 8619
rect 19061 8579 19119 8585
rect 19426 8576 19432 8628
rect 19484 8616 19490 8628
rect 20622 8616 20628 8628
rect 19484 8588 20628 8616
rect 19484 8576 19490 8588
rect 17586 8548 17592 8560
rect 17328 8520 17592 8548
rect 17586 8508 17592 8520
rect 17644 8508 17650 8560
rect 16850 8480 16856 8492
rect 14139 8452 15976 8480
rect 16408 8452 16856 8480
rect 14139 8449 14151 8452
rect 14093 8443 14151 8449
rect 1394 8372 1400 8424
rect 1452 8412 1458 8424
rect 15948 8421 15976 8452
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 19720 8489 19748 8588
rect 20622 8576 20628 8588
rect 20680 8576 20686 8628
rect 20990 8576 20996 8628
rect 21048 8616 21054 8628
rect 21453 8619 21511 8625
rect 21453 8616 21465 8619
rect 21048 8588 21465 8616
rect 21048 8576 21054 8588
rect 21453 8585 21465 8588
rect 21499 8585 21511 8619
rect 21453 8579 21511 8585
rect 22097 8619 22155 8625
rect 22097 8585 22109 8619
rect 22143 8616 22155 8619
rect 22370 8616 22376 8628
rect 22143 8588 22376 8616
rect 22143 8585 22155 8588
rect 22097 8579 22155 8585
rect 22370 8576 22376 8588
rect 22428 8576 22434 8628
rect 22738 8576 22744 8628
rect 22796 8616 22802 8628
rect 24121 8619 24179 8625
rect 24121 8616 24133 8619
rect 22796 8588 24133 8616
rect 22796 8576 22802 8588
rect 24121 8585 24133 8588
rect 24167 8585 24179 8619
rect 24121 8579 24179 8585
rect 24486 8576 24492 8628
rect 24544 8576 24550 8628
rect 25498 8576 25504 8628
rect 25556 8576 25562 8628
rect 25869 8619 25927 8625
rect 25869 8585 25881 8619
rect 25915 8616 25927 8619
rect 26050 8616 26056 8628
rect 25915 8588 26056 8616
rect 25915 8585 25927 8588
rect 25869 8579 25927 8585
rect 26050 8576 26056 8588
rect 26108 8576 26114 8628
rect 27614 8576 27620 8628
rect 27672 8616 27678 8628
rect 28353 8619 28411 8625
rect 28353 8616 28365 8619
rect 27672 8588 28365 8616
rect 27672 8576 27678 8588
rect 28353 8585 28365 8588
rect 28399 8585 28411 8619
rect 29454 8616 29460 8628
rect 28353 8579 28411 8585
rect 28552 8588 29460 8616
rect 20438 8508 20444 8560
rect 20496 8508 20502 8560
rect 23658 8508 23664 8560
rect 23716 8508 23722 8560
rect 19705 8483 19763 8489
rect 19705 8449 19717 8483
rect 19751 8449 19763 8483
rect 19705 8443 19763 8449
rect 24857 8483 24915 8489
rect 24857 8449 24869 8483
rect 24903 8480 24915 8483
rect 25038 8480 25044 8492
rect 24903 8452 25044 8480
rect 24903 8449 24915 8452
rect 24857 8443 24915 8449
rect 25038 8440 25044 8452
rect 25096 8440 25102 8492
rect 26418 8440 26424 8492
rect 26476 8480 26482 8492
rect 27709 8483 27767 8489
rect 27709 8480 27721 8483
rect 26476 8452 27721 8480
rect 26476 8440 26482 8452
rect 27709 8449 27721 8452
rect 27755 8480 27767 8483
rect 28552 8480 28580 8588
rect 29454 8576 29460 8588
rect 29512 8576 29518 8628
rect 31018 8576 31024 8628
rect 31076 8576 31082 8628
rect 31294 8576 31300 8628
rect 31352 8616 31358 8628
rect 31481 8619 31539 8625
rect 31481 8616 31493 8619
rect 31352 8588 31493 8616
rect 31352 8576 31358 8588
rect 31481 8585 31493 8588
rect 31527 8585 31539 8619
rect 33870 8616 33876 8628
rect 31481 8579 31539 8585
rect 32324 8588 33876 8616
rect 29086 8548 29092 8560
rect 28828 8520 29092 8548
rect 28828 8489 28856 8520
rect 29086 8508 29092 8520
rect 29144 8508 29150 8560
rect 30374 8508 30380 8560
rect 30432 8508 30438 8560
rect 30742 8508 30748 8560
rect 30800 8548 30806 8560
rect 32324 8548 32352 8588
rect 33870 8576 33876 8588
rect 33928 8576 33934 8628
rect 34238 8576 34244 8628
rect 34296 8616 34302 8628
rect 34333 8619 34391 8625
rect 34333 8616 34345 8619
rect 34296 8588 34345 8616
rect 34296 8576 34302 8588
rect 34333 8585 34345 8588
rect 34379 8585 34391 8619
rect 34333 8579 34391 8585
rect 34606 8576 34612 8628
rect 34664 8576 34670 8628
rect 34885 8619 34943 8625
rect 34885 8585 34897 8619
rect 34931 8585 34943 8619
rect 34885 8579 34943 8585
rect 34624 8548 34652 8576
rect 30800 8520 32352 8548
rect 33810 8520 34652 8548
rect 34900 8548 34928 8579
rect 35342 8576 35348 8628
rect 35400 8576 35406 8628
rect 38933 8619 38991 8625
rect 38933 8585 38945 8619
rect 38979 8616 38991 8619
rect 44818 8616 44824 8628
rect 38979 8588 44824 8616
rect 38979 8585 38991 8588
rect 38933 8579 38991 8585
rect 44818 8576 44824 8588
rect 44876 8576 44882 8628
rect 34900 8520 39160 8548
rect 30800 8508 30806 8520
rect 27755 8452 28580 8480
rect 28813 8483 28871 8489
rect 27755 8449 27767 8452
rect 27709 8443 27767 8449
rect 28813 8449 28825 8483
rect 28859 8449 28871 8483
rect 30392 8480 30420 8508
rect 30222 8452 30788 8480
rect 28813 8443 28871 8449
rect 30760 8424 30788 8452
rect 31386 8440 31392 8492
rect 31444 8440 31450 8492
rect 32324 8489 32352 8520
rect 32309 8483 32367 8489
rect 32309 8449 32321 8483
rect 32355 8449 32367 8483
rect 32309 8443 32367 8449
rect 35250 8440 35256 8492
rect 35308 8440 35314 8492
rect 36722 8480 36728 8492
rect 35360 8452 36728 8480
rect 1581 8415 1639 8421
rect 1581 8412 1593 8415
rect 1452 8384 1593 8412
rect 1452 8372 1458 8384
rect 1581 8381 1593 8384
rect 1627 8381 1639 8415
rect 1581 8375 1639 8381
rect 15933 8415 15991 8421
rect 15933 8381 15945 8415
rect 15979 8381 15991 8415
rect 15933 8375 15991 8381
rect 16114 8372 16120 8424
rect 16172 8412 16178 8424
rect 18874 8412 18880 8424
rect 16172 8384 18880 8412
rect 16172 8372 16178 8384
rect 18874 8372 18880 8384
rect 18932 8372 18938 8424
rect 19981 8415 20039 8421
rect 19981 8381 19993 8415
rect 20027 8412 20039 8415
rect 21450 8412 21456 8424
rect 20027 8384 21456 8412
rect 20027 8381 20039 8384
rect 19981 8375 20039 8381
rect 21450 8372 21456 8384
rect 21508 8372 21514 8424
rect 21542 8372 21548 8424
rect 21600 8412 21606 8424
rect 21821 8415 21879 8421
rect 21821 8412 21833 8415
rect 21600 8384 21833 8412
rect 21600 8372 21606 8384
rect 21821 8381 21833 8384
rect 21867 8381 21879 8415
rect 21821 8375 21879 8381
rect 22094 8372 22100 8424
rect 22152 8412 22158 8424
rect 22373 8415 22431 8421
rect 22373 8412 22385 8415
rect 22152 8384 22385 8412
rect 22152 8372 22158 8384
rect 22373 8381 22385 8384
rect 22419 8381 22431 8415
rect 22373 8375 22431 8381
rect 22649 8415 22707 8421
rect 22649 8381 22661 8415
rect 22695 8412 22707 8415
rect 25222 8412 25228 8424
rect 22695 8384 25228 8412
rect 22695 8381 22707 8384
rect 22649 8375 22707 8381
rect 25222 8372 25228 8384
rect 25280 8372 25286 8424
rect 29089 8415 29147 8421
rect 29089 8381 29101 8415
rect 29135 8412 29147 8415
rect 30374 8412 30380 8424
rect 29135 8384 30380 8412
rect 29135 8381 29147 8384
rect 29089 8375 29147 8381
rect 30374 8372 30380 8384
rect 30432 8372 30438 8424
rect 30742 8372 30748 8424
rect 30800 8372 30806 8424
rect 31662 8372 31668 8424
rect 31720 8372 31726 8424
rect 32585 8415 32643 8421
rect 32585 8381 32597 8415
rect 32631 8412 32643 8415
rect 35360 8412 35388 8452
rect 36722 8440 36728 8452
rect 36780 8440 36786 8492
rect 39132 8489 39160 8520
rect 39574 8508 39580 8560
rect 39632 8548 39638 8560
rect 44177 8551 44235 8557
rect 44177 8548 44189 8551
rect 39632 8520 44189 8548
rect 39632 8508 39638 8520
rect 44177 8517 44189 8520
rect 44223 8517 44235 8551
rect 44177 8511 44235 8517
rect 44361 8551 44419 8557
rect 44361 8517 44373 8551
rect 44407 8548 44419 8551
rect 47670 8548 47676 8560
rect 44407 8520 47676 8548
rect 44407 8517 44419 8520
rect 44361 8511 44419 8517
rect 47670 8508 47676 8520
rect 47728 8508 47734 8560
rect 49142 8508 49148 8560
rect 49200 8508 49206 8560
rect 37645 8483 37703 8489
rect 37645 8449 37657 8483
rect 37691 8449 37703 8483
rect 37645 8443 37703 8449
rect 39117 8483 39175 8489
rect 39117 8449 39129 8483
rect 39163 8449 39175 8483
rect 39117 8443 39175 8449
rect 40313 8483 40371 8489
rect 40313 8449 40325 8483
rect 40359 8480 40371 8483
rect 40865 8483 40923 8489
rect 40865 8480 40877 8483
rect 40359 8452 40877 8480
rect 40359 8449 40371 8452
rect 40313 8443 40371 8449
rect 40865 8449 40877 8452
rect 40911 8480 40923 8483
rect 41322 8480 41328 8492
rect 40911 8452 41328 8480
rect 40911 8449 40923 8452
rect 40865 8443 40923 8449
rect 32631 8384 35388 8412
rect 35437 8415 35495 8421
rect 32631 8381 32643 8384
rect 32585 8375 32643 8381
rect 35437 8381 35449 8415
rect 35483 8381 35495 8415
rect 35437 8375 35495 8381
rect 18598 8304 18604 8356
rect 18656 8304 18662 8356
rect 26050 8304 26056 8356
rect 26108 8304 26114 8356
rect 30561 8347 30619 8353
rect 30561 8313 30573 8347
rect 30607 8344 30619 8347
rect 32214 8344 32220 8356
rect 30607 8316 32220 8344
rect 30607 8313 30619 8316
rect 30561 8307 30619 8313
rect 32214 8304 32220 8316
rect 32272 8304 32278 8356
rect 34054 8304 34060 8356
rect 34112 8344 34118 8356
rect 35452 8344 35480 8375
rect 35802 8372 35808 8424
rect 35860 8412 35866 8424
rect 37660 8412 37688 8443
rect 41322 8440 41328 8452
rect 41380 8440 41386 8492
rect 45830 8440 45836 8492
rect 45888 8440 45894 8492
rect 46750 8440 46756 8492
rect 46808 8480 46814 8492
rect 47949 8483 48007 8489
rect 47949 8480 47961 8483
rect 46808 8452 47961 8480
rect 46808 8440 46814 8452
rect 47949 8449 47961 8452
rect 47995 8449 48007 8483
rect 47949 8443 48007 8449
rect 35860 8384 37688 8412
rect 40497 8415 40555 8421
rect 35860 8372 35866 8384
rect 40497 8381 40509 8415
rect 40543 8412 40555 8415
rect 40543 8384 45554 8412
rect 40543 8381 40555 8384
rect 40497 8375 40555 8381
rect 34112 8316 35480 8344
rect 37461 8347 37519 8353
rect 34112 8304 34118 8316
rect 37461 8313 37473 8347
rect 37507 8344 37519 8347
rect 41414 8344 41420 8356
rect 37507 8316 41420 8344
rect 37507 8313 37519 8316
rect 37461 8307 37519 8313
rect 41414 8304 41420 8316
rect 41472 8304 41478 8356
rect 45526 8344 45554 8384
rect 46842 8372 46848 8424
rect 46900 8372 46906 8424
rect 47578 8344 47584 8356
rect 45526 8316 47584 8344
rect 47578 8304 47584 8316
rect 47636 8304 47642 8356
rect 15378 8236 15384 8288
rect 15436 8236 15442 8288
rect 16390 8236 16396 8288
rect 16448 8236 16454 8288
rect 27798 8236 27804 8288
rect 27856 8276 27862 8288
rect 32766 8276 32772 8288
rect 27856 8248 32772 8276
rect 27856 8236 27862 8248
rect 32766 8236 32772 8248
rect 32824 8276 32830 8288
rect 34422 8276 34428 8288
rect 32824 8248 34428 8276
rect 32824 8236 32830 8248
rect 34422 8236 34428 8248
rect 34480 8236 34486 8288
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 2133 8075 2191 8081
rect 2133 8072 2145 8075
rect 1452 8044 2145 8072
rect 1452 8032 1458 8044
rect 2133 8041 2145 8044
rect 2179 8041 2191 8075
rect 2133 8035 2191 8041
rect 16574 8032 16580 8084
rect 16632 8032 16638 8084
rect 17126 8032 17132 8084
rect 17184 8072 17190 8084
rect 17497 8075 17555 8081
rect 17497 8072 17509 8075
rect 17184 8044 17509 8072
rect 17184 8032 17190 8044
rect 17497 8041 17509 8044
rect 17543 8041 17555 8075
rect 17497 8035 17555 8041
rect 17957 8075 18015 8081
rect 17957 8041 17969 8075
rect 18003 8072 18015 8075
rect 18690 8072 18696 8084
rect 18003 8044 18696 8072
rect 18003 8041 18015 8044
rect 17957 8035 18015 8041
rect 18690 8032 18696 8044
rect 18748 8032 18754 8084
rect 20346 8032 20352 8084
rect 20404 8072 20410 8084
rect 20441 8075 20499 8081
rect 20441 8072 20453 8075
rect 20404 8044 20453 8072
rect 20404 8032 20410 8044
rect 20441 8041 20453 8044
rect 20487 8041 20499 8075
rect 20441 8035 20499 8041
rect 15381 8007 15439 8013
rect 15381 7973 15393 8007
rect 15427 8004 15439 8007
rect 17862 8004 17868 8016
rect 15427 7976 17868 8004
rect 15427 7973 15439 7976
rect 15381 7967 15439 7973
rect 17862 7964 17868 7976
rect 17920 7964 17926 8016
rect 20456 8004 20484 8035
rect 20806 8032 20812 8084
rect 20864 8072 20870 8084
rect 21818 8072 21824 8084
rect 20864 8044 21824 8072
rect 20864 8032 20870 8044
rect 21818 8032 21824 8044
rect 21876 8072 21882 8084
rect 23109 8075 23167 8081
rect 23109 8072 23121 8075
rect 21876 8044 23121 8072
rect 21876 8032 21882 8044
rect 23109 8041 23121 8044
rect 23155 8041 23167 8075
rect 23109 8035 23167 8041
rect 25222 8032 25228 8084
rect 25280 8032 25286 8084
rect 30374 8032 30380 8084
rect 30432 8032 30438 8084
rect 31021 8075 31079 8081
rect 31021 8041 31033 8075
rect 31067 8072 31079 8075
rect 35250 8072 35256 8084
rect 31067 8044 35256 8072
rect 31067 8041 31079 8044
rect 31021 8035 31079 8041
rect 35250 8032 35256 8044
rect 35308 8032 35314 8084
rect 20901 8007 20959 8013
rect 20901 8004 20913 8007
rect 18340 7976 19932 8004
rect 20456 7976 20913 8004
rect 14826 7896 14832 7948
rect 14884 7936 14890 7948
rect 15841 7939 15899 7945
rect 15841 7936 15853 7939
rect 14884 7908 15853 7936
rect 14884 7896 14890 7908
rect 15841 7905 15853 7908
rect 15887 7905 15899 7939
rect 15841 7899 15899 7905
rect 16022 7896 16028 7948
rect 16080 7896 16086 7948
rect 18340 7936 18368 7976
rect 16776 7908 18368 7936
rect 1302 7828 1308 7880
rect 1360 7868 1366 7880
rect 1581 7871 1639 7877
rect 1581 7868 1593 7871
rect 1360 7840 1593 7868
rect 1360 7828 1366 7840
rect 1581 7837 1593 7840
rect 1627 7868 1639 7871
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 1627 7840 2329 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 2317 7837 2329 7840
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 15378 7828 15384 7880
rect 15436 7868 15442 7880
rect 15749 7871 15807 7877
rect 15749 7868 15761 7871
rect 15436 7840 15761 7868
rect 15436 7828 15442 7840
rect 15749 7837 15761 7840
rect 15795 7837 15807 7871
rect 15749 7831 15807 7837
rect 10686 7800 10692 7812
rect 1780 7772 10692 7800
rect 1780 7741 1808 7772
rect 10686 7760 10692 7772
rect 10744 7760 10750 7812
rect 14366 7760 14372 7812
rect 14424 7800 14430 7812
rect 16776 7800 16804 7908
rect 18414 7896 18420 7948
rect 18472 7896 18478 7948
rect 18506 7896 18512 7948
rect 18564 7896 18570 7948
rect 19904 7945 19932 7976
rect 20901 7973 20913 7976
rect 20947 7973 20959 8007
rect 20901 7967 20959 7973
rect 30650 7964 30656 8016
rect 30708 8004 30714 8016
rect 32861 8007 32919 8013
rect 32861 8004 32873 8007
rect 30708 7976 32873 8004
rect 30708 7964 30714 7976
rect 32861 7973 32873 7976
rect 32907 7973 32919 8007
rect 32861 7967 32919 7973
rect 19889 7939 19947 7945
rect 19889 7905 19901 7939
rect 19935 7905 19947 7939
rect 19889 7899 19947 7905
rect 19981 7939 20039 7945
rect 19981 7905 19993 7939
rect 20027 7905 20039 7939
rect 19981 7899 20039 7905
rect 16853 7871 16911 7877
rect 16853 7837 16865 7871
rect 16899 7868 16911 7871
rect 18598 7868 18604 7880
rect 16899 7840 18604 7868
rect 16899 7837 16911 7840
rect 16853 7831 16911 7837
rect 18598 7828 18604 7840
rect 18656 7868 18662 7880
rect 19996 7868 20024 7899
rect 20714 7896 20720 7948
rect 20772 7936 20778 7948
rect 21361 7939 21419 7945
rect 21361 7936 21373 7939
rect 20772 7908 21373 7936
rect 20772 7896 20778 7908
rect 21361 7905 21373 7908
rect 21407 7936 21419 7939
rect 22002 7936 22008 7948
rect 21407 7908 22008 7936
rect 21407 7905 21419 7908
rect 21361 7899 21419 7905
rect 22002 7896 22008 7908
rect 22060 7896 22066 7948
rect 28994 7896 29000 7948
rect 29052 7896 29058 7948
rect 31110 7896 31116 7948
rect 31168 7936 31174 7948
rect 31481 7939 31539 7945
rect 31481 7936 31493 7939
rect 31168 7908 31493 7936
rect 31168 7896 31174 7908
rect 31481 7905 31493 7908
rect 31527 7905 31539 7939
rect 31481 7899 31539 7905
rect 31665 7939 31723 7945
rect 31665 7905 31677 7939
rect 31711 7936 31723 7939
rect 32674 7936 32680 7948
rect 31711 7908 32680 7936
rect 31711 7905 31723 7908
rect 31665 7899 31723 7905
rect 32674 7896 32680 7908
rect 32732 7896 32738 7948
rect 49145 7939 49203 7945
rect 49145 7905 49157 7939
rect 49191 7936 49203 7939
rect 49234 7936 49240 7948
rect 49191 7908 49240 7936
rect 49191 7905 49203 7908
rect 49145 7899 49203 7905
rect 49234 7896 49240 7908
rect 49292 7896 49298 7948
rect 18656 7840 20024 7868
rect 18656 7828 18662 7840
rect 23842 7828 23848 7880
rect 23900 7868 23906 7880
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 23900 7840 24593 7868
rect 23900 7828 23906 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 29733 7871 29791 7877
rect 29733 7837 29745 7871
rect 29779 7868 29791 7871
rect 29822 7868 29828 7880
rect 29779 7840 29828 7868
rect 29779 7837 29791 7840
rect 29733 7831 29791 7837
rect 29822 7828 29828 7840
rect 29880 7828 29886 7880
rect 32214 7828 32220 7880
rect 32272 7828 32278 7880
rect 34422 7828 34428 7880
rect 34480 7868 34486 7880
rect 38749 7871 38807 7877
rect 38749 7868 38761 7871
rect 34480 7840 38761 7868
rect 34480 7828 34486 7840
rect 38749 7837 38761 7840
rect 38795 7868 38807 7871
rect 39209 7871 39267 7877
rect 39209 7868 39221 7871
rect 38795 7840 39221 7868
rect 38795 7837 38807 7840
rect 38749 7831 38807 7837
rect 39209 7837 39221 7840
rect 39255 7837 39267 7871
rect 39209 7831 39267 7837
rect 47026 7828 47032 7880
rect 47084 7868 47090 7880
rect 47949 7871 48007 7877
rect 47949 7868 47961 7871
rect 47084 7840 47961 7868
rect 47084 7828 47090 7840
rect 47949 7837 47961 7840
rect 47995 7837 48007 7871
rect 47949 7831 48007 7837
rect 20717 7803 20775 7809
rect 20717 7800 20729 7803
rect 14424 7772 16804 7800
rect 18340 7772 20729 7800
rect 14424 7760 14430 7772
rect 1765 7735 1823 7741
rect 1765 7701 1777 7735
rect 1811 7701 1823 7735
rect 1765 7695 1823 7701
rect 15102 7692 15108 7744
rect 15160 7692 15166 7744
rect 17770 7692 17776 7744
rect 17828 7732 17834 7744
rect 18340 7741 18368 7772
rect 20717 7769 20729 7772
rect 20763 7800 20775 7803
rect 21266 7800 21272 7812
rect 20763 7772 21272 7800
rect 20763 7769 20775 7772
rect 20717 7763 20775 7769
rect 21266 7760 21272 7772
rect 21324 7760 21330 7812
rect 21637 7803 21695 7809
rect 21637 7769 21649 7803
rect 21683 7769 21695 7803
rect 22862 7772 23520 7800
rect 21637 7763 21695 7769
rect 18325 7735 18383 7741
rect 18325 7732 18337 7735
rect 17828 7704 18337 7732
rect 17828 7692 17834 7704
rect 18325 7701 18337 7704
rect 18371 7701 18383 7735
rect 18325 7695 18383 7701
rect 18598 7692 18604 7744
rect 18656 7732 18662 7744
rect 18969 7735 19027 7741
rect 18969 7732 18981 7735
rect 18656 7704 18981 7732
rect 18656 7692 18662 7704
rect 18969 7701 18981 7704
rect 19015 7701 19027 7735
rect 18969 7695 19027 7701
rect 19426 7692 19432 7744
rect 19484 7692 19490 7744
rect 19794 7692 19800 7744
rect 19852 7692 19858 7744
rect 20898 7692 20904 7744
rect 20956 7732 20962 7744
rect 20993 7735 21051 7741
rect 20993 7732 21005 7735
rect 20956 7704 21005 7732
rect 20956 7692 20962 7704
rect 20993 7701 21005 7704
rect 21039 7701 21051 7735
rect 21652 7732 21680 7763
rect 23290 7732 23296 7744
rect 21652 7704 23296 7732
rect 20993 7695 21051 7701
rect 23290 7692 23296 7704
rect 23348 7692 23354 7744
rect 23492 7741 23520 7772
rect 28350 7760 28356 7812
rect 28408 7800 28414 7812
rect 31389 7803 31447 7809
rect 28408 7772 30880 7800
rect 28408 7760 28414 7772
rect 23477 7735 23535 7741
rect 23477 7701 23489 7735
rect 23523 7732 23535 7735
rect 23658 7732 23664 7744
rect 23523 7704 23664 7732
rect 23523 7701 23535 7704
rect 23477 7695 23535 7701
rect 23658 7692 23664 7704
rect 23716 7732 23722 7744
rect 24121 7735 24179 7741
rect 24121 7732 24133 7735
rect 23716 7704 24133 7732
rect 23716 7692 23722 7704
rect 24121 7701 24133 7704
rect 24167 7701 24179 7735
rect 24121 7695 24179 7701
rect 27798 7692 27804 7744
rect 27856 7732 27862 7744
rect 27985 7735 28043 7741
rect 27985 7732 27997 7735
rect 27856 7704 27997 7732
rect 27856 7692 27862 7704
rect 27985 7701 27997 7704
rect 28031 7701 28043 7735
rect 27985 7695 28043 7701
rect 30742 7692 30748 7744
rect 30800 7692 30806 7744
rect 30852 7732 30880 7772
rect 31389 7769 31401 7803
rect 31435 7800 31447 7803
rect 33321 7803 33379 7809
rect 33321 7800 33333 7803
rect 31435 7772 33333 7800
rect 31435 7769 31447 7772
rect 31389 7763 31447 7769
rect 33321 7769 33333 7772
rect 33367 7769 33379 7803
rect 38013 7803 38071 7809
rect 38013 7800 38025 7803
rect 33321 7763 33379 7769
rect 37568 7772 38025 7800
rect 37568 7741 37596 7772
rect 38013 7769 38025 7772
rect 38059 7769 38071 7803
rect 38013 7763 38071 7769
rect 38933 7803 38991 7809
rect 38933 7769 38945 7803
rect 38979 7800 38991 7803
rect 40586 7800 40592 7812
rect 38979 7772 40592 7800
rect 38979 7769 38991 7772
rect 38933 7763 38991 7769
rect 40586 7760 40592 7772
rect 40644 7760 40650 7812
rect 37553 7735 37611 7741
rect 37553 7732 37565 7735
rect 30852 7704 37565 7732
rect 37553 7701 37565 7704
rect 37599 7701 37611 7735
rect 37553 7695 37611 7701
rect 38105 7735 38163 7741
rect 38105 7701 38117 7735
rect 38151 7732 38163 7735
rect 38654 7732 38660 7744
rect 38151 7704 38660 7732
rect 38151 7701 38163 7704
rect 38105 7695 38163 7701
rect 38654 7692 38660 7704
rect 38712 7692 38718 7744
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 16298 7488 16304 7540
rect 16356 7528 16362 7540
rect 17497 7531 17555 7537
rect 17497 7528 17509 7531
rect 16356 7500 17509 7528
rect 16356 7488 16362 7500
rect 17497 7497 17509 7500
rect 17543 7497 17555 7531
rect 17497 7491 17555 7497
rect 18233 7531 18291 7537
rect 18233 7497 18245 7531
rect 18279 7497 18291 7531
rect 18233 7491 18291 7497
rect 16022 7420 16028 7472
rect 16080 7460 16086 7472
rect 18248 7460 18276 7491
rect 18322 7488 18328 7540
rect 18380 7528 18386 7540
rect 18601 7531 18659 7537
rect 18601 7528 18613 7531
rect 18380 7500 18613 7528
rect 18380 7488 18386 7500
rect 18601 7497 18613 7500
rect 18647 7497 18659 7531
rect 18601 7491 18659 7497
rect 18690 7488 18696 7540
rect 18748 7488 18754 7540
rect 19242 7488 19248 7540
rect 19300 7528 19306 7540
rect 20073 7531 20131 7537
rect 20073 7528 20085 7531
rect 19300 7500 20085 7528
rect 19300 7488 19306 7500
rect 20073 7497 20085 7500
rect 20119 7497 20131 7531
rect 20073 7491 20131 7497
rect 20346 7488 20352 7540
rect 20404 7488 20410 7540
rect 21450 7488 21456 7540
rect 21508 7488 21514 7540
rect 22278 7488 22284 7540
rect 22336 7528 22342 7540
rect 22649 7531 22707 7537
rect 22649 7528 22661 7531
rect 22336 7500 22661 7528
rect 22336 7488 22342 7500
rect 22649 7497 22661 7500
rect 22695 7497 22707 7531
rect 22649 7491 22707 7497
rect 23290 7488 23296 7540
rect 23348 7528 23354 7540
rect 23753 7531 23811 7537
rect 23753 7528 23765 7531
rect 23348 7500 23765 7528
rect 23348 7488 23354 7500
rect 23753 7497 23765 7500
rect 23799 7497 23811 7531
rect 23753 7491 23811 7497
rect 29638 7488 29644 7540
rect 29696 7488 29702 7540
rect 31386 7488 31392 7540
rect 31444 7488 31450 7540
rect 32858 7488 32864 7540
rect 32916 7528 32922 7540
rect 32953 7531 33011 7537
rect 32953 7528 32965 7531
rect 32916 7500 32965 7528
rect 32916 7488 32922 7500
rect 32953 7497 32965 7500
rect 32999 7497 33011 7531
rect 32953 7491 33011 7497
rect 37366 7488 37372 7540
rect 37424 7488 37430 7540
rect 19794 7460 19800 7472
rect 16080 7432 16896 7460
rect 18248 7432 19800 7460
rect 16080 7420 16086 7432
rect 1302 7352 1308 7404
rect 1360 7392 1366 7404
rect 1581 7395 1639 7401
rect 1581 7392 1593 7395
rect 1360 7364 1593 7392
rect 1360 7352 1366 7364
rect 1581 7361 1593 7364
rect 1627 7392 1639 7395
rect 2133 7395 2191 7401
rect 2133 7392 2145 7395
rect 1627 7364 2145 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 2133 7361 2145 7364
rect 2179 7361 2191 7395
rect 2133 7355 2191 7361
rect 14090 7352 14096 7404
rect 14148 7392 14154 7404
rect 16868 7401 16896 7432
rect 19794 7420 19800 7432
rect 19852 7420 19858 7472
rect 20898 7420 20904 7472
rect 20956 7460 20962 7472
rect 22462 7460 22468 7472
rect 20956 7432 22468 7460
rect 20956 7420 20962 7432
rect 22462 7420 22468 7432
rect 22520 7420 22526 7472
rect 29546 7420 29552 7472
rect 29604 7460 29610 7472
rect 30929 7463 30987 7469
rect 30929 7460 30941 7463
rect 29604 7432 30941 7460
rect 29604 7420 29610 7432
rect 30929 7429 30941 7432
rect 30975 7429 30987 7463
rect 37384 7460 37412 7488
rect 37829 7463 37887 7469
rect 37829 7460 37841 7463
rect 37384 7432 37841 7460
rect 30929 7423 30987 7429
rect 37829 7429 37841 7432
rect 37875 7429 37887 7463
rect 37829 7423 37887 7429
rect 44818 7420 44824 7472
rect 44876 7420 44882 7472
rect 49145 7463 49203 7469
rect 49145 7429 49157 7463
rect 49191 7460 49203 7463
rect 49326 7460 49332 7472
rect 49191 7432 49332 7460
rect 49191 7429 49203 7432
rect 49145 7423 49203 7429
rect 49326 7420 49332 7432
rect 49384 7420 49390 7472
rect 16209 7395 16267 7401
rect 16209 7392 16221 7395
rect 14148 7364 16221 7392
rect 14148 7352 14154 7364
rect 16209 7361 16221 7364
rect 16255 7361 16267 7395
rect 16209 7355 16267 7361
rect 16853 7395 16911 7401
rect 16853 7361 16865 7395
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 19429 7395 19487 7401
rect 19429 7361 19441 7395
rect 19475 7361 19487 7395
rect 19429 7355 19487 7361
rect 17310 7324 17316 7336
rect 12406 7296 17316 7324
rect 1765 7259 1823 7265
rect 1765 7225 1777 7259
rect 1811 7256 1823 7259
rect 12406 7256 12434 7296
rect 17310 7284 17316 7296
rect 17368 7284 17374 7336
rect 18877 7327 18935 7333
rect 18877 7293 18889 7327
rect 18923 7324 18935 7327
rect 18966 7324 18972 7336
rect 18923 7296 18972 7324
rect 18923 7293 18935 7296
rect 18877 7287 18935 7293
rect 18966 7284 18972 7296
rect 19024 7284 19030 7336
rect 19444 7324 19472 7355
rect 20806 7352 20812 7404
rect 20864 7352 20870 7404
rect 21726 7352 21732 7404
rect 21784 7392 21790 7404
rect 22005 7395 22063 7401
rect 22005 7392 22017 7395
rect 21784 7364 22017 7392
rect 21784 7352 21790 7364
rect 22005 7361 22017 7364
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 22738 7352 22744 7404
rect 22796 7392 22802 7404
rect 23109 7395 23167 7401
rect 23109 7392 23121 7395
rect 22796 7364 23121 7392
rect 22796 7352 22802 7364
rect 23109 7361 23121 7364
rect 23155 7361 23167 7395
rect 23109 7355 23167 7361
rect 30285 7395 30343 7401
rect 30285 7361 30297 7395
rect 30331 7392 30343 7395
rect 31478 7392 31484 7404
rect 30331 7364 31484 7392
rect 30331 7361 30343 7364
rect 30285 7355 30343 7361
rect 31478 7352 31484 7364
rect 31536 7352 31542 7404
rect 32309 7395 32367 7401
rect 32309 7361 32321 7395
rect 32355 7392 32367 7395
rect 34054 7392 34060 7404
rect 32355 7364 34060 7392
rect 32355 7361 32367 7364
rect 32309 7355 32367 7361
rect 34054 7352 34060 7364
rect 34112 7352 34118 7404
rect 38565 7395 38623 7401
rect 38565 7361 38577 7395
rect 38611 7392 38623 7395
rect 39025 7395 39083 7401
rect 39025 7392 39037 7395
rect 38611 7364 39037 7392
rect 38611 7361 38623 7364
rect 38565 7355 38623 7361
rect 39025 7361 39037 7364
rect 39071 7361 39083 7395
rect 39025 7355 39083 7361
rect 21634 7324 21640 7336
rect 19444 7296 21640 7324
rect 21634 7284 21640 7296
rect 21692 7284 21698 7336
rect 29730 7284 29736 7336
rect 29788 7324 29794 7336
rect 38580 7324 38608 7355
rect 46934 7352 46940 7404
rect 46992 7392 46998 7404
rect 47949 7395 48007 7401
rect 47949 7392 47961 7395
rect 46992 7364 47961 7392
rect 46992 7352 46998 7364
rect 47949 7361 47961 7364
rect 47995 7361 48007 7395
rect 47949 7355 48007 7361
rect 29788 7296 38608 7324
rect 29788 7284 29794 7296
rect 38654 7284 38660 7336
rect 38712 7324 38718 7336
rect 47026 7324 47032 7336
rect 38712 7296 47032 7324
rect 38712 7284 38718 7296
rect 47026 7284 47032 7296
rect 47084 7284 47090 7336
rect 1811 7228 12434 7256
rect 16025 7259 16083 7265
rect 1811 7225 1823 7228
rect 1765 7219 1823 7225
rect 16025 7225 16037 7259
rect 16071 7256 16083 7259
rect 19518 7256 19524 7268
rect 16071 7228 19524 7256
rect 16071 7225 16083 7228
rect 16025 7219 16083 7225
rect 19518 7216 19524 7228
rect 19576 7216 19582 7268
rect 38749 7259 38807 7265
rect 38749 7225 38761 7259
rect 38795 7256 38807 7259
rect 45005 7259 45063 7265
rect 38795 7228 42104 7256
rect 38795 7225 38807 7228
rect 38749 7219 38807 7225
rect 15102 7148 15108 7200
rect 15160 7188 15166 7200
rect 15749 7191 15807 7197
rect 15749 7188 15761 7191
rect 15160 7160 15761 7188
rect 15160 7148 15166 7160
rect 15749 7157 15761 7160
rect 15795 7188 15807 7191
rect 16390 7188 16396 7200
rect 15795 7160 16396 7188
rect 15795 7157 15807 7160
rect 15749 7151 15807 7157
rect 16390 7148 16396 7160
rect 16448 7188 16454 7200
rect 17957 7191 18015 7197
rect 17957 7188 17969 7191
rect 16448 7160 17969 7188
rect 16448 7148 16454 7160
rect 17957 7157 17969 7160
rect 18003 7188 18015 7191
rect 18690 7188 18696 7200
rect 18003 7160 18696 7188
rect 18003 7157 18015 7160
rect 17957 7151 18015 7157
rect 18690 7148 18696 7160
rect 18748 7148 18754 7200
rect 37918 7148 37924 7200
rect 37976 7148 37982 7200
rect 42076 7188 42104 7228
rect 45005 7225 45017 7259
rect 45051 7256 45063 7259
rect 47210 7256 47216 7268
rect 45051 7228 47216 7256
rect 45051 7225 45063 7228
rect 45005 7219 45063 7225
rect 47210 7216 47216 7228
rect 47268 7216 47274 7268
rect 45738 7188 45744 7200
rect 42076 7160 45744 7188
rect 45738 7148 45744 7160
rect 45796 7148 45802 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 18690 6944 18696 6996
rect 18748 6984 18754 6996
rect 19889 6987 19947 6993
rect 19889 6984 19901 6987
rect 18748 6956 19901 6984
rect 18748 6944 18754 6956
rect 19889 6953 19901 6956
rect 19935 6984 19947 6987
rect 20346 6984 20352 6996
rect 19935 6956 20352 6984
rect 19935 6953 19947 6956
rect 19889 6947 19947 6953
rect 20346 6944 20352 6956
rect 20404 6944 20410 6996
rect 31110 6944 31116 6996
rect 31168 6984 31174 6996
rect 31297 6987 31355 6993
rect 31297 6984 31309 6987
rect 31168 6956 31309 6984
rect 31168 6944 31174 6956
rect 31297 6953 31309 6956
rect 31343 6953 31355 6987
rect 31297 6947 31355 6953
rect 37918 6876 37924 6928
rect 37976 6916 37982 6928
rect 47118 6916 47124 6928
rect 37976 6888 47124 6916
rect 37976 6876 37982 6888
rect 47118 6876 47124 6888
rect 47176 6876 47182 6928
rect 17402 6808 17408 6860
rect 17460 6848 17466 6860
rect 18877 6851 18935 6857
rect 18877 6848 18889 6851
rect 17460 6820 18889 6848
rect 17460 6808 17466 6820
rect 18877 6817 18889 6820
rect 18923 6817 18935 6851
rect 18877 6811 18935 6817
rect 19702 6808 19708 6860
rect 19760 6848 19766 6860
rect 20993 6851 21051 6857
rect 20993 6848 21005 6851
rect 19760 6820 21005 6848
rect 19760 6808 19766 6820
rect 20993 6817 21005 6820
rect 21039 6817 21051 6851
rect 20993 6811 21051 6817
rect 21358 6808 21364 6860
rect 21416 6848 21422 6860
rect 22189 6851 22247 6857
rect 22189 6848 22201 6851
rect 21416 6820 22201 6848
rect 21416 6808 21422 6820
rect 22189 6817 22201 6820
rect 22235 6817 22247 6851
rect 22189 6811 22247 6817
rect 30006 6808 30012 6860
rect 30064 6848 30070 6860
rect 31021 6851 31079 6857
rect 31021 6848 31033 6851
rect 30064 6820 31033 6848
rect 30064 6808 30070 6820
rect 31021 6817 31033 6820
rect 31067 6817 31079 6851
rect 31021 6811 31079 6817
rect 49142 6808 49148 6860
rect 49200 6808 49206 6860
rect 1302 6740 1308 6792
rect 1360 6780 1366 6792
rect 2501 6783 2559 6789
rect 2501 6780 2513 6783
rect 1360 6752 2513 6780
rect 1360 6740 1366 6752
rect 2501 6749 2513 6752
rect 2547 6780 2559 6783
rect 2777 6783 2835 6789
rect 2777 6780 2789 6783
rect 2547 6752 2789 6780
rect 2547 6749 2559 6752
rect 2501 6743 2559 6749
rect 2777 6749 2789 6752
rect 2823 6749 2835 6783
rect 18233 6783 18291 6789
rect 2777 6743 2835 6749
rect 9646 6752 18000 6780
rect 1210 6672 1216 6724
rect 1268 6712 1274 6724
rect 1673 6715 1731 6721
rect 1673 6712 1685 6715
rect 1268 6684 1685 6712
rect 1268 6672 1274 6684
rect 1673 6681 1685 6684
rect 1719 6681 1731 6715
rect 1673 6675 1731 6681
rect 1857 6715 1915 6721
rect 1857 6681 1869 6715
rect 1903 6712 1915 6715
rect 9646 6712 9674 6752
rect 1903 6684 9674 6712
rect 17972 6712 18000 6752
rect 18233 6749 18245 6783
rect 18279 6780 18291 6783
rect 19058 6780 19064 6792
rect 18279 6752 19064 6780
rect 18279 6749 18291 6752
rect 18233 6743 18291 6749
rect 19058 6740 19064 6752
rect 19116 6740 19122 6792
rect 20070 6740 20076 6792
rect 20128 6780 20134 6792
rect 20349 6783 20407 6789
rect 20349 6780 20361 6783
rect 20128 6752 20361 6780
rect 20128 6740 20134 6752
rect 20349 6749 20361 6752
rect 20395 6749 20407 6783
rect 20349 6743 20407 6749
rect 21174 6740 21180 6792
rect 21232 6780 21238 6792
rect 21545 6783 21603 6789
rect 21545 6780 21557 6783
rect 21232 6752 21557 6780
rect 21232 6740 21238 6752
rect 21545 6749 21557 6752
rect 21591 6749 21603 6783
rect 21545 6743 21603 6749
rect 30377 6783 30435 6789
rect 30377 6749 30389 6783
rect 30423 6780 30435 6783
rect 30466 6780 30472 6792
rect 30423 6752 30472 6780
rect 30423 6749 30435 6752
rect 30377 6743 30435 6749
rect 30466 6740 30472 6752
rect 30524 6740 30530 6792
rect 40586 6740 40592 6792
rect 40644 6780 40650 6792
rect 46109 6783 46167 6789
rect 46109 6780 46121 6783
rect 40644 6752 46121 6780
rect 40644 6740 40650 6752
rect 46109 6749 46121 6752
rect 46155 6749 46167 6783
rect 46109 6743 46167 6749
rect 47670 6740 47676 6792
rect 47728 6780 47734 6792
rect 47949 6783 48007 6789
rect 47949 6780 47961 6783
rect 47728 6752 47961 6780
rect 47728 6740 47734 6752
rect 47949 6749 47961 6752
rect 47995 6749 48007 6783
rect 47949 6743 48007 6749
rect 27798 6712 27804 6724
rect 17972 6684 27804 6712
rect 1903 6681 1915 6684
rect 1857 6675 1915 6681
rect 27798 6672 27804 6684
rect 27856 6672 27862 6724
rect 47305 6715 47363 6721
rect 47305 6681 47317 6715
rect 47351 6712 47363 6715
rect 48866 6712 48872 6724
rect 47351 6684 48872 6712
rect 47351 6681 47363 6684
rect 47305 6675 47363 6681
rect 48866 6672 48872 6684
rect 48924 6672 48930 6724
rect 2317 6647 2375 6653
rect 2317 6613 2329 6647
rect 2363 6644 2375 6647
rect 2406 6644 2412 6656
rect 2363 6616 2412 6644
rect 2363 6613 2375 6616
rect 2317 6607 2375 6613
rect 2406 6604 2412 6616
rect 2464 6604 2470 6656
rect 16390 6604 16396 6656
rect 16448 6604 16454 6656
rect 17770 6604 17776 6656
rect 17828 6604 17834 6656
rect 18874 6604 18880 6656
rect 18932 6644 18938 6656
rect 19429 6647 19487 6653
rect 19429 6644 19441 6647
rect 18932 6616 19441 6644
rect 18932 6604 18938 6616
rect 19429 6613 19441 6616
rect 19475 6613 19487 6647
rect 19429 6607 19487 6613
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 1210 6400 1216 6452
rect 1268 6440 1274 6452
rect 2133 6443 2191 6449
rect 2133 6440 2145 6443
rect 1268 6412 2145 6440
rect 1268 6400 1274 6412
rect 2133 6409 2145 6412
rect 2179 6409 2191 6443
rect 2133 6403 2191 6409
rect 18690 6400 18696 6452
rect 18748 6400 18754 6452
rect 19610 6400 19616 6452
rect 19668 6440 19674 6452
rect 19889 6443 19947 6449
rect 19889 6440 19901 6443
rect 19668 6412 19901 6440
rect 19668 6400 19674 6412
rect 19889 6409 19901 6412
rect 19935 6409 19947 6443
rect 19889 6403 19947 6409
rect 34146 6332 34152 6384
rect 34204 6372 34210 6384
rect 37553 6375 37611 6381
rect 37553 6372 37565 6375
rect 34204 6344 37565 6372
rect 34204 6332 34210 6344
rect 37553 6341 37565 6344
rect 37599 6372 37611 6375
rect 38013 6375 38071 6381
rect 38013 6372 38025 6375
rect 37599 6344 38025 6372
rect 37599 6341 37611 6344
rect 37553 6335 37611 6341
rect 38013 6341 38025 6344
rect 38059 6341 38071 6375
rect 38013 6335 38071 6341
rect 41414 6332 41420 6384
rect 41472 6372 41478 6384
rect 43993 6375 44051 6381
rect 43993 6372 44005 6375
rect 41472 6344 44005 6372
rect 41472 6332 41478 6344
rect 43993 6341 44005 6344
rect 44039 6341 44051 6375
rect 43993 6335 44051 6341
rect 49145 6375 49203 6381
rect 49145 6341 49157 6375
rect 49191 6372 49203 6375
rect 49326 6372 49332 6384
rect 49191 6344 49332 6372
rect 49191 6341 49203 6344
rect 49145 6335 49203 6341
rect 49326 6332 49332 6344
rect 49384 6332 49390 6384
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 1581 6307 1639 6313
rect 1581 6304 1593 6307
rect 1360 6276 1593 6304
rect 1360 6264 1366 6276
rect 1581 6273 1593 6276
rect 1627 6304 1639 6307
rect 2317 6307 2375 6313
rect 2317 6304 2329 6307
rect 1627 6276 2329 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 2317 6273 2329 6276
rect 2363 6273 2375 6307
rect 2317 6267 2375 6273
rect 17862 6264 17868 6316
rect 17920 6304 17926 6316
rect 18325 6307 18383 6313
rect 18325 6304 18337 6307
rect 17920 6276 18337 6304
rect 17920 6264 17926 6276
rect 18325 6273 18337 6276
rect 18371 6273 18383 6307
rect 18325 6267 18383 6273
rect 18782 6264 18788 6316
rect 18840 6304 18846 6316
rect 19245 6307 19303 6313
rect 19245 6304 19257 6307
rect 18840 6276 19257 6304
rect 18840 6264 18846 6276
rect 19245 6273 19257 6276
rect 19291 6273 19303 6307
rect 19245 6267 19303 6273
rect 19426 6264 19432 6316
rect 19484 6304 19490 6316
rect 20533 6307 20591 6313
rect 20533 6304 20545 6307
rect 19484 6276 20545 6304
rect 19484 6264 19490 6276
rect 20533 6273 20545 6276
rect 20579 6273 20591 6307
rect 20533 6267 20591 6273
rect 42702 6264 42708 6316
rect 42760 6304 42766 6316
rect 47949 6307 48007 6313
rect 47949 6304 47961 6307
rect 42760 6276 47961 6304
rect 42760 6264 42766 6276
rect 47949 6273 47961 6276
rect 47995 6273 48007 6307
rect 47949 6267 48007 6273
rect 28442 6196 28448 6248
rect 28500 6236 28506 6248
rect 36906 6236 36912 6248
rect 28500 6208 36912 6236
rect 28500 6196 28506 6208
rect 36906 6196 36912 6208
rect 36964 6196 36970 6248
rect 1765 6171 1823 6177
rect 1765 6137 1777 6171
rect 1811 6168 1823 6171
rect 10042 6168 10048 6180
rect 1811 6140 10048 6168
rect 1811 6137 1823 6140
rect 1765 6131 1823 6137
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 18141 6171 18199 6177
rect 18141 6137 18153 6171
rect 18187 6168 18199 6171
rect 21174 6168 21180 6180
rect 18187 6140 21180 6168
rect 18187 6137 18199 6140
rect 18141 6131 18199 6137
rect 21174 6128 21180 6140
rect 21232 6128 21238 6180
rect 26050 6128 26056 6180
rect 26108 6168 26114 6180
rect 35802 6168 35808 6180
rect 26108 6140 35808 6168
rect 26108 6128 26114 6140
rect 35802 6128 35808 6140
rect 35860 6128 35866 6180
rect 44177 6171 44235 6177
rect 44177 6137 44189 6171
rect 44223 6168 44235 6171
rect 46934 6168 46940 6180
rect 44223 6140 46940 6168
rect 44223 6137 44235 6140
rect 44177 6131 44235 6137
rect 46934 6128 46940 6140
rect 46992 6128 46998 6180
rect 20349 6103 20407 6109
rect 20349 6069 20361 6103
rect 20395 6100 20407 6103
rect 22738 6100 22744 6112
rect 20395 6072 22744 6100
rect 20395 6069 20407 6072
rect 20349 6063 20407 6069
rect 22738 6060 22744 6072
rect 22796 6060 22802 6112
rect 37642 6060 37648 6112
rect 37700 6060 37706 6112
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 37642 5856 37648 5908
rect 37700 5896 37706 5908
rect 47302 5896 47308 5908
rect 37700 5868 47308 5896
rect 37700 5856 37706 5868
rect 47302 5856 47308 5868
rect 47360 5856 47366 5908
rect 1765 5831 1823 5837
rect 1765 5797 1777 5831
rect 1811 5828 1823 5831
rect 13446 5828 13452 5840
rect 1811 5800 13452 5828
rect 1811 5797 1823 5800
rect 1765 5791 1823 5797
rect 13446 5788 13452 5800
rect 13504 5788 13510 5840
rect 3053 5763 3111 5769
rect 3053 5760 3065 5763
rect 1596 5732 3065 5760
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 1596 5701 1624 5732
rect 3053 5729 3065 5732
rect 3099 5729 3111 5763
rect 3053 5723 3111 5729
rect 49145 5763 49203 5769
rect 49145 5729 49157 5763
rect 49191 5760 49203 5763
rect 49234 5760 49240 5772
rect 49191 5732 49240 5760
rect 49191 5729 49203 5732
rect 49145 5723 49203 5729
rect 49234 5720 49240 5732
rect 49292 5720 49298 5772
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1360 5664 1593 5692
rect 1360 5652 1366 5664
rect 1581 5661 1593 5664
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5692 2375 5695
rect 2774 5692 2780 5704
rect 2363 5664 2780 5692
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 2774 5652 2780 5664
rect 2832 5692 2838 5704
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 2832 5664 2881 5692
rect 2832 5652 2838 5664
rect 2869 5661 2881 5664
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 40034 5652 40040 5704
rect 40092 5692 40098 5704
rect 43717 5695 43775 5701
rect 43717 5692 43729 5695
rect 40092 5664 43729 5692
rect 40092 5652 40098 5664
rect 43717 5661 43729 5664
rect 43763 5661 43775 5695
rect 43717 5655 43775 5661
rect 47578 5652 47584 5704
rect 47636 5692 47642 5704
rect 47949 5695 48007 5701
rect 47949 5692 47961 5695
rect 47636 5664 47961 5692
rect 47636 5652 47642 5664
rect 47949 5661 47961 5664
rect 47995 5661 48007 5695
rect 47949 5655 48007 5661
rect 15470 5624 15476 5636
rect 2516 5596 15476 5624
rect 2516 5565 2544 5596
rect 15470 5584 15476 5596
rect 15528 5584 15534 5636
rect 43901 5627 43959 5633
rect 43901 5593 43913 5627
rect 43947 5624 43959 5627
rect 45830 5624 45836 5636
rect 43947 5596 45836 5624
rect 43947 5593 43959 5596
rect 43901 5587 43959 5593
rect 45830 5584 45836 5596
rect 45888 5584 45894 5636
rect 2501 5559 2559 5565
rect 2501 5525 2513 5559
rect 2547 5525 2559 5559
rect 2501 5519 2559 5525
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 24026 5556 24032 5568
rect 19392 5528 24032 5556
rect 19392 5516 19398 5528
rect 24026 5516 24032 5528
rect 24084 5516 24090 5568
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 37274 5312 37280 5364
rect 37332 5352 37338 5364
rect 37369 5355 37427 5361
rect 37369 5352 37381 5355
rect 37332 5324 37381 5352
rect 37332 5312 37338 5324
rect 37369 5321 37381 5324
rect 37415 5321 37427 5355
rect 37369 5315 37427 5321
rect 31294 5244 31300 5296
rect 31352 5284 31358 5296
rect 38565 5287 38623 5293
rect 38565 5284 38577 5287
rect 31352 5256 38577 5284
rect 31352 5244 31358 5256
rect 38565 5253 38577 5256
rect 38611 5284 38623 5287
rect 39025 5287 39083 5293
rect 39025 5284 39037 5287
rect 38611 5256 39037 5284
rect 38611 5253 38623 5256
rect 38565 5247 38623 5253
rect 39025 5253 39037 5256
rect 39071 5253 39083 5287
rect 39025 5247 39083 5253
rect 49142 5244 49148 5296
rect 49200 5244 49206 5296
rect 37274 5176 37280 5228
rect 37332 5216 37338 5228
rect 37829 5219 37887 5225
rect 37829 5216 37841 5219
rect 37332 5188 37841 5216
rect 37332 5176 37338 5188
rect 37829 5185 37841 5188
rect 37875 5185 37887 5219
rect 37829 5179 37887 5185
rect 45738 5176 45744 5228
rect 45796 5216 45802 5228
rect 45833 5219 45891 5225
rect 45833 5216 45845 5219
rect 45796 5188 45845 5216
rect 45796 5176 45802 5188
rect 45833 5185 45845 5188
rect 45879 5185 45891 5219
rect 45833 5179 45891 5185
rect 47210 5176 47216 5228
rect 47268 5216 47274 5228
rect 47949 5219 48007 5225
rect 47949 5216 47961 5219
rect 47268 5188 47961 5216
rect 47268 5176 47274 5188
rect 47949 5185 47961 5188
rect 47995 5185 48007 5219
rect 47949 5179 48007 5185
rect 1302 5108 1308 5160
rect 1360 5148 1366 5160
rect 1581 5151 1639 5157
rect 1581 5148 1593 5151
rect 1360 5120 1593 5148
rect 1360 5108 1366 5120
rect 1581 5117 1593 5120
rect 1627 5117 1639 5151
rect 1581 5111 1639 5117
rect 1857 5151 1915 5157
rect 1857 5117 1869 5151
rect 1903 5148 1915 5151
rect 10778 5148 10784 5160
rect 1903 5120 10784 5148
rect 1903 5117 1915 5120
rect 1857 5111 1915 5117
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 46845 5151 46903 5157
rect 46845 5117 46857 5151
rect 46891 5148 46903 5151
rect 48314 5148 48320 5160
rect 46891 5120 48320 5148
rect 46891 5117 46903 5120
rect 46845 5111 46903 5117
rect 48314 5108 48320 5120
rect 48372 5108 48378 5160
rect 38749 5083 38807 5089
rect 38749 5049 38761 5083
rect 38795 5080 38807 5083
rect 40034 5080 40040 5092
rect 38795 5052 40040 5080
rect 38795 5049 38807 5052
rect 38749 5043 38807 5049
rect 40034 5040 40040 5052
rect 40092 5040 40098 5092
rect 37918 4972 37924 5024
rect 37976 4972 37982 5024
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 1302 4768 1308 4820
rect 1360 4808 1366 4820
rect 2133 4811 2191 4817
rect 2133 4808 2145 4811
rect 1360 4780 2145 4808
rect 1360 4768 1366 4780
rect 2133 4777 2145 4780
rect 2179 4777 2191 4811
rect 2133 4771 2191 4777
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 22370 4808 22376 4820
rect 5592 4780 22376 4808
rect 5592 4768 5598 4780
rect 22370 4768 22376 4780
rect 22428 4768 22434 4820
rect 36906 4768 36912 4820
rect 36964 4768 36970 4820
rect 37918 4768 37924 4820
rect 37976 4808 37982 4820
rect 47210 4808 47216 4820
rect 37976 4780 47216 4808
rect 37976 4768 37982 4780
rect 47210 4768 47216 4780
rect 47268 4768 47274 4820
rect 31662 4740 31668 4752
rect 25240 4712 31668 4740
rect 25240 4681 25268 4712
rect 31662 4700 31668 4712
rect 31720 4700 31726 4752
rect 25225 4675 25283 4681
rect 25225 4641 25237 4675
rect 25271 4641 25283 4675
rect 25225 4635 25283 4641
rect 26234 4632 26240 4684
rect 26292 4632 26298 4684
rect 49145 4675 49203 4681
rect 49145 4641 49157 4675
rect 49191 4672 49203 4675
rect 49418 4672 49424 4684
rect 49191 4644 49424 4672
rect 49191 4641 49203 4644
rect 49145 4635 49203 4641
rect 49418 4632 49424 4644
rect 49476 4632 49482 4684
rect 1302 4564 1308 4616
rect 1360 4604 1366 4616
rect 1581 4607 1639 4613
rect 1581 4604 1593 4607
rect 1360 4576 1593 4604
rect 1360 4564 1366 4576
rect 1581 4573 1593 4576
rect 1627 4604 1639 4607
rect 2317 4607 2375 4613
rect 2317 4604 2329 4607
rect 1627 4576 2329 4604
rect 1627 4573 1639 4576
rect 1581 4567 1639 4573
rect 2317 4573 2329 4576
rect 2363 4573 2375 4607
rect 2317 4567 2375 4573
rect 22240 4607 22298 4613
rect 22240 4573 22252 4607
rect 22286 4604 22298 4607
rect 22462 4604 22468 4616
rect 22286 4576 22468 4604
rect 22286 4573 22298 4576
rect 22240 4567 22298 4573
rect 22462 4564 22468 4576
rect 22520 4564 22526 4616
rect 22646 4564 22652 4616
rect 22704 4604 22710 4616
rect 22868 4607 22926 4613
rect 22868 4604 22880 4607
rect 22704 4576 22880 4604
rect 22704 4564 22710 4576
rect 22868 4573 22880 4576
rect 22914 4573 22926 4607
rect 22868 4567 22926 4573
rect 23290 4564 23296 4616
rect 23348 4604 23354 4616
rect 23696 4607 23754 4613
rect 23696 4604 23708 4607
rect 23348 4576 23708 4604
rect 23348 4564 23354 4576
rect 23696 4573 23708 4576
rect 23742 4573 23754 4607
rect 23696 4567 23754 4573
rect 27062 4564 27068 4616
rect 27120 4604 27126 4616
rect 38105 4607 38163 4613
rect 38105 4604 38117 4607
rect 27120 4576 38117 4604
rect 27120 4564 27126 4576
rect 38105 4573 38117 4576
rect 38151 4604 38163 4607
rect 38565 4607 38623 4613
rect 38565 4604 38577 4607
rect 38151 4576 38577 4604
rect 38151 4573 38163 4576
rect 38105 4567 38163 4573
rect 38565 4573 38577 4576
rect 38611 4573 38623 4607
rect 38565 4567 38623 4573
rect 47026 4564 47032 4616
rect 47084 4604 47090 4616
rect 47949 4607 48007 4613
rect 47949 4604 47961 4607
rect 47084 4576 47961 4604
rect 47084 4564 47090 4576
rect 47949 4573 47961 4576
rect 47995 4573 48007 4607
rect 47949 4567 48007 4573
rect 22327 4539 22385 4545
rect 1780 4508 6914 4536
rect 1780 4477 1808 4508
rect 1765 4471 1823 4477
rect 1765 4437 1777 4471
rect 1811 4437 1823 4471
rect 6886 4468 6914 4508
rect 22327 4505 22339 4539
rect 22373 4536 22385 4539
rect 23566 4536 23572 4548
rect 22373 4508 23572 4536
rect 22373 4505 22385 4508
rect 22327 4499 22385 4505
rect 23566 4496 23572 4508
rect 23624 4496 23630 4548
rect 23799 4539 23857 4545
rect 23799 4505 23811 4539
rect 23845 4536 23857 4539
rect 25409 4539 25467 4545
rect 25409 4536 25421 4539
rect 23845 4508 25421 4536
rect 23845 4505 23857 4508
rect 23799 4499 23857 4505
rect 25409 4505 25421 4508
rect 25455 4505 25467 4539
rect 25409 4499 25467 4505
rect 36906 4496 36912 4548
rect 36964 4536 36970 4548
rect 37369 4539 37427 4545
rect 37369 4536 37381 4539
rect 36964 4508 37381 4536
rect 36964 4496 36970 4508
rect 37369 4505 37381 4508
rect 37415 4505 37427 4539
rect 37369 4499 37427 4505
rect 38289 4539 38347 4545
rect 38289 4505 38301 4539
rect 38335 4536 38347 4539
rect 38335 4508 41414 4536
rect 38335 4505 38347 4508
rect 38289 4499 38347 4505
rect 19334 4468 19340 4480
rect 6886 4440 19340 4468
rect 1765 4431 1823 4437
rect 19334 4428 19340 4440
rect 19392 4428 19398 4480
rect 22971 4471 23029 4477
rect 22971 4437 22983 4471
rect 23017 4468 23029 4471
rect 24026 4468 24032 4480
rect 23017 4440 24032 4468
rect 23017 4437 23029 4440
rect 22971 4431 23029 4437
rect 24026 4428 24032 4440
rect 24084 4428 24090 4480
rect 24213 4471 24271 4477
rect 24213 4437 24225 4471
rect 24259 4468 24271 4471
rect 24762 4468 24768 4480
rect 24259 4440 24768 4468
rect 24259 4437 24271 4440
rect 24213 4431 24271 4437
rect 24762 4428 24768 4440
rect 24820 4428 24826 4480
rect 37461 4471 37519 4477
rect 37461 4437 37473 4471
rect 37507 4468 37519 4471
rect 39390 4468 39396 4480
rect 37507 4440 39396 4468
rect 37507 4437 37519 4440
rect 37461 4431 37519 4437
rect 39390 4428 39396 4440
rect 39448 4428 39454 4480
rect 41386 4468 41414 4508
rect 44450 4468 44456 4480
rect 41386 4440 44456 4468
rect 44450 4428 44456 4440
rect 44508 4428 44514 4480
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 23658 4264 23664 4276
rect 23584 4236 23664 4264
rect 1394 4156 1400 4208
rect 1452 4196 1458 4208
rect 1673 4199 1731 4205
rect 1673 4196 1685 4199
rect 1452 4168 1685 4196
rect 1452 4156 1458 4168
rect 1673 4165 1685 4168
rect 1719 4196 1731 4199
rect 23584 4196 23612 4236
rect 23658 4224 23664 4236
rect 23716 4264 23722 4276
rect 24762 4264 24768 4276
rect 23716 4236 24768 4264
rect 23716 4224 23722 4236
rect 24762 4224 24768 4236
rect 24820 4224 24826 4276
rect 1719 4168 2452 4196
rect 23506 4168 23612 4196
rect 1719 4165 1731 4168
rect 1673 4159 1731 4165
rect 1302 4088 1308 4140
rect 1360 4128 1366 4140
rect 2317 4131 2375 4137
rect 2317 4128 2329 4131
rect 1360 4100 2329 4128
rect 1360 4088 1366 4100
rect 2317 4097 2329 4100
rect 2363 4097 2375 4131
rect 2424 4128 2452 4168
rect 24026 4156 24032 4208
rect 24084 4196 24090 4208
rect 24489 4199 24547 4205
rect 24489 4196 24501 4199
rect 24084 4168 24501 4196
rect 24084 4156 24090 4168
rect 24489 4165 24501 4168
rect 24535 4165 24547 4199
rect 24489 4159 24547 4165
rect 27338 4156 27344 4208
rect 27396 4156 27402 4208
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 2424 4100 3065 4128
rect 2317 4091 2375 4097
rect 3053 4097 3065 4100
rect 3099 4097 3111 4131
rect 3053 4091 3111 4097
rect 2332 4060 2360 4091
rect 16482 4088 16488 4140
rect 16540 4128 16546 4140
rect 18325 4131 18383 4137
rect 18325 4128 18337 4131
rect 16540 4100 18337 4128
rect 16540 4088 16546 4100
rect 18325 4097 18337 4100
rect 18371 4097 18383 4131
rect 18325 4091 18383 4097
rect 27154 4088 27160 4140
rect 27212 4088 27218 4140
rect 34238 4088 34244 4140
rect 34296 4128 34302 4140
rect 39206 4128 39212 4140
rect 34296 4100 39212 4128
rect 34296 4088 34302 4100
rect 39206 4088 39212 4100
rect 39264 4088 39270 4140
rect 39298 4088 39304 4140
rect 39356 4128 39362 4140
rect 45833 4131 45891 4137
rect 45833 4128 45845 4131
rect 39356 4100 45845 4128
rect 39356 4088 39362 4100
rect 45833 4097 45845 4100
rect 45879 4097 45891 4131
rect 45833 4091 45891 4097
rect 47118 4088 47124 4140
rect 47176 4128 47182 4140
rect 47949 4131 48007 4137
rect 47949 4128 47961 4131
rect 47176 4100 47961 4128
rect 47176 4088 47182 4100
rect 47949 4097 47961 4100
rect 47995 4097 48007 4131
rect 47949 4091 48007 4097
rect 49145 4131 49203 4137
rect 49145 4097 49157 4131
rect 49191 4128 49203 4131
rect 49326 4128 49332 4140
rect 49191 4100 49332 4128
rect 49191 4097 49203 4100
rect 49145 4091 49203 4097
rect 49326 4088 49332 4100
rect 49384 4088 49390 4140
rect 2869 4063 2927 4069
rect 2869 4060 2881 4063
rect 2332 4032 2881 4060
rect 2869 4029 2881 4032
rect 2915 4029 2927 4063
rect 17770 4060 17776 4072
rect 2869 4023 2927 4029
rect 6886 4032 17776 4060
rect 2501 3995 2559 4001
rect 2501 3961 2513 3995
rect 2547 3992 2559 3995
rect 6886 3992 6914 4032
rect 17770 4020 17776 4032
rect 17828 4020 17834 4072
rect 18509 4063 18567 4069
rect 18509 4029 18521 4063
rect 18555 4029 18567 4063
rect 18509 4023 18567 4029
rect 2547 3964 6914 3992
rect 2547 3961 2559 3964
rect 2501 3955 2559 3961
rect 16482 3952 16488 4004
rect 16540 3992 16546 4004
rect 18524 3992 18552 4023
rect 20162 4020 20168 4072
rect 20220 4020 20226 4072
rect 22002 4020 22008 4072
rect 22060 4020 22066 4072
rect 22278 4020 22284 4072
rect 22336 4020 22342 4072
rect 24305 4063 24363 4069
rect 24305 4029 24317 4063
rect 24351 4029 24363 4063
rect 24305 4023 24363 4029
rect 16540 3964 22094 3992
rect 16540 3952 16546 3964
rect 1765 3927 1823 3933
rect 1765 3893 1777 3927
rect 1811 3924 1823 3927
rect 5534 3924 5540 3936
rect 1811 3896 5540 3924
rect 1811 3893 1823 3896
rect 1765 3887 1823 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 20714 3924 20720 3936
rect 7524 3896 20720 3924
rect 7524 3884 7530 3896
rect 20714 3884 20720 3896
rect 20772 3884 20778 3936
rect 22066 3924 22094 3964
rect 22462 3924 22468 3936
rect 22066 3896 22468 3924
rect 22462 3884 22468 3896
rect 22520 3884 22526 3936
rect 23658 3884 23664 3936
rect 23716 3924 23722 3936
rect 23753 3927 23811 3933
rect 23753 3924 23765 3927
rect 23716 3896 23765 3924
rect 23716 3884 23722 3896
rect 23753 3893 23765 3896
rect 23799 3893 23811 3927
rect 24320 3924 24348 4023
rect 24486 4020 24492 4072
rect 24544 4060 24550 4072
rect 25682 4060 25688 4072
rect 24544 4032 25688 4060
rect 24544 4020 24550 4032
rect 25682 4020 25688 4032
rect 25740 4020 25746 4072
rect 27617 4063 27675 4069
rect 27617 4060 27629 4063
rect 25792 4032 27629 4060
rect 24394 3952 24400 4004
rect 24452 3992 24458 4004
rect 25792 3992 25820 4032
rect 27617 4029 27629 4032
rect 27663 4029 27675 4063
rect 27617 4023 27675 4029
rect 46658 4020 46664 4072
rect 46716 4020 46722 4072
rect 24452 3964 25820 3992
rect 24452 3952 24458 3964
rect 27154 3952 27160 4004
rect 27212 3992 27218 4004
rect 33594 3992 33600 4004
rect 27212 3964 33600 3992
rect 27212 3952 27218 3964
rect 33594 3952 33600 3964
rect 33652 3952 33658 4004
rect 30650 3924 30656 3936
rect 24320 3896 30656 3924
rect 23753 3887 23811 3893
rect 30650 3884 30656 3896
rect 30708 3884 30714 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 5350 3680 5356 3732
rect 5408 3720 5414 3732
rect 20073 3723 20131 3729
rect 5408 3692 17724 3720
rect 5408 3680 5414 3692
rect 15378 3612 15384 3664
rect 15436 3652 15442 3664
rect 17589 3655 17647 3661
rect 17589 3652 17601 3655
rect 15436 3624 17601 3652
rect 15436 3612 15442 3624
rect 17589 3621 17601 3624
rect 17635 3621 17647 3655
rect 17589 3615 17647 3621
rect 1118 3544 1124 3596
rect 1176 3584 1182 3596
rect 17218 3584 17224 3596
rect 1176 3556 17224 3584
rect 1176 3544 1182 3556
rect 17218 3544 17224 3556
rect 17276 3544 17282 3596
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1581 3519 1639 3525
rect 1581 3516 1593 3519
rect 1360 3488 1593 3516
rect 1360 3476 1366 3488
rect 1581 3485 1593 3488
rect 1627 3485 1639 3519
rect 1581 3479 1639 3485
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 7558 3516 7564 3528
rect 1903 3488 7564 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 7558 3476 7564 3488
rect 7616 3476 7622 3528
rect 16482 3476 16488 3528
rect 16540 3476 16546 3528
rect 17696 3448 17724 3692
rect 20073 3689 20085 3723
rect 20119 3720 20131 3723
rect 22278 3720 22284 3732
rect 20119 3692 22284 3720
rect 20119 3689 20131 3692
rect 20073 3683 20131 3689
rect 22278 3680 22284 3692
rect 22336 3680 22342 3732
rect 23983 3723 24041 3729
rect 23983 3689 23995 3723
rect 24029 3720 24041 3723
rect 27338 3720 27344 3732
rect 24029 3692 27344 3720
rect 24029 3689 24041 3692
rect 23983 3683 24041 3689
rect 27338 3680 27344 3692
rect 27396 3680 27402 3732
rect 36541 3723 36599 3729
rect 36541 3689 36553 3723
rect 36587 3720 36599 3723
rect 39298 3720 39304 3732
rect 36587 3692 39304 3720
rect 36587 3689 36599 3692
rect 36541 3683 36599 3689
rect 39298 3680 39304 3692
rect 39356 3680 39362 3732
rect 20714 3612 20720 3664
rect 20772 3652 20778 3664
rect 21910 3652 21916 3664
rect 20772 3624 21916 3652
rect 20772 3612 20778 3624
rect 21910 3612 21916 3624
rect 21968 3652 21974 3664
rect 21968 3624 25084 3652
rect 21968 3612 21974 3624
rect 19794 3584 19800 3596
rect 17788 3556 19800 3584
rect 17788 3525 17816 3556
rect 19794 3544 19800 3556
rect 19852 3544 19858 3596
rect 21174 3544 21180 3596
rect 21232 3544 21238 3596
rect 21361 3587 21419 3593
rect 21361 3553 21373 3587
rect 21407 3584 21419 3587
rect 22094 3584 22100 3596
rect 21407 3556 22100 3584
rect 21407 3553 21419 3556
rect 21361 3547 21419 3553
rect 22094 3544 22100 3556
rect 22152 3584 22158 3596
rect 23290 3584 23296 3596
rect 22152 3556 23296 3584
rect 22152 3544 22158 3556
rect 23290 3544 23296 3556
rect 23348 3544 23354 3596
rect 23566 3544 23572 3596
rect 23624 3584 23630 3596
rect 25056 3593 25084 3624
rect 36998 3612 37004 3664
rect 37056 3652 37062 3664
rect 45554 3652 45560 3664
rect 37056 3624 45560 3652
rect 37056 3612 37062 3624
rect 45554 3612 45560 3624
rect 45612 3612 45618 3664
rect 24765 3587 24823 3593
rect 24765 3584 24777 3587
rect 23624 3556 24777 3584
rect 23624 3544 23630 3556
rect 24765 3553 24777 3556
rect 24811 3553 24823 3587
rect 24765 3547 24823 3553
rect 25041 3587 25099 3593
rect 25041 3553 25053 3587
rect 25087 3553 25099 3587
rect 25041 3547 25099 3553
rect 34514 3544 34520 3596
rect 34572 3584 34578 3596
rect 47670 3584 47676 3596
rect 34572 3556 47676 3584
rect 34572 3544 34578 3556
rect 47670 3544 47676 3556
rect 47728 3544 47734 3596
rect 49142 3544 49148 3596
rect 49200 3544 49206 3596
rect 17773 3519 17831 3525
rect 17773 3485 17785 3519
rect 17819 3485 17831 3519
rect 17773 3479 17831 3485
rect 19426 3476 19432 3528
rect 19484 3476 19490 3528
rect 22922 3476 22928 3528
rect 22980 3516 22986 3528
rect 23880 3519 23938 3525
rect 23880 3516 23892 3519
rect 22980 3488 23892 3516
rect 22980 3476 22986 3488
rect 23880 3485 23892 3488
rect 23926 3485 23938 3519
rect 23880 3479 23938 3485
rect 24581 3519 24639 3525
rect 24581 3485 24593 3519
rect 24627 3485 24639 3519
rect 24581 3479 24639 3485
rect 23017 3451 23075 3457
rect 17696 3420 22094 3448
rect 12526 3340 12532 3392
rect 12584 3380 12590 3392
rect 16577 3383 16635 3389
rect 16577 3380 16589 3383
rect 12584 3352 16589 3380
rect 12584 3340 12590 3352
rect 16577 3349 16589 3352
rect 16623 3349 16635 3383
rect 22066 3380 22094 3420
rect 23017 3417 23029 3451
rect 23063 3448 23075 3451
rect 24394 3448 24400 3460
rect 23063 3420 24400 3448
rect 23063 3417 23075 3420
rect 23017 3411 23075 3417
rect 24394 3408 24400 3420
rect 24452 3408 24458 3460
rect 24486 3380 24492 3392
rect 22066 3352 24492 3380
rect 16577 3343 16635 3349
rect 24486 3340 24492 3352
rect 24544 3340 24550 3392
rect 24596 3380 24624 3479
rect 35802 3476 35808 3528
rect 35860 3516 35866 3528
rect 36449 3519 36507 3525
rect 36449 3516 36461 3519
rect 35860 3488 36461 3516
rect 35860 3476 35866 3488
rect 36449 3485 36461 3488
rect 36495 3516 36507 3519
rect 36909 3519 36967 3525
rect 36909 3516 36921 3519
rect 36495 3488 36921 3516
rect 36495 3485 36507 3488
rect 36449 3479 36507 3485
rect 36909 3485 36921 3488
rect 36955 3485 36967 3519
rect 36909 3479 36967 3485
rect 40034 3476 40040 3528
rect 40092 3516 40098 3528
rect 46109 3519 46167 3525
rect 46109 3516 46121 3519
rect 40092 3488 46121 3516
rect 40092 3476 40098 3488
rect 46109 3485 46121 3488
rect 46155 3485 46167 3519
rect 46109 3479 46167 3485
rect 46934 3476 46940 3528
rect 46992 3516 46998 3528
rect 47949 3519 48007 3525
rect 47949 3516 47961 3519
rect 46992 3488 47961 3516
rect 46992 3476 46998 3488
rect 47949 3485 47961 3488
rect 47995 3485 48007 3519
rect 47949 3479 48007 3485
rect 40862 3408 40868 3460
rect 40920 3448 40926 3460
rect 43438 3448 43444 3460
rect 40920 3420 43444 3448
rect 40920 3408 40926 3420
rect 43438 3408 43444 3420
rect 43496 3408 43502 3460
rect 47305 3451 47363 3457
rect 47305 3417 47317 3451
rect 47351 3448 47363 3451
rect 48682 3448 48688 3460
rect 47351 3420 48688 3448
rect 47351 3417 47363 3420
rect 47305 3411 47363 3417
rect 48682 3408 48688 3420
rect 48740 3408 48746 3460
rect 25866 3380 25872 3392
rect 24596 3352 25872 3380
rect 25866 3340 25872 3352
rect 25924 3340 25930 3392
rect 40954 3340 40960 3392
rect 41012 3380 41018 3392
rect 49786 3380 49792 3392
rect 41012 3352 49792 3380
rect 41012 3340 41018 3352
rect 49786 3340 49792 3352
rect 49844 3340 49850 3392
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 1302 3136 1308 3188
rect 1360 3176 1366 3188
rect 2133 3179 2191 3185
rect 2133 3176 2145 3179
rect 1360 3148 2145 3176
rect 1360 3136 1366 3148
rect 2133 3145 2145 3148
rect 2179 3145 2191 3179
rect 2133 3139 2191 3145
rect 17218 3136 17224 3188
rect 17276 3176 17282 3188
rect 24210 3176 24216 3188
rect 17276 3148 24216 3176
rect 17276 3136 17282 3148
rect 24210 3136 24216 3148
rect 24268 3136 24274 3188
rect 30742 3176 30748 3188
rect 29748 3148 30748 3176
rect 16114 3068 16120 3120
rect 16172 3108 16178 3120
rect 22094 3108 22100 3120
rect 16172 3080 17356 3108
rect 16172 3068 16178 3080
rect 1302 3000 1308 3052
rect 1360 3040 1366 3052
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 1360 3012 1593 3040
rect 1360 3000 1366 3012
rect 1581 3009 1593 3012
rect 1627 3040 1639 3043
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 1627 3012 2513 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 14274 3000 14280 3052
rect 14332 3040 14338 3052
rect 14553 3043 14611 3049
rect 14553 3040 14565 3043
rect 14332 3012 14565 3040
rect 14332 3000 14338 3012
rect 14553 3009 14565 3012
rect 14599 3009 14611 3043
rect 16390 3040 16396 3052
rect 15962 3012 16396 3040
rect 14553 3003 14611 3009
rect 16390 3000 16396 3012
rect 16448 3000 16454 3052
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 11054 2932 11060 2984
rect 11112 2972 11118 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 11112 2944 14841 2972
rect 11112 2932 11118 2944
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 1765 2907 1823 2913
rect 1765 2873 1777 2907
rect 1811 2904 1823 2907
rect 11238 2904 11244 2916
rect 1811 2876 11244 2904
rect 1811 2873 1823 2876
rect 1765 2867 1823 2873
rect 11238 2864 11244 2876
rect 11296 2864 11302 2916
rect 17052 2904 17080 3003
rect 17328 2981 17356 3080
rect 19076 3080 22100 3108
rect 19076 3049 19104 3080
rect 22094 3068 22100 3080
rect 22152 3068 22158 3120
rect 22922 3068 22928 3120
rect 22980 3068 22986 3120
rect 23658 3068 23664 3120
rect 23716 3108 23722 3120
rect 23716 3080 25084 3108
rect 23716 3068 23722 3080
rect 19061 3043 19119 3049
rect 19061 3009 19073 3043
rect 19107 3009 19119 3043
rect 19061 3003 19119 3009
rect 19518 3000 19524 3052
rect 19576 3040 19582 3052
rect 19613 3043 19671 3049
rect 19613 3040 19625 3043
rect 19576 3012 19625 3040
rect 19576 3000 19582 3012
rect 19613 3009 19625 3012
rect 19659 3009 19671 3043
rect 19613 3003 19671 3009
rect 22738 3000 22744 3052
rect 22796 3000 22802 3052
rect 25056 3049 25084 3080
rect 27706 3068 27712 3120
rect 27764 3108 27770 3120
rect 29748 3108 29776 3148
rect 30742 3136 30748 3148
rect 30800 3176 30806 3188
rect 31205 3179 31263 3185
rect 31205 3176 31217 3179
rect 30800 3148 31217 3176
rect 30800 3136 30806 3148
rect 31205 3145 31217 3148
rect 31251 3145 31263 3179
rect 31205 3139 31263 3145
rect 49145 3111 49203 3117
rect 27764 3080 29854 3108
rect 27764 3068 27770 3080
rect 49145 3077 49157 3111
rect 49191 3108 49203 3111
rect 49234 3108 49240 3120
rect 49191 3080 49240 3108
rect 49191 3077 49203 3080
rect 49145 3071 49203 3077
rect 49234 3068 49240 3080
rect 49292 3068 49298 3120
rect 25041 3043 25099 3049
rect 25041 3009 25053 3043
rect 25087 3009 25099 3043
rect 25041 3003 25099 3009
rect 27614 3000 27620 3052
rect 27672 3040 27678 3052
rect 27893 3043 27951 3049
rect 27893 3040 27905 3043
rect 27672 3012 27905 3040
rect 27672 3000 27678 3012
rect 27893 3009 27905 3012
rect 27939 3009 27951 3043
rect 27893 3003 27951 3009
rect 29086 3000 29092 3052
rect 29144 3000 29150 3052
rect 39390 3000 39396 3052
rect 39448 3040 39454 3052
rect 43993 3043 44051 3049
rect 43993 3040 44005 3043
rect 39448 3012 44005 3040
rect 39448 3000 39454 3012
rect 43993 3009 44005 3012
rect 44039 3009 44051 3043
rect 43993 3003 44051 3009
rect 45830 3000 45836 3052
rect 45888 3000 45894 3052
rect 47302 3000 47308 3052
rect 47360 3040 47366 3052
rect 47949 3043 48007 3049
rect 47949 3040 47961 3043
rect 47360 3012 47961 3040
rect 47360 3000 47366 3012
rect 47949 3009 47961 3012
rect 47995 3009 48007 3043
rect 47949 3003 48007 3009
rect 17313 2975 17371 2981
rect 17313 2941 17325 2975
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 19794 2932 19800 2984
rect 19852 2932 19858 2984
rect 21453 2975 21511 2981
rect 21453 2941 21465 2975
rect 21499 2972 21511 2975
rect 22278 2972 22284 2984
rect 21499 2944 22284 2972
rect 21499 2941 21511 2944
rect 21453 2935 21511 2941
rect 22278 2932 22284 2944
rect 22336 2932 22342 2984
rect 24581 2975 24639 2981
rect 24581 2941 24593 2975
rect 24627 2972 24639 2975
rect 26510 2972 26516 2984
rect 24627 2944 26516 2972
rect 24627 2941 24639 2944
rect 24581 2935 24639 2941
rect 26510 2932 26516 2944
rect 26568 2932 26574 2984
rect 28537 2975 28595 2981
rect 28537 2941 28549 2975
rect 28583 2972 28595 2975
rect 29365 2975 29423 2981
rect 29365 2972 29377 2975
rect 28583 2944 29377 2972
rect 28583 2941 28595 2944
rect 28537 2935 28595 2941
rect 29365 2941 29377 2944
rect 29411 2941 29423 2975
rect 29365 2935 29423 2941
rect 45189 2975 45247 2981
rect 45189 2941 45201 2975
rect 45235 2972 45247 2975
rect 46750 2972 46756 2984
rect 45235 2944 46756 2972
rect 45235 2941 45247 2944
rect 45189 2935 45247 2941
rect 46750 2932 46756 2944
rect 46808 2932 46814 2984
rect 46842 2932 46848 2984
rect 46900 2932 46906 2984
rect 18877 2907 18935 2913
rect 18877 2904 18889 2907
rect 17052 2876 18889 2904
rect 18877 2873 18889 2876
rect 18923 2873 18935 2907
rect 19812 2904 19840 2932
rect 22646 2904 22652 2916
rect 19812 2876 22652 2904
rect 18877 2867 18935 2873
rect 22646 2864 22652 2876
rect 22704 2904 22710 2916
rect 23382 2904 23388 2916
rect 22704 2876 23388 2904
rect 22704 2864 22710 2876
rect 23382 2864 23388 2876
rect 23440 2864 23446 2916
rect 2314 2796 2320 2848
rect 2372 2796 2378 2848
rect 2774 2796 2780 2848
rect 2832 2796 2838 2848
rect 3326 2796 3332 2848
rect 3384 2836 3390 2848
rect 8846 2836 8852 2848
rect 3384 2808 8852 2836
rect 3384 2796 3390 2808
rect 8846 2796 8852 2808
rect 8904 2796 8910 2848
rect 16301 2839 16359 2845
rect 16301 2805 16313 2839
rect 16347 2836 16359 2839
rect 19426 2836 19432 2848
rect 16347 2808 19432 2836
rect 16347 2805 16359 2808
rect 16301 2799 16359 2805
rect 19426 2796 19432 2808
rect 19484 2836 19490 2848
rect 20990 2836 20996 2848
rect 19484 2808 20996 2836
rect 19484 2796 19490 2808
rect 20990 2796 20996 2808
rect 21048 2796 21054 2848
rect 24854 2796 24860 2848
rect 24912 2836 24918 2848
rect 25685 2839 25743 2845
rect 25685 2836 25697 2839
rect 24912 2808 25697 2836
rect 24912 2796 24918 2808
rect 25685 2805 25697 2808
rect 25731 2805 25743 2839
rect 25685 2799 25743 2805
rect 30834 2796 30840 2848
rect 30892 2796 30898 2848
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 3053 2635 3111 2641
rect 3053 2601 3065 2635
rect 3099 2632 3111 2635
rect 9490 2632 9496 2644
rect 3099 2604 9496 2632
rect 3099 2601 3111 2604
rect 3053 2595 3111 2601
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 9677 2635 9735 2641
rect 9677 2601 9689 2635
rect 9723 2632 9735 2635
rect 11054 2632 11060 2644
rect 9723 2604 11060 2632
rect 9723 2601 9735 2604
rect 9677 2595 9735 2601
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 16390 2592 16396 2644
rect 16448 2592 16454 2644
rect 20990 2592 20996 2644
rect 21048 2592 21054 2644
rect 22741 2635 22799 2641
rect 22741 2601 22753 2635
rect 22787 2632 22799 2635
rect 23658 2632 23664 2644
rect 22787 2604 23664 2632
rect 22787 2601 22799 2604
rect 22741 2595 22799 2601
rect 23658 2592 23664 2604
rect 23716 2592 23722 2644
rect 23753 2635 23811 2641
rect 23753 2601 23765 2635
rect 23799 2632 23811 2635
rect 26329 2635 26387 2641
rect 26329 2632 26341 2635
rect 23799 2604 26341 2632
rect 23799 2601 23811 2604
rect 23753 2595 23811 2601
rect 26329 2601 26341 2604
rect 26375 2632 26387 2635
rect 27614 2632 27620 2644
rect 26375 2604 27620 2632
rect 26375 2601 26387 2604
rect 26329 2595 26387 2601
rect 27614 2592 27620 2604
rect 27672 2592 27678 2644
rect 27893 2635 27951 2641
rect 27893 2601 27905 2635
rect 27939 2601 27951 2635
rect 27893 2595 27951 2601
rect 2501 2567 2559 2573
rect 2501 2533 2513 2567
rect 2547 2564 2559 2567
rect 20898 2564 20904 2576
rect 2547 2536 6914 2564
rect 2547 2533 2559 2536
rect 2501 2527 2559 2533
rect 2774 2496 2780 2508
rect 1596 2468 2780 2496
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1596 2437 1624 2468
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 6886 2496 6914 2536
rect 9692 2536 20904 2564
rect 9692 2496 9720 2536
rect 20898 2524 20904 2536
rect 20956 2524 20962 2576
rect 21361 2567 21419 2573
rect 21361 2533 21373 2567
rect 21407 2564 21419 2567
rect 22830 2564 22836 2576
rect 21407 2536 22836 2564
rect 21407 2533 21419 2536
rect 21361 2527 21419 2533
rect 6886 2468 9720 2496
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 12253 2499 12311 2505
rect 12253 2496 12265 2499
rect 11756 2468 12265 2496
rect 11756 2456 11762 2468
rect 12253 2465 12265 2468
rect 12299 2465 12311 2499
rect 12253 2459 12311 2465
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 13872 2468 14749 2496
rect 13872 2456 13878 2468
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 21376 2496 21404 2527
rect 22830 2524 22836 2536
rect 22888 2524 22894 2576
rect 22925 2567 22983 2573
rect 22925 2533 22937 2567
rect 22971 2564 22983 2567
rect 23290 2564 23296 2576
rect 22971 2536 23296 2564
rect 22971 2533 22983 2536
rect 22925 2527 22983 2533
rect 23290 2524 23296 2536
rect 23348 2524 23354 2576
rect 23382 2524 23388 2576
rect 23440 2564 23446 2576
rect 23937 2567 23995 2573
rect 23937 2564 23949 2567
rect 23440 2536 23949 2564
rect 23440 2524 23446 2536
rect 23937 2533 23949 2536
rect 23983 2533 23995 2567
rect 23937 2527 23995 2533
rect 25866 2524 25872 2576
rect 25924 2564 25930 2576
rect 27430 2564 27436 2576
rect 25924 2536 27436 2564
rect 25924 2524 25930 2536
rect 27430 2524 27436 2536
rect 27488 2524 27494 2576
rect 27706 2564 27712 2576
rect 27540 2536 27712 2564
rect 14737 2459 14795 2465
rect 20456 2468 21404 2496
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 1360 2400 1593 2428
rect 1360 2388 1366 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 2314 2428 2320 2440
rect 1581 2391 1639 2397
rect 1688 2400 2320 2428
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 1688 2360 1716 2400
rect 2314 2388 2320 2400
rect 2372 2388 2378 2440
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3513 2431 3571 2437
rect 3513 2428 3525 2431
rect 3292 2400 3525 2428
rect 3292 2388 3298 2400
rect 3513 2397 3525 2400
rect 3559 2397 3571 2431
rect 3513 2391 3571 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9732 2400 9873 2428
rect 9732 2388 9738 2400
rect 9861 2397 9873 2400
rect 9907 2428 9919 2431
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 9907 2400 10149 2428
rect 9907 2397 9919 2400
rect 9861 2391 9919 2397
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 10137 2391 10195 2397
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2428 12035 2431
rect 12526 2428 12532 2440
rect 12023 2400 12532 2428
rect 12023 2397 12035 2400
rect 11977 2391 12035 2397
rect 12526 2388 12532 2400
rect 12584 2388 12590 2440
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2428 14519 2431
rect 15378 2428 15384 2440
rect 14507 2400 15384 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 15378 2388 15384 2400
rect 15436 2388 15442 2440
rect 20456 2437 20484 2468
rect 22002 2456 22008 2508
rect 22060 2496 22066 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 22060 2468 24593 2496
rect 22060 2456 22066 2468
rect 24581 2465 24593 2468
rect 24627 2465 24639 2499
rect 24581 2459 24639 2465
rect 24854 2456 24860 2508
rect 24912 2456 24918 2508
rect 24946 2456 24952 2508
rect 25004 2496 25010 2508
rect 26697 2499 26755 2505
rect 26697 2496 26709 2499
rect 25004 2468 26709 2496
rect 25004 2456 25010 2468
rect 26697 2465 26709 2468
rect 26743 2496 26755 2499
rect 27540 2496 27568 2536
rect 27706 2524 27712 2536
rect 27764 2524 27770 2576
rect 27908 2564 27936 2595
rect 31662 2592 31668 2644
rect 31720 2632 31726 2644
rect 32953 2635 33011 2641
rect 32953 2632 32965 2635
rect 31720 2604 32965 2632
rect 31720 2592 31726 2604
rect 32953 2601 32965 2604
rect 32999 2601 33011 2635
rect 32953 2595 33011 2601
rect 33594 2592 33600 2644
rect 33652 2632 33658 2644
rect 35069 2635 35127 2641
rect 35069 2632 35081 2635
rect 33652 2604 35081 2632
rect 33652 2592 33658 2604
rect 35069 2601 35081 2604
rect 35115 2601 35127 2635
rect 35069 2595 35127 2601
rect 30834 2564 30840 2576
rect 27908 2536 30840 2564
rect 30834 2524 30840 2536
rect 30892 2564 30898 2576
rect 30892 2536 40724 2564
rect 30892 2524 30898 2536
rect 37737 2499 37795 2505
rect 37737 2496 37749 2499
rect 26743 2468 27568 2496
rect 27632 2468 37749 2496
rect 26743 2465 26755 2468
rect 26697 2459 26755 2465
rect 27632 2437 27660 2468
rect 37737 2465 37749 2468
rect 37783 2465 37795 2499
rect 37737 2459 37795 2465
rect 17681 2431 17739 2437
rect 17681 2397 17693 2431
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 20441 2431 20499 2437
rect 20441 2397 20453 2431
rect 20487 2397 20499 2431
rect 20441 2391 20499 2397
rect 20901 2431 20959 2437
rect 20901 2397 20913 2431
rect 20947 2428 20959 2431
rect 22465 2431 22523 2437
rect 22465 2428 22477 2431
rect 20947 2400 22477 2428
rect 20947 2397 20959 2400
rect 20901 2391 20959 2397
rect 22465 2397 22477 2400
rect 22511 2428 22523 2431
rect 23477 2431 23535 2437
rect 23477 2428 23489 2431
rect 22511 2400 23489 2428
rect 22511 2397 22523 2400
rect 22465 2391 22523 2397
rect 23477 2397 23489 2400
rect 23523 2428 23535 2431
rect 27617 2431 27675 2437
rect 27617 2428 27629 2431
rect 23523 2400 24072 2428
rect 23523 2397 23535 2400
rect 23477 2391 23535 2397
rect 10594 2360 10600 2372
rect 1268 2332 1716 2360
rect 1780 2332 10600 2360
rect 1268 2320 1274 2332
rect 1780 2301 1808 2332
rect 10594 2320 10600 2332
rect 10652 2320 10658 2372
rect 1765 2295 1823 2301
rect 1765 2261 1777 2295
rect 1811 2261 1823 2295
rect 1765 2255 1823 2261
rect 9490 2252 9496 2304
rect 9548 2292 9554 2304
rect 12342 2292 12348 2304
rect 9548 2264 12348 2292
rect 9548 2252 9554 2264
rect 12342 2252 12348 2264
rect 12400 2252 12406 2304
rect 17696 2292 17724 2391
rect 18322 2320 18328 2372
rect 18380 2360 18386 2372
rect 18417 2363 18475 2369
rect 18417 2360 18429 2363
rect 18380 2332 18429 2360
rect 18380 2320 18386 2332
rect 18417 2329 18429 2332
rect 18463 2329 18475 2363
rect 18417 2323 18475 2329
rect 20257 2295 20315 2301
rect 20257 2292 20269 2295
rect 17696 2264 20269 2292
rect 20257 2261 20269 2264
rect 20303 2261 20315 2295
rect 24044 2292 24072 2400
rect 26206 2400 27629 2428
rect 24854 2320 24860 2372
rect 24912 2360 24918 2372
rect 26206 2360 26234 2400
rect 27617 2397 27629 2400
rect 27663 2397 27675 2431
rect 27617 2391 27675 2397
rect 28626 2388 28632 2440
rect 28684 2428 28690 2440
rect 28905 2431 28963 2437
rect 28905 2428 28917 2431
rect 28684 2400 28917 2428
rect 28684 2388 28690 2400
rect 28905 2397 28917 2400
rect 28951 2428 28963 2431
rect 29181 2431 29239 2437
rect 29181 2428 29193 2431
rect 28951 2400 29193 2428
rect 28951 2397 28963 2400
rect 28905 2391 28963 2397
rect 29181 2397 29193 2400
rect 29227 2397 29239 2431
rect 29181 2391 29239 2397
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30800 2400 31033 2428
rect 30800 2388 30806 2400
rect 31021 2397 31033 2400
rect 31067 2428 31079 2431
rect 31297 2431 31355 2437
rect 31297 2428 31309 2431
rect 31067 2400 31309 2428
rect 31067 2397 31079 2400
rect 31021 2391 31079 2397
rect 31297 2397 31309 2400
rect 31343 2397 31355 2431
rect 31297 2391 31355 2397
rect 33134 2388 33140 2440
rect 33192 2428 33198 2440
rect 33413 2431 33471 2437
rect 33413 2428 33425 2431
rect 33192 2400 33425 2428
rect 33192 2388 33198 2400
rect 33413 2397 33425 2400
rect 33459 2397 33471 2431
rect 33413 2391 33471 2397
rect 34974 2388 34980 2440
rect 35032 2428 35038 2440
rect 40696 2437 40724 2536
rect 41322 2456 41328 2508
rect 41380 2496 41386 2508
rect 41417 2499 41475 2505
rect 41417 2496 41429 2499
rect 41380 2468 41429 2496
rect 41380 2456 41386 2468
rect 41417 2465 41429 2468
rect 41463 2465 41475 2499
rect 41417 2459 41475 2465
rect 49142 2456 49148 2508
rect 49200 2456 49206 2508
rect 35253 2431 35311 2437
rect 35253 2428 35265 2431
rect 35032 2400 35265 2428
rect 35032 2388 35038 2400
rect 35253 2397 35265 2400
rect 35299 2428 35311 2431
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 35299 2400 35541 2428
rect 35299 2397 35311 2400
rect 35253 2391 35311 2397
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 35529 2391 35587 2397
rect 37108 2400 37473 2428
rect 24912 2332 25346 2360
rect 26160 2332 26234 2360
rect 24912 2320 24918 2332
rect 26160 2292 26188 2332
rect 27430 2320 27436 2372
rect 27488 2360 27494 2372
rect 27488 2332 28764 2360
rect 27488 2320 27494 2332
rect 24044 2264 26188 2292
rect 20257 2255 20315 2261
rect 27154 2252 27160 2304
rect 27212 2292 27218 2304
rect 28736 2301 28764 2332
rect 37108 2304 37136 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 40681 2431 40739 2437
rect 40681 2397 40693 2431
rect 40727 2397 40739 2431
rect 40681 2391 40739 2397
rect 44450 2388 44456 2440
rect 44508 2428 44514 2440
rect 45833 2431 45891 2437
rect 45833 2428 45845 2431
rect 44508 2400 45845 2428
rect 44508 2388 44514 2400
rect 45833 2397 45845 2400
rect 45879 2397 45891 2431
rect 45833 2391 45891 2397
rect 47210 2388 47216 2440
rect 47268 2428 47274 2440
rect 47949 2431 48007 2437
rect 47949 2428 47961 2431
rect 47268 2400 47961 2428
rect 47268 2388 47274 2400
rect 47949 2397 47961 2400
rect 47995 2397 48007 2431
rect 47949 2391 48007 2397
rect 47029 2363 47087 2369
rect 47029 2329 47041 2363
rect 47075 2360 47087 2363
rect 48498 2360 48504 2372
rect 47075 2332 48504 2360
rect 47075 2329 47087 2332
rect 47029 2323 47087 2329
rect 48498 2320 48504 2332
rect 48556 2320 48562 2372
rect 28077 2295 28135 2301
rect 28077 2292 28089 2295
rect 27212 2264 28089 2292
rect 27212 2252 27218 2264
rect 28077 2261 28089 2264
rect 28123 2261 28135 2295
rect 28077 2255 28135 2261
rect 28721 2295 28779 2301
rect 28721 2261 28733 2295
rect 28767 2261 28779 2295
rect 28721 2255 28779 2261
rect 30650 2252 30656 2304
rect 30708 2292 30714 2304
rect 30837 2295 30895 2301
rect 30837 2292 30849 2295
rect 30708 2264 30849 2292
rect 30708 2252 30714 2264
rect 30837 2261 30849 2264
rect 30883 2261 30895 2295
rect 30837 2255 30895 2261
rect 37090 2252 37096 2304
rect 37148 2252 37154 2304
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
rect 1302 2048 1308 2100
rect 1360 2088 1366 2100
rect 3234 2088 3240 2100
rect 1360 2060 3240 2088
rect 1360 2048 1366 2060
rect 3234 2048 3240 2060
rect 3292 2048 3298 2100
rect 22462 2048 22468 2100
rect 22520 2088 22526 2100
rect 27154 2088 27160 2100
rect 22520 2060 27160 2088
rect 22520 2048 22526 2060
rect 27154 2048 27160 2060
rect 27212 2048 27218 2100
<< via1 >>
rect 24676 26324 24728 26376
rect 43904 26324 43956 26376
rect 28908 26256 28960 26308
rect 45100 26256 45152 26308
rect 27528 26188 27580 26240
rect 40040 26188 40092 26240
rect 33416 26120 33468 26172
rect 45284 26120 45336 26172
rect 34428 26052 34480 26104
rect 45836 26052 45888 26104
rect 33784 25984 33836 26036
rect 44640 25984 44692 26036
rect 37004 25916 37056 25968
rect 46020 25916 46072 25968
rect 25228 25712 25280 25764
rect 38660 25712 38712 25764
rect 31852 25644 31904 25696
rect 38936 25644 38988 25696
rect 25872 25576 25924 25628
rect 40592 25576 40644 25628
rect 24032 25508 24084 25560
rect 42616 25508 42668 25560
rect 29828 25440 29880 25492
rect 43352 25440 43404 25492
rect 31576 25372 31628 25424
rect 48412 25372 48464 25424
rect 22468 25304 22520 25356
rect 48780 25304 48832 25356
rect 28632 25236 28684 25288
rect 38844 25236 38896 25288
rect 38936 25236 38988 25288
rect 43444 25236 43496 25288
rect 37740 25168 37792 25220
rect 48964 25168 49016 25220
rect 35992 25100 36044 25152
rect 42524 25100 42576 25152
rect 35808 25032 35860 25084
rect 44364 25032 44416 25084
rect 33324 24964 33376 25016
rect 42340 24964 42392 25016
rect 37648 24896 37700 24948
rect 44456 24896 44508 24948
rect 3056 24828 3108 24880
rect 9864 24828 9916 24880
rect 36728 24828 36780 24880
rect 43996 24828 44048 24880
rect 3424 24760 3476 24812
rect 7196 24760 7248 24812
rect 19432 24760 19484 24812
rect 25504 24760 25556 24812
rect 34244 24760 34296 24812
rect 38752 24760 38804 24812
rect 40224 24760 40276 24812
rect 45652 24760 45704 24812
rect 20536 24692 20588 24744
rect 28356 24692 28408 24744
rect 34060 24692 34112 24744
rect 39672 24692 39724 24744
rect 43812 24692 43864 24744
rect 46572 24692 46624 24744
rect 11796 24624 11848 24676
rect 25412 24624 25464 24676
rect 36544 24624 36596 24676
rect 40316 24624 40368 24676
rect 42432 24624 42484 24676
rect 47584 24624 47636 24676
rect 2136 24556 2188 24608
rect 10968 24556 11020 24608
rect 19616 24556 19668 24608
rect 25780 24556 25832 24608
rect 30288 24556 30340 24608
rect 35808 24556 35860 24608
rect 36728 24556 36780 24608
rect 39212 24556 39264 24608
rect 43628 24556 43680 24608
rect 47952 24556 48004 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 2780 24352 2832 24404
rect 6184 24352 6236 24404
rect 3516 24216 3568 24268
rect 6460 24216 6512 24268
rect 13452 24352 13504 24404
rect 21732 24352 21784 24404
rect 22284 24352 22336 24404
rect 2320 24148 2372 24200
rect 4896 24148 4948 24200
rect 5264 24148 5316 24200
rect 8668 24216 8720 24268
rect 7380 24191 7432 24200
rect 7380 24157 7389 24191
rect 7389 24157 7423 24191
rect 7423 24157 7432 24191
rect 7380 24148 7432 24157
rect 9680 24148 9732 24200
rect 10784 24148 10836 24200
rect 11612 24148 11664 24200
rect 14280 24284 14332 24336
rect 14464 24216 14516 24268
rect 18328 24216 18380 24268
rect 19248 24216 19300 24268
rect 19432 24327 19484 24336
rect 19432 24293 19441 24327
rect 19441 24293 19475 24327
rect 19475 24293 19484 24327
rect 19432 24284 19484 24293
rect 22376 24284 22428 24336
rect 5908 24080 5960 24132
rect 12532 24080 12584 24132
rect 17132 24148 17184 24200
rect 17776 24148 17828 24200
rect 19616 24191 19668 24200
rect 19616 24157 19625 24191
rect 19625 24157 19659 24191
rect 19659 24157 19668 24191
rect 19616 24148 19668 24157
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 23388 24216 23440 24268
rect 24860 24395 24912 24404
rect 24860 24361 24869 24395
rect 24869 24361 24903 24395
rect 24903 24361 24912 24395
rect 24860 24352 24912 24361
rect 25136 24352 25188 24404
rect 30196 24352 30248 24404
rect 36268 24352 36320 24404
rect 39396 24352 39448 24404
rect 27620 24284 27672 24336
rect 29644 24284 29696 24336
rect 30288 24284 30340 24336
rect 3976 24055 4028 24064
rect 3976 24021 3985 24055
rect 3985 24021 4019 24055
rect 4019 24021 4028 24055
rect 3976 24012 4028 24021
rect 8852 24012 8904 24064
rect 12440 24012 12492 24064
rect 15016 24012 15068 24064
rect 17408 24012 17460 24064
rect 19156 24012 19208 24064
rect 22560 24148 22612 24200
rect 20260 24080 20312 24132
rect 24032 24191 24084 24200
rect 24032 24157 24041 24191
rect 24041 24157 24075 24191
rect 24075 24157 24084 24191
rect 24032 24148 24084 24157
rect 34060 24259 34112 24268
rect 34060 24225 34069 24259
rect 34069 24225 34103 24259
rect 34103 24225 34112 24259
rect 34060 24216 34112 24225
rect 34244 24259 34296 24268
rect 34244 24225 34253 24259
rect 34253 24225 34287 24259
rect 34287 24225 34296 24259
rect 34244 24216 34296 24225
rect 35256 24284 35308 24336
rect 40040 24352 40092 24404
rect 41144 24352 41196 24404
rect 47952 24395 48004 24404
rect 47952 24361 47961 24395
rect 47961 24361 47995 24395
rect 47995 24361 48004 24395
rect 47952 24352 48004 24361
rect 44732 24284 44784 24336
rect 44824 24284 44876 24336
rect 47216 24284 47268 24336
rect 35348 24259 35400 24268
rect 35348 24225 35357 24259
rect 35357 24225 35391 24259
rect 35391 24225 35400 24259
rect 35348 24216 35400 24225
rect 35808 24216 35860 24268
rect 36544 24259 36596 24268
rect 36544 24225 36553 24259
rect 36553 24225 36587 24259
rect 36587 24225 36596 24259
rect 36544 24216 36596 24225
rect 36728 24259 36780 24268
rect 36728 24225 36737 24259
rect 36737 24225 36771 24259
rect 36771 24225 36780 24259
rect 36728 24216 36780 24225
rect 37924 24259 37976 24268
rect 37924 24225 37933 24259
rect 37933 24225 37967 24259
rect 37967 24225 37976 24259
rect 37924 24216 37976 24225
rect 38384 24216 38436 24268
rect 39488 24216 39540 24268
rect 26608 24148 26660 24200
rect 27344 24148 27396 24200
rect 28356 24191 28408 24200
rect 28356 24157 28365 24191
rect 28365 24157 28399 24191
rect 28399 24157 28408 24191
rect 28356 24148 28408 24157
rect 30288 24148 30340 24200
rect 31484 24148 31536 24200
rect 35072 24148 35124 24200
rect 37832 24191 37884 24200
rect 37832 24157 37841 24191
rect 37841 24157 37875 24191
rect 37875 24157 37884 24191
rect 37832 24148 37884 24157
rect 22744 24080 22796 24132
rect 26884 24080 26936 24132
rect 29368 24080 29420 24132
rect 31116 24080 31168 24132
rect 31300 24080 31352 24132
rect 33876 24080 33928 24132
rect 25964 24012 26016 24064
rect 26516 24055 26568 24064
rect 26516 24021 26525 24055
rect 26525 24021 26559 24055
rect 26559 24021 26568 24055
rect 26516 24012 26568 24021
rect 26792 24012 26844 24064
rect 29644 24012 29696 24064
rect 29920 24055 29972 24064
rect 29920 24021 29929 24055
rect 29929 24021 29963 24055
rect 29963 24021 29972 24055
rect 29920 24012 29972 24021
rect 31668 24012 31720 24064
rect 32128 24055 32180 24064
rect 32128 24021 32137 24055
rect 32137 24021 32171 24055
rect 32171 24021 32180 24055
rect 32128 24012 32180 24021
rect 33600 24055 33652 24064
rect 33600 24021 33609 24055
rect 33609 24021 33643 24055
rect 33643 24021 33652 24055
rect 33600 24012 33652 24021
rect 35164 24012 35216 24064
rect 35532 24080 35584 24132
rect 39120 24148 39172 24200
rect 39396 24148 39448 24200
rect 40224 24148 40276 24200
rect 38292 24080 38344 24132
rect 35348 24012 35400 24064
rect 36084 24055 36136 24064
rect 36084 24021 36093 24055
rect 36093 24021 36127 24055
rect 36127 24021 36136 24055
rect 36084 24012 36136 24021
rect 36176 24012 36228 24064
rect 39948 24012 40000 24064
rect 41144 24259 41196 24268
rect 41144 24225 41153 24259
rect 41153 24225 41187 24259
rect 41187 24225 41196 24259
rect 41144 24216 41196 24225
rect 41420 24259 41472 24268
rect 41420 24225 41429 24259
rect 41429 24225 41463 24259
rect 41463 24225 41472 24259
rect 41420 24216 41472 24225
rect 45468 24259 45520 24268
rect 45468 24225 45477 24259
rect 45477 24225 45511 24259
rect 45511 24225 45520 24259
rect 45468 24216 45520 24225
rect 46296 24216 46348 24268
rect 45192 24191 45244 24200
rect 45192 24157 45201 24191
rect 45201 24157 45235 24191
rect 45235 24157 45244 24191
rect 45192 24148 45244 24157
rect 48228 24216 48280 24268
rect 48780 24259 48832 24268
rect 48780 24225 48789 24259
rect 48789 24225 48823 24259
rect 48823 24225 48832 24259
rect 48780 24216 48832 24225
rect 42156 24080 42208 24132
rect 41788 24012 41840 24064
rect 42432 24012 42484 24064
rect 44180 24012 44232 24064
rect 44732 24055 44784 24064
rect 44732 24021 44741 24055
rect 44741 24021 44775 24055
rect 44775 24021 44784 24055
rect 44732 24012 44784 24021
rect 45008 24012 45060 24064
rect 46756 24080 46808 24132
rect 47124 24080 47176 24132
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 1860 23808 1912 23860
rect 15568 23808 15620 23860
rect 2136 23783 2188 23792
rect 2136 23749 2145 23783
rect 2145 23749 2179 23783
rect 2179 23749 2188 23783
rect 2136 23740 2188 23749
rect 3976 23740 4028 23792
rect 3332 23672 3384 23724
rect 4804 23715 4856 23724
rect 4804 23681 4813 23715
rect 4813 23681 4847 23715
rect 4847 23681 4856 23715
rect 4804 23672 4856 23681
rect 6828 23715 6880 23724
rect 6828 23681 6837 23715
rect 6837 23681 6871 23715
rect 6871 23681 6880 23715
rect 6828 23672 6880 23681
rect 9312 23740 9364 23792
rect 10692 23783 10744 23792
rect 10692 23749 10701 23783
rect 10701 23749 10735 23783
rect 10735 23749 10744 23783
rect 10692 23740 10744 23749
rect 10784 23740 10836 23792
rect 10048 23672 10100 23724
rect 11796 23715 11848 23724
rect 11796 23681 11805 23715
rect 11805 23681 11839 23715
rect 11839 23681 11848 23715
rect 11796 23672 11848 23681
rect 4160 23604 4212 23656
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 9128 23604 9180 23656
rect 14740 23740 14792 23792
rect 12072 23715 12124 23724
rect 12072 23681 12081 23715
rect 12081 23681 12115 23715
rect 12115 23681 12124 23715
rect 12072 23672 12124 23681
rect 15292 23740 15344 23792
rect 17040 23740 17092 23792
rect 19708 23808 19760 23860
rect 20536 23851 20588 23860
rect 20536 23817 20545 23851
rect 20545 23817 20579 23851
rect 20579 23817 20588 23851
rect 20536 23808 20588 23817
rect 22284 23808 22336 23860
rect 22376 23851 22428 23860
rect 22376 23817 22385 23851
rect 22385 23817 22419 23851
rect 22419 23817 22428 23851
rect 22376 23808 22428 23817
rect 22468 23851 22520 23860
rect 22468 23817 22477 23851
rect 22477 23817 22511 23851
rect 22511 23817 22520 23851
rect 22468 23808 22520 23817
rect 23572 23808 23624 23860
rect 24676 23808 24728 23860
rect 18972 23740 19024 23792
rect 20352 23740 20404 23792
rect 20996 23740 21048 23792
rect 21272 23783 21324 23792
rect 21272 23749 21281 23783
rect 21281 23749 21315 23783
rect 21315 23749 21324 23783
rect 21272 23740 21324 23749
rect 21640 23740 21692 23792
rect 26792 23808 26844 23860
rect 29368 23851 29420 23860
rect 29368 23817 29377 23851
rect 29377 23817 29411 23851
rect 29411 23817 29420 23851
rect 29368 23808 29420 23817
rect 26516 23740 26568 23792
rect 28540 23740 28592 23792
rect 14740 23604 14792 23656
rect 9680 23536 9732 23588
rect 16764 23604 16816 23656
rect 17224 23672 17276 23724
rect 18328 23604 18380 23656
rect 18788 23715 18840 23724
rect 18788 23681 18797 23715
rect 18797 23681 18831 23715
rect 18831 23681 18840 23715
rect 18788 23672 18840 23681
rect 24124 23672 24176 23724
rect 27436 23672 27488 23724
rect 28172 23672 28224 23724
rect 30564 23740 30616 23792
rect 30932 23740 30984 23792
rect 32680 23715 32732 23724
rect 32680 23681 32689 23715
rect 32689 23681 32723 23715
rect 32723 23681 32732 23715
rect 32680 23672 32732 23681
rect 19156 23604 19208 23656
rect 15292 23536 15344 23588
rect 22560 23647 22612 23656
rect 22560 23613 22569 23647
rect 22569 23613 22603 23647
rect 22603 23613 22612 23647
rect 22560 23604 22612 23613
rect 23664 23604 23716 23656
rect 24860 23647 24912 23656
rect 24860 23613 24869 23647
rect 24869 23613 24903 23647
rect 24903 23613 24912 23647
rect 24860 23604 24912 23613
rect 29736 23604 29788 23656
rect 3424 23468 3476 23520
rect 6644 23468 6696 23520
rect 17224 23468 17276 23520
rect 20628 23468 20680 23520
rect 23296 23511 23348 23520
rect 23296 23477 23305 23511
rect 23305 23477 23339 23511
rect 23339 23477 23348 23511
rect 23296 23468 23348 23477
rect 29000 23536 29052 23588
rect 32588 23604 32640 23656
rect 35532 23808 35584 23860
rect 35624 23851 35676 23860
rect 35624 23817 35633 23851
rect 35633 23817 35667 23851
rect 35667 23817 35676 23851
rect 35624 23808 35676 23817
rect 35992 23808 36044 23860
rect 38936 23808 38988 23860
rect 33784 23783 33836 23792
rect 33784 23749 33793 23783
rect 33793 23749 33827 23783
rect 33827 23749 33836 23783
rect 33784 23740 33836 23749
rect 34244 23740 34296 23792
rect 35164 23740 35216 23792
rect 38568 23740 38620 23792
rect 35532 23672 35584 23724
rect 26608 23511 26660 23520
rect 26608 23477 26617 23511
rect 26617 23477 26651 23511
rect 26651 23477 26660 23511
rect 26608 23468 26660 23477
rect 27528 23468 27580 23520
rect 27804 23511 27856 23520
rect 27804 23477 27813 23511
rect 27813 23477 27847 23511
rect 27847 23477 27856 23511
rect 27804 23468 27856 23477
rect 30288 23468 30340 23520
rect 33508 23647 33560 23656
rect 33508 23613 33517 23647
rect 33517 23613 33551 23647
rect 33551 23613 33560 23647
rect 33508 23604 33560 23613
rect 35164 23604 35216 23656
rect 36452 23647 36504 23656
rect 36452 23613 36461 23647
rect 36461 23613 36495 23647
rect 36495 23613 36504 23647
rect 36452 23604 36504 23613
rect 35348 23468 35400 23520
rect 35624 23468 35676 23520
rect 36268 23468 36320 23520
rect 36912 23511 36964 23520
rect 36912 23477 36921 23511
rect 36921 23477 36955 23511
rect 36955 23477 36964 23511
rect 36912 23468 36964 23477
rect 39488 23672 39540 23724
rect 39764 23672 39816 23724
rect 39396 23647 39448 23656
rect 39396 23613 39405 23647
rect 39405 23613 39439 23647
rect 39439 23613 39448 23647
rect 39396 23604 39448 23613
rect 39856 23604 39908 23656
rect 44732 23808 44784 23860
rect 45100 23740 45152 23792
rect 42800 23672 42852 23724
rect 44272 23672 44324 23724
rect 45560 23672 45612 23724
rect 46204 23672 46256 23724
rect 46940 23740 46992 23792
rect 47492 23740 47544 23792
rect 41144 23647 41196 23656
rect 41144 23613 41153 23647
rect 41153 23613 41187 23647
rect 41187 23613 41196 23647
rect 41144 23604 41196 23613
rect 42892 23647 42944 23656
rect 42892 23613 42901 23647
rect 42901 23613 42935 23647
rect 42935 23613 42944 23647
rect 42892 23604 42944 23613
rect 43904 23647 43956 23656
rect 43904 23613 43913 23647
rect 43913 23613 43947 23647
rect 43947 23613 43956 23647
rect 43904 23604 43956 23613
rect 45100 23604 45152 23656
rect 43812 23536 43864 23588
rect 47952 23672 48004 23724
rect 45560 23536 45612 23588
rect 40040 23468 40092 23520
rect 40132 23468 40184 23520
rect 41880 23468 41932 23520
rect 41972 23468 42024 23520
rect 47584 23468 47636 23520
rect 49056 23511 49108 23520
rect 49056 23477 49065 23511
rect 49065 23477 49099 23511
rect 49099 23477 49108 23511
rect 49056 23468 49108 23477
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 6828 23264 6880 23316
rect 13268 23264 13320 23316
rect 17132 23264 17184 23316
rect 17592 23264 17644 23316
rect 19616 23264 19668 23316
rect 19708 23307 19760 23316
rect 19708 23273 19717 23307
rect 19717 23273 19751 23307
rect 19751 23273 19760 23307
rect 19708 23264 19760 23273
rect 8576 23196 8628 23248
rect 5264 23128 5316 23180
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 9404 23171 9456 23180
rect 9404 23137 9413 23171
rect 9413 23137 9447 23171
rect 9447 23137 9456 23171
rect 9404 23128 9456 23137
rect 11244 23171 11296 23180
rect 11244 23137 11253 23171
rect 11253 23137 11287 23171
rect 11287 23137 11296 23171
rect 11244 23128 11296 23137
rect 13360 23171 13412 23180
rect 13360 23137 13369 23171
rect 13369 23137 13403 23171
rect 13403 23137 13412 23171
rect 13360 23128 13412 23137
rect 14280 23171 14332 23180
rect 14280 23137 14289 23171
rect 14289 23137 14323 23171
rect 14323 23137 14332 23171
rect 14280 23128 14332 23137
rect 14556 23128 14608 23180
rect 16396 23171 16448 23180
rect 16396 23137 16405 23171
rect 16405 23137 16439 23171
rect 16439 23137 16448 23171
rect 16396 23128 16448 23137
rect 18604 23196 18656 23248
rect 22560 23264 22612 23316
rect 18788 23128 18840 23180
rect 21180 23128 21232 23180
rect 29828 23264 29880 23316
rect 33784 23264 33836 23316
rect 35348 23264 35400 23316
rect 35808 23264 35860 23316
rect 23388 23196 23440 23248
rect 23112 23171 23164 23180
rect 23112 23137 23121 23171
rect 23121 23137 23155 23171
rect 23155 23137 23164 23171
rect 23112 23128 23164 23137
rect 2780 23035 2832 23044
rect 2780 23001 2789 23035
rect 2789 23001 2823 23035
rect 2823 23001 2832 23035
rect 2780 22992 2832 23001
rect 3976 23103 4028 23112
rect 3976 23069 3985 23103
rect 3985 23069 4019 23103
rect 4019 23069 4028 23103
rect 3976 23060 4028 23069
rect 4436 23060 4488 23112
rect 7104 23060 7156 23112
rect 9220 23060 9272 23112
rect 4344 22992 4396 23044
rect 12440 23103 12492 23112
rect 12440 23069 12449 23103
rect 12449 23069 12483 23103
rect 12483 23069 12492 23103
rect 12440 23060 12492 23069
rect 16672 23060 16724 23112
rect 17132 23103 17184 23112
rect 17132 23069 17141 23103
rect 17141 23069 17175 23103
rect 17175 23069 17184 23103
rect 17132 23060 17184 23069
rect 19892 23103 19944 23112
rect 19892 23069 19901 23103
rect 19901 23069 19935 23103
rect 19935 23069 19944 23103
rect 19892 23060 19944 23069
rect 22008 23060 22060 23112
rect 23664 23128 23716 23180
rect 25964 23171 26016 23180
rect 25964 23137 25973 23171
rect 25973 23137 26007 23171
rect 26007 23137 26016 23171
rect 25964 23128 26016 23137
rect 23848 23103 23900 23112
rect 23848 23069 23857 23103
rect 23857 23069 23891 23103
rect 23891 23069 23900 23103
rect 23848 23060 23900 23069
rect 25596 23060 25648 23112
rect 26976 23060 27028 23112
rect 30012 23196 30064 23248
rect 30932 23239 30984 23248
rect 30932 23205 30941 23239
rect 30941 23205 30975 23239
rect 30975 23205 30984 23239
rect 30932 23196 30984 23205
rect 38752 23264 38804 23316
rect 39764 23264 39816 23316
rect 40040 23307 40092 23316
rect 40040 23273 40049 23307
rect 40049 23273 40083 23307
rect 40083 23273 40092 23307
rect 40040 23264 40092 23273
rect 41052 23307 41104 23316
rect 41052 23273 41061 23307
rect 41061 23273 41095 23307
rect 41095 23273 41104 23307
rect 41052 23264 41104 23273
rect 43260 23264 43312 23316
rect 43536 23264 43588 23316
rect 43904 23307 43956 23316
rect 39396 23196 39448 23248
rect 39488 23239 39540 23248
rect 39488 23205 39497 23239
rect 39497 23205 39531 23239
rect 39531 23205 39540 23239
rect 39488 23196 39540 23205
rect 40132 23196 40184 23248
rect 40408 23196 40460 23248
rect 42892 23196 42944 23248
rect 43628 23196 43680 23248
rect 27620 23128 27672 23180
rect 28356 23171 28408 23180
rect 28356 23137 28365 23171
rect 28365 23137 28399 23171
rect 28399 23137 28408 23171
rect 28356 23128 28408 23137
rect 14096 22992 14148 23044
rect 14648 23035 14700 23044
rect 14648 23001 14657 23035
rect 14657 23001 14691 23035
rect 14691 23001 14700 23035
rect 14648 22992 14700 23001
rect 17500 22992 17552 23044
rect 18420 22992 18472 23044
rect 14280 22924 14332 22976
rect 17592 22924 17644 22976
rect 17776 22924 17828 22976
rect 20628 23035 20680 23044
rect 20628 23001 20637 23035
rect 20637 23001 20671 23035
rect 20671 23001 20680 23035
rect 20628 22992 20680 23001
rect 20720 22992 20772 23044
rect 21088 22992 21140 23044
rect 24032 22992 24084 23044
rect 24216 22992 24268 23044
rect 22100 22967 22152 22976
rect 22100 22933 22109 22967
rect 22109 22933 22143 22967
rect 22143 22933 22152 22967
rect 22100 22924 22152 22933
rect 22468 22924 22520 22976
rect 23756 22924 23808 22976
rect 25320 22924 25372 22976
rect 28172 22992 28224 23044
rect 30196 23171 30248 23180
rect 30196 23137 30205 23171
rect 30205 23137 30239 23171
rect 30239 23137 30248 23171
rect 30196 23128 30248 23137
rect 30288 23171 30340 23180
rect 30288 23137 30297 23171
rect 30297 23137 30331 23171
rect 30331 23137 30340 23171
rect 30288 23128 30340 23137
rect 31668 23171 31720 23180
rect 31668 23137 31677 23171
rect 31677 23137 31711 23171
rect 31711 23137 31720 23171
rect 31668 23128 31720 23137
rect 32864 23128 32916 23180
rect 34888 23128 34940 23180
rect 37464 23128 37516 23180
rect 39028 23128 39080 23180
rect 39304 23128 39356 23180
rect 39764 23128 39816 23180
rect 27436 22967 27488 22976
rect 27436 22933 27445 22967
rect 27445 22933 27479 22967
rect 27479 22933 27488 22967
rect 27436 22924 27488 22933
rect 31024 23060 31076 23112
rect 31208 23060 31260 23112
rect 33968 23060 34020 23112
rect 41512 23171 41564 23180
rect 41512 23137 41521 23171
rect 41521 23137 41555 23171
rect 41555 23137 41564 23171
rect 41512 23128 41564 23137
rect 40776 23060 40828 23112
rect 43076 23060 43128 23112
rect 43904 23273 43913 23307
rect 43913 23273 43947 23307
rect 43947 23273 43956 23307
rect 43904 23264 43956 23273
rect 44180 23264 44232 23316
rect 44824 23307 44876 23316
rect 44824 23273 44833 23307
rect 44833 23273 44867 23307
rect 44867 23273 44876 23307
rect 44824 23264 44876 23273
rect 45100 23264 45152 23316
rect 45284 23264 45336 23316
rect 47584 23307 47636 23316
rect 47584 23273 47593 23307
rect 47593 23273 47627 23307
rect 47627 23273 47636 23307
rect 47584 23264 47636 23273
rect 47768 23264 47820 23316
rect 48504 23307 48556 23316
rect 48504 23273 48513 23307
rect 48513 23273 48547 23307
rect 48547 23273 48556 23307
rect 48504 23264 48556 23273
rect 48964 23264 49016 23316
rect 44088 23196 44140 23248
rect 43904 23128 43956 23180
rect 45560 23128 45612 23180
rect 44088 23060 44140 23112
rect 44548 23060 44600 23112
rect 28724 22992 28776 23044
rect 30840 22992 30892 23044
rect 30932 22992 30984 23044
rect 32128 22992 32180 23044
rect 35256 23035 35308 23044
rect 35256 23001 35265 23035
rect 35265 23001 35299 23035
rect 35299 23001 35308 23035
rect 35256 22992 35308 23001
rect 35992 22992 36044 23044
rect 29092 22924 29144 22976
rect 29276 22924 29328 22976
rect 29368 22967 29420 22976
rect 29368 22933 29377 22967
rect 29377 22933 29411 22967
rect 29411 22933 29420 22967
rect 29368 22924 29420 22933
rect 30104 22967 30156 22976
rect 30104 22933 30113 22967
rect 30113 22933 30147 22967
rect 30147 22933 30156 22967
rect 30104 22924 30156 22933
rect 30656 22924 30708 22976
rect 31484 22924 31536 22976
rect 35900 22924 35952 22976
rect 36728 22967 36780 22976
rect 36728 22933 36737 22967
rect 36737 22933 36771 22967
rect 36771 22933 36780 22967
rect 36728 22924 36780 22933
rect 39488 22992 39540 23044
rect 40500 23035 40552 23044
rect 40500 23001 40509 23035
rect 40509 23001 40543 23035
rect 40543 23001 40552 23035
rect 40500 22992 40552 23001
rect 38292 22924 38344 22976
rect 39304 22967 39356 22976
rect 39304 22933 39313 22967
rect 39313 22933 39347 22967
rect 39347 22933 39356 22967
rect 39304 22924 39356 22933
rect 39764 22924 39816 22976
rect 41696 22992 41748 23044
rect 43628 22992 43680 23044
rect 44640 22992 44692 23044
rect 44824 22992 44876 23044
rect 48320 23103 48372 23112
rect 48320 23069 48329 23103
rect 48329 23069 48363 23103
rect 48363 23069 48372 23103
rect 48320 23060 48372 23069
rect 47308 22992 47360 23044
rect 43720 22924 43772 22976
rect 43996 22924 44048 22976
rect 46480 22924 46532 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 3148 22720 3200 22772
rect 6736 22720 6788 22772
rect 6828 22720 6880 22772
rect 2872 22652 2924 22704
rect 4252 22652 4304 22704
rect 14464 22652 14516 22704
rect 1860 22584 1912 22636
rect 3884 22584 3936 22636
rect 4068 22584 4120 22636
rect 5816 22584 5868 22636
rect 6920 22584 6972 22636
rect 9772 22627 9824 22636
rect 9772 22593 9781 22627
rect 9781 22593 9815 22627
rect 9815 22593 9824 22627
rect 9772 22584 9824 22593
rect 16580 22720 16632 22772
rect 16672 22720 16724 22772
rect 15844 22695 15896 22704
rect 15844 22661 15853 22695
rect 15853 22661 15887 22695
rect 15887 22661 15896 22695
rect 15844 22652 15896 22661
rect 2872 22516 2924 22568
rect 4160 22559 4212 22568
rect 4160 22525 4169 22559
rect 4169 22525 4203 22559
rect 4203 22525 4212 22559
rect 4160 22516 4212 22525
rect 5080 22559 5132 22568
rect 5080 22525 5089 22559
rect 5089 22525 5123 22559
rect 5123 22525 5132 22559
rect 5080 22516 5132 22525
rect 7656 22516 7708 22568
rect 9680 22516 9732 22568
rect 9956 22516 10008 22568
rect 3424 22448 3476 22500
rect 5632 22448 5684 22500
rect 11612 22516 11664 22568
rect 11796 22516 11848 22568
rect 11980 22559 12032 22568
rect 11980 22525 11989 22559
rect 11989 22525 12023 22559
rect 12023 22525 12032 22559
rect 11980 22516 12032 22525
rect 13820 22559 13872 22568
rect 13820 22525 13829 22559
rect 13829 22525 13863 22559
rect 13863 22525 13872 22559
rect 13820 22516 13872 22525
rect 10416 22448 10468 22500
rect 18420 22652 18472 22704
rect 18604 22763 18656 22772
rect 18604 22729 18613 22763
rect 18613 22729 18647 22763
rect 18647 22729 18656 22763
rect 18604 22720 18656 22729
rect 19064 22763 19116 22772
rect 19064 22729 19073 22763
rect 19073 22729 19107 22763
rect 19107 22729 19116 22763
rect 19064 22720 19116 22729
rect 19524 22652 19576 22704
rect 20352 22652 20404 22704
rect 21088 22652 21140 22704
rect 21824 22652 21876 22704
rect 25136 22720 25188 22772
rect 23296 22652 23348 22704
rect 23572 22652 23624 22704
rect 24400 22652 24452 22704
rect 26424 22720 26476 22772
rect 26884 22720 26936 22772
rect 27436 22720 27488 22772
rect 16856 22627 16908 22636
rect 16856 22593 16865 22627
rect 16865 22593 16899 22627
rect 16899 22593 16908 22627
rect 16856 22584 16908 22593
rect 21180 22584 21232 22636
rect 22008 22627 22060 22636
rect 22008 22593 22017 22627
rect 22017 22593 22051 22627
rect 22051 22593 22060 22627
rect 22008 22584 22060 22593
rect 26516 22652 26568 22704
rect 26976 22652 27028 22704
rect 27712 22652 27764 22704
rect 28632 22652 28684 22704
rect 30012 22652 30064 22704
rect 5724 22380 5776 22432
rect 9404 22380 9456 22432
rect 13268 22380 13320 22432
rect 13360 22380 13412 22432
rect 18788 22448 18840 22500
rect 19432 22516 19484 22568
rect 22652 22516 22704 22568
rect 24124 22516 24176 22568
rect 24308 22516 24360 22568
rect 16856 22380 16908 22432
rect 17132 22380 17184 22432
rect 17868 22380 17920 22432
rect 22100 22380 22152 22432
rect 22744 22380 22796 22432
rect 24860 22627 24912 22636
rect 24860 22593 24869 22627
rect 24869 22593 24903 22627
rect 24903 22593 24912 22627
rect 24860 22584 24912 22593
rect 27436 22584 27488 22636
rect 24584 22516 24636 22568
rect 24584 22423 24636 22432
rect 24584 22389 24593 22423
rect 24593 22389 24627 22423
rect 24627 22389 24636 22423
rect 24584 22380 24636 22389
rect 27804 22516 27856 22568
rect 26148 22448 26200 22500
rect 26516 22448 26568 22500
rect 27252 22448 27304 22500
rect 30380 22516 30432 22568
rect 30840 22720 30892 22772
rect 31760 22720 31812 22772
rect 33416 22763 33468 22772
rect 33416 22729 33425 22763
rect 33425 22729 33459 22763
rect 33459 22729 33468 22763
rect 33416 22720 33468 22729
rect 33508 22720 33560 22772
rect 33600 22652 33652 22704
rect 32496 22584 32548 22636
rect 34888 22720 34940 22772
rect 35624 22720 35676 22772
rect 33876 22652 33928 22704
rect 34244 22652 34296 22704
rect 41696 22720 41748 22772
rect 44272 22720 44324 22772
rect 46940 22763 46992 22772
rect 46940 22729 46949 22763
rect 46949 22729 46983 22763
rect 46983 22729 46992 22763
rect 46940 22720 46992 22729
rect 47308 22720 47360 22772
rect 48504 22763 48556 22772
rect 48504 22729 48513 22763
rect 48513 22729 48547 22763
rect 48547 22729 48556 22763
rect 48504 22720 48556 22729
rect 49148 22720 49200 22772
rect 39488 22652 39540 22704
rect 39580 22652 39632 22704
rect 31668 22516 31720 22568
rect 26240 22380 26292 22432
rect 26608 22423 26660 22432
rect 26608 22389 26617 22423
rect 26617 22389 26651 22423
rect 26651 22389 26660 22423
rect 26608 22380 26660 22389
rect 31208 22448 31260 22500
rect 32772 22559 32824 22568
rect 32772 22525 32781 22559
rect 32781 22525 32815 22559
rect 32815 22525 32824 22559
rect 32772 22516 32824 22525
rect 29736 22380 29788 22432
rect 29920 22380 29972 22432
rect 30288 22423 30340 22432
rect 30288 22389 30297 22423
rect 30297 22389 30331 22423
rect 30331 22389 30340 22423
rect 30288 22380 30340 22389
rect 37096 22584 37148 22636
rect 37464 22627 37516 22636
rect 37464 22593 37473 22627
rect 37473 22593 37507 22627
rect 37507 22593 37516 22627
rect 37464 22584 37516 22593
rect 40040 22627 40092 22636
rect 40040 22593 40049 22627
rect 40049 22593 40083 22627
rect 40083 22593 40092 22627
rect 40040 22584 40092 22593
rect 34428 22516 34480 22568
rect 34612 22516 34664 22568
rect 33692 22448 33744 22500
rect 35532 22448 35584 22500
rect 40132 22559 40184 22568
rect 40132 22525 40141 22559
rect 40141 22525 40175 22559
rect 40175 22525 40184 22559
rect 40132 22516 40184 22525
rect 40224 22559 40276 22568
rect 40224 22525 40233 22559
rect 40233 22525 40267 22559
rect 40267 22525 40276 22559
rect 40224 22516 40276 22525
rect 40500 22652 40552 22704
rect 41328 22652 41380 22704
rect 41880 22695 41932 22704
rect 41880 22661 41889 22695
rect 41889 22661 41923 22695
rect 41923 22661 41932 22695
rect 41880 22652 41932 22661
rect 42156 22652 42208 22704
rect 43076 22652 43128 22704
rect 46480 22652 46532 22704
rect 41052 22584 41104 22636
rect 43352 22584 43404 22636
rect 43536 22627 43588 22636
rect 43536 22593 43545 22627
rect 43545 22593 43579 22627
rect 43579 22593 43588 22627
rect 43536 22584 43588 22593
rect 44364 22584 44416 22636
rect 45836 22627 45888 22636
rect 45836 22593 45845 22627
rect 45845 22593 45879 22627
rect 45879 22593 45888 22627
rect 45836 22584 45888 22593
rect 40408 22448 40460 22500
rect 34704 22380 34756 22432
rect 35900 22380 35952 22432
rect 36728 22380 36780 22432
rect 38752 22380 38804 22432
rect 39672 22423 39724 22432
rect 39672 22389 39681 22423
rect 39681 22389 39715 22423
rect 39715 22389 39724 22423
rect 39672 22380 39724 22389
rect 42616 22491 42668 22500
rect 42616 22457 42625 22491
rect 42625 22457 42659 22491
rect 42659 22457 42668 22491
rect 42616 22448 42668 22457
rect 44088 22516 44140 22568
rect 44732 22516 44784 22568
rect 45008 22516 45060 22568
rect 46112 22559 46164 22568
rect 46112 22525 46121 22559
rect 46121 22525 46155 22559
rect 46155 22525 46164 22559
rect 46112 22516 46164 22525
rect 46848 22584 46900 22636
rect 47768 22584 47820 22636
rect 49332 22584 49384 22636
rect 46848 22448 46900 22500
rect 49148 22448 49200 22500
rect 48320 22380 48372 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 1584 22176 1636 22228
rect 4620 22176 4672 22228
rect 13912 22176 13964 22228
rect 16856 22176 16908 22228
rect 18420 22176 18472 22228
rect 21640 22176 21692 22228
rect 21824 22176 21876 22228
rect 2228 22108 2280 22160
rect 4528 22108 4580 22160
rect 1308 22040 1360 22092
rect 3792 22040 3844 22092
rect 6736 22083 6788 22092
rect 6736 22049 6745 22083
rect 6745 22049 6779 22083
rect 6779 22049 6788 22083
rect 6736 22040 6788 22049
rect 8576 22083 8628 22092
rect 8576 22049 8585 22083
rect 8585 22049 8619 22083
rect 8619 22049 8628 22083
rect 8576 22040 8628 22049
rect 9864 22083 9916 22092
rect 9864 22049 9873 22083
rect 9873 22049 9907 22083
rect 9907 22049 9916 22083
rect 9864 22040 9916 22049
rect 10048 22040 10100 22092
rect 1768 22015 1820 22024
rect 1768 21981 1777 22015
rect 1777 21981 1811 22015
rect 1811 21981 1820 22015
rect 1768 21972 1820 21981
rect 7656 21972 7708 22024
rect 7932 22015 7984 22024
rect 7932 21981 7941 22015
rect 7941 21981 7975 22015
rect 7975 21981 7984 22015
rect 7932 21972 7984 21981
rect 9128 22015 9180 22024
rect 9128 21981 9137 22015
rect 9137 21981 9171 22015
rect 9171 21981 9180 22015
rect 9128 21972 9180 21981
rect 11796 22108 11848 22160
rect 11888 22108 11940 22160
rect 11704 22083 11756 22092
rect 11704 22049 11713 22083
rect 11713 22049 11747 22083
rect 11747 22049 11756 22083
rect 11704 22040 11756 22049
rect 13636 22108 13688 22160
rect 14280 22040 14332 22092
rect 14740 22083 14792 22092
rect 14740 22049 14749 22083
rect 14749 22049 14783 22083
rect 14783 22049 14792 22083
rect 14740 22040 14792 22049
rect 17132 22108 17184 22160
rect 11796 21972 11848 22024
rect 15200 22015 15252 22024
rect 15200 21981 15209 22015
rect 15209 21981 15243 22015
rect 15243 21981 15252 22015
rect 15200 21972 15252 21981
rect 17500 22015 17552 22024
rect 17500 21981 17509 22015
rect 17509 21981 17543 22015
rect 17543 21981 17552 22015
rect 17500 21972 17552 21981
rect 11060 21947 11112 21956
rect 11060 21913 11069 21947
rect 11069 21913 11103 21947
rect 11103 21913 11112 21947
rect 11060 21904 11112 21913
rect 14372 21904 14424 21956
rect 14832 21904 14884 21956
rect 16856 21904 16908 21956
rect 9404 21836 9456 21888
rect 14188 21879 14240 21888
rect 14188 21845 14197 21879
rect 14197 21845 14231 21879
rect 14231 21845 14240 21879
rect 14188 21836 14240 21845
rect 15292 21836 15344 21888
rect 17040 21836 17092 21888
rect 17776 21836 17828 21888
rect 20352 22040 20404 22092
rect 20444 22040 20496 22092
rect 20628 22040 20680 22092
rect 22468 22040 22520 22092
rect 18052 21972 18104 22024
rect 19340 21972 19392 22024
rect 19432 21972 19484 22024
rect 20076 21972 20128 22024
rect 21180 22015 21232 22024
rect 21180 21981 21189 22015
rect 21189 21981 21223 22015
rect 21223 21981 21232 22015
rect 21180 21972 21232 21981
rect 23756 22176 23808 22228
rect 25136 22176 25188 22228
rect 27252 22176 27304 22228
rect 27344 22176 27396 22228
rect 22652 22108 22704 22160
rect 22744 22040 22796 22092
rect 25780 22108 25832 22160
rect 23204 21972 23256 22024
rect 23296 21972 23348 22024
rect 24216 22040 24268 22092
rect 25412 22040 25464 22092
rect 26148 22040 26200 22092
rect 26608 22108 26660 22160
rect 26700 22108 26752 22160
rect 27620 22108 27672 22160
rect 29368 22176 29420 22228
rect 30288 22176 30340 22228
rect 30380 22219 30432 22228
rect 30380 22185 30389 22219
rect 30389 22185 30423 22219
rect 30423 22185 30432 22219
rect 30380 22176 30432 22185
rect 29920 22108 29972 22160
rect 25044 22015 25096 22024
rect 25044 21981 25053 22015
rect 25053 21981 25087 22015
rect 25087 21981 25096 22015
rect 25044 21972 25096 21981
rect 26884 21972 26936 22024
rect 18144 21904 18196 21956
rect 20168 21904 20220 21956
rect 20720 21904 20772 21956
rect 19432 21836 19484 21888
rect 19984 21879 20036 21888
rect 19984 21845 19993 21879
rect 19993 21845 20027 21879
rect 20027 21845 20036 21879
rect 19984 21836 20036 21845
rect 23020 21836 23072 21888
rect 24308 21836 24360 21888
rect 25412 21836 25464 21888
rect 28908 22040 28960 22092
rect 28816 21972 28868 22024
rect 29644 21972 29696 22024
rect 31668 22176 31720 22228
rect 32496 22176 32548 22228
rect 34244 22176 34296 22228
rect 32588 22151 32640 22160
rect 32588 22117 32597 22151
rect 32597 22117 32631 22151
rect 32631 22117 32640 22151
rect 32588 22108 32640 22117
rect 31208 22040 31260 22092
rect 32312 22040 32364 22092
rect 33324 22040 33376 22092
rect 29368 21904 29420 21956
rect 31208 21904 31260 21956
rect 31392 21904 31444 21956
rect 32128 21904 32180 21956
rect 33508 22083 33560 22092
rect 33508 22049 33517 22083
rect 33517 22049 33551 22083
rect 33551 22049 33560 22083
rect 33508 22040 33560 22049
rect 33784 22108 33836 22160
rect 34336 22108 34388 22160
rect 33876 22040 33928 22092
rect 38568 22176 38620 22228
rect 38844 22176 38896 22228
rect 39764 22176 39816 22228
rect 40040 22176 40092 22228
rect 35900 21972 35952 22024
rect 38752 22108 38804 22160
rect 38292 22040 38344 22092
rect 38568 22040 38620 22092
rect 40776 22108 40828 22160
rect 41052 22108 41104 22160
rect 43628 22176 43680 22228
rect 45560 22176 45612 22228
rect 45652 22176 45704 22228
rect 40868 22040 40920 22092
rect 41420 22040 41472 22092
rect 42340 22040 42392 22092
rect 37188 21972 37240 22024
rect 39396 21972 39448 22024
rect 42892 22151 42944 22160
rect 42892 22117 42901 22151
rect 42901 22117 42935 22151
rect 42935 22117 42944 22151
rect 42892 22108 42944 22117
rect 43536 22083 43588 22092
rect 43536 22049 43545 22083
rect 43545 22049 43579 22083
rect 43579 22049 43588 22083
rect 43536 22040 43588 22049
rect 43352 21972 43404 22024
rect 43720 21972 43772 22024
rect 26332 21879 26384 21888
rect 26332 21845 26341 21879
rect 26341 21845 26375 21879
rect 26375 21845 26384 21879
rect 26332 21836 26384 21845
rect 26700 21836 26752 21888
rect 27344 21836 27396 21888
rect 28632 21836 28684 21888
rect 31760 21836 31812 21888
rect 32680 21836 32732 21888
rect 33140 21836 33192 21888
rect 34520 21879 34572 21888
rect 34520 21845 34529 21879
rect 34529 21845 34563 21879
rect 34563 21845 34572 21879
rect 34520 21836 34572 21845
rect 35164 21836 35216 21888
rect 35256 21879 35308 21888
rect 35256 21845 35265 21879
rect 35265 21845 35299 21879
rect 35299 21845 35308 21879
rect 35256 21836 35308 21845
rect 36176 21836 36228 21888
rect 36452 21879 36504 21888
rect 36452 21845 36461 21879
rect 36461 21845 36495 21879
rect 36495 21845 36504 21879
rect 36452 21836 36504 21845
rect 36544 21879 36596 21888
rect 36544 21845 36553 21879
rect 36553 21845 36587 21879
rect 36587 21845 36596 21879
rect 36544 21836 36596 21845
rect 37464 21904 37516 21956
rect 37556 21904 37608 21956
rect 39580 21947 39632 21956
rect 39580 21913 39589 21947
rect 39589 21913 39623 21947
rect 39623 21913 39632 21947
rect 39580 21904 39632 21913
rect 40592 21904 40644 21956
rect 44548 21904 44600 21956
rect 46020 22108 46072 22160
rect 47308 22176 47360 22228
rect 49240 22176 49292 22228
rect 48596 22040 48648 22092
rect 45284 21972 45336 22024
rect 45652 21972 45704 22024
rect 45744 21972 45796 22024
rect 47308 22015 47360 22024
rect 47308 21981 47317 22015
rect 47317 21981 47351 22015
rect 47351 21981 47360 22015
rect 47308 21972 47360 21981
rect 49056 21972 49108 22024
rect 37280 21836 37332 21888
rect 40040 21879 40092 21888
rect 40040 21845 40049 21879
rect 40049 21845 40083 21879
rect 40083 21845 40092 21879
rect 40040 21836 40092 21845
rect 40500 21879 40552 21888
rect 40500 21845 40509 21879
rect 40509 21845 40543 21879
rect 40543 21845 40552 21879
rect 40500 21836 40552 21845
rect 41512 21836 41564 21888
rect 41696 21879 41748 21888
rect 41696 21845 41705 21879
rect 41705 21845 41739 21879
rect 41739 21845 41748 21879
rect 41696 21836 41748 21845
rect 43444 21836 43496 21888
rect 45468 21904 45520 21956
rect 49148 21947 49200 21956
rect 49148 21913 49157 21947
rect 49157 21913 49191 21947
rect 49191 21913 49200 21947
rect 49148 21904 49200 21913
rect 49424 21904 49476 21956
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 9220 21632 9272 21684
rect 11796 21675 11848 21684
rect 11796 21641 11805 21675
rect 11805 21641 11839 21675
rect 11839 21641 11848 21675
rect 11796 21632 11848 21641
rect 13360 21632 13412 21684
rect 14740 21675 14792 21684
rect 14740 21641 14749 21675
rect 14749 21641 14783 21675
rect 14783 21641 14792 21675
rect 14740 21632 14792 21641
rect 15108 21675 15160 21684
rect 15108 21641 15117 21675
rect 15117 21641 15151 21675
rect 15151 21641 15160 21675
rect 15108 21632 15160 21641
rect 15568 21632 15620 21684
rect 20628 21632 20680 21684
rect 22284 21632 22336 21684
rect 25136 21675 25188 21684
rect 25136 21641 25145 21675
rect 25145 21641 25179 21675
rect 25179 21641 25188 21675
rect 25136 21632 25188 21641
rect 27160 21675 27212 21684
rect 27160 21641 27169 21675
rect 27169 21641 27203 21675
rect 27203 21641 27212 21675
rect 27160 21632 27212 21641
rect 28540 21632 28592 21684
rect 28724 21675 28776 21684
rect 28724 21641 28733 21675
rect 28733 21641 28767 21675
rect 28767 21641 28776 21675
rect 28724 21632 28776 21641
rect 31760 21632 31812 21684
rect 32128 21632 32180 21684
rect 32404 21632 32456 21684
rect 35808 21632 35860 21684
rect 40040 21632 40092 21684
rect 40132 21632 40184 21684
rect 1768 21564 1820 21616
rect 3976 21564 4028 21616
rect 4252 21564 4304 21616
rect 5356 21564 5408 21616
rect 3424 21496 3476 21548
rect 5080 21496 5132 21548
rect 5172 21496 5224 21548
rect 7748 21564 7800 21616
rect 10324 21564 10376 21616
rect 7288 21496 7340 21548
rect 17040 21564 17092 21616
rect 17132 21564 17184 21616
rect 1400 21428 1452 21480
rect 4344 21428 4396 21480
rect 6644 21428 6696 21480
rect 7840 21428 7892 21480
rect 5448 21403 5500 21412
rect 5448 21369 5457 21403
rect 5457 21369 5491 21403
rect 5491 21369 5500 21403
rect 5448 21360 5500 21369
rect 3608 21292 3660 21344
rect 11980 21539 12032 21548
rect 11980 21505 11989 21539
rect 11989 21505 12023 21539
rect 12023 21505 12032 21539
rect 11980 21496 12032 21505
rect 9772 21428 9824 21480
rect 10324 21428 10376 21480
rect 11152 21471 11204 21480
rect 11152 21437 11161 21471
rect 11161 21437 11195 21471
rect 11195 21437 11204 21471
rect 11152 21428 11204 21437
rect 13636 21539 13688 21548
rect 13636 21505 13645 21539
rect 13645 21505 13679 21539
rect 13679 21505 13688 21539
rect 13636 21496 13688 21505
rect 14924 21496 14976 21548
rect 16120 21539 16172 21548
rect 16120 21505 16129 21539
rect 16129 21505 16163 21539
rect 16163 21505 16172 21539
rect 16120 21496 16172 21505
rect 17224 21539 17276 21548
rect 17224 21505 17233 21539
rect 17233 21505 17267 21539
rect 17267 21505 17276 21539
rect 17224 21496 17276 21505
rect 15016 21428 15068 21480
rect 15292 21471 15344 21480
rect 15292 21437 15301 21471
rect 15301 21437 15335 21471
rect 15335 21437 15344 21471
rect 15292 21428 15344 21437
rect 20076 21564 20128 21616
rect 20444 21564 20496 21616
rect 23020 21564 23072 21616
rect 23388 21564 23440 21616
rect 28172 21564 28224 21616
rect 28632 21564 28684 21616
rect 29276 21564 29328 21616
rect 30196 21564 30248 21616
rect 34244 21564 34296 21616
rect 34980 21564 35032 21616
rect 35992 21564 36044 21616
rect 36912 21607 36964 21616
rect 36912 21573 36921 21607
rect 36921 21573 36955 21607
rect 36955 21573 36964 21607
rect 36912 21564 36964 21573
rect 37556 21564 37608 21616
rect 38568 21564 38620 21616
rect 38752 21564 38804 21616
rect 21272 21496 21324 21548
rect 17960 21428 18012 21480
rect 9588 21292 9640 21344
rect 20168 21428 20220 21480
rect 20628 21428 20680 21480
rect 21548 21496 21600 21548
rect 21916 21539 21968 21548
rect 21916 21505 21925 21539
rect 21925 21505 21959 21539
rect 21959 21505 21968 21539
rect 21916 21496 21968 21505
rect 22008 21496 22060 21548
rect 23296 21428 23348 21480
rect 25228 21471 25280 21480
rect 25228 21437 25237 21471
rect 25237 21437 25271 21471
rect 25271 21437 25280 21471
rect 25228 21428 25280 21437
rect 25964 21539 26016 21548
rect 25964 21505 25973 21539
rect 25973 21505 26007 21539
rect 26007 21505 26016 21539
rect 25964 21496 26016 21505
rect 26608 21539 26660 21548
rect 26608 21505 26617 21539
rect 26617 21505 26651 21539
rect 26651 21505 26660 21539
rect 26608 21496 26660 21505
rect 29092 21496 29144 21548
rect 29552 21496 29604 21548
rect 28172 21428 28224 21480
rect 28632 21428 28684 21480
rect 28816 21471 28868 21480
rect 28816 21437 28825 21471
rect 28825 21437 28859 21471
rect 28859 21437 28868 21471
rect 28816 21428 28868 21437
rect 28908 21471 28960 21480
rect 28908 21437 28917 21471
rect 28917 21437 28951 21471
rect 28951 21437 28960 21471
rect 28908 21428 28960 21437
rect 29460 21428 29512 21480
rect 30748 21428 30800 21480
rect 31300 21471 31352 21480
rect 31300 21437 31309 21471
rect 31309 21437 31343 21471
rect 31343 21437 31352 21471
rect 31300 21428 31352 21437
rect 32036 21428 32088 21480
rect 32496 21428 32548 21480
rect 33048 21428 33100 21480
rect 33600 21539 33652 21548
rect 33600 21505 33609 21539
rect 33609 21505 33643 21539
rect 33643 21505 33652 21539
rect 33600 21496 33652 21505
rect 33692 21471 33744 21480
rect 33692 21437 33701 21471
rect 33701 21437 33735 21471
rect 33735 21437 33744 21471
rect 33692 21428 33744 21437
rect 20076 21360 20128 21412
rect 15752 21292 15804 21344
rect 16856 21335 16908 21344
rect 16856 21301 16865 21335
rect 16865 21301 16899 21335
rect 16899 21301 16908 21335
rect 16856 21292 16908 21301
rect 17500 21292 17552 21344
rect 20352 21335 20404 21344
rect 20352 21301 20361 21335
rect 20361 21301 20395 21335
rect 20395 21301 20404 21335
rect 20352 21292 20404 21301
rect 20536 21292 20588 21344
rect 22376 21360 22428 21412
rect 21916 21292 21968 21344
rect 22100 21335 22152 21344
rect 22100 21301 22109 21335
rect 22109 21301 22143 21335
rect 22143 21301 22152 21335
rect 22100 21292 22152 21301
rect 24768 21335 24820 21344
rect 24768 21301 24777 21335
rect 24777 21301 24811 21335
rect 24811 21301 24820 21335
rect 24768 21292 24820 21301
rect 26148 21360 26200 21412
rect 30840 21360 30892 21412
rect 29368 21292 29420 21344
rect 30196 21292 30248 21344
rect 30472 21292 30524 21344
rect 31760 21292 31812 21344
rect 32496 21292 32548 21344
rect 32588 21292 32640 21344
rect 34428 21496 34480 21548
rect 34796 21539 34848 21548
rect 34796 21505 34805 21539
rect 34805 21505 34839 21539
rect 34839 21505 34848 21539
rect 34796 21496 34848 21505
rect 35164 21360 35216 21412
rect 36176 21471 36228 21480
rect 36176 21437 36185 21471
rect 36185 21437 36219 21471
rect 36219 21437 36228 21471
rect 36176 21428 36228 21437
rect 36636 21428 36688 21480
rect 37648 21428 37700 21480
rect 37740 21360 37792 21412
rect 35440 21292 35492 21344
rect 35716 21335 35768 21344
rect 35716 21301 35725 21335
rect 35725 21301 35759 21335
rect 35759 21301 35768 21335
rect 35716 21292 35768 21301
rect 36360 21292 36412 21344
rect 36820 21335 36872 21344
rect 36820 21301 36829 21335
rect 36829 21301 36863 21335
rect 36863 21301 36872 21335
rect 36820 21292 36872 21301
rect 37372 21335 37424 21344
rect 37372 21301 37381 21335
rect 37381 21301 37415 21335
rect 37415 21301 37424 21335
rect 37372 21292 37424 21301
rect 37556 21292 37608 21344
rect 38384 21428 38436 21480
rect 39028 21428 39080 21480
rect 39304 21428 39356 21480
rect 42248 21632 42300 21684
rect 42892 21632 42944 21684
rect 43260 21632 43312 21684
rect 45284 21632 45336 21684
rect 45560 21632 45612 21684
rect 47400 21632 47452 21684
rect 48228 21632 48280 21684
rect 41512 21564 41564 21616
rect 40684 21471 40736 21480
rect 39396 21360 39448 21412
rect 40684 21437 40693 21471
rect 40693 21437 40727 21471
rect 40727 21437 40736 21471
rect 40684 21428 40736 21437
rect 40776 21471 40828 21480
rect 40776 21437 40785 21471
rect 40785 21437 40819 21471
rect 40819 21437 40828 21471
rect 40776 21428 40828 21437
rect 41512 21428 41564 21480
rect 42248 21428 42300 21480
rect 43904 21539 43956 21548
rect 43904 21505 43913 21539
rect 43913 21505 43947 21539
rect 43947 21505 43956 21539
rect 43904 21496 43956 21505
rect 44272 21564 44324 21616
rect 44824 21564 44876 21616
rect 44548 21539 44600 21548
rect 44548 21505 44557 21539
rect 44557 21505 44591 21539
rect 44591 21505 44600 21539
rect 44548 21496 44600 21505
rect 44732 21496 44784 21548
rect 45008 21496 45060 21548
rect 45836 21539 45888 21548
rect 45836 21505 45845 21539
rect 45845 21505 45879 21539
rect 45879 21505 45888 21539
rect 45836 21496 45888 21505
rect 45928 21496 45980 21548
rect 48596 21564 48648 21616
rect 46848 21496 46900 21548
rect 48504 21496 48556 21548
rect 47584 21428 47636 21480
rect 45560 21360 45612 21412
rect 38292 21292 38344 21344
rect 40592 21292 40644 21344
rect 42064 21335 42116 21344
rect 42064 21301 42073 21335
rect 42073 21301 42107 21335
rect 42107 21301 42116 21335
rect 42064 21292 42116 21301
rect 42340 21292 42392 21344
rect 43720 21335 43772 21344
rect 43720 21301 43729 21335
rect 43729 21301 43763 21335
rect 43763 21301 43772 21335
rect 43720 21292 43772 21301
rect 44364 21335 44416 21344
rect 44364 21301 44373 21335
rect 44373 21301 44407 21335
rect 44407 21301 44416 21335
rect 44364 21292 44416 21301
rect 45008 21335 45060 21344
rect 45008 21301 45017 21335
rect 45017 21301 45051 21335
rect 45051 21301 45060 21335
rect 45008 21292 45060 21301
rect 45192 21292 45244 21344
rect 45744 21292 45796 21344
rect 48872 21292 48924 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 3424 21088 3476 21140
rect 6460 21088 6512 21140
rect 7656 21131 7708 21140
rect 7656 21097 7665 21131
rect 7665 21097 7699 21131
rect 7699 21097 7708 21131
rect 7656 21088 7708 21097
rect 9680 21088 9732 21140
rect 10416 21088 10468 21140
rect 3976 21020 4028 21072
rect 8024 21020 8076 21072
rect 9036 21063 9088 21072
rect 9036 21029 9045 21063
rect 9045 21029 9079 21063
rect 9079 21029 9088 21063
rect 9036 21020 9088 21029
rect 9588 21020 9640 21072
rect 2780 20859 2832 20868
rect 2780 20825 2789 20859
rect 2789 20825 2823 20859
rect 2823 20825 2832 20859
rect 2780 20816 2832 20825
rect 4160 20952 4212 21004
rect 5632 20952 5684 21004
rect 7012 20884 7064 20936
rect 8300 20952 8352 21004
rect 7840 20927 7892 20936
rect 7840 20893 7849 20927
rect 7849 20893 7883 20927
rect 7883 20893 7892 20927
rect 7840 20884 7892 20893
rect 9496 20884 9548 20936
rect 15292 21088 15344 21140
rect 16948 21131 17000 21140
rect 16948 21097 16957 21131
rect 16957 21097 16991 21131
rect 16991 21097 17000 21131
rect 16948 21088 17000 21097
rect 17224 21088 17276 21140
rect 20536 21088 20588 21140
rect 20628 21088 20680 21140
rect 21548 21088 21600 21140
rect 22284 21088 22336 21140
rect 24768 21088 24820 21140
rect 26240 21088 26292 21140
rect 30104 21088 30156 21140
rect 30564 21088 30616 21140
rect 12900 20952 12952 21004
rect 12532 20884 12584 20936
rect 13268 20952 13320 21004
rect 14188 20952 14240 21004
rect 14372 20995 14424 21004
rect 14372 20961 14381 20995
rect 14381 20961 14415 20995
rect 14415 20961 14424 20995
rect 14372 20952 14424 20961
rect 15016 20952 15068 21004
rect 18328 21020 18380 21072
rect 22836 21063 22888 21072
rect 22836 21029 22845 21063
rect 22845 21029 22879 21063
rect 22879 21029 22888 21063
rect 22836 21020 22888 21029
rect 13452 20884 13504 20936
rect 13820 20884 13872 20936
rect 15936 20884 15988 20936
rect 16764 20884 16816 20936
rect 17500 20995 17552 21004
rect 17500 20961 17509 20995
rect 17509 20961 17543 20995
rect 17543 20961 17552 20995
rect 17500 20952 17552 20961
rect 9956 20816 10008 20868
rect 12808 20816 12860 20868
rect 13084 20816 13136 20868
rect 13176 20816 13228 20868
rect 18788 20952 18840 21004
rect 21180 20952 21232 21004
rect 21732 20952 21784 21004
rect 21916 20952 21968 21004
rect 22744 20952 22796 21004
rect 23756 20995 23808 21004
rect 23756 20961 23765 20995
rect 23765 20961 23799 20995
rect 23799 20961 23808 20995
rect 23756 20952 23808 20961
rect 23848 20995 23900 21004
rect 23848 20961 23857 20995
rect 23857 20961 23891 20995
rect 23891 20961 23900 20995
rect 23848 20952 23900 20961
rect 26332 20995 26384 21004
rect 26332 20961 26341 20995
rect 26341 20961 26375 20995
rect 26375 20961 26384 20995
rect 26332 20952 26384 20961
rect 27528 20995 27580 21004
rect 27528 20961 27537 20995
rect 27537 20961 27571 20995
rect 27571 20961 27580 20995
rect 27528 20952 27580 20961
rect 29736 21063 29788 21072
rect 29736 21029 29745 21063
rect 29745 21029 29779 21063
rect 29779 21029 29788 21063
rect 29736 21020 29788 21029
rect 29000 20952 29052 21004
rect 30104 20952 30156 21004
rect 30748 20952 30800 21004
rect 35716 21088 35768 21140
rect 36912 21131 36964 21140
rect 36912 21097 36921 21131
rect 36921 21097 36955 21131
rect 36955 21097 36964 21131
rect 36912 21088 36964 21097
rect 37188 21088 37240 21140
rect 31760 21020 31812 21072
rect 32404 21020 32456 21072
rect 39212 21088 39264 21140
rect 40316 21088 40368 21140
rect 40500 21088 40552 21140
rect 44272 21088 44324 21140
rect 44916 21088 44968 21140
rect 45836 21131 45888 21140
rect 45836 21097 45845 21131
rect 45845 21097 45879 21131
rect 45879 21097 45888 21131
rect 45836 21088 45888 21097
rect 46020 21131 46072 21140
rect 46020 21097 46029 21131
rect 46029 21097 46063 21131
rect 46063 21097 46072 21131
rect 46020 21088 46072 21097
rect 46572 21088 46624 21140
rect 47584 21088 47636 21140
rect 48320 21088 48372 21140
rect 39304 21020 39356 21072
rect 8024 20748 8076 20800
rect 12256 20748 12308 20800
rect 12624 20748 12676 20800
rect 13728 20748 13780 20800
rect 14464 20748 14516 20800
rect 17960 20859 18012 20868
rect 17960 20825 17969 20859
rect 17969 20825 18003 20859
rect 18003 20825 18012 20859
rect 17960 20816 18012 20825
rect 20260 20816 20312 20868
rect 16396 20791 16448 20800
rect 16396 20757 16405 20791
rect 16405 20757 16439 20791
rect 16439 20757 16448 20791
rect 16396 20748 16448 20757
rect 17316 20791 17368 20800
rect 17316 20757 17325 20791
rect 17325 20757 17359 20791
rect 17359 20757 17368 20791
rect 17316 20748 17368 20757
rect 18604 20791 18656 20800
rect 18604 20757 18613 20791
rect 18613 20757 18647 20791
rect 18647 20757 18656 20791
rect 18604 20748 18656 20757
rect 22836 20884 22888 20936
rect 24768 20884 24820 20936
rect 28540 20884 28592 20936
rect 29920 20927 29972 20936
rect 29920 20893 29929 20927
rect 29929 20893 29963 20927
rect 29963 20893 29972 20927
rect 29920 20884 29972 20893
rect 22744 20816 22796 20868
rect 22560 20748 22612 20800
rect 23296 20748 23348 20800
rect 23664 20791 23716 20800
rect 23664 20757 23673 20791
rect 23673 20757 23707 20791
rect 23707 20757 23716 20791
rect 23664 20748 23716 20757
rect 25136 20748 25188 20800
rect 26792 20816 26844 20868
rect 27620 20816 27672 20868
rect 27804 20816 27856 20868
rect 31300 20884 31352 20936
rect 31852 20884 31904 20936
rect 30564 20816 30616 20868
rect 31576 20816 31628 20868
rect 26148 20791 26200 20800
rect 26148 20757 26157 20791
rect 26157 20757 26191 20791
rect 26191 20757 26200 20791
rect 26148 20748 26200 20757
rect 26332 20748 26384 20800
rect 28724 20791 28776 20800
rect 28724 20757 28733 20791
rect 28733 20757 28767 20791
rect 28767 20757 28776 20791
rect 28724 20748 28776 20757
rect 28908 20748 28960 20800
rect 30104 20748 30156 20800
rect 31300 20748 31352 20800
rect 31852 20748 31904 20800
rect 32864 20952 32916 21004
rect 33140 20952 33192 21004
rect 32312 20884 32364 20936
rect 33048 20816 33100 20868
rect 34888 20995 34940 21004
rect 34888 20961 34897 20995
rect 34897 20961 34931 20995
rect 34931 20961 34940 20995
rect 34888 20952 34940 20961
rect 36728 20952 36780 21004
rect 42340 21020 42392 21072
rect 42800 21020 42852 21072
rect 39948 20952 40000 21004
rect 40592 20995 40644 21004
rect 40592 20961 40601 20995
rect 40601 20961 40635 20995
rect 40635 20961 40644 20995
rect 40592 20952 40644 20961
rect 37648 20927 37700 20936
rect 37648 20893 37657 20927
rect 37657 20893 37691 20927
rect 37691 20893 37700 20927
rect 37648 20884 37700 20893
rect 39212 20884 39264 20936
rect 42432 20995 42484 21004
rect 42432 20961 42441 20995
rect 42441 20961 42475 20995
rect 42475 20961 42484 20995
rect 42432 20952 42484 20961
rect 42708 20995 42760 21004
rect 42708 20961 42717 20995
rect 42717 20961 42751 20995
rect 42751 20961 42760 20995
rect 42708 20952 42760 20961
rect 48780 20952 48832 21004
rect 42892 20884 42944 20936
rect 43812 20884 43864 20936
rect 44456 20884 44508 20936
rect 45100 20884 45152 20936
rect 46388 20884 46440 20936
rect 47032 20884 47084 20936
rect 47676 20884 47728 20936
rect 48228 20884 48280 20936
rect 49056 20927 49108 20936
rect 49056 20893 49065 20927
rect 49065 20893 49099 20927
rect 49099 20893 49108 20927
rect 49056 20884 49108 20893
rect 33784 20748 33836 20800
rect 34152 20748 34204 20800
rect 36636 20791 36688 20800
rect 36636 20757 36645 20791
rect 36645 20757 36679 20791
rect 36679 20757 36688 20791
rect 36636 20748 36688 20757
rect 37280 20791 37332 20800
rect 37280 20757 37289 20791
rect 37289 20757 37323 20791
rect 37323 20757 37332 20791
rect 37280 20748 37332 20757
rect 38568 20816 38620 20868
rect 40776 20748 40828 20800
rect 41328 20816 41380 20868
rect 42984 20816 43036 20868
rect 42800 20748 42852 20800
rect 44272 20748 44324 20800
rect 49240 20791 49292 20800
rect 49240 20757 49249 20791
rect 49249 20757 49283 20791
rect 49283 20757 49292 20791
rect 49240 20748 49292 20757
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 7288 20544 7340 20596
rect 1860 20408 1912 20460
rect 3608 20451 3660 20460
rect 3608 20417 3617 20451
rect 3617 20417 3651 20451
rect 3651 20417 3660 20451
rect 3608 20408 3660 20417
rect 2872 20340 2924 20392
rect 3884 20383 3936 20392
rect 3884 20349 3893 20383
rect 3893 20349 3927 20383
rect 3927 20349 3936 20383
rect 3884 20340 3936 20349
rect 5908 20408 5960 20460
rect 8852 20408 8904 20460
rect 9128 20451 9180 20460
rect 9128 20417 9137 20451
rect 9137 20417 9171 20451
rect 9171 20417 9180 20451
rect 9128 20408 9180 20417
rect 7196 20383 7248 20392
rect 7196 20349 7205 20383
rect 7205 20349 7239 20383
rect 7239 20349 7248 20383
rect 7196 20340 7248 20349
rect 8300 20340 8352 20392
rect 9404 20340 9456 20392
rect 10232 20408 10284 20460
rect 10508 20451 10560 20460
rect 10508 20417 10517 20451
rect 10517 20417 10551 20451
rect 10551 20417 10560 20451
rect 10508 20408 10560 20417
rect 11704 20519 11756 20528
rect 11704 20485 11713 20519
rect 11713 20485 11747 20519
rect 11747 20485 11756 20519
rect 11704 20476 11756 20485
rect 12256 20519 12308 20528
rect 12256 20485 12265 20519
rect 12265 20485 12299 20519
rect 12299 20485 12308 20519
rect 12256 20476 12308 20485
rect 13912 20544 13964 20596
rect 15108 20544 15160 20596
rect 15384 20544 15436 20596
rect 19064 20544 19116 20596
rect 15936 20476 15988 20528
rect 20444 20544 20496 20596
rect 20720 20587 20772 20596
rect 20720 20553 20729 20587
rect 20729 20553 20763 20587
rect 20763 20553 20772 20587
rect 20720 20544 20772 20553
rect 22008 20587 22060 20596
rect 22008 20553 22017 20587
rect 22017 20553 22051 20587
rect 22051 20553 22060 20587
rect 22008 20544 22060 20553
rect 22744 20587 22796 20596
rect 22744 20553 22753 20587
rect 22753 20553 22787 20587
rect 22787 20553 22796 20587
rect 22744 20544 22796 20553
rect 20076 20476 20128 20528
rect 20352 20476 20404 20528
rect 22468 20476 22520 20528
rect 12072 20451 12124 20460
rect 12072 20417 12081 20451
rect 12081 20417 12115 20451
rect 12115 20417 12124 20451
rect 12072 20408 12124 20417
rect 12716 20451 12768 20460
rect 12716 20417 12725 20451
rect 12725 20417 12759 20451
rect 12759 20417 12768 20451
rect 12716 20408 12768 20417
rect 15200 20408 15252 20460
rect 16120 20451 16172 20460
rect 16120 20417 16129 20451
rect 16129 20417 16163 20451
rect 16163 20417 16172 20451
rect 16120 20408 16172 20417
rect 16764 20408 16816 20460
rect 17408 20451 17460 20460
rect 17408 20417 17417 20451
rect 17417 20417 17451 20451
rect 17451 20417 17460 20451
rect 17408 20408 17460 20417
rect 18420 20408 18472 20460
rect 21088 20451 21140 20460
rect 21088 20417 21097 20451
rect 21097 20417 21131 20451
rect 21131 20417 21140 20451
rect 21088 20408 21140 20417
rect 22836 20408 22888 20460
rect 11612 20340 11664 20392
rect 12348 20340 12400 20392
rect 12624 20340 12676 20392
rect 11520 20272 11572 20324
rect 13084 20272 13136 20324
rect 13820 20383 13872 20392
rect 13820 20349 13829 20383
rect 13829 20349 13863 20383
rect 13863 20349 13872 20383
rect 13820 20340 13872 20349
rect 14188 20340 14240 20392
rect 17040 20340 17092 20392
rect 17776 20340 17828 20392
rect 15476 20272 15528 20324
rect 19800 20340 19852 20392
rect 21180 20383 21232 20392
rect 21180 20349 21189 20383
rect 21189 20349 21223 20383
rect 21223 20349 21232 20383
rect 21180 20340 21232 20349
rect 11152 20247 11204 20256
rect 11152 20213 11161 20247
rect 11161 20213 11195 20247
rect 11195 20213 11204 20247
rect 11152 20204 11204 20213
rect 12440 20204 12492 20256
rect 13636 20204 13688 20256
rect 16212 20247 16264 20256
rect 16212 20213 16221 20247
rect 16221 20213 16255 20247
rect 16255 20213 16264 20247
rect 16212 20204 16264 20213
rect 16764 20247 16816 20256
rect 16764 20213 16773 20247
rect 16773 20213 16807 20247
rect 16807 20213 16816 20247
rect 16764 20204 16816 20213
rect 16856 20204 16908 20256
rect 18328 20204 18380 20256
rect 25964 20544 26016 20596
rect 26056 20544 26108 20596
rect 27344 20544 27396 20596
rect 23480 20451 23532 20460
rect 23480 20417 23489 20451
rect 23489 20417 23523 20451
rect 23523 20417 23532 20451
rect 24400 20476 24452 20528
rect 24584 20476 24636 20528
rect 25504 20476 25556 20528
rect 27620 20476 27672 20528
rect 23480 20408 23532 20417
rect 26056 20408 26108 20460
rect 26240 20451 26292 20460
rect 26240 20417 26249 20451
rect 26249 20417 26283 20451
rect 26283 20417 26292 20451
rect 26240 20408 26292 20417
rect 27252 20451 27304 20460
rect 27252 20417 27261 20451
rect 27261 20417 27295 20451
rect 27295 20417 27304 20451
rect 27252 20408 27304 20417
rect 29644 20544 29696 20596
rect 29828 20544 29880 20596
rect 30104 20544 30156 20596
rect 29276 20476 29328 20528
rect 30012 20476 30064 20528
rect 30380 20476 30432 20528
rect 31208 20476 31260 20528
rect 33048 20476 33100 20528
rect 33968 20544 34020 20596
rect 35808 20544 35860 20596
rect 36176 20544 36228 20596
rect 36268 20476 36320 20528
rect 23388 20340 23440 20392
rect 23756 20340 23808 20392
rect 24124 20383 24176 20392
rect 24124 20349 24133 20383
rect 24133 20349 24167 20383
rect 24167 20349 24176 20383
rect 24124 20340 24176 20349
rect 24584 20340 24636 20392
rect 25412 20340 25464 20392
rect 25596 20383 25648 20392
rect 25596 20349 25605 20383
rect 25605 20349 25639 20383
rect 25639 20349 25648 20383
rect 25596 20340 25648 20349
rect 28540 20340 28592 20392
rect 29276 20340 29328 20392
rect 29736 20340 29788 20392
rect 30196 20340 30248 20392
rect 20352 20204 20404 20256
rect 21088 20204 21140 20256
rect 23848 20204 23900 20256
rect 27252 20272 27304 20324
rect 30380 20272 30432 20324
rect 34704 20408 34756 20460
rect 35256 20451 35308 20460
rect 35256 20417 35265 20451
rect 35265 20417 35299 20451
rect 35299 20417 35308 20451
rect 35256 20408 35308 20417
rect 35624 20408 35676 20460
rect 35808 20408 35860 20460
rect 37280 20544 37332 20596
rect 37924 20544 37976 20596
rect 42064 20544 42116 20596
rect 42156 20587 42208 20596
rect 42156 20553 42165 20587
rect 42165 20553 42199 20587
rect 42199 20553 42208 20587
rect 42156 20544 42208 20553
rect 42708 20544 42760 20596
rect 43812 20587 43864 20596
rect 43812 20553 43821 20587
rect 43821 20553 43855 20587
rect 43855 20553 43864 20587
rect 43812 20544 43864 20553
rect 44456 20544 44508 20596
rect 44732 20544 44784 20596
rect 44824 20587 44876 20596
rect 44824 20553 44833 20587
rect 44833 20553 44867 20587
rect 44867 20553 44876 20587
rect 44824 20544 44876 20553
rect 46756 20544 46808 20596
rect 47124 20544 47176 20596
rect 47676 20544 47728 20596
rect 38752 20476 38804 20528
rect 39764 20476 39816 20528
rect 40316 20519 40368 20528
rect 40316 20485 40325 20519
rect 40325 20485 40359 20519
rect 40359 20485 40368 20519
rect 40316 20476 40368 20485
rect 31208 20383 31260 20392
rect 31208 20349 31217 20383
rect 31217 20349 31251 20383
rect 31251 20349 31260 20383
rect 31208 20340 31260 20349
rect 32312 20383 32364 20392
rect 32312 20349 32321 20383
rect 32321 20349 32355 20383
rect 32355 20349 32364 20383
rect 32312 20340 32364 20349
rect 32680 20340 32732 20392
rect 31116 20272 31168 20324
rect 25780 20204 25832 20256
rect 27068 20204 27120 20256
rect 27712 20204 27764 20256
rect 29184 20204 29236 20256
rect 30288 20204 30340 20256
rect 30656 20247 30708 20256
rect 30656 20213 30665 20247
rect 30665 20213 30699 20247
rect 30699 20213 30708 20247
rect 30656 20204 30708 20213
rect 30932 20204 30984 20256
rect 33692 20272 33744 20324
rect 35716 20340 35768 20392
rect 36820 20408 36872 20460
rect 37188 20408 37240 20460
rect 43904 20476 43956 20528
rect 46388 20476 46440 20528
rect 49332 20476 49384 20528
rect 36728 20383 36780 20392
rect 36728 20349 36737 20383
rect 36737 20349 36771 20383
rect 36771 20349 36780 20383
rect 36728 20340 36780 20349
rect 37740 20383 37792 20392
rect 37740 20349 37749 20383
rect 37749 20349 37783 20383
rect 37783 20349 37792 20383
rect 37740 20340 37792 20349
rect 40960 20408 41012 20460
rect 36452 20272 36504 20324
rect 39028 20272 39080 20324
rect 41052 20340 41104 20392
rect 34060 20204 34112 20256
rect 35532 20204 35584 20256
rect 36084 20204 36136 20256
rect 39764 20204 39816 20256
rect 39948 20247 40000 20256
rect 39948 20213 39957 20247
rect 39957 20213 39991 20247
rect 39991 20213 40000 20247
rect 39948 20204 40000 20213
rect 41144 20272 41196 20324
rect 44088 20408 44140 20460
rect 47032 20408 47084 20460
rect 48596 20451 48648 20460
rect 48596 20417 48605 20451
rect 48605 20417 48639 20451
rect 48639 20417 48648 20451
rect 48596 20408 48648 20417
rect 49056 20451 49108 20460
rect 49056 20417 49065 20451
rect 49065 20417 49099 20451
rect 49099 20417 49108 20451
rect 49056 20408 49108 20417
rect 41512 20340 41564 20392
rect 42616 20340 42668 20392
rect 42984 20340 43036 20392
rect 45560 20340 45612 20392
rect 41972 20272 42024 20324
rect 43260 20272 43312 20324
rect 41788 20247 41840 20256
rect 41788 20213 41797 20247
rect 41797 20213 41831 20247
rect 41831 20213 41840 20247
rect 41788 20204 41840 20213
rect 48320 20204 48372 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 3608 20000 3660 20052
rect 11152 20000 11204 20052
rect 12348 20000 12400 20052
rect 12440 20000 12492 20052
rect 12624 20000 12676 20052
rect 15384 20000 15436 20052
rect 15476 20043 15528 20052
rect 15476 20009 15485 20043
rect 15485 20009 15519 20043
rect 15519 20009 15528 20043
rect 15476 20000 15528 20009
rect 16948 20000 17000 20052
rect 19524 20000 19576 20052
rect 21272 20000 21324 20052
rect 26700 20000 26752 20052
rect 26792 20043 26844 20052
rect 26792 20009 26801 20043
rect 26801 20009 26835 20043
rect 26835 20009 26844 20043
rect 26792 20000 26844 20009
rect 27712 20000 27764 20052
rect 28816 20000 28868 20052
rect 29276 20043 29328 20052
rect 29276 20009 29285 20043
rect 29285 20009 29319 20043
rect 29319 20009 29328 20043
rect 29276 20000 29328 20009
rect 29368 20000 29420 20052
rect 5264 19932 5316 19984
rect 10416 19932 10468 19984
rect 4528 19907 4580 19916
rect 4528 19873 4537 19907
rect 4537 19873 4571 19907
rect 4571 19873 4580 19907
rect 4528 19864 4580 19873
rect 6184 19864 6236 19916
rect 6368 19864 6420 19916
rect 9956 19864 10008 19916
rect 12348 19864 12400 19916
rect 1768 19839 1820 19848
rect 1768 19805 1777 19839
rect 1777 19805 1811 19839
rect 1811 19805 1820 19839
rect 1768 19796 1820 19805
rect 5724 19796 5776 19848
rect 6000 19839 6052 19848
rect 6000 19805 6009 19839
rect 6009 19805 6043 19839
rect 6043 19805 6052 19839
rect 6000 19796 6052 19805
rect 7840 19839 7892 19848
rect 7840 19805 7849 19839
rect 7849 19805 7883 19839
rect 7883 19805 7892 19839
rect 7840 19796 7892 19805
rect 7932 19796 7984 19848
rect 2780 19771 2832 19780
rect 2780 19737 2789 19771
rect 2789 19737 2823 19771
rect 2823 19737 2832 19771
rect 2780 19728 2832 19737
rect 4252 19728 4304 19780
rect 7656 19703 7708 19712
rect 7656 19669 7665 19703
rect 7665 19669 7699 19703
rect 7699 19669 7708 19703
rect 7656 19660 7708 19669
rect 10140 19728 10192 19780
rect 11704 19796 11756 19848
rect 14372 19975 14424 19984
rect 14372 19941 14381 19975
rect 14381 19941 14415 19975
rect 14415 19941 14424 19975
rect 14372 19932 14424 19941
rect 15200 19932 15252 19984
rect 15844 19932 15896 19984
rect 19800 19932 19852 19984
rect 21824 19932 21876 19984
rect 13820 19864 13872 19916
rect 17776 19864 17828 19916
rect 17868 19864 17920 19916
rect 13636 19796 13688 19848
rect 14096 19796 14148 19848
rect 15936 19839 15988 19848
rect 15936 19805 15945 19839
rect 15945 19805 15979 19839
rect 15979 19805 15988 19839
rect 15936 19796 15988 19805
rect 16948 19796 17000 19848
rect 18420 19796 18472 19848
rect 9220 19703 9272 19712
rect 9220 19669 9229 19703
rect 9229 19669 9263 19703
rect 9263 19669 9272 19703
rect 9220 19660 9272 19669
rect 16304 19728 16356 19780
rect 18604 19728 18656 19780
rect 10600 19660 10652 19712
rect 10784 19660 10836 19712
rect 12440 19660 12492 19712
rect 12532 19660 12584 19712
rect 13636 19660 13688 19712
rect 15108 19660 15160 19712
rect 17592 19660 17644 19712
rect 19892 19728 19944 19780
rect 23940 19932 23992 19984
rect 24124 19932 24176 19984
rect 23756 19907 23808 19916
rect 23756 19873 23765 19907
rect 23765 19873 23799 19907
rect 23799 19873 23808 19907
rect 23756 19864 23808 19873
rect 20444 19839 20496 19848
rect 20444 19805 20453 19839
rect 20453 19805 20487 19839
rect 20487 19805 20496 19839
rect 20444 19796 20496 19805
rect 21732 19796 21784 19848
rect 22468 19796 22520 19848
rect 25228 19864 25280 19916
rect 28632 19907 28684 19916
rect 28632 19873 28641 19907
rect 28641 19873 28675 19907
rect 28675 19873 28684 19907
rect 28632 19864 28684 19873
rect 28908 19932 28960 19984
rect 33508 20000 33560 20052
rect 33968 20000 34020 20052
rect 29460 19864 29512 19916
rect 29644 19864 29696 19916
rect 31392 19907 31444 19916
rect 31392 19873 31401 19907
rect 31401 19873 31435 19907
rect 31435 19873 31444 19907
rect 31392 19864 31444 19873
rect 31484 19907 31536 19916
rect 31484 19873 31493 19907
rect 31493 19873 31527 19907
rect 31527 19873 31536 19907
rect 31484 19864 31536 19873
rect 24676 19839 24728 19848
rect 24676 19805 24685 19839
rect 24685 19805 24719 19839
rect 24719 19805 24728 19839
rect 24676 19796 24728 19805
rect 27528 19796 27580 19848
rect 28816 19796 28868 19848
rect 30196 19839 30248 19848
rect 30196 19805 30205 19839
rect 30205 19805 30239 19839
rect 30239 19805 30248 19839
rect 30196 19796 30248 19805
rect 30380 19796 30432 19848
rect 31024 19796 31076 19848
rect 31300 19839 31352 19848
rect 31300 19805 31309 19839
rect 31309 19805 31343 19839
rect 31343 19805 31352 19839
rect 31300 19796 31352 19805
rect 20996 19728 21048 19780
rect 22100 19728 22152 19780
rect 23296 19728 23348 19780
rect 21732 19660 21784 19712
rect 22008 19660 22060 19712
rect 22468 19703 22520 19712
rect 22468 19669 22477 19703
rect 22477 19669 22511 19703
rect 22511 19669 22520 19703
rect 22468 19660 22520 19669
rect 23572 19703 23624 19712
rect 23572 19669 23581 19703
rect 23581 19669 23615 19703
rect 23615 19669 23624 19703
rect 23572 19660 23624 19669
rect 24492 19703 24544 19712
rect 24492 19669 24501 19703
rect 24501 19669 24535 19703
rect 24535 19669 24544 19703
rect 24492 19660 24544 19669
rect 24952 19703 25004 19712
rect 24952 19669 24961 19703
rect 24961 19669 24995 19703
rect 24995 19669 25004 19703
rect 24952 19660 25004 19669
rect 25044 19660 25096 19712
rect 25780 19660 25832 19712
rect 26240 19660 26292 19712
rect 27068 19660 27120 19712
rect 27252 19703 27304 19712
rect 27252 19669 27261 19703
rect 27261 19669 27295 19703
rect 27295 19669 27304 19703
rect 27252 19660 27304 19669
rect 31208 19728 31260 19780
rect 34428 19932 34480 19984
rect 34704 20000 34756 20052
rect 35348 20000 35400 20052
rect 37188 20000 37240 20052
rect 37280 20043 37332 20052
rect 37280 20009 37289 20043
rect 37289 20009 37323 20043
rect 37323 20009 37332 20043
rect 37280 20000 37332 20009
rect 35624 19932 35676 19984
rect 38752 19932 38804 19984
rect 40776 19932 40828 19984
rect 41512 19932 41564 19984
rect 41972 19932 42024 19984
rect 42616 20043 42668 20052
rect 42616 20009 42625 20043
rect 42625 20009 42659 20043
rect 42659 20009 42668 20043
rect 42616 20000 42668 20009
rect 43352 20043 43404 20052
rect 43352 20009 43361 20043
rect 43361 20009 43395 20043
rect 43395 20009 43404 20043
rect 43352 20000 43404 20009
rect 46204 20000 46256 20052
rect 47492 20043 47544 20052
rect 47492 20009 47501 20043
rect 47501 20009 47535 20043
rect 47535 20009 47544 20043
rect 47492 20000 47544 20009
rect 48964 20000 49016 20052
rect 43720 19932 43772 19984
rect 48780 19932 48832 19984
rect 32220 19864 32272 19916
rect 32864 19864 32916 19916
rect 32956 19864 33008 19916
rect 33876 19907 33928 19916
rect 33876 19873 33885 19907
rect 33885 19873 33919 19907
rect 33919 19873 33928 19907
rect 33876 19864 33928 19873
rect 34060 19907 34112 19916
rect 34060 19873 34069 19907
rect 34069 19873 34103 19907
rect 34103 19873 34112 19907
rect 34060 19864 34112 19873
rect 36084 19864 36136 19916
rect 37372 19864 37424 19916
rect 37464 19864 37516 19916
rect 37924 19864 37976 19916
rect 39028 19864 39080 19916
rect 39580 19864 39632 19916
rect 40132 19864 40184 19916
rect 32496 19839 32548 19848
rect 32496 19805 32505 19839
rect 32505 19805 32539 19839
rect 32539 19805 32548 19839
rect 32496 19796 32548 19805
rect 32772 19796 32824 19848
rect 35900 19796 35952 19848
rect 38844 19839 38896 19848
rect 38844 19805 38853 19839
rect 38853 19805 38887 19839
rect 38887 19805 38896 19839
rect 38844 19796 38896 19805
rect 29276 19660 29328 19712
rect 29460 19660 29512 19712
rect 30104 19703 30156 19712
rect 30104 19669 30113 19703
rect 30113 19669 30147 19703
rect 30147 19669 30156 19703
rect 30104 19660 30156 19669
rect 32128 19703 32180 19712
rect 32128 19669 32137 19703
rect 32137 19669 32171 19703
rect 32171 19669 32180 19703
rect 32128 19660 32180 19669
rect 32404 19660 32456 19712
rect 33048 19660 33100 19712
rect 34704 19728 34756 19780
rect 37280 19728 37332 19780
rect 40316 19796 40368 19848
rect 40500 19839 40552 19848
rect 40500 19805 40509 19839
rect 40509 19805 40543 19839
rect 40543 19805 40552 19839
rect 40500 19796 40552 19805
rect 43444 19796 43496 19848
rect 48688 19796 48740 19848
rect 35072 19660 35124 19712
rect 35348 19703 35400 19712
rect 35348 19669 35357 19703
rect 35357 19669 35391 19703
rect 35391 19669 35400 19703
rect 35348 19660 35400 19669
rect 35808 19660 35860 19712
rect 35900 19660 35952 19712
rect 36452 19703 36504 19712
rect 36452 19669 36461 19703
rect 36461 19669 36495 19703
rect 36495 19669 36504 19703
rect 36452 19660 36504 19669
rect 37648 19703 37700 19712
rect 37648 19669 37657 19703
rect 37657 19669 37691 19703
rect 37691 19669 37700 19703
rect 37648 19660 37700 19669
rect 38384 19660 38436 19712
rect 38568 19660 38620 19712
rect 38660 19660 38712 19712
rect 39856 19660 39908 19712
rect 40040 19703 40092 19712
rect 40040 19669 40049 19703
rect 40049 19669 40083 19703
rect 40083 19669 40092 19703
rect 40040 19660 40092 19669
rect 42340 19728 42392 19780
rect 44640 19728 44692 19780
rect 49332 19728 49384 19780
rect 40684 19660 40736 19712
rect 40960 19660 41012 19712
rect 45284 19660 45336 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 6276 19456 6328 19508
rect 7932 19456 7984 19508
rect 4620 19431 4672 19440
rect 4620 19397 4629 19431
rect 4629 19397 4663 19431
rect 4663 19397 4672 19431
rect 4620 19388 4672 19397
rect 6092 19388 6144 19440
rect 9864 19499 9916 19508
rect 9864 19465 9873 19499
rect 9873 19465 9907 19499
rect 9907 19465 9916 19499
rect 9864 19456 9916 19465
rect 9956 19456 10008 19508
rect 13360 19456 13412 19508
rect 16304 19499 16356 19508
rect 16304 19465 16313 19499
rect 16313 19465 16347 19499
rect 16347 19465 16356 19499
rect 16304 19456 16356 19465
rect 16672 19456 16724 19508
rect 21272 19456 21324 19508
rect 21732 19456 21784 19508
rect 23572 19456 23624 19508
rect 26148 19456 26200 19508
rect 28356 19456 28408 19508
rect 28724 19456 28776 19508
rect 32036 19456 32088 19508
rect 32220 19456 32272 19508
rect 32772 19456 32824 19508
rect 34612 19456 34664 19508
rect 34704 19499 34756 19508
rect 34704 19465 34713 19499
rect 34713 19465 34747 19499
rect 34747 19465 34756 19499
rect 34704 19456 34756 19465
rect 35164 19499 35216 19508
rect 35164 19465 35173 19499
rect 35173 19465 35207 19499
rect 35207 19465 35216 19499
rect 35164 19456 35216 19465
rect 36452 19456 36504 19508
rect 40500 19499 40552 19508
rect 40500 19465 40509 19499
rect 40509 19465 40543 19499
rect 40543 19465 40552 19499
rect 40500 19456 40552 19465
rect 40684 19456 40736 19508
rect 2872 19320 2924 19372
rect 5264 19320 5316 19372
rect 6828 19295 6880 19304
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 5264 19184 5316 19236
rect 7748 19320 7800 19372
rect 7932 19320 7984 19372
rect 8760 19363 8812 19372
rect 8760 19329 8769 19363
rect 8769 19329 8803 19363
rect 8803 19329 8812 19363
rect 8760 19320 8812 19329
rect 7012 19252 7064 19304
rect 2320 19116 2372 19168
rect 6184 19159 6236 19168
rect 6184 19125 6193 19159
rect 6193 19125 6227 19159
rect 6227 19125 6236 19159
rect 6184 19116 6236 19125
rect 6552 19116 6604 19168
rect 6644 19159 6696 19168
rect 6644 19125 6653 19159
rect 6653 19125 6687 19159
rect 6687 19125 6696 19159
rect 6644 19116 6696 19125
rect 7840 19184 7892 19236
rect 7932 19184 7984 19236
rect 8944 19184 8996 19236
rect 10324 19388 10376 19440
rect 11336 19388 11388 19440
rect 12072 19388 12124 19440
rect 9312 19320 9364 19372
rect 10140 19320 10192 19372
rect 9496 19252 9548 19304
rect 11796 19363 11848 19372
rect 11796 19329 11805 19363
rect 11805 19329 11839 19363
rect 11839 19329 11848 19363
rect 11796 19320 11848 19329
rect 15568 19388 15620 19440
rect 14556 19363 14608 19372
rect 14556 19329 14565 19363
rect 14565 19329 14599 19363
rect 14599 19329 14608 19363
rect 14556 19320 14608 19329
rect 17868 19388 17920 19440
rect 17224 19363 17276 19372
rect 17224 19329 17233 19363
rect 17233 19329 17267 19363
rect 17267 19329 17276 19363
rect 17224 19320 17276 19329
rect 17776 19320 17828 19372
rect 18604 19388 18656 19440
rect 20536 19388 20588 19440
rect 24032 19388 24084 19440
rect 24400 19388 24452 19440
rect 25780 19388 25832 19440
rect 29276 19388 29328 19440
rect 19432 19320 19484 19372
rect 20720 19320 20772 19372
rect 21824 19320 21876 19372
rect 22100 19320 22152 19372
rect 22468 19363 22520 19372
rect 22468 19329 22477 19363
rect 22477 19329 22511 19363
rect 22511 19329 22520 19363
rect 22468 19320 22520 19329
rect 23388 19320 23440 19372
rect 11152 19184 11204 19236
rect 13452 19252 13504 19304
rect 14004 19252 14056 19304
rect 16028 19252 16080 19304
rect 16948 19252 17000 19304
rect 17592 19252 17644 19304
rect 20076 19252 20128 19304
rect 20996 19252 21048 19304
rect 22008 19252 22060 19304
rect 22652 19295 22704 19304
rect 22652 19261 22661 19295
rect 22661 19261 22695 19295
rect 22695 19261 22704 19295
rect 22652 19252 22704 19261
rect 25320 19252 25372 19304
rect 10508 19116 10560 19168
rect 11796 19116 11848 19168
rect 12440 19159 12492 19168
rect 12440 19125 12449 19159
rect 12449 19125 12483 19159
rect 12483 19125 12492 19159
rect 12440 19116 12492 19125
rect 14372 19116 14424 19168
rect 14924 19116 14976 19168
rect 17684 19116 17736 19168
rect 22376 19184 22428 19236
rect 23480 19116 23532 19168
rect 25964 19320 26016 19372
rect 25688 19252 25740 19304
rect 25504 19227 25556 19236
rect 25504 19193 25513 19227
rect 25513 19193 25547 19227
rect 25547 19193 25556 19227
rect 25504 19184 25556 19193
rect 25872 19184 25924 19236
rect 26700 19320 26752 19372
rect 28632 19320 28684 19372
rect 28724 19320 28776 19372
rect 27620 19252 27672 19304
rect 27160 19116 27212 19168
rect 27252 19159 27304 19168
rect 27252 19125 27261 19159
rect 27261 19125 27295 19159
rect 27295 19125 27304 19159
rect 27252 19116 27304 19125
rect 27896 19252 27948 19304
rect 29644 19363 29696 19372
rect 29644 19329 29653 19363
rect 29653 19329 29687 19363
rect 29687 19329 29696 19363
rect 29644 19320 29696 19329
rect 30288 19363 30340 19372
rect 30288 19329 30297 19363
rect 30297 19329 30331 19363
rect 30331 19329 30340 19363
rect 30288 19320 30340 19329
rect 30840 19388 30892 19440
rect 35624 19388 35676 19440
rect 38476 19388 38528 19440
rect 38752 19388 38804 19440
rect 39856 19388 39908 19440
rect 30932 19320 30984 19372
rect 31208 19320 31260 19372
rect 31760 19320 31812 19372
rect 31852 19320 31904 19372
rect 32220 19320 32272 19372
rect 32312 19320 32364 19372
rect 32956 19320 33008 19372
rect 33048 19320 33100 19372
rect 28080 19184 28132 19236
rect 31576 19184 31628 19236
rect 33232 19252 33284 19304
rect 33508 19252 33560 19304
rect 33876 19363 33928 19372
rect 33876 19329 33885 19363
rect 33885 19329 33919 19363
rect 33919 19329 33928 19363
rect 33876 19320 33928 19329
rect 33968 19363 34020 19372
rect 33968 19329 33977 19363
rect 33977 19329 34011 19363
rect 34011 19329 34020 19363
rect 33968 19320 34020 19329
rect 34520 19320 34572 19372
rect 35164 19320 35216 19372
rect 35716 19320 35768 19372
rect 35992 19320 36044 19372
rect 34152 19295 34204 19304
rect 34152 19261 34161 19295
rect 34161 19261 34195 19295
rect 34195 19261 34204 19295
rect 34152 19252 34204 19261
rect 32036 19116 32088 19168
rect 32956 19184 33008 19236
rect 33968 19184 34020 19236
rect 34980 19252 35032 19304
rect 35808 19252 35860 19304
rect 37004 19252 37056 19304
rect 37188 19320 37240 19372
rect 37740 19320 37792 19372
rect 42156 19456 42208 19508
rect 42708 19499 42760 19508
rect 42708 19465 42717 19499
rect 42717 19465 42751 19499
rect 42751 19465 42760 19499
rect 42708 19456 42760 19465
rect 37832 19252 37884 19304
rect 40684 19252 40736 19304
rect 37188 19184 37240 19236
rect 39764 19184 39816 19236
rect 41972 19363 42024 19372
rect 41972 19329 41981 19363
rect 41981 19329 42015 19363
rect 42015 19329 42024 19363
rect 41972 19320 42024 19329
rect 48872 19456 48924 19508
rect 49148 19363 49200 19372
rect 49148 19329 49157 19363
rect 49157 19329 49191 19363
rect 49191 19329 49200 19363
rect 49148 19320 49200 19329
rect 47768 19252 47820 19304
rect 48412 19295 48464 19304
rect 48412 19261 48421 19295
rect 48421 19261 48455 19295
rect 48455 19261 48464 19295
rect 48412 19252 48464 19261
rect 47216 19184 47268 19236
rect 36636 19116 36688 19168
rect 36912 19159 36964 19168
rect 36912 19125 36921 19159
rect 36921 19125 36955 19159
rect 36955 19125 36964 19159
rect 36912 19116 36964 19125
rect 38752 19116 38804 19168
rect 39672 19159 39724 19168
rect 39672 19125 39681 19159
rect 39681 19125 39715 19159
rect 39715 19125 39724 19159
rect 39672 19116 39724 19125
rect 42432 19159 42484 19168
rect 42432 19125 42441 19159
rect 42441 19125 42475 19159
rect 42475 19125 42484 19159
rect 42432 19116 42484 19125
rect 48504 19116 48556 19168
rect 49056 19116 49108 19168
rect 49240 19159 49292 19168
rect 49240 19125 49249 19159
rect 49249 19125 49283 19159
rect 49283 19125 49292 19159
rect 49240 19116 49292 19125
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 6000 18912 6052 18964
rect 7196 18912 7248 18964
rect 12440 18912 12492 18964
rect 12532 18912 12584 18964
rect 14556 18912 14608 18964
rect 16120 18912 16172 18964
rect 16304 18912 16356 18964
rect 17316 18912 17368 18964
rect 19984 18912 20036 18964
rect 22376 18912 22428 18964
rect 6644 18844 6696 18896
rect 7748 18844 7800 18896
rect 10324 18844 10376 18896
rect 11796 18844 11848 18896
rect 13544 18844 13596 18896
rect 16396 18844 16448 18896
rect 3516 18776 3568 18828
rect 6184 18776 6236 18828
rect 9036 18776 9088 18828
rect 9680 18776 9732 18828
rect 13820 18776 13872 18828
rect 15292 18776 15344 18828
rect 17040 18819 17092 18828
rect 17040 18785 17049 18819
rect 17049 18785 17083 18819
rect 17083 18785 17092 18819
rect 17040 18776 17092 18785
rect 17684 18887 17736 18896
rect 17684 18853 17693 18887
rect 17693 18853 17727 18887
rect 17727 18853 17736 18887
rect 17684 18844 17736 18853
rect 19892 18844 19944 18896
rect 24032 18912 24084 18964
rect 25136 18912 25188 18964
rect 4252 18708 4304 18760
rect 2780 18683 2832 18692
rect 2780 18649 2789 18683
rect 2789 18649 2823 18683
rect 2823 18649 2832 18683
rect 2780 18640 2832 18649
rect 7380 18708 7432 18760
rect 5264 18572 5316 18624
rect 6552 18572 6604 18624
rect 8300 18640 8352 18692
rect 8484 18640 8536 18692
rect 9496 18640 9548 18692
rect 8668 18572 8720 18624
rect 9864 18572 9916 18624
rect 10048 18751 10100 18760
rect 10048 18717 10057 18751
rect 10057 18717 10091 18751
rect 10091 18717 10100 18751
rect 10048 18708 10100 18717
rect 12440 18708 12492 18760
rect 14188 18708 14240 18760
rect 14280 18751 14332 18760
rect 14280 18717 14289 18751
rect 14289 18717 14323 18751
rect 14323 18717 14332 18751
rect 14280 18708 14332 18717
rect 17132 18708 17184 18760
rect 19248 18708 19300 18760
rect 19432 18751 19484 18760
rect 19432 18717 19441 18751
rect 19441 18717 19475 18751
rect 19475 18717 19484 18751
rect 19432 18708 19484 18717
rect 19616 18751 19668 18760
rect 19616 18717 19625 18751
rect 19625 18717 19659 18751
rect 19659 18717 19668 18751
rect 19616 18708 19668 18717
rect 20628 18776 20680 18828
rect 21916 18776 21968 18828
rect 21272 18708 21324 18760
rect 25044 18776 25096 18828
rect 26516 18912 26568 18964
rect 28540 18912 28592 18964
rect 29552 18912 29604 18964
rect 30104 18912 30156 18964
rect 30748 18955 30800 18964
rect 30748 18921 30757 18955
rect 30757 18921 30791 18955
rect 30791 18921 30800 18955
rect 30748 18912 30800 18921
rect 27528 18844 27580 18896
rect 32036 18844 32088 18896
rect 33140 18912 33192 18964
rect 36544 18912 36596 18964
rect 40132 18912 40184 18964
rect 41052 18912 41104 18964
rect 42156 18912 42208 18964
rect 49240 18912 49292 18964
rect 22284 18751 22336 18760
rect 22284 18717 22293 18751
rect 22293 18717 22327 18751
rect 22327 18717 22336 18751
rect 22284 18708 22336 18717
rect 23572 18708 23624 18760
rect 23940 18708 23992 18760
rect 24032 18708 24084 18760
rect 26608 18776 26660 18828
rect 27160 18776 27212 18828
rect 10784 18683 10836 18692
rect 10784 18649 10793 18683
rect 10793 18649 10827 18683
rect 10827 18649 10836 18683
rect 10784 18640 10836 18649
rect 15844 18640 15896 18692
rect 16488 18640 16540 18692
rect 15200 18572 15252 18624
rect 15292 18572 15344 18624
rect 16304 18572 16356 18624
rect 16948 18615 17000 18624
rect 16948 18581 16957 18615
rect 16957 18581 16991 18615
rect 16991 18581 17000 18615
rect 16948 18572 17000 18581
rect 17868 18640 17920 18692
rect 19248 18572 19300 18624
rect 19340 18615 19392 18624
rect 19340 18581 19349 18615
rect 19349 18581 19383 18615
rect 19383 18581 19392 18615
rect 19340 18572 19392 18581
rect 20812 18572 20864 18624
rect 21456 18615 21508 18624
rect 21456 18581 21465 18615
rect 21465 18581 21499 18615
rect 21499 18581 21508 18615
rect 21456 18572 21508 18581
rect 21732 18572 21784 18624
rect 22560 18572 22612 18624
rect 23388 18572 23440 18624
rect 26148 18640 26200 18692
rect 26608 18640 26660 18692
rect 29644 18776 29696 18828
rect 29828 18776 29880 18828
rect 30748 18776 30800 18828
rect 32220 18776 32272 18828
rect 35348 18844 35400 18896
rect 37556 18844 37608 18896
rect 38200 18844 38252 18896
rect 33508 18776 33560 18828
rect 33876 18776 33928 18828
rect 35256 18776 35308 18828
rect 35624 18819 35676 18828
rect 35624 18785 35633 18819
rect 35633 18785 35667 18819
rect 35667 18785 35676 18819
rect 35624 18776 35676 18785
rect 38476 18776 38528 18828
rect 42248 18844 42300 18896
rect 42340 18776 42392 18828
rect 27528 18708 27580 18760
rect 28632 18708 28684 18760
rect 29184 18751 29236 18760
rect 29184 18717 29193 18751
rect 29193 18717 29227 18751
rect 29227 18717 29236 18751
rect 29184 18708 29236 18717
rect 29368 18708 29420 18760
rect 31208 18708 31260 18760
rect 37188 18708 37240 18760
rect 29460 18640 29512 18692
rect 31392 18640 31444 18692
rect 35900 18640 35952 18692
rect 36636 18640 36688 18692
rect 37832 18640 37884 18692
rect 41696 18708 41748 18760
rect 41604 18640 41656 18692
rect 48780 18708 48832 18760
rect 49148 18708 49200 18760
rect 42616 18640 42668 18692
rect 24032 18615 24084 18624
rect 24032 18581 24041 18615
rect 24041 18581 24075 18615
rect 24075 18581 24084 18615
rect 24032 18572 24084 18581
rect 24676 18572 24728 18624
rect 25412 18572 25464 18624
rect 26424 18572 26476 18624
rect 28540 18572 28592 18624
rect 29092 18615 29144 18624
rect 29092 18581 29101 18615
rect 29101 18581 29135 18615
rect 29135 18581 29144 18615
rect 29092 18572 29144 18581
rect 30012 18572 30064 18624
rect 30104 18615 30156 18624
rect 30104 18581 30113 18615
rect 30113 18581 30147 18615
rect 30147 18581 30156 18615
rect 30104 18572 30156 18581
rect 31300 18572 31352 18624
rect 32036 18572 32088 18624
rect 33600 18572 33652 18624
rect 33968 18572 34020 18624
rect 35808 18572 35860 18624
rect 36912 18572 36964 18624
rect 37740 18572 37792 18624
rect 38476 18615 38528 18624
rect 38476 18581 38485 18615
rect 38485 18581 38519 18615
rect 38519 18581 38528 18615
rect 38476 18572 38528 18581
rect 39212 18615 39264 18624
rect 39212 18581 39221 18615
rect 39221 18581 39255 18615
rect 39255 18581 39264 18615
rect 39212 18572 39264 18581
rect 42800 18572 42852 18624
rect 48412 18615 48464 18624
rect 48412 18581 48421 18615
rect 48421 18581 48455 18615
rect 48455 18581 48464 18615
rect 48412 18572 48464 18581
rect 48872 18572 48924 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 7288 18368 7340 18420
rect 4068 18300 4120 18352
rect 6368 18300 6420 18352
rect 6460 18300 6512 18352
rect 1768 18275 1820 18284
rect 1768 18241 1777 18275
rect 1777 18241 1811 18275
rect 1811 18241 1820 18275
rect 1768 18232 1820 18241
rect 3516 18275 3568 18284
rect 3516 18241 3525 18275
rect 3525 18241 3559 18275
rect 3559 18241 3568 18275
rect 3516 18232 3568 18241
rect 4712 18275 4764 18284
rect 4712 18241 4721 18275
rect 4721 18241 4755 18275
rect 4755 18241 4764 18275
rect 4712 18232 4764 18241
rect 2780 18207 2832 18216
rect 2780 18173 2789 18207
rect 2789 18173 2823 18207
rect 2823 18173 2832 18207
rect 2780 18164 2832 18173
rect 5172 18139 5224 18148
rect 5172 18105 5181 18139
rect 5181 18105 5215 18139
rect 5215 18105 5224 18139
rect 5172 18096 5224 18105
rect 7196 18275 7248 18284
rect 7196 18241 7205 18275
rect 7205 18241 7239 18275
rect 7239 18241 7248 18275
rect 7196 18232 7248 18241
rect 7748 18343 7800 18352
rect 7748 18309 7757 18343
rect 7757 18309 7791 18343
rect 7791 18309 7800 18343
rect 7748 18300 7800 18309
rect 6092 18096 6144 18148
rect 8668 18300 8720 18352
rect 10324 18368 10376 18420
rect 12808 18368 12860 18420
rect 15200 18411 15252 18420
rect 15200 18377 15209 18411
rect 15209 18377 15243 18411
rect 15243 18377 15252 18411
rect 15200 18368 15252 18377
rect 16212 18411 16264 18420
rect 16212 18377 16221 18411
rect 16221 18377 16255 18411
rect 16255 18377 16264 18411
rect 16212 18368 16264 18377
rect 17132 18411 17184 18420
rect 17132 18377 17141 18411
rect 17141 18377 17175 18411
rect 17175 18377 17184 18411
rect 17132 18368 17184 18377
rect 17868 18411 17920 18420
rect 17868 18377 17877 18411
rect 17877 18377 17911 18411
rect 17911 18377 17920 18411
rect 17868 18368 17920 18377
rect 9956 18232 10008 18284
rect 6460 18028 6512 18080
rect 7012 18071 7064 18080
rect 7012 18037 7021 18071
rect 7021 18037 7055 18071
rect 7055 18037 7064 18071
rect 7012 18028 7064 18037
rect 8300 18028 8352 18080
rect 8576 18028 8628 18080
rect 9588 18164 9640 18216
rect 11152 18232 11204 18284
rect 11796 18232 11848 18284
rect 14004 18232 14056 18284
rect 14188 18232 14240 18284
rect 10416 18139 10468 18148
rect 10416 18105 10425 18139
rect 10425 18105 10459 18139
rect 10459 18105 10468 18139
rect 10416 18096 10468 18105
rect 10784 18028 10836 18080
rect 11060 18028 11112 18080
rect 11244 18028 11296 18080
rect 12072 18096 12124 18148
rect 12348 18164 12400 18216
rect 12532 18096 12584 18148
rect 12440 18028 12492 18080
rect 13360 18164 13412 18216
rect 13452 18164 13504 18216
rect 15476 18232 15528 18284
rect 18420 18232 18472 18284
rect 19984 18300 20036 18352
rect 20168 18300 20220 18352
rect 19248 18275 19300 18284
rect 19248 18241 19257 18275
rect 19257 18241 19291 18275
rect 19291 18241 19300 18275
rect 19248 18232 19300 18241
rect 14004 18096 14056 18148
rect 16028 18164 16080 18216
rect 16764 18164 16816 18216
rect 17684 18164 17736 18216
rect 18604 18164 18656 18216
rect 19892 18207 19944 18216
rect 19892 18173 19901 18207
rect 19901 18173 19935 18207
rect 19935 18173 19944 18207
rect 19892 18164 19944 18173
rect 14280 18028 14332 18080
rect 16488 18096 16540 18148
rect 17040 18096 17092 18148
rect 21456 18368 21508 18420
rect 25136 18411 25188 18420
rect 25136 18377 25145 18411
rect 25145 18377 25179 18411
rect 25179 18377 25188 18411
rect 25136 18368 25188 18377
rect 25504 18368 25556 18420
rect 27252 18368 27304 18420
rect 21272 18300 21324 18352
rect 23204 18300 23256 18352
rect 23388 18343 23440 18352
rect 23388 18309 23397 18343
rect 23397 18309 23431 18343
rect 23431 18309 23440 18343
rect 23388 18300 23440 18309
rect 23848 18300 23900 18352
rect 27712 18368 27764 18420
rect 23296 18232 23348 18284
rect 24860 18232 24912 18284
rect 24584 18096 24636 18148
rect 15844 18028 15896 18080
rect 16580 18028 16632 18080
rect 17408 18071 17460 18080
rect 17408 18037 17417 18071
rect 17417 18037 17451 18071
rect 17451 18037 17460 18071
rect 17408 18028 17460 18037
rect 21732 18028 21784 18080
rect 22008 18071 22060 18080
rect 22008 18037 22017 18071
rect 22017 18037 22051 18071
rect 22051 18037 22060 18071
rect 22008 18028 22060 18037
rect 23204 18028 23256 18080
rect 30104 18368 30156 18420
rect 30380 18368 30432 18420
rect 31116 18368 31168 18420
rect 31760 18300 31812 18352
rect 25044 18275 25096 18284
rect 25044 18241 25053 18275
rect 25053 18241 25087 18275
rect 25087 18241 25096 18275
rect 25044 18232 25096 18241
rect 26516 18232 26568 18284
rect 28632 18232 28684 18284
rect 25228 18207 25280 18216
rect 25228 18173 25237 18207
rect 25237 18173 25271 18207
rect 25271 18173 25280 18207
rect 25228 18164 25280 18173
rect 26424 18207 26476 18216
rect 26424 18173 26433 18207
rect 26433 18173 26467 18207
rect 26467 18173 26476 18207
rect 26424 18164 26476 18173
rect 26792 18164 26844 18216
rect 30104 18275 30156 18284
rect 30104 18241 30113 18275
rect 30113 18241 30147 18275
rect 30147 18241 30156 18275
rect 33416 18368 33468 18420
rect 38476 18368 38528 18420
rect 39764 18411 39816 18420
rect 33600 18300 33652 18352
rect 34152 18300 34204 18352
rect 30104 18232 30156 18241
rect 28816 18164 28868 18216
rect 28908 18207 28960 18216
rect 28908 18173 28917 18207
rect 28917 18173 28951 18207
rect 28951 18173 28960 18207
rect 28908 18164 28960 18173
rect 29552 18164 29604 18216
rect 30564 18164 30616 18216
rect 31392 18207 31444 18216
rect 31392 18173 31401 18207
rect 31401 18173 31435 18207
rect 31435 18173 31444 18207
rect 31392 18164 31444 18173
rect 31576 18207 31628 18216
rect 31576 18173 31585 18207
rect 31585 18173 31619 18207
rect 31619 18173 31628 18207
rect 31576 18164 31628 18173
rect 32312 18164 32364 18216
rect 33140 18232 33192 18284
rect 32864 18207 32916 18216
rect 32864 18173 32873 18207
rect 32873 18173 32907 18207
rect 32907 18173 32916 18207
rect 32864 18164 32916 18173
rect 30472 18096 30524 18148
rect 32496 18096 32548 18148
rect 33876 18207 33928 18216
rect 33876 18173 33885 18207
rect 33885 18173 33919 18207
rect 33919 18173 33928 18207
rect 37372 18300 37424 18352
rect 37464 18300 37516 18352
rect 39764 18377 39773 18411
rect 39773 18377 39807 18411
rect 39807 18377 39816 18411
rect 39764 18368 39816 18377
rect 40040 18368 40092 18420
rect 42156 18411 42208 18420
rect 42156 18377 42165 18411
rect 42165 18377 42199 18411
rect 42199 18377 42208 18411
rect 42156 18368 42208 18377
rect 48780 18411 48832 18420
rect 48780 18377 48789 18411
rect 48789 18377 48823 18411
rect 48823 18377 48832 18411
rect 48780 18368 48832 18377
rect 38844 18300 38896 18352
rect 48412 18300 48464 18352
rect 37280 18232 37332 18284
rect 37924 18232 37976 18284
rect 39672 18232 39724 18284
rect 33876 18164 33928 18173
rect 36820 18164 36872 18216
rect 36912 18207 36964 18216
rect 36912 18173 36921 18207
rect 36921 18173 36955 18207
rect 36955 18173 36964 18207
rect 36912 18164 36964 18173
rect 37740 18164 37792 18216
rect 35716 18096 35768 18148
rect 37832 18096 37884 18148
rect 38292 18207 38344 18216
rect 38292 18173 38301 18207
rect 38301 18173 38335 18207
rect 38335 18173 38344 18207
rect 38292 18164 38344 18173
rect 38384 18164 38436 18216
rect 41696 18232 41748 18284
rect 41880 18232 41932 18284
rect 49056 18275 49108 18284
rect 41052 18164 41104 18216
rect 49056 18241 49065 18275
rect 49065 18241 49099 18275
rect 49099 18241 49108 18275
rect 49056 18232 49108 18241
rect 41604 18139 41656 18148
rect 41604 18105 41613 18139
rect 41613 18105 41647 18139
rect 41647 18105 41656 18139
rect 41604 18096 41656 18105
rect 25044 18028 25096 18080
rect 27160 18071 27212 18080
rect 27160 18037 27169 18071
rect 27169 18037 27203 18071
rect 27203 18037 27212 18071
rect 27160 18028 27212 18037
rect 27620 18028 27672 18080
rect 28632 18028 28684 18080
rect 29092 18028 29144 18080
rect 30932 18028 30984 18080
rect 31576 18028 31628 18080
rect 34520 18028 34572 18080
rect 35348 18071 35400 18080
rect 35348 18037 35357 18071
rect 35357 18037 35391 18071
rect 35391 18037 35400 18071
rect 35348 18028 35400 18037
rect 37188 18028 37240 18080
rect 37464 18028 37516 18080
rect 38844 18028 38896 18080
rect 41512 18028 41564 18080
rect 43352 18028 43404 18080
rect 48320 18028 48372 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 8392 17867 8444 17876
rect 8392 17833 8401 17867
rect 8401 17833 8435 17867
rect 8435 17833 8444 17867
rect 8392 17824 8444 17833
rect 11152 17824 11204 17876
rect 11428 17824 11480 17876
rect 14924 17824 14976 17876
rect 1768 17756 1820 17808
rect 8484 17756 8536 17808
rect 8852 17756 8904 17808
rect 9956 17756 10008 17808
rect 13360 17756 13412 17808
rect 16028 17867 16080 17876
rect 16028 17833 16037 17867
rect 16037 17833 16071 17867
rect 16071 17833 16080 17867
rect 16028 17824 16080 17833
rect 19892 17824 19944 17876
rect 20260 17824 20312 17876
rect 24492 17824 24544 17876
rect 24584 17867 24636 17876
rect 24584 17833 24593 17867
rect 24593 17833 24627 17867
rect 24627 17833 24636 17867
rect 24584 17824 24636 17833
rect 22836 17756 22888 17808
rect 30288 17824 30340 17876
rect 30380 17824 30432 17876
rect 30840 17824 30892 17876
rect 31944 17824 31996 17876
rect 32588 17824 32640 17876
rect 32864 17824 32916 17876
rect 33784 17867 33836 17876
rect 33784 17833 33793 17867
rect 33793 17833 33827 17867
rect 33827 17833 33836 17867
rect 33784 17824 33836 17833
rect 34704 17824 34756 17876
rect 24768 17756 24820 17808
rect 1216 17688 1268 17740
rect 3332 17688 3384 17740
rect 7012 17688 7064 17740
rect 4344 17620 4396 17672
rect 4896 17620 4948 17672
rect 8576 17663 8628 17672
rect 8576 17629 8585 17663
rect 8585 17629 8619 17663
rect 8619 17629 8628 17663
rect 8576 17620 8628 17629
rect 9404 17663 9456 17672
rect 9404 17629 9413 17663
rect 9413 17629 9447 17663
rect 9447 17629 9456 17663
rect 9404 17620 9456 17629
rect 4988 17484 5040 17536
rect 9680 17484 9732 17536
rect 9864 17527 9916 17536
rect 9864 17493 9873 17527
rect 9873 17493 9907 17527
rect 9907 17493 9916 17527
rect 9864 17484 9916 17493
rect 10324 17527 10376 17536
rect 10324 17493 10333 17527
rect 10333 17493 10367 17527
rect 10367 17493 10376 17527
rect 10324 17484 10376 17493
rect 10508 17731 10560 17740
rect 10508 17697 10517 17731
rect 10517 17697 10551 17731
rect 10551 17697 10560 17731
rect 10508 17688 10560 17697
rect 10784 17620 10836 17672
rect 12348 17688 12400 17740
rect 12716 17688 12768 17740
rect 14280 17731 14332 17740
rect 14280 17697 14289 17731
rect 14289 17697 14323 17731
rect 14323 17697 14332 17731
rect 14280 17688 14332 17697
rect 15108 17688 15160 17740
rect 15200 17688 15252 17740
rect 16672 17688 16724 17740
rect 12440 17620 12492 17672
rect 13544 17663 13596 17672
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 13544 17620 13596 17629
rect 15844 17620 15896 17672
rect 11336 17595 11388 17604
rect 11336 17561 11345 17595
rect 11345 17561 11379 17595
rect 11379 17561 11388 17595
rect 11336 17552 11388 17561
rect 14556 17595 14608 17604
rect 14556 17561 14565 17595
rect 14565 17561 14599 17595
rect 14599 17561 14608 17595
rect 14556 17552 14608 17561
rect 17868 17620 17920 17672
rect 18328 17688 18380 17740
rect 18512 17688 18564 17740
rect 18604 17688 18656 17740
rect 19340 17688 19392 17740
rect 20444 17688 20496 17740
rect 21088 17688 21140 17740
rect 22284 17688 22336 17740
rect 25044 17731 25096 17740
rect 25044 17697 25053 17731
rect 25053 17697 25087 17731
rect 25087 17697 25096 17731
rect 25044 17688 25096 17697
rect 28816 17756 28868 17808
rect 29000 17756 29052 17808
rect 33968 17756 34020 17808
rect 37372 17756 37424 17808
rect 25596 17688 25648 17740
rect 26608 17688 26660 17740
rect 19524 17620 19576 17672
rect 11520 17484 11572 17536
rect 11704 17484 11756 17536
rect 12256 17484 12308 17536
rect 13452 17484 13504 17536
rect 14372 17484 14424 17536
rect 18328 17552 18380 17604
rect 15936 17484 15988 17536
rect 16580 17484 16632 17536
rect 18972 17484 19024 17536
rect 22008 17620 22060 17672
rect 24952 17620 25004 17672
rect 25228 17620 25280 17672
rect 25780 17620 25832 17672
rect 20352 17552 20404 17604
rect 20904 17552 20956 17604
rect 23296 17552 23348 17604
rect 21364 17484 21416 17536
rect 21916 17527 21968 17536
rect 21916 17493 21925 17527
rect 21925 17493 21959 17527
rect 21959 17493 21968 17527
rect 21916 17484 21968 17493
rect 25044 17484 25096 17536
rect 26056 17484 26108 17536
rect 28356 17688 28408 17740
rect 28816 17620 28868 17672
rect 30380 17620 30432 17672
rect 31668 17688 31720 17740
rect 33232 17731 33284 17740
rect 33232 17697 33241 17731
rect 33241 17697 33275 17731
rect 33275 17697 33284 17731
rect 33232 17688 33284 17697
rect 33692 17688 33744 17740
rect 34060 17688 34112 17740
rect 31024 17620 31076 17672
rect 31944 17620 31996 17672
rect 34612 17688 34664 17740
rect 34888 17688 34940 17740
rect 35716 17688 35768 17740
rect 36084 17731 36136 17740
rect 36084 17697 36093 17731
rect 36093 17697 36127 17731
rect 36127 17697 36136 17731
rect 36084 17688 36136 17697
rect 36636 17688 36688 17740
rect 32496 17552 32548 17604
rect 35624 17620 35676 17672
rect 37188 17620 37240 17672
rect 37464 17620 37516 17672
rect 38568 17824 38620 17876
rect 42340 17867 42392 17876
rect 42340 17833 42349 17867
rect 42349 17833 42383 17867
rect 42383 17833 42392 17867
rect 42340 17824 42392 17833
rect 42616 17867 42668 17876
rect 42616 17833 42625 17867
rect 42625 17833 42659 17867
rect 42659 17833 42668 17867
rect 42616 17824 42668 17833
rect 39764 17756 39816 17808
rect 38568 17731 38620 17740
rect 38568 17697 38577 17731
rect 38577 17697 38611 17731
rect 38611 17697 38620 17731
rect 38568 17688 38620 17697
rect 39212 17731 39264 17740
rect 39212 17697 39221 17731
rect 39221 17697 39255 17731
rect 39255 17697 39264 17731
rect 39212 17688 39264 17697
rect 39948 17688 40000 17740
rect 28908 17484 28960 17536
rect 29276 17527 29328 17536
rect 29276 17493 29285 17527
rect 29285 17493 29319 17527
rect 29319 17493 29328 17527
rect 29276 17484 29328 17493
rect 34520 17552 34572 17604
rect 34980 17552 35032 17604
rect 32772 17527 32824 17536
rect 32772 17493 32781 17527
rect 32781 17493 32815 17527
rect 32815 17493 32824 17527
rect 32772 17484 32824 17493
rect 33784 17484 33836 17536
rect 34704 17484 34756 17536
rect 35348 17527 35400 17536
rect 35348 17493 35357 17527
rect 35357 17493 35391 17527
rect 35391 17493 35400 17527
rect 35348 17484 35400 17493
rect 40316 17552 40368 17604
rect 37832 17484 37884 17536
rect 38844 17484 38896 17536
rect 40224 17484 40276 17536
rect 40592 17620 40644 17672
rect 41880 17756 41932 17808
rect 49056 17663 49108 17672
rect 49056 17629 49065 17663
rect 49065 17629 49099 17663
rect 49099 17629 49108 17663
rect 49056 17620 49108 17629
rect 48412 17552 48464 17604
rect 42064 17484 42116 17536
rect 49148 17484 49200 17536
rect 49240 17527 49292 17536
rect 49240 17493 49249 17527
rect 49249 17493 49283 17527
rect 49283 17493 49292 17527
rect 49240 17484 49292 17493
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 4436 17280 4488 17332
rect 4804 17323 4856 17332
rect 4804 17289 4813 17323
rect 4813 17289 4847 17323
rect 4847 17289 4856 17323
rect 4804 17280 4856 17289
rect 5080 17280 5132 17332
rect 8300 17280 8352 17332
rect 8760 17280 8812 17332
rect 9956 17280 10008 17332
rect 12532 17280 12584 17332
rect 14004 17323 14056 17332
rect 14004 17289 14013 17323
rect 14013 17289 14047 17323
rect 14047 17289 14056 17323
rect 14004 17280 14056 17289
rect 15384 17280 15436 17332
rect 17684 17280 17736 17332
rect 18972 17280 19024 17332
rect 24216 17280 24268 17332
rect 24768 17280 24820 17332
rect 24860 17323 24912 17332
rect 24860 17289 24869 17323
rect 24869 17289 24903 17323
rect 24903 17289 24912 17323
rect 24860 17280 24912 17289
rect 27804 17323 27856 17332
rect 27804 17289 27813 17323
rect 27813 17289 27847 17323
rect 27847 17289 27856 17323
rect 27804 17280 27856 17289
rect 29092 17323 29144 17332
rect 29092 17289 29101 17323
rect 29101 17289 29135 17323
rect 29135 17289 29144 17323
rect 29092 17280 29144 17289
rect 29920 17280 29972 17332
rect 32036 17280 32088 17332
rect 32772 17280 32824 17332
rect 36268 17280 36320 17332
rect 37648 17280 37700 17332
rect 38384 17280 38436 17332
rect 1308 17076 1360 17128
rect 4988 17187 5040 17196
rect 4988 17153 4997 17187
rect 4997 17153 5031 17187
rect 5031 17153 5040 17187
rect 4988 17144 5040 17153
rect 5632 17187 5684 17196
rect 5632 17153 5641 17187
rect 5641 17153 5675 17187
rect 5675 17153 5684 17187
rect 5632 17144 5684 17153
rect 6552 17187 6604 17196
rect 6552 17153 6561 17187
rect 6561 17153 6595 17187
rect 6595 17153 6604 17187
rect 6552 17144 6604 17153
rect 7104 17144 7156 17196
rect 9864 17212 9916 17264
rect 12440 17212 12492 17264
rect 20168 17212 20220 17264
rect 20904 17212 20956 17264
rect 26516 17255 26568 17264
rect 26516 17221 26525 17255
rect 26525 17221 26559 17255
rect 26559 17221 26568 17255
rect 26516 17212 26568 17221
rect 27068 17212 27120 17264
rect 27988 17212 28040 17264
rect 30104 17212 30156 17264
rect 30748 17212 30800 17264
rect 6644 17076 6696 17128
rect 9312 17187 9364 17196
rect 9312 17153 9321 17187
rect 9321 17153 9355 17187
rect 9355 17153 9364 17187
rect 9312 17144 9364 17153
rect 9956 17187 10008 17196
rect 9956 17153 9965 17187
rect 9965 17153 9999 17187
rect 9999 17153 10008 17187
rect 9956 17144 10008 17153
rect 11428 17144 11480 17196
rect 12164 17144 12216 17196
rect 12624 17144 12676 17196
rect 15384 17144 15436 17196
rect 4160 16940 4212 16992
rect 8024 16940 8076 16992
rect 10600 17076 10652 17128
rect 10876 17119 10928 17128
rect 10876 17085 10885 17119
rect 10885 17085 10919 17119
rect 10919 17085 10928 17119
rect 10876 17076 10928 17085
rect 9128 17051 9180 17060
rect 9128 17017 9137 17051
rect 9137 17017 9171 17051
rect 9171 17017 9180 17051
rect 9128 17008 9180 17017
rect 12164 17008 12216 17060
rect 12440 17051 12492 17060
rect 12440 17017 12449 17051
rect 12449 17017 12483 17051
rect 12483 17017 12492 17051
rect 15476 17076 15528 17128
rect 16580 17144 16632 17196
rect 18512 17144 18564 17196
rect 19340 17187 19392 17196
rect 19340 17153 19349 17187
rect 19349 17153 19383 17187
rect 19383 17153 19392 17187
rect 19340 17144 19392 17153
rect 22192 17187 22244 17196
rect 22192 17153 22201 17187
rect 22201 17153 22235 17187
rect 22235 17153 22244 17187
rect 22192 17144 22244 17153
rect 22284 17144 22336 17196
rect 24032 17144 24084 17196
rect 24952 17144 25004 17196
rect 16120 17119 16172 17128
rect 16120 17085 16129 17119
rect 16129 17085 16163 17119
rect 16163 17085 16172 17119
rect 16120 17076 16172 17085
rect 12440 17008 12492 17017
rect 12532 16940 12584 16992
rect 13452 16940 13504 16992
rect 14832 17008 14884 17060
rect 14740 16940 14792 16992
rect 15016 16940 15068 16992
rect 15568 17051 15620 17060
rect 15568 17017 15577 17051
rect 15577 17017 15611 17051
rect 15611 17017 15620 17051
rect 15568 17008 15620 17017
rect 17040 17008 17092 17060
rect 16948 16940 17000 16992
rect 17408 17119 17460 17128
rect 17408 17085 17417 17119
rect 17417 17085 17451 17119
rect 17451 17085 17460 17119
rect 17408 17076 17460 17085
rect 17868 17076 17920 17128
rect 18604 16940 18656 16992
rect 20076 17076 20128 17128
rect 22376 17076 22428 17128
rect 25504 17119 25556 17128
rect 25504 17085 25513 17119
rect 25513 17085 25547 17119
rect 25547 17085 25556 17119
rect 25504 17076 25556 17085
rect 27804 17144 27856 17196
rect 29368 17144 29420 17196
rect 32496 17212 32548 17264
rect 32588 17255 32640 17264
rect 32588 17221 32597 17255
rect 32597 17221 32631 17255
rect 32631 17221 32640 17255
rect 32588 17212 32640 17221
rect 34152 17212 34204 17264
rect 35808 17212 35860 17264
rect 41604 17280 41656 17332
rect 42616 17280 42668 17332
rect 48412 17323 48464 17332
rect 48412 17289 48421 17323
rect 48421 17289 48455 17323
rect 48455 17289 48464 17323
rect 48412 17280 48464 17289
rect 34612 17187 34664 17196
rect 34612 17153 34621 17187
rect 34621 17153 34655 17187
rect 34655 17153 34664 17187
rect 34612 17144 34664 17153
rect 36360 17187 36412 17196
rect 36360 17153 36369 17187
rect 36369 17153 36403 17187
rect 36403 17153 36412 17187
rect 36360 17144 36412 17153
rect 38384 17144 38436 17196
rect 38568 17144 38620 17196
rect 41052 17187 41104 17196
rect 41052 17153 41061 17187
rect 41061 17153 41095 17187
rect 41095 17153 41104 17187
rect 41052 17144 41104 17153
rect 48780 17144 48832 17196
rect 49240 17144 49292 17196
rect 22008 17051 22060 17060
rect 22008 17017 22017 17051
rect 22017 17017 22051 17051
rect 22051 17017 22060 17051
rect 22008 17008 22060 17017
rect 24492 17008 24544 17060
rect 20168 16940 20220 16992
rect 26608 16940 26660 16992
rect 27896 17008 27948 17060
rect 28080 17076 28132 17128
rect 29092 17076 29144 17128
rect 29644 17076 29696 17128
rect 30748 17076 30800 17128
rect 29000 16940 29052 16992
rect 29460 16940 29512 16992
rect 30564 16940 30616 16992
rect 31208 16940 31260 16992
rect 31392 16940 31444 16992
rect 31760 16940 31812 16992
rect 31944 16940 31996 16992
rect 33232 17076 33284 17128
rect 34244 17076 34296 17128
rect 34888 17076 34940 17128
rect 35440 17076 35492 17128
rect 36544 17119 36596 17128
rect 36544 17085 36553 17119
rect 36553 17085 36587 17119
rect 36587 17085 36596 17119
rect 36544 17076 36596 17085
rect 38752 17076 38804 17128
rect 33692 17008 33744 17060
rect 34980 17008 35032 17060
rect 33876 16940 33928 16992
rect 34244 16940 34296 16992
rect 37740 17008 37792 17060
rect 43352 17076 43404 17128
rect 37096 16940 37148 16992
rect 37372 16940 37424 16992
rect 38568 16940 38620 16992
rect 40592 16983 40644 16992
rect 40592 16949 40601 16983
rect 40601 16949 40635 16983
rect 40635 16949 40644 16983
rect 40592 16940 40644 16949
rect 48688 16940 48740 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 5816 16736 5868 16788
rect 8576 16736 8628 16788
rect 8668 16736 8720 16788
rect 10232 16736 10284 16788
rect 10876 16736 10928 16788
rect 14464 16736 14516 16788
rect 14740 16736 14792 16788
rect 16212 16736 16264 16788
rect 5632 16668 5684 16720
rect 8484 16668 8536 16720
rect 16028 16668 16080 16720
rect 16488 16668 16540 16720
rect 16948 16736 17000 16788
rect 17592 16736 17644 16788
rect 19248 16736 19300 16788
rect 23296 16736 23348 16788
rect 29368 16736 29420 16788
rect 32128 16736 32180 16788
rect 33508 16736 33560 16788
rect 34152 16736 34204 16788
rect 34796 16736 34848 16788
rect 35900 16736 35952 16788
rect 36360 16736 36412 16788
rect 37004 16736 37056 16788
rect 41052 16736 41104 16788
rect 48780 16779 48832 16788
rect 48780 16745 48789 16779
rect 48789 16745 48823 16779
rect 48823 16745 48832 16779
rect 48780 16736 48832 16745
rect 17408 16668 17460 16720
rect 8300 16643 8352 16652
rect 8300 16609 8309 16643
rect 8309 16609 8343 16643
rect 8343 16609 8352 16643
rect 8300 16600 8352 16609
rect 8944 16600 8996 16652
rect 10140 16600 10192 16652
rect 10416 16600 10468 16652
rect 13452 16643 13504 16652
rect 13452 16609 13461 16643
rect 13461 16609 13495 16643
rect 13495 16609 13504 16643
rect 13452 16600 13504 16609
rect 14004 16600 14056 16652
rect 14096 16643 14148 16652
rect 14096 16609 14105 16643
rect 14105 16609 14139 16643
rect 14139 16609 14148 16643
rect 14096 16600 14148 16609
rect 14372 16600 14424 16652
rect 4068 16532 4120 16584
rect 4160 16575 4212 16584
rect 4160 16541 4169 16575
rect 4169 16541 4203 16575
rect 4203 16541 4212 16575
rect 4160 16532 4212 16541
rect 4804 16575 4856 16584
rect 4804 16541 4813 16575
rect 4813 16541 4847 16575
rect 4847 16541 4856 16575
rect 4804 16532 4856 16541
rect 6368 16532 6420 16584
rect 6460 16532 6512 16584
rect 8024 16532 8076 16584
rect 10048 16575 10100 16584
rect 10048 16541 10057 16575
rect 10057 16541 10091 16575
rect 10091 16541 10100 16575
rect 10048 16532 10100 16541
rect 1308 16464 1360 16516
rect 9404 16507 9456 16516
rect 9404 16473 9413 16507
rect 9413 16473 9447 16507
rect 9447 16473 9456 16507
rect 9404 16464 9456 16473
rect 9588 16464 9640 16516
rect 3976 16439 4028 16448
rect 3976 16405 3985 16439
rect 3985 16405 4019 16439
rect 4019 16405 4028 16439
rect 3976 16396 4028 16405
rect 5356 16396 5408 16448
rect 6920 16396 6972 16448
rect 8852 16396 8904 16448
rect 8944 16396 8996 16448
rect 11244 16532 11296 16584
rect 11336 16532 11388 16584
rect 12440 16532 12492 16584
rect 13636 16532 13688 16584
rect 14832 16575 14884 16584
rect 14832 16541 14841 16575
rect 14841 16541 14875 16575
rect 14875 16541 14884 16575
rect 14832 16532 14884 16541
rect 11888 16464 11940 16516
rect 12072 16464 12124 16516
rect 15108 16600 15160 16652
rect 20168 16668 20220 16720
rect 20904 16668 20956 16720
rect 21088 16643 21140 16652
rect 21088 16609 21097 16643
rect 21097 16609 21131 16643
rect 21131 16609 21140 16643
rect 21088 16600 21140 16609
rect 22744 16600 22796 16652
rect 23940 16668 23992 16720
rect 24032 16668 24084 16720
rect 29000 16668 29052 16720
rect 30380 16668 30432 16720
rect 30472 16668 30524 16720
rect 31024 16668 31076 16720
rect 32864 16668 32916 16720
rect 34612 16668 34664 16720
rect 15752 16575 15804 16584
rect 15752 16541 15761 16575
rect 15761 16541 15795 16575
rect 15795 16541 15804 16575
rect 15752 16532 15804 16541
rect 16672 16464 16724 16516
rect 11520 16439 11572 16448
rect 11520 16405 11529 16439
rect 11529 16405 11563 16439
rect 11563 16405 11572 16439
rect 11520 16396 11572 16405
rect 11612 16439 11664 16448
rect 11612 16405 11621 16439
rect 11621 16405 11655 16439
rect 11655 16405 11664 16439
rect 11612 16396 11664 16405
rect 11980 16396 12032 16448
rect 12992 16439 13044 16448
rect 12992 16405 13001 16439
rect 13001 16405 13035 16439
rect 13035 16405 13044 16439
rect 12992 16396 13044 16405
rect 14464 16439 14516 16448
rect 14464 16405 14473 16439
rect 14473 16405 14507 16439
rect 14507 16405 14516 16439
rect 14464 16396 14516 16405
rect 18328 16464 18380 16516
rect 19248 16464 19300 16516
rect 20720 16464 20772 16516
rect 19340 16396 19392 16448
rect 19432 16439 19484 16448
rect 19432 16405 19441 16439
rect 19441 16405 19475 16439
rect 19475 16405 19484 16439
rect 19432 16396 19484 16405
rect 19800 16439 19852 16448
rect 19800 16405 19809 16439
rect 19809 16405 19843 16439
rect 19843 16405 19852 16439
rect 19800 16396 19852 16405
rect 20904 16464 20956 16516
rect 23756 16464 23808 16516
rect 24860 16600 24912 16652
rect 28356 16600 28408 16652
rect 29184 16600 29236 16652
rect 28448 16532 28500 16584
rect 22376 16396 22428 16448
rect 22836 16439 22888 16448
rect 22836 16405 22845 16439
rect 22845 16405 22879 16439
rect 22879 16405 22888 16439
rect 22836 16396 22888 16405
rect 23296 16439 23348 16448
rect 23296 16405 23305 16439
rect 23305 16405 23339 16439
rect 23339 16405 23348 16439
rect 23296 16396 23348 16405
rect 23480 16396 23532 16448
rect 24308 16396 24360 16448
rect 25780 16464 25832 16516
rect 26608 16464 26660 16516
rect 27528 16464 27580 16516
rect 28908 16532 28960 16584
rect 29736 16532 29788 16584
rect 29920 16600 29972 16652
rect 31392 16600 31444 16652
rect 32496 16600 32548 16652
rect 32956 16600 33008 16652
rect 34796 16600 34848 16652
rect 33600 16532 33652 16584
rect 37372 16668 37424 16720
rect 35716 16643 35768 16652
rect 35716 16609 35725 16643
rect 35725 16609 35759 16643
rect 35759 16609 35768 16643
rect 35716 16600 35768 16609
rect 36728 16575 36780 16584
rect 36728 16541 36737 16575
rect 36737 16541 36771 16575
rect 36771 16541 36780 16575
rect 36728 16532 36780 16541
rect 37004 16532 37056 16584
rect 30380 16464 30432 16516
rect 31668 16464 31720 16516
rect 31760 16507 31812 16516
rect 31760 16473 31769 16507
rect 31769 16473 31803 16507
rect 31803 16473 31812 16507
rect 31760 16464 31812 16473
rect 27436 16396 27488 16448
rect 29184 16439 29236 16448
rect 29184 16405 29193 16439
rect 29193 16405 29227 16439
rect 29227 16405 29236 16439
rect 29184 16396 29236 16405
rect 29736 16439 29788 16448
rect 29736 16405 29745 16439
rect 29745 16405 29779 16439
rect 29779 16405 29788 16439
rect 29736 16396 29788 16405
rect 30196 16396 30248 16448
rect 30288 16396 30340 16448
rect 34152 16464 34204 16516
rect 34244 16396 34296 16448
rect 34980 16396 35032 16448
rect 36636 16439 36688 16448
rect 36636 16405 36645 16439
rect 36645 16405 36679 16439
rect 36679 16405 36688 16439
rect 36636 16396 36688 16405
rect 36912 16464 36964 16516
rect 40592 16600 40644 16652
rect 37188 16532 37240 16584
rect 37464 16532 37516 16584
rect 37740 16575 37792 16584
rect 37740 16541 37749 16575
rect 37749 16541 37783 16575
rect 37783 16541 37792 16575
rect 37740 16532 37792 16541
rect 38476 16464 38528 16516
rect 40316 16532 40368 16584
rect 41328 16532 41380 16584
rect 49148 16532 49200 16584
rect 40684 16507 40736 16516
rect 40684 16473 40693 16507
rect 40693 16473 40727 16507
rect 40727 16473 40736 16507
rect 40684 16464 40736 16473
rect 39672 16396 39724 16448
rect 42156 16396 42208 16448
rect 49240 16439 49292 16448
rect 49240 16405 49249 16439
rect 49249 16405 49283 16439
rect 49283 16405 49292 16439
rect 49240 16396 49292 16405
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 3976 16192 4028 16244
rect 5908 16192 5960 16244
rect 6368 16192 6420 16244
rect 9128 16192 9180 16244
rect 10140 16235 10192 16244
rect 10140 16201 10149 16235
rect 10149 16201 10183 16235
rect 10183 16201 10192 16235
rect 10140 16192 10192 16201
rect 4068 16124 4120 16176
rect 8944 16124 8996 16176
rect 9864 16167 9916 16176
rect 9864 16133 9873 16167
rect 9873 16133 9907 16167
rect 9907 16133 9916 16167
rect 9864 16124 9916 16133
rect 11428 16192 11480 16244
rect 11612 16192 11664 16244
rect 14464 16192 14516 16244
rect 15660 16192 15712 16244
rect 16028 16235 16080 16244
rect 16028 16201 16037 16235
rect 16037 16201 16071 16235
rect 16071 16201 16080 16235
rect 16028 16192 16080 16201
rect 17224 16192 17276 16244
rect 19248 16192 19300 16244
rect 20076 16192 20128 16244
rect 22836 16192 22888 16244
rect 25044 16192 25096 16244
rect 10600 16167 10652 16176
rect 10600 16133 10609 16167
rect 10609 16133 10643 16167
rect 10643 16133 10652 16167
rect 10600 16124 10652 16133
rect 10968 16124 11020 16176
rect 12072 16124 12124 16176
rect 12992 16124 13044 16176
rect 15016 16124 15068 16176
rect 20904 16124 20956 16176
rect 21548 16167 21600 16176
rect 21548 16133 21557 16167
rect 21557 16133 21591 16167
rect 21591 16133 21600 16167
rect 21548 16124 21600 16133
rect 23664 16124 23716 16176
rect 5448 16056 5500 16108
rect 8300 16056 8352 16108
rect 11980 16056 12032 16108
rect 12348 16099 12400 16108
rect 12348 16065 12357 16099
rect 12357 16065 12391 16099
rect 12391 16065 12400 16099
rect 12348 16056 12400 16065
rect 1308 15988 1360 16040
rect 4344 15988 4396 16040
rect 8668 16031 8720 16040
rect 8668 15997 8677 16031
rect 8677 15997 8711 16031
rect 8711 15997 8720 16031
rect 8668 15988 8720 15997
rect 9680 15988 9732 16040
rect 9864 15920 9916 15972
rect 10048 15988 10100 16040
rect 12624 16031 12676 16040
rect 12624 15997 12633 16031
rect 12633 15997 12667 16031
rect 12667 15997 12676 16031
rect 12624 15988 12676 15997
rect 13728 16031 13780 16040
rect 13728 15997 13737 16031
rect 13737 15997 13771 16031
rect 13771 15997 13780 16031
rect 13728 15988 13780 15997
rect 14832 16099 14884 16108
rect 14832 16065 14841 16099
rect 14841 16065 14875 16099
rect 14875 16065 14884 16099
rect 14832 16056 14884 16065
rect 15936 16099 15988 16108
rect 15936 16065 15945 16099
rect 15945 16065 15979 16099
rect 15979 16065 15988 16099
rect 15936 16056 15988 16065
rect 14004 15988 14056 16040
rect 16304 15988 16356 16040
rect 17684 16099 17736 16108
rect 17684 16065 17693 16099
rect 17693 16065 17727 16099
rect 17727 16065 17736 16099
rect 17684 16056 17736 16065
rect 18604 16056 18656 16108
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 24768 16124 24820 16176
rect 25872 16192 25924 16244
rect 26424 16192 26476 16244
rect 26608 16235 26660 16244
rect 26608 16201 26617 16235
rect 26617 16201 26651 16235
rect 26651 16201 26660 16235
rect 26608 16192 26660 16201
rect 27344 16192 27396 16244
rect 27528 16192 27580 16244
rect 27160 16124 27212 16176
rect 28908 16124 28960 16176
rect 29276 16192 29328 16244
rect 30380 16192 30432 16244
rect 30656 16192 30708 16244
rect 31944 16192 31996 16244
rect 32680 16192 32732 16244
rect 33968 16235 34020 16244
rect 33968 16201 33977 16235
rect 33977 16201 34011 16235
rect 34011 16201 34020 16235
rect 33968 16192 34020 16201
rect 34980 16192 35032 16244
rect 35348 16192 35400 16244
rect 36912 16192 36964 16244
rect 37372 16192 37424 16244
rect 38660 16192 38712 16244
rect 41604 16235 41656 16244
rect 41604 16201 41613 16235
rect 41613 16201 41647 16235
rect 41647 16201 41656 16235
rect 41604 16192 41656 16201
rect 30288 16124 30340 16176
rect 30932 16167 30984 16176
rect 30932 16133 30941 16167
rect 30941 16133 30975 16167
rect 30975 16133 30984 16167
rect 30932 16124 30984 16133
rect 34796 16167 34848 16176
rect 34796 16133 34805 16167
rect 34805 16133 34839 16167
rect 34839 16133 34848 16167
rect 34796 16124 34848 16133
rect 36728 16124 36780 16176
rect 38568 16124 38620 16176
rect 38752 16124 38804 16176
rect 48964 16124 49016 16176
rect 27436 16056 27488 16108
rect 28356 16099 28408 16108
rect 28356 16065 28365 16099
rect 28365 16065 28399 16099
rect 28399 16065 28408 16099
rect 28356 16056 28408 16065
rect 30196 16056 30248 16108
rect 6276 15852 6328 15904
rect 9496 15852 9548 15904
rect 11152 15895 11204 15904
rect 11152 15861 11161 15895
rect 11161 15861 11195 15895
rect 11195 15861 11204 15895
rect 11152 15852 11204 15861
rect 12072 15852 12124 15904
rect 14832 15852 14884 15904
rect 15844 15852 15896 15904
rect 18604 15920 18656 15972
rect 17224 15852 17276 15904
rect 17868 15852 17920 15904
rect 17960 15852 18012 15904
rect 18512 15852 18564 15904
rect 19340 15988 19392 16040
rect 23572 16031 23624 16040
rect 23572 15997 23581 16031
rect 23581 15997 23615 16031
rect 23615 15997 23624 16031
rect 23572 15988 23624 15997
rect 26424 15988 26476 16040
rect 20996 15852 21048 15904
rect 22284 15852 22336 15904
rect 22560 15852 22612 15904
rect 22652 15895 22704 15904
rect 22652 15861 22661 15895
rect 22661 15861 22695 15895
rect 22695 15861 22704 15895
rect 22652 15852 22704 15861
rect 23940 15852 23992 15904
rect 24400 15852 24452 15904
rect 27344 15920 27396 15972
rect 28724 15988 28776 16040
rect 30840 15988 30892 16040
rect 30380 15920 30432 15972
rect 31116 15920 31168 15972
rect 33876 16099 33928 16108
rect 33876 16065 33885 16099
rect 33885 16065 33919 16099
rect 33919 16065 33928 16099
rect 33876 16056 33928 16065
rect 36360 16056 36412 16108
rect 37188 16056 37240 16108
rect 39764 16056 39816 16108
rect 42248 16056 42300 16108
rect 49056 16099 49108 16108
rect 32956 16031 33008 16040
rect 32956 15997 32965 16031
rect 32965 15997 32999 16031
rect 32999 15997 33008 16031
rect 32956 15988 33008 15997
rect 34152 16031 34204 16040
rect 34152 15997 34161 16031
rect 34161 15997 34195 16031
rect 34195 15997 34204 16031
rect 34152 15988 34204 15997
rect 34888 15988 34940 16040
rect 35348 16031 35400 16040
rect 35348 15997 35357 16031
rect 35357 15997 35391 16031
rect 35391 15997 35400 16031
rect 35348 15988 35400 15997
rect 35440 15988 35492 16040
rect 37004 15988 37056 16040
rect 37464 15988 37516 16040
rect 41052 16031 41104 16040
rect 41052 15997 41061 16031
rect 41061 15997 41095 16031
rect 41095 15997 41104 16031
rect 41052 15988 41104 15997
rect 33784 15920 33836 15972
rect 33416 15852 33468 15904
rect 33508 15895 33560 15904
rect 33508 15861 33517 15895
rect 33517 15861 33551 15895
rect 33551 15861 33560 15895
rect 33508 15852 33560 15861
rect 36360 15920 36412 15972
rect 37648 15920 37700 15972
rect 39856 15920 39908 15972
rect 49056 16065 49065 16099
rect 49065 16065 49099 16099
rect 49099 16065 49108 16099
rect 49056 16056 49108 16065
rect 38568 15852 38620 15904
rect 39580 15852 39632 15904
rect 42340 15852 42392 15904
rect 48596 15852 48648 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 3516 15648 3568 15700
rect 11244 15648 11296 15700
rect 11520 15648 11572 15700
rect 14556 15648 14608 15700
rect 15752 15648 15804 15700
rect 9772 15580 9824 15632
rect 10140 15580 10192 15632
rect 12348 15580 12400 15632
rect 1308 15512 1360 15564
rect 10784 15555 10836 15564
rect 10784 15521 10793 15555
rect 10793 15521 10827 15555
rect 10827 15521 10836 15555
rect 10784 15512 10836 15521
rect 9680 15444 9732 15496
rect 10692 15444 10744 15496
rect 12624 15512 12676 15564
rect 15108 15512 15160 15564
rect 15844 15555 15896 15564
rect 15844 15521 15853 15555
rect 15853 15521 15887 15555
rect 15887 15521 15896 15555
rect 15844 15512 15896 15521
rect 17960 15580 18012 15632
rect 17500 15555 17552 15564
rect 17500 15521 17509 15555
rect 17509 15521 17543 15555
rect 17543 15521 17552 15555
rect 17500 15512 17552 15521
rect 18420 15648 18472 15700
rect 18604 15648 18656 15700
rect 20812 15648 20864 15700
rect 22652 15648 22704 15700
rect 26148 15648 26200 15700
rect 21916 15580 21968 15632
rect 22008 15580 22060 15632
rect 22376 15623 22428 15632
rect 22376 15589 22385 15623
rect 22385 15589 22419 15623
rect 22419 15589 22428 15623
rect 22376 15580 22428 15589
rect 22560 15580 22612 15632
rect 24584 15580 24636 15632
rect 19340 15555 19392 15564
rect 19340 15521 19349 15555
rect 19349 15521 19383 15555
rect 19383 15521 19392 15555
rect 19340 15512 19392 15521
rect 20352 15555 20404 15564
rect 20352 15521 20361 15555
rect 20361 15521 20395 15555
rect 20395 15521 20404 15555
rect 20352 15512 20404 15521
rect 20904 15555 20956 15564
rect 20904 15521 20913 15555
rect 20913 15521 20947 15555
rect 20947 15521 20956 15555
rect 20904 15512 20956 15521
rect 21732 15555 21784 15564
rect 21732 15521 21741 15555
rect 21741 15521 21775 15555
rect 21775 15521 21784 15555
rect 21732 15512 21784 15521
rect 13728 15444 13780 15496
rect 14280 15487 14332 15496
rect 14280 15453 14289 15487
rect 14289 15453 14323 15487
rect 14323 15453 14332 15487
rect 14280 15444 14332 15453
rect 17132 15444 17184 15496
rect 17684 15444 17736 15496
rect 18972 15444 19024 15496
rect 22560 15487 22612 15496
rect 22560 15453 22569 15487
rect 22569 15453 22603 15487
rect 22603 15453 22612 15487
rect 22560 15444 22612 15453
rect 6920 15376 6972 15428
rect 7656 15376 7708 15428
rect 9404 15419 9456 15428
rect 9404 15385 9413 15419
rect 9413 15385 9447 15419
rect 9447 15385 9456 15419
rect 9404 15376 9456 15385
rect 11152 15376 11204 15428
rect 11520 15376 11572 15428
rect 15568 15376 15620 15428
rect 18420 15376 18472 15428
rect 19248 15376 19300 15428
rect 6644 15351 6696 15360
rect 6644 15317 6653 15351
rect 6653 15317 6687 15351
rect 6687 15317 6696 15351
rect 6644 15308 6696 15317
rect 8668 15351 8720 15360
rect 8668 15317 8677 15351
rect 8677 15317 8711 15351
rect 8711 15317 8720 15351
rect 9036 15351 9088 15360
rect 8668 15308 8720 15317
rect 9036 15317 9045 15351
rect 9045 15317 9079 15351
rect 9079 15317 9088 15351
rect 9036 15308 9088 15317
rect 9496 15351 9548 15360
rect 9496 15317 9505 15351
rect 9505 15317 9539 15351
rect 9539 15317 9548 15351
rect 9496 15308 9548 15317
rect 10232 15308 10284 15360
rect 12072 15308 12124 15360
rect 14556 15308 14608 15360
rect 16856 15308 16908 15360
rect 17592 15308 17644 15360
rect 19892 15308 19944 15360
rect 20536 15308 20588 15360
rect 21272 15308 21324 15360
rect 21548 15351 21600 15360
rect 21548 15317 21557 15351
rect 21557 15317 21591 15351
rect 21591 15317 21600 15351
rect 21548 15308 21600 15317
rect 21640 15351 21692 15360
rect 21640 15317 21649 15351
rect 21649 15317 21683 15351
rect 21683 15317 21692 15351
rect 21640 15308 21692 15317
rect 23388 15512 23440 15564
rect 24768 15580 24820 15632
rect 23848 15444 23900 15496
rect 25136 15555 25188 15564
rect 25136 15521 25145 15555
rect 25145 15521 25179 15555
rect 25179 15521 25188 15555
rect 25136 15512 25188 15521
rect 26792 15648 26844 15700
rect 26976 15691 27028 15700
rect 26976 15657 26985 15691
rect 26985 15657 27019 15691
rect 27019 15657 27028 15691
rect 26976 15648 27028 15657
rect 27528 15648 27580 15700
rect 31852 15648 31904 15700
rect 34152 15648 34204 15700
rect 34244 15648 34296 15700
rect 27068 15580 27120 15632
rect 27436 15580 27488 15632
rect 28632 15580 28684 15632
rect 26424 15555 26476 15564
rect 26424 15521 26433 15555
rect 26433 15521 26467 15555
rect 26467 15521 26476 15555
rect 26424 15512 26476 15521
rect 26608 15512 26660 15564
rect 28540 15512 28592 15564
rect 28908 15580 28960 15632
rect 32312 15580 32364 15632
rect 33048 15580 33100 15632
rect 29184 15512 29236 15564
rect 32864 15512 32916 15564
rect 34336 15512 34388 15564
rect 27712 15444 27764 15496
rect 28724 15444 28776 15496
rect 30288 15444 30340 15496
rect 32036 15444 32088 15496
rect 32772 15444 32824 15496
rect 37648 15648 37700 15700
rect 42156 15648 42208 15700
rect 48964 15648 49016 15700
rect 37188 15623 37240 15632
rect 35164 15555 35216 15564
rect 35164 15521 35173 15555
rect 35173 15521 35207 15555
rect 35207 15521 35216 15555
rect 35164 15512 35216 15521
rect 34888 15487 34940 15496
rect 34888 15453 34897 15487
rect 34897 15453 34931 15487
rect 34931 15453 34940 15487
rect 34888 15444 34940 15453
rect 36176 15444 36228 15496
rect 37188 15589 37197 15623
rect 37197 15589 37231 15623
rect 37231 15589 37240 15623
rect 37188 15580 37240 15589
rect 39488 15623 39540 15632
rect 39488 15589 39497 15623
rect 39497 15589 39531 15623
rect 39531 15589 39540 15623
rect 39488 15580 39540 15589
rect 41328 15580 41380 15632
rect 25412 15308 25464 15360
rect 25872 15351 25924 15360
rect 25872 15317 25881 15351
rect 25881 15317 25915 15351
rect 25915 15317 25924 15351
rect 25872 15308 25924 15317
rect 26240 15351 26292 15360
rect 26240 15317 26249 15351
rect 26249 15317 26283 15351
rect 26283 15317 26292 15351
rect 26240 15308 26292 15317
rect 26700 15376 26752 15428
rect 31024 15376 31076 15428
rect 34244 15376 34296 15428
rect 26792 15308 26844 15360
rect 26976 15308 27028 15360
rect 27436 15351 27488 15360
rect 27436 15317 27445 15351
rect 27445 15317 27479 15351
rect 27479 15317 27488 15351
rect 27436 15308 27488 15317
rect 31116 15308 31168 15360
rect 32772 15308 32824 15360
rect 33048 15351 33100 15360
rect 33048 15317 33057 15351
rect 33057 15317 33091 15351
rect 33091 15317 33100 15351
rect 33048 15308 33100 15317
rect 35256 15308 35308 15360
rect 36084 15308 36136 15360
rect 37464 15444 37516 15496
rect 42340 15512 42392 15564
rect 42248 15487 42300 15496
rect 42248 15453 42257 15487
rect 42257 15453 42291 15487
rect 42291 15453 42300 15487
rect 42248 15444 42300 15453
rect 49332 15487 49384 15496
rect 49332 15453 49341 15487
rect 49341 15453 49375 15487
rect 49375 15453 49384 15487
rect 49332 15444 49384 15453
rect 38476 15376 38528 15428
rect 36912 15351 36964 15360
rect 36912 15317 36921 15351
rect 36921 15317 36955 15351
rect 36955 15317 36964 15351
rect 36912 15308 36964 15317
rect 38384 15308 38436 15360
rect 40316 15376 40368 15428
rect 41604 15376 41656 15428
rect 40040 15308 40092 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 9864 15147 9916 15156
rect 9864 15113 9873 15147
rect 9873 15113 9907 15147
rect 9907 15113 9916 15147
rect 9864 15104 9916 15113
rect 10324 15104 10376 15156
rect 12072 15104 12124 15156
rect 12808 15104 12860 15156
rect 14832 15104 14884 15156
rect 14924 15104 14976 15156
rect 8852 15036 8904 15088
rect 11980 15036 12032 15088
rect 12532 15036 12584 15088
rect 13912 15036 13964 15088
rect 6644 14968 6696 15020
rect 10968 15011 11020 15020
rect 10968 14977 10977 15011
rect 10977 14977 11011 15011
rect 11011 14977 11020 15011
rect 10968 14968 11020 14977
rect 11152 14968 11204 15020
rect 12716 14968 12768 15020
rect 1308 14900 1360 14952
rect 12256 14900 12308 14952
rect 12532 14900 12584 14952
rect 16764 15104 16816 15156
rect 17132 15104 17184 15156
rect 15292 15036 15344 15088
rect 17316 15079 17368 15088
rect 17316 15045 17325 15079
rect 17325 15045 17359 15079
rect 17359 15045 17368 15079
rect 17316 15036 17368 15045
rect 18696 15147 18748 15156
rect 18696 15113 18705 15147
rect 18705 15113 18739 15147
rect 18739 15113 18748 15147
rect 18696 15104 18748 15113
rect 19800 15104 19852 15156
rect 20720 15147 20772 15156
rect 20720 15113 20729 15147
rect 20729 15113 20763 15147
rect 20763 15113 20772 15147
rect 20720 15104 20772 15113
rect 21180 15104 21232 15156
rect 21640 15104 21692 15156
rect 23480 15104 23532 15156
rect 26056 15104 26108 15156
rect 27068 15147 27120 15156
rect 27068 15113 27077 15147
rect 27077 15113 27111 15147
rect 27111 15113 27120 15147
rect 27068 15104 27120 15113
rect 27252 15104 27304 15156
rect 21732 15036 21784 15088
rect 19800 14968 19852 15020
rect 20536 14968 20588 15020
rect 21456 14968 21508 15020
rect 17132 14900 17184 14952
rect 10416 14764 10468 14816
rect 10692 14764 10744 14816
rect 11060 14807 11112 14816
rect 11060 14773 11069 14807
rect 11069 14773 11103 14807
rect 11103 14773 11112 14807
rect 11060 14764 11112 14773
rect 14280 14832 14332 14884
rect 17868 14900 17920 14952
rect 18788 14943 18840 14952
rect 18788 14909 18797 14943
rect 18797 14909 18831 14943
rect 18831 14909 18840 14943
rect 18788 14900 18840 14909
rect 18880 14943 18932 14952
rect 18880 14909 18889 14943
rect 18889 14909 18923 14943
rect 18923 14909 18932 14943
rect 18880 14900 18932 14909
rect 19984 14943 20036 14952
rect 19984 14909 19993 14943
rect 19993 14909 20027 14943
rect 20027 14909 20036 14943
rect 19984 14900 20036 14909
rect 20076 14943 20128 14952
rect 20076 14909 20085 14943
rect 20085 14909 20119 14943
rect 20119 14909 20128 14943
rect 20076 14900 20128 14909
rect 20904 14900 20956 14952
rect 21272 14943 21324 14952
rect 21272 14909 21281 14943
rect 21281 14909 21315 14943
rect 21315 14909 21324 14943
rect 21272 14900 21324 14909
rect 25780 15036 25832 15088
rect 24492 15011 24544 15020
rect 24492 14977 24501 15011
rect 24501 14977 24535 15011
rect 24535 14977 24544 15011
rect 24492 14968 24544 14977
rect 25688 14968 25740 15020
rect 27252 15011 27304 15020
rect 18420 14832 18472 14884
rect 13452 14764 13504 14816
rect 15292 14807 15344 14816
rect 15292 14773 15301 14807
rect 15301 14773 15335 14807
rect 15335 14773 15344 14807
rect 15292 14764 15344 14773
rect 16488 14764 16540 14816
rect 16856 14764 16908 14816
rect 17316 14764 17368 14816
rect 17500 14764 17552 14816
rect 20444 14764 20496 14816
rect 21456 14764 21508 14816
rect 24584 14943 24636 14952
rect 24584 14909 24593 14943
rect 24593 14909 24627 14943
rect 24627 14909 24636 14943
rect 24584 14900 24636 14909
rect 24124 14832 24176 14884
rect 24768 14900 24820 14952
rect 27252 14977 27261 15011
rect 27261 14977 27295 15011
rect 27295 14977 27304 15011
rect 27252 14968 27304 14977
rect 28724 15104 28776 15156
rect 29092 15104 29144 15156
rect 28356 15036 28408 15088
rect 28448 15036 28500 15088
rect 29828 15036 29880 15088
rect 23756 14764 23808 14816
rect 24492 14764 24544 14816
rect 25136 14764 25188 14816
rect 25412 14764 25464 14816
rect 25596 14764 25648 14816
rect 26240 14764 26292 14816
rect 28908 14900 28960 14952
rect 27160 14832 27212 14884
rect 28080 14832 28132 14884
rect 26792 14764 26844 14816
rect 28816 14764 28868 14816
rect 30104 14900 30156 14952
rect 30104 14764 30156 14816
rect 30748 14943 30800 14952
rect 30748 14909 30757 14943
rect 30757 14909 30791 14943
rect 30791 14909 30800 14943
rect 30748 14900 30800 14909
rect 33784 15104 33836 15156
rect 34520 15104 34572 15156
rect 34704 15104 34756 15156
rect 36268 15147 36320 15156
rect 36268 15113 36277 15147
rect 36277 15113 36311 15147
rect 36311 15113 36320 15147
rect 36268 15104 36320 15113
rect 40132 15104 40184 15156
rect 41604 15104 41656 15156
rect 38476 15036 38528 15088
rect 48412 15036 48464 15088
rect 32680 15011 32732 15020
rect 32680 14977 32689 15011
rect 32689 14977 32723 15011
rect 32723 14977 32732 15011
rect 32680 14968 32732 14977
rect 31024 14900 31076 14952
rect 32588 14900 32640 14952
rect 33324 14900 33376 14952
rect 30932 14832 30984 14884
rect 34152 14943 34204 14952
rect 34152 14909 34161 14943
rect 34161 14909 34195 14943
rect 34195 14909 34204 14943
rect 34152 14900 34204 14909
rect 35992 14968 36044 15020
rect 39856 14968 39908 15020
rect 40316 14968 40368 15020
rect 42064 14968 42116 15020
rect 49056 15011 49108 15020
rect 49056 14977 49065 15011
rect 49065 14977 49099 15011
rect 49099 14977 49108 15011
rect 49056 14968 49108 14977
rect 33232 14764 33284 14816
rect 35072 14764 35124 14816
rect 35532 14900 35584 14952
rect 36636 14900 36688 14952
rect 37464 14943 37516 14952
rect 37464 14909 37473 14943
rect 37473 14909 37507 14943
rect 37507 14909 37516 14943
rect 37464 14900 37516 14909
rect 40040 14900 40092 14952
rect 35808 14832 35860 14884
rect 37372 14832 37424 14884
rect 39948 14832 40000 14884
rect 48320 14832 48372 14884
rect 36268 14764 36320 14816
rect 37096 14764 37148 14816
rect 38200 14764 38252 14816
rect 38292 14764 38344 14816
rect 41144 14764 41196 14816
rect 45836 14764 45888 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 9680 14560 9732 14612
rect 10508 14560 10560 14612
rect 16028 14560 16080 14612
rect 16396 14560 16448 14612
rect 16948 14560 17000 14612
rect 18696 14560 18748 14612
rect 21732 14560 21784 14612
rect 23480 14560 23532 14612
rect 23756 14603 23808 14612
rect 23756 14569 23765 14603
rect 23765 14569 23799 14603
rect 23799 14569 23808 14603
rect 23756 14560 23808 14569
rect 24584 14560 24636 14612
rect 29092 14560 29144 14612
rect 30840 14560 30892 14612
rect 33876 14560 33928 14612
rect 33968 14560 34020 14612
rect 37740 14560 37792 14612
rect 41604 14560 41656 14612
rect 5448 14492 5500 14544
rect 11060 14492 11112 14544
rect 12348 14492 12400 14544
rect 1308 14424 1360 14476
rect 13360 14424 13412 14476
rect 13544 14467 13596 14476
rect 13544 14433 13553 14467
rect 13553 14433 13587 14467
rect 13587 14433 13596 14467
rect 13544 14424 13596 14433
rect 13820 14424 13872 14476
rect 9588 14331 9640 14340
rect 9588 14297 9597 14331
rect 9597 14297 9631 14331
rect 9631 14297 9640 14331
rect 9588 14288 9640 14297
rect 10324 14331 10376 14340
rect 10324 14297 10333 14331
rect 10333 14297 10367 14331
rect 10367 14297 10376 14331
rect 10324 14288 10376 14297
rect 11428 14356 11480 14408
rect 11980 14356 12032 14408
rect 16212 14467 16264 14476
rect 16212 14433 16221 14467
rect 16221 14433 16255 14467
rect 16255 14433 16264 14467
rect 16212 14424 16264 14433
rect 18420 14492 18472 14544
rect 19800 14492 19852 14544
rect 16672 14424 16724 14476
rect 17040 14424 17092 14476
rect 17408 14467 17460 14476
rect 17408 14433 17417 14467
rect 17417 14433 17451 14467
rect 17451 14433 17460 14467
rect 17408 14424 17460 14433
rect 18604 14467 18656 14476
rect 16948 14356 17000 14408
rect 17224 14399 17276 14408
rect 17224 14365 17233 14399
rect 17233 14365 17267 14399
rect 17267 14365 17276 14399
rect 17224 14356 17276 14365
rect 17316 14356 17368 14408
rect 18604 14433 18613 14467
rect 18613 14433 18647 14467
rect 18647 14433 18656 14467
rect 18604 14424 18656 14433
rect 18696 14467 18748 14476
rect 18696 14433 18705 14467
rect 18705 14433 18739 14467
rect 18739 14433 18748 14467
rect 18696 14424 18748 14433
rect 19064 14424 19116 14476
rect 21088 14467 21140 14476
rect 21088 14433 21097 14467
rect 21097 14433 21131 14467
rect 21131 14433 21140 14467
rect 21088 14424 21140 14433
rect 22652 14492 22704 14544
rect 25596 14492 25648 14544
rect 21732 14424 21784 14476
rect 22744 14424 22796 14476
rect 24400 14424 24452 14476
rect 24676 14424 24728 14476
rect 24860 14424 24912 14476
rect 27160 14424 27212 14476
rect 17684 14356 17736 14408
rect 20352 14356 20404 14408
rect 20996 14356 21048 14408
rect 23940 14399 23992 14408
rect 12256 14331 12308 14340
rect 12256 14297 12265 14331
rect 12265 14297 12299 14331
rect 12299 14297 12308 14331
rect 12256 14288 12308 14297
rect 11244 14263 11296 14272
rect 11244 14229 11253 14263
rect 11253 14229 11287 14263
rect 11287 14229 11296 14263
rect 11244 14220 11296 14229
rect 11336 14220 11388 14272
rect 13912 14220 13964 14272
rect 14188 14220 14240 14272
rect 14832 14331 14884 14340
rect 14832 14297 14841 14331
rect 14841 14297 14875 14331
rect 14875 14297 14884 14331
rect 14832 14288 14884 14297
rect 14924 14263 14976 14272
rect 14924 14229 14933 14263
rect 14933 14229 14967 14263
rect 14967 14229 14976 14263
rect 14924 14220 14976 14229
rect 17868 14288 17920 14340
rect 16028 14263 16080 14272
rect 16028 14229 16037 14263
rect 16037 14229 16071 14263
rect 16071 14229 16080 14263
rect 16028 14220 16080 14229
rect 16120 14263 16172 14272
rect 16120 14229 16129 14263
rect 16129 14229 16163 14263
rect 16163 14229 16172 14263
rect 16120 14220 16172 14229
rect 16212 14220 16264 14272
rect 17132 14220 17184 14272
rect 17408 14220 17460 14272
rect 21916 14288 21968 14340
rect 23020 14288 23072 14340
rect 23940 14365 23949 14399
rect 23949 14365 23983 14399
rect 23983 14365 23992 14399
rect 23940 14356 23992 14365
rect 24032 14356 24084 14408
rect 27068 14356 27120 14408
rect 28724 14492 28776 14544
rect 28540 14467 28592 14476
rect 28540 14433 28549 14467
rect 28549 14433 28583 14467
rect 28583 14433 28592 14467
rect 32036 14492 32088 14544
rect 32864 14492 32916 14544
rect 34796 14492 34848 14544
rect 36544 14492 36596 14544
rect 28540 14424 28592 14433
rect 30380 14424 30432 14476
rect 30748 14424 30800 14476
rect 31668 14424 31720 14476
rect 32956 14424 33008 14476
rect 33600 14424 33652 14476
rect 34152 14424 34204 14476
rect 34888 14467 34940 14476
rect 34888 14433 34897 14467
rect 34897 14433 34931 14467
rect 34931 14433 34940 14467
rect 34888 14424 34940 14433
rect 37464 14424 37516 14476
rect 37832 14424 37884 14476
rect 39856 14492 39908 14544
rect 45560 14492 45612 14544
rect 48596 14492 48648 14544
rect 38936 14424 38988 14476
rect 39948 14424 40000 14476
rect 23480 14288 23532 14340
rect 26240 14288 26292 14340
rect 31024 14356 31076 14408
rect 31116 14356 31168 14408
rect 31484 14356 31536 14408
rect 19156 14220 19208 14272
rect 19708 14220 19760 14272
rect 20076 14263 20128 14272
rect 20076 14229 20085 14263
rect 20085 14229 20119 14263
rect 20119 14229 20128 14263
rect 20076 14220 20128 14229
rect 20904 14220 20956 14272
rect 21732 14220 21784 14272
rect 23296 14220 23348 14272
rect 23848 14220 23900 14272
rect 24216 14220 24268 14272
rect 25504 14220 25556 14272
rect 28632 14220 28684 14272
rect 29276 14263 29328 14272
rect 29276 14229 29285 14263
rect 29285 14229 29319 14263
rect 29319 14229 29328 14263
rect 29276 14220 29328 14229
rect 29460 14220 29512 14272
rect 30196 14263 30248 14272
rect 30196 14229 30205 14263
rect 30205 14229 30239 14263
rect 30239 14229 30248 14263
rect 30196 14220 30248 14229
rect 30472 14220 30524 14272
rect 32036 14220 32088 14272
rect 33140 14288 33192 14340
rect 33416 14356 33468 14408
rect 38476 14356 38528 14408
rect 39488 14399 39540 14408
rect 39488 14365 39497 14399
rect 39497 14365 39531 14399
rect 39531 14365 39540 14399
rect 39488 14356 39540 14365
rect 41144 14399 41196 14408
rect 41144 14365 41153 14399
rect 41153 14365 41187 14399
rect 41187 14365 41196 14399
rect 41144 14356 41196 14365
rect 49056 14399 49108 14408
rect 49056 14365 49065 14399
rect 49065 14365 49099 14399
rect 49099 14365 49108 14399
rect 49056 14356 49108 14365
rect 35164 14331 35216 14340
rect 35164 14297 35173 14331
rect 35173 14297 35207 14331
rect 35207 14297 35216 14331
rect 35164 14288 35216 14297
rect 35440 14288 35492 14340
rect 36176 14288 36228 14340
rect 32588 14220 32640 14272
rect 36084 14220 36136 14272
rect 38936 14220 38988 14272
rect 39304 14263 39356 14272
rect 39304 14229 39313 14263
rect 39313 14229 39347 14263
rect 39347 14229 39356 14263
rect 39304 14220 39356 14229
rect 40684 14263 40736 14272
rect 40684 14229 40693 14263
rect 40693 14229 40727 14263
rect 40727 14229 40736 14263
rect 40684 14220 40736 14229
rect 41420 14220 41472 14272
rect 44180 14220 44232 14272
rect 48320 14220 48372 14272
rect 49240 14263 49292 14272
rect 49240 14229 49249 14263
rect 49249 14229 49283 14263
rect 49283 14229 49292 14263
rect 49240 14220 49292 14229
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 9772 14016 9824 14068
rect 9864 14059 9916 14068
rect 9864 14025 9873 14059
rect 9873 14025 9907 14059
rect 9907 14025 9916 14059
rect 9864 14016 9916 14025
rect 11244 13948 11296 14000
rect 11520 14016 11572 14068
rect 15108 14059 15160 14068
rect 15108 14025 15117 14059
rect 15117 14025 15151 14059
rect 15151 14025 15160 14059
rect 15108 14016 15160 14025
rect 12532 13948 12584 14000
rect 13360 13948 13412 14000
rect 13912 13948 13964 14000
rect 14188 13948 14240 14000
rect 16120 14016 16172 14068
rect 17408 14016 17460 14068
rect 17776 14016 17828 14068
rect 20720 14016 20772 14068
rect 20996 14016 21048 14068
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 4068 13880 4120 13932
rect 10232 13880 10284 13932
rect 940 13812 992 13864
rect 7380 13812 7432 13864
rect 9588 13855 9640 13864
rect 9588 13821 9597 13855
rect 9597 13821 9631 13855
rect 9631 13821 9640 13855
rect 9588 13812 9640 13821
rect 10324 13812 10376 13864
rect 12716 13880 12768 13932
rect 12348 13744 12400 13796
rect 12256 13676 12308 13728
rect 12624 13812 12676 13864
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 17684 13948 17736 14000
rect 18512 13948 18564 14000
rect 17132 13880 17184 13932
rect 17316 13880 17368 13932
rect 19524 13880 19576 13932
rect 21088 13880 21140 13932
rect 23296 14016 23348 14068
rect 24032 14016 24084 14068
rect 26424 14016 26476 14068
rect 28448 14016 28500 14068
rect 22284 13991 22336 14000
rect 22284 13957 22293 13991
rect 22293 13957 22327 13991
rect 22327 13957 22336 13991
rect 22284 13948 22336 13957
rect 25228 13948 25280 14000
rect 26792 13948 26844 14000
rect 27068 13948 27120 14000
rect 29276 13948 29328 14000
rect 30380 14016 30432 14068
rect 32772 14016 32824 14068
rect 35072 14016 35124 14068
rect 35624 14016 35676 14068
rect 35716 14059 35768 14068
rect 35716 14025 35725 14059
rect 35725 14025 35759 14059
rect 35759 14025 35768 14059
rect 35716 14016 35768 14025
rect 15936 13812 15988 13864
rect 14648 13744 14700 13796
rect 16396 13744 16448 13796
rect 16488 13744 16540 13796
rect 18144 13812 18196 13864
rect 19616 13812 19668 13864
rect 19708 13855 19760 13864
rect 19708 13821 19717 13855
rect 19717 13821 19751 13855
rect 19751 13821 19760 13855
rect 19708 13812 19760 13821
rect 21916 13812 21968 13864
rect 23020 13812 23072 13864
rect 24860 13923 24912 13932
rect 24860 13889 24869 13923
rect 24869 13889 24903 13923
rect 24903 13889 24912 13923
rect 24860 13880 24912 13889
rect 29000 13880 29052 13932
rect 33692 13880 33744 13932
rect 34428 13880 34480 13932
rect 37188 14016 37240 14068
rect 37280 14016 37332 14068
rect 37740 14016 37792 14068
rect 39120 14016 39172 14068
rect 36360 13948 36412 14000
rect 36728 13948 36780 14000
rect 41420 14016 41472 14068
rect 41512 14016 41564 14068
rect 47860 14016 47912 14068
rect 48412 14059 48464 14068
rect 48412 14025 48421 14059
rect 48421 14025 48455 14059
rect 48455 14025 48464 14059
rect 48412 14016 48464 14025
rect 48504 14016 48556 14068
rect 39304 13948 39356 14000
rect 49148 13991 49200 14000
rect 49148 13957 49157 13991
rect 49157 13957 49191 13991
rect 49191 13957 49200 13991
rect 49148 13948 49200 13957
rect 23480 13812 23532 13864
rect 25136 13855 25188 13864
rect 25136 13821 25145 13855
rect 25145 13821 25179 13855
rect 25179 13821 25188 13855
rect 25136 13812 25188 13821
rect 14004 13676 14056 13728
rect 16304 13676 16356 13728
rect 16948 13719 17000 13728
rect 16948 13685 16957 13719
rect 16957 13685 16991 13719
rect 16991 13685 17000 13719
rect 16948 13676 17000 13685
rect 30840 13812 30892 13864
rect 32220 13812 32272 13864
rect 32588 13855 32640 13864
rect 32588 13821 32597 13855
rect 32597 13821 32631 13855
rect 32631 13821 32640 13855
rect 32588 13812 32640 13821
rect 33140 13812 33192 13864
rect 33600 13812 33652 13864
rect 31852 13744 31904 13796
rect 34060 13855 34112 13864
rect 34060 13821 34069 13855
rect 34069 13821 34103 13855
rect 34103 13821 34112 13855
rect 34060 13812 34112 13821
rect 34520 13812 34572 13864
rect 36544 13880 36596 13932
rect 37740 13880 37792 13932
rect 36084 13744 36136 13796
rect 37096 13812 37148 13864
rect 39212 13880 39264 13932
rect 37924 13855 37976 13864
rect 37924 13821 37933 13855
rect 37933 13821 37967 13855
rect 37967 13821 37976 13855
rect 37924 13812 37976 13821
rect 20076 13676 20128 13728
rect 28540 13676 28592 13728
rect 29368 13676 29420 13728
rect 30288 13676 30340 13728
rect 31300 13676 31352 13728
rect 33968 13676 34020 13728
rect 34980 13676 35032 13728
rect 35072 13676 35124 13728
rect 36176 13676 36228 13728
rect 37188 13676 37240 13728
rect 38292 13812 38344 13864
rect 39856 13923 39908 13932
rect 39856 13889 39865 13923
rect 39865 13889 39899 13923
rect 39899 13889 39908 13923
rect 39856 13880 39908 13889
rect 40868 13923 40920 13932
rect 40868 13889 40877 13923
rect 40877 13889 40911 13923
rect 40911 13889 40920 13923
rect 40868 13880 40920 13889
rect 40960 13923 41012 13932
rect 40960 13889 40969 13923
rect 40969 13889 41003 13923
rect 41003 13889 41012 13923
rect 40960 13880 41012 13889
rect 45836 13923 45888 13932
rect 45836 13889 45845 13923
rect 45845 13889 45879 13923
rect 45879 13889 45888 13923
rect 45836 13880 45888 13889
rect 48228 13880 48280 13932
rect 38200 13744 38252 13796
rect 46572 13812 46624 13864
rect 41144 13744 41196 13796
rect 41052 13676 41104 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 9036 13472 9088 13524
rect 13820 13472 13872 13524
rect 14464 13515 14516 13524
rect 14464 13481 14473 13515
rect 14473 13481 14507 13515
rect 14507 13481 14516 13515
rect 14464 13472 14516 13481
rect 15200 13515 15252 13524
rect 15200 13481 15209 13515
rect 15209 13481 15243 13515
rect 15243 13481 15252 13515
rect 15200 13472 15252 13481
rect 15568 13472 15620 13524
rect 19248 13472 19300 13524
rect 19892 13472 19944 13524
rect 19984 13472 20036 13524
rect 21364 13472 21416 13524
rect 12440 13404 12492 13456
rect 12808 13404 12860 13456
rect 14188 13404 14240 13456
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 2780 13336 2832 13345
rect 9864 13336 9916 13388
rect 11520 13336 11572 13388
rect 12532 13336 12584 13388
rect 13544 13336 13596 13388
rect 15660 13379 15712 13388
rect 15660 13345 15669 13379
rect 15669 13345 15703 13379
rect 15703 13345 15712 13379
rect 15660 13336 15712 13345
rect 18144 13404 18196 13456
rect 18604 13404 18656 13456
rect 19064 13404 19116 13456
rect 1768 13311 1820 13320
rect 1768 13277 1777 13311
rect 1777 13277 1811 13311
rect 1811 13277 1820 13311
rect 1768 13268 1820 13277
rect 6920 13268 6972 13320
rect 9956 13243 10008 13252
rect 9956 13209 9965 13243
rect 9965 13209 9999 13243
rect 9999 13209 10008 13243
rect 9956 13200 10008 13209
rect 10876 13311 10928 13320
rect 10876 13277 10885 13311
rect 10885 13277 10919 13311
rect 10919 13277 10928 13311
rect 10876 13268 10928 13277
rect 13360 13268 13412 13320
rect 13728 13268 13780 13320
rect 16212 13268 16264 13320
rect 11060 13200 11112 13252
rect 11612 13200 11664 13252
rect 14280 13200 14332 13252
rect 14372 13243 14424 13252
rect 14372 13209 14381 13243
rect 14381 13209 14415 13243
rect 14415 13209 14424 13243
rect 14372 13200 14424 13209
rect 15384 13200 15436 13252
rect 16488 13268 16540 13320
rect 17316 13336 17368 13388
rect 17500 13336 17552 13388
rect 19800 13336 19852 13388
rect 17960 13311 18012 13320
rect 17960 13277 17969 13311
rect 17969 13277 18003 13311
rect 18003 13277 18012 13311
rect 17960 13268 18012 13277
rect 18420 13268 18472 13320
rect 19616 13268 19668 13320
rect 21364 13379 21416 13388
rect 21364 13345 21373 13379
rect 21373 13345 21407 13379
rect 21407 13345 21416 13379
rect 23112 13447 23164 13456
rect 23112 13413 23121 13447
rect 23121 13413 23155 13447
rect 23155 13413 23164 13447
rect 23112 13404 23164 13413
rect 23848 13472 23900 13524
rect 24952 13472 25004 13524
rect 25136 13472 25188 13524
rect 29092 13472 29144 13524
rect 29460 13472 29512 13524
rect 27436 13404 27488 13456
rect 27620 13404 27672 13456
rect 34428 13472 34480 13524
rect 34520 13472 34572 13524
rect 21364 13336 21416 13345
rect 21272 13268 21324 13320
rect 22100 13268 22152 13320
rect 16580 13200 16632 13252
rect 12072 13132 12124 13184
rect 14832 13175 14884 13184
rect 14832 13141 14841 13175
rect 14841 13141 14875 13175
rect 14875 13141 14884 13175
rect 14832 13132 14884 13141
rect 14924 13132 14976 13184
rect 17592 13175 17644 13184
rect 17592 13141 17601 13175
rect 17601 13141 17635 13175
rect 17635 13141 17644 13175
rect 17592 13132 17644 13141
rect 19064 13200 19116 13252
rect 23756 13379 23808 13388
rect 23756 13345 23765 13379
rect 23765 13345 23799 13379
rect 23799 13345 23808 13379
rect 23756 13336 23808 13345
rect 27804 13336 27856 13388
rect 30840 13404 30892 13456
rect 32956 13404 33008 13456
rect 24952 13268 25004 13320
rect 25228 13311 25280 13320
rect 25228 13277 25237 13311
rect 25237 13277 25271 13311
rect 25271 13277 25280 13311
rect 25228 13268 25280 13277
rect 25504 13268 25556 13320
rect 27068 13268 27120 13320
rect 30196 13336 30248 13388
rect 32220 13336 32272 13388
rect 33968 13379 34020 13388
rect 33968 13345 33977 13379
rect 33977 13345 34011 13379
rect 34011 13345 34020 13379
rect 33968 13336 34020 13345
rect 35716 13404 35768 13456
rect 34152 13336 34204 13388
rect 30104 13311 30156 13320
rect 30104 13277 30113 13311
rect 30113 13277 30147 13311
rect 30147 13277 30156 13311
rect 30104 13268 30156 13277
rect 32864 13268 32916 13320
rect 34612 13268 34664 13320
rect 22744 13200 22796 13252
rect 25872 13200 25924 13252
rect 20076 13132 20128 13184
rect 20260 13132 20312 13184
rect 21640 13132 21692 13184
rect 22284 13175 22336 13184
rect 22284 13141 22293 13175
rect 22293 13141 22327 13175
rect 22327 13141 22336 13175
rect 22284 13132 22336 13141
rect 23204 13132 23256 13184
rect 24492 13175 24544 13184
rect 24492 13141 24501 13175
rect 24501 13141 24535 13175
rect 24535 13141 24544 13175
rect 24492 13132 24544 13141
rect 26056 13132 26108 13184
rect 26976 13132 27028 13184
rect 30012 13132 30064 13184
rect 30472 13132 30524 13184
rect 31484 13243 31536 13252
rect 31484 13209 31493 13243
rect 31493 13209 31527 13243
rect 31527 13209 31536 13243
rect 31484 13200 31536 13209
rect 31944 13200 31996 13252
rect 33324 13200 33376 13252
rect 33600 13200 33652 13252
rect 35716 13311 35768 13320
rect 35716 13277 35725 13311
rect 35725 13277 35759 13311
rect 35759 13277 35768 13311
rect 35716 13268 35768 13277
rect 35808 13200 35860 13252
rect 32128 13132 32180 13184
rect 32312 13132 32364 13184
rect 35348 13132 35400 13184
rect 36176 13447 36228 13456
rect 36176 13413 36185 13447
rect 36185 13413 36219 13447
rect 36219 13413 36228 13447
rect 36176 13404 36228 13413
rect 36728 13379 36780 13388
rect 36728 13345 36737 13379
rect 36737 13345 36771 13379
rect 36771 13345 36780 13379
rect 36728 13336 36780 13345
rect 36452 13311 36504 13320
rect 36452 13277 36461 13311
rect 36461 13277 36495 13311
rect 36495 13277 36504 13311
rect 36452 13268 36504 13277
rect 38200 13515 38252 13524
rect 38200 13481 38209 13515
rect 38209 13481 38243 13515
rect 38243 13481 38252 13515
rect 38200 13472 38252 13481
rect 38568 13336 38620 13388
rect 41144 13311 41196 13320
rect 41144 13277 41153 13311
rect 41153 13277 41187 13311
rect 41187 13277 41196 13311
rect 41144 13268 41196 13277
rect 46572 13268 46624 13320
rect 49148 13311 49200 13320
rect 49148 13277 49157 13311
rect 49157 13277 49191 13311
rect 49191 13277 49200 13311
rect 49148 13268 49200 13277
rect 37188 13200 37240 13252
rect 38752 13200 38804 13252
rect 39028 13132 39080 13184
rect 39304 13175 39356 13184
rect 39304 13141 39313 13175
rect 39313 13141 39347 13175
rect 39347 13141 39356 13175
rect 39304 13132 39356 13141
rect 39580 13175 39632 13184
rect 39580 13141 39589 13175
rect 39589 13141 39623 13175
rect 39623 13141 39632 13175
rect 39580 13132 39632 13141
rect 41788 13175 41840 13184
rect 41788 13141 41797 13175
rect 41797 13141 41831 13175
rect 41831 13141 41840 13175
rect 41788 13132 41840 13141
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 5632 12928 5684 12980
rect 9864 12971 9916 12980
rect 9864 12937 9873 12971
rect 9873 12937 9907 12971
rect 9907 12937 9916 12971
rect 9864 12928 9916 12937
rect 10416 12928 10468 12980
rect 11060 12928 11112 12980
rect 1308 12792 1360 12844
rect 11336 12792 11388 12844
rect 12072 12971 12124 12980
rect 12072 12937 12081 12971
rect 12081 12937 12115 12971
rect 12115 12937 12124 12971
rect 12072 12928 12124 12937
rect 12256 12928 12308 12980
rect 15936 12971 15988 12980
rect 15936 12937 15945 12971
rect 15945 12937 15979 12971
rect 15979 12937 15988 12971
rect 15936 12928 15988 12937
rect 16856 12928 16908 12980
rect 19708 12928 19760 12980
rect 22652 12928 22704 12980
rect 23572 12928 23624 12980
rect 23756 12928 23808 12980
rect 27068 12928 27120 12980
rect 27160 12928 27212 12980
rect 29368 12928 29420 12980
rect 12256 12792 12308 12844
rect 1216 12724 1268 12776
rect 9496 12724 9548 12776
rect 10968 12767 11020 12776
rect 10968 12733 10977 12767
rect 10977 12733 11011 12767
rect 11011 12733 11020 12767
rect 10968 12724 11020 12733
rect 12532 12792 12584 12844
rect 13360 12860 13412 12912
rect 14372 12860 14424 12912
rect 16580 12860 16632 12912
rect 17040 12860 17092 12912
rect 12808 12724 12860 12776
rect 16028 12835 16080 12844
rect 16028 12801 16037 12835
rect 16037 12801 16071 12835
rect 16071 12801 16080 12835
rect 16028 12792 16080 12801
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 18236 12792 18288 12844
rect 15292 12724 15344 12776
rect 2780 12656 2832 12708
rect 10048 12656 10100 12708
rect 10416 12631 10468 12640
rect 10416 12597 10425 12631
rect 10425 12597 10459 12631
rect 10459 12597 10468 12631
rect 10416 12588 10468 12597
rect 11428 12588 11480 12640
rect 12808 12631 12860 12640
rect 12808 12597 12817 12631
rect 12817 12597 12851 12631
rect 12851 12597 12860 12631
rect 12808 12588 12860 12597
rect 16488 12724 16540 12776
rect 21180 12860 21232 12912
rect 21548 12860 21600 12912
rect 23848 12860 23900 12912
rect 24124 12860 24176 12912
rect 24216 12903 24268 12912
rect 24216 12869 24225 12903
rect 24225 12869 24259 12903
rect 24259 12869 24268 12903
rect 24216 12860 24268 12869
rect 26792 12903 26844 12912
rect 26792 12869 26801 12903
rect 26801 12869 26835 12903
rect 26835 12869 26844 12903
rect 26792 12860 26844 12869
rect 19524 12835 19576 12844
rect 19524 12801 19533 12835
rect 19533 12801 19567 12835
rect 19567 12801 19576 12835
rect 19524 12792 19576 12801
rect 21916 12792 21968 12844
rect 22376 12792 22428 12844
rect 22836 12792 22888 12844
rect 23480 12792 23532 12844
rect 27712 12860 27764 12912
rect 28172 12860 28224 12912
rect 29000 12860 29052 12912
rect 29736 12860 29788 12912
rect 30288 12860 30340 12912
rect 18604 12767 18656 12776
rect 18604 12733 18613 12767
rect 18613 12733 18647 12767
rect 18647 12733 18656 12767
rect 18604 12724 18656 12733
rect 18880 12724 18932 12776
rect 19616 12767 19668 12776
rect 19616 12733 19625 12767
rect 19625 12733 19659 12767
rect 19659 12733 19668 12767
rect 19616 12724 19668 12733
rect 16580 12656 16632 12708
rect 19156 12699 19208 12708
rect 19156 12665 19165 12699
rect 19165 12665 19199 12699
rect 19199 12665 19208 12699
rect 19156 12656 19208 12665
rect 20628 12699 20680 12708
rect 20628 12665 20637 12699
rect 20637 12665 20671 12699
rect 20671 12665 20680 12699
rect 20628 12656 20680 12665
rect 18420 12588 18472 12640
rect 20260 12631 20312 12640
rect 20260 12597 20269 12631
rect 20269 12597 20303 12631
rect 20303 12597 20312 12631
rect 20260 12588 20312 12597
rect 21180 12767 21232 12776
rect 21180 12733 21189 12767
rect 21189 12733 21223 12767
rect 21223 12733 21232 12767
rect 21180 12724 21232 12733
rect 22008 12767 22060 12776
rect 22008 12733 22017 12767
rect 22017 12733 22051 12767
rect 22051 12733 22060 12767
rect 22008 12724 22060 12733
rect 22100 12724 22152 12776
rect 25964 12724 26016 12776
rect 29276 12792 29328 12844
rect 29552 12792 29604 12844
rect 32312 12928 32364 12980
rect 35716 12928 35768 12980
rect 35808 12928 35860 12980
rect 31392 12835 31444 12844
rect 31392 12801 31401 12835
rect 31401 12801 31435 12835
rect 31435 12801 31444 12835
rect 31392 12792 31444 12801
rect 32220 12792 32272 12844
rect 32496 12860 32548 12912
rect 34612 12860 34664 12912
rect 34796 12860 34848 12912
rect 36452 12860 36504 12912
rect 41788 12928 41840 12980
rect 33692 12792 33744 12844
rect 34428 12792 34480 12844
rect 38476 12860 38528 12912
rect 39856 12860 39908 12912
rect 39028 12792 39080 12844
rect 41604 12835 41656 12844
rect 41604 12801 41613 12835
rect 41613 12801 41647 12835
rect 41647 12801 41656 12835
rect 41604 12792 41656 12801
rect 44180 12792 44232 12844
rect 47860 12792 47912 12844
rect 49148 12835 49200 12844
rect 49148 12801 49157 12835
rect 49157 12801 49191 12835
rect 49191 12801 49200 12835
rect 49148 12792 49200 12801
rect 21272 12656 21324 12708
rect 21824 12588 21876 12640
rect 22468 12588 22520 12640
rect 22836 12588 22888 12640
rect 25228 12656 25280 12708
rect 25412 12656 25464 12708
rect 28540 12656 28592 12708
rect 31576 12724 31628 12776
rect 29460 12588 29512 12640
rect 30104 12588 30156 12640
rect 31024 12631 31076 12640
rect 31024 12597 31033 12631
rect 31033 12597 31067 12631
rect 31067 12597 31076 12631
rect 31024 12588 31076 12597
rect 33324 12724 33376 12776
rect 34888 12724 34940 12776
rect 36452 12767 36504 12776
rect 36452 12733 36461 12767
rect 36461 12733 36495 12767
rect 36495 12733 36504 12767
rect 36452 12724 36504 12733
rect 33968 12656 34020 12708
rect 34152 12656 34204 12708
rect 35440 12656 35492 12708
rect 44180 12656 44232 12708
rect 35164 12588 35216 12640
rect 38476 12588 38528 12640
rect 38752 12588 38804 12640
rect 47952 12588 48004 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 2780 12427 2832 12436
rect 2780 12393 2789 12427
rect 2789 12393 2823 12427
rect 2823 12393 2832 12427
rect 2780 12384 2832 12393
rect 5264 12248 5316 12300
rect 1308 12180 1360 12232
rect 7564 12044 7616 12096
rect 13084 12384 13136 12436
rect 12256 12248 12308 12300
rect 18604 12384 18656 12436
rect 21640 12384 21692 12436
rect 22560 12384 22612 12436
rect 23664 12316 23716 12368
rect 13912 12248 13964 12300
rect 16948 12248 17000 12300
rect 17684 12248 17736 12300
rect 19708 12248 19760 12300
rect 20812 12248 20864 12300
rect 22744 12291 22796 12300
rect 22744 12257 22753 12291
rect 22753 12257 22787 12291
rect 22787 12257 22796 12291
rect 22744 12248 22796 12257
rect 25596 12384 25648 12436
rect 26056 12384 26108 12436
rect 27620 12384 27672 12436
rect 29736 12384 29788 12436
rect 26332 12359 26384 12368
rect 26332 12325 26341 12359
rect 26341 12325 26375 12359
rect 26375 12325 26384 12359
rect 26332 12316 26384 12325
rect 27344 12316 27396 12368
rect 31392 12316 31444 12368
rect 36452 12384 36504 12436
rect 36636 12427 36688 12436
rect 36636 12393 36645 12427
rect 36645 12393 36679 12427
rect 36679 12393 36688 12427
rect 36636 12384 36688 12393
rect 37096 12427 37148 12436
rect 37096 12393 37105 12427
rect 37105 12393 37139 12427
rect 37139 12393 37148 12427
rect 37096 12384 37148 12393
rect 38200 12384 38252 12436
rect 39580 12427 39632 12436
rect 39580 12393 39589 12427
rect 39589 12393 39623 12427
rect 39623 12393 39632 12427
rect 39580 12384 39632 12393
rect 34060 12316 34112 12368
rect 37188 12316 37240 12368
rect 37280 12316 37332 12368
rect 38936 12316 38988 12368
rect 10232 12087 10284 12096
rect 10232 12053 10241 12087
rect 10241 12053 10275 12087
rect 10275 12053 10284 12087
rect 10232 12044 10284 12053
rect 13728 12180 13780 12232
rect 14280 12180 14332 12232
rect 16488 12180 16540 12232
rect 18328 12180 18380 12232
rect 21272 12223 21324 12232
rect 21272 12189 21281 12223
rect 21281 12189 21315 12223
rect 21315 12189 21324 12223
rect 21272 12180 21324 12189
rect 26976 12248 27028 12300
rect 27528 12291 27580 12300
rect 27528 12257 27537 12291
rect 27537 12257 27571 12291
rect 27571 12257 27580 12291
rect 27528 12248 27580 12257
rect 28816 12248 28868 12300
rect 30012 12291 30064 12300
rect 30012 12257 30021 12291
rect 30021 12257 30055 12291
rect 30055 12257 30064 12291
rect 30012 12248 30064 12257
rect 32220 12291 32272 12300
rect 32220 12257 32229 12291
rect 32229 12257 32263 12291
rect 32263 12257 32272 12291
rect 32220 12248 32272 12257
rect 34152 12248 34204 12300
rect 34704 12248 34756 12300
rect 35716 12248 35768 12300
rect 36176 12248 36228 12300
rect 10876 12112 10928 12164
rect 11612 12112 11664 12164
rect 13084 12112 13136 12164
rect 13452 12112 13504 12164
rect 15292 12112 15344 12164
rect 11060 12044 11112 12096
rect 12256 12044 12308 12096
rect 15936 12044 15988 12096
rect 16028 12044 16080 12096
rect 17500 12112 17552 12164
rect 17868 12112 17920 12164
rect 19432 12155 19484 12164
rect 19432 12121 19441 12155
rect 19441 12121 19475 12155
rect 19475 12121 19484 12155
rect 19432 12112 19484 12121
rect 21180 12112 21232 12164
rect 21640 12112 21692 12164
rect 17132 12087 17184 12096
rect 17132 12053 17141 12087
rect 17141 12053 17175 12087
rect 17175 12053 17184 12087
rect 17132 12044 17184 12053
rect 17224 12087 17276 12096
rect 17224 12053 17233 12087
rect 17233 12053 17267 12087
rect 17267 12053 17276 12087
rect 17224 12044 17276 12053
rect 21272 12044 21324 12096
rect 21456 12044 21508 12096
rect 24492 12180 24544 12232
rect 25964 12180 26016 12232
rect 26792 12180 26844 12232
rect 27160 12180 27212 12232
rect 29092 12180 29144 12232
rect 29368 12180 29420 12232
rect 34244 12180 34296 12232
rect 36728 12248 36780 12300
rect 37556 12291 37608 12300
rect 37556 12257 37565 12291
rect 37565 12257 37599 12291
rect 37599 12257 37608 12291
rect 37556 12248 37608 12257
rect 37740 12291 37792 12300
rect 37740 12257 37749 12291
rect 37749 12257 37783 12291
rect 37783 12257 37792 12291
rect 37740 12248 37792 12257
rect 22468 12087 22520 12096
rect 22468 12053 22477 12087
rect 22477 12053 22511 12087
rect 22511 12053 22520 12087
rect 22468 12044 22520 12053
rect 22560 12087 22612 12096
rect 22560 12053 22569 12087
rect 22569 12053 22603 12087
rect 22603 12053 22612 12087
rect 22560 12044 22612 12053
rect 24676 12044 24728 12096
rect 26240 12044 26292 12096
rect 30288 12112 30340 12164
rect 30472 12112 30524 12164
rect 33232 12112 33284 12164
rect 37464 12223 37516 12232
rect 37464 12189 37473 12223
rect 37473 12189 37507 12223
rect 37507 12189 37516 12223
rect 37464 12180 37516 12189
rect 27344 12087 27396 12096
rect 27344 12053 27353 12087
rect 27353 12053 27387 12087
rect 27387 12053 27396 12087
rect 27344 12044 27396 12053
rect 27620 12044 27672 12096
rect 28356 12044 28408 12096
rect 28448 12087 28500 12096
rect 28448 12053 28457 12087
rect 28457 12053 28491 12087
rect 28491 12053 28500 12087
rect 28448 12044 28500 12053
rect 30380 12044 30432 12096
rect 35440 12112 35492 12164
rect 34520 12044 34572 12096
rect 38476 12180 38528 12232
rect 41604 12223 41656 12232
rect 41604 12189 41613 12223
rect 41613 12189 41647 12223
rect 41647 12189 41656 12223
rect 41604 12180 41656 12189
rect 49148 12291 49200 12300
rect 49148 12257 49157 12291
rect 49157 12257 49191 12291
rect 49191 12257 49200 12291
rect 49148 12248 49200 12257
rect 47952 12223 48004 12232
rect 47952 12189 47961 12223
rect 47961 12189 47995 12223
rect 47995 12189 48004 12223
rect 47952 12180 48004 12189
rect 40132 12155 40184 12164
rect 40132 12121 40141 12155
rect 40141 12121 40175 12155
rect 40175 12121 40184 12155
rect 40132 12112 40184 12121
rect 47216 12112 47268 12164
rect 38936 12087 38988 12096
rect 38936 12053 38945 12087
rect 38945 12053 38979 12087
rect 38979 12053 38988 12087
rect 38936 12044 38988 12053
rect 40776 12087 40828 12096
rect 40776 12053 40785 12087
rect 40785 12053 40819 12087
rect 40819 12053 40828 12087
rect 40776 12044 40828 12053
rect 45928 12087 45980 12096
rect 45928 12053 45937 12087
rect 45937 12053 45971 12087
rect 45971 12053 45980 12087
rect 45928 12044 45980 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 4344 11840 4396 11892
rect 9864 11840 9916 11892
rect 10876 11840 10928 11892
rect 1216 11704 1268 11756
rect 1308 11636 1360 11688
rect 10600 11772 10652 11824
rect 13360 11840 13412 11892
rect 15476 11840 15528 11892
rect 16488 11883 16540 11892
rect 16488 11849 16497 11883
rect 16497 11849 16531 11883
rect 16531 11849 16540 11883
rect 16488 11840 16540 11849
rect 16580 11840 16632 11892
rect 20076 11840 20128 11892
rect 20536 11840 20588 11892
rect 22008 11840 22060 11892
rect 22376 11840 22428 11892
rect 25596 11840 25648 11892
rect 25964 11883 26016 11892
rect 25964 11849 25973 11883
rect 25973 11849 26007 11883
rect 26007 11849 26016 11883
rect 25964 11840 26016 11849
rect 27344 11840 27396 11892
rect 28448 11840 28500 11892
rect 14188 11772 14240 11824
rect 14280 11772 14332 11824
rect 14004 11704 14056 11756
rect 14740 11704 14792 11756
rect 15476 11747 15528 11756
rect 15476 11713 15485 11747
rect 15485 11713 15519 11747
rect 15519 11713 15528 11747
rect 15476 11704 15528 11713
rect 20812 11772 20864 11824
rect 22100 11815 22152 11824
rect 22100 11781 22109 11815
rect 22109 11781 22143 11815
rect 22143 11781 22152 11815
rect 22100 11772 22152 11781
rect 23388 11815 23440 11824
rect 23388 11781 23397 11815
rect 23397 11781 23431 11815
rect 23431 11781 23440 11815
rect 23388 11772 23440 11781
rect 16856 11747 16908 11756
rect 12164 11636 12216 11688
rect 12624 11679 12676 11688
rect 12624 11645 12633 11679
rect 12633 11645 12667 11679
rect 12667 11645 12676 11679
rect 12624 11636 12676 11645
rect 12072 11500 12124 11552
rect 13636 11500 13688 11552
rect 14740 11568 14792 11620
rect 14832 11543 14884 11552
rect 14832 11509 14841 11543
rect 14841 11509 14875 11543
rect 14875 11509 14884 11543
rect 14832 11500 14884 11509
rect 15016 11500 15068 11552
rect 15476 11500 15528 11552
rect 16212 11543 16264 11552
rect 16212 11509 16221 11543
rect 16221 11509 16255 11543
rect 16255 11509 16264 11543
rect 16212 11500 16264 11509
rect 16856 11713 16865 11747
rect 16865 11713 16899 11747
rect 16899 11713 16908 11747
rect 16856 11704 16908 11713
rect 18236 11704 18288 11756
rect 19248 11636 19300 11688
rect 22652 11704 22704 11756
rect 24492 11772 24544 11824
rect 27344 11704 27396 11756
rect 28448 11704 28500 11756
rect 29092 11772 29144 11824
rect 29460 11772 29512 11824
rect 30288 11840 30340 11892
rect 31300 11883 31352 11892
rect 31300 11849 31309 11883
rect 31309 11849 31343 11883
rect 31343 11849 31352 11883
rect 31300 11840 31352 11849
rect 32680 11840 32732 11892
rect 30104 11704 30156 11756
rect 37280 11840 37332 11892
rect 34796 11772 34848 11824
rect 36728 11772 36780 11824
rect 37372 11772 37424 11824
rect 19892 11636 19944 11688
rect 18328 11568 18380 11620
rect 20168 11636 20220 11688
rect 21272 11636 21324 11688
rect 21364 11679 21416 11688
rect 21364 11645 21373 11679
rect 21373 11645 21407 11679
rect 21407 11645 21416 11679
rect 21364 11636 21416 11645
rect 20076 11568 20128 11620
rect 22744 11636 22796 11688
rect 26332 11636 26384 11688
rect 27436 11636 27488 11688
rect 22560 11568 22612 11620
rect 27160 11611 27212 11620
rect 27160 11577 27169 11611
rect 27169 11577 27203 11611
rect 27203 11577 27212 11611
rect 27160 11568 27212 11577
rect 19340 11500 19392 11552
rect 19708 11500 19760 11552
rect 22100 11500 22152 11552
rect 28816 11679 28868 11688
rect 28816 11645 28825 11679
rect 28825 11645 28859 11679
rect 28859 11645 28868 11679
rect 28816 11636 28868 11645
rect 29368 11636 29420 11688
rect 31944 11636 31996 11688
rect 32312 11636 32364 11688
rect 32772 11679 32824 11688
rect 32772 11645 32781 11679
rect 32781 11645 32815 11679
rect 32815 11645 32824 11679
rect 32772 11636 32824 11645
rect 29828 11568 29880 11620
rect 30748 11568 30800 11620
rect 34520 11636 34572 11688
rect 34888 11636 34940 11688
rect 38384 11704 38436 11756
rect 40776 11772 40828 11824
rect 49148 11815 49200 11824
rect 49148 11781 49157 11815
rect 49157 11781 49191 11815
rect 49191 11781 49200 11815
rect 49148 11772 49200 11781
rect 45928 11704 45980 11756
rect 35072 11568 35124 11620
rect 29276 11500 29328 11552
rect 29552 11500 29604 11552
rect 31760 11500 31812 11552
rect 32312 11500 32364 11552
rect 33600 11500 33652 11552
rect 33876 11500 33928 11552
rect 35164 11500 35216 11552
rect 39120 11679 39172 11688
rect 39120 11645 39129 11679
rect 39129 11645 39163 11679
rect 39163 11645 39172 11679
rect 39120 11636 39172 11645
rect 39212 11679 39264 11688
rect 39212 11645 39221 11679
rect 39221 11645 39255 11679
rect 39255 11645 39264 11679
rect 39212 11636 39264 11645
rect 40132 11636 40184 11688
rect 37372 11568 37424 11620
rect 41604 11568 41656 11620
rect 46664 11568 46716 11620
rect 35624 11500 35676 11552
rect 35992 11500 36044 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 1216 11296 1268 11348
rect 9864 11296 9916 11348
rect 10784 11296 10836 11348
rect 1768 11271 1820 11280
rect 1768 11237 1777 11271
rect 1777 11237 1811 11271
rect 1811 11237 1820 11271
rect 1768 11228 1820 11237
rect 10232 11228 10284 11280
rect 10876 11160 10928 11212
rect 13912 11271 13964 11280
rect 13912 11237 13921 11271
rect 13921 11237 13955 11271
rect 13955 11237 13964 11271
rect 13912 11228 13964 11237
rect 14556 11339 14608 11348
rect 14556 11305 14565 11339
rect 14565 11305 14599 11339
rect 14599 11305 14608 11339
rect 14556 11296 14608 11305
rect 16212 11296 16264 11348
rect 16488 11296 16540 11348
rect 16948 11339 17000 11348
rect 16948 11305 16957 11339
rect 16957 11305 16991 11339
rect 16991 11305 17000 11339
rect 16948 11296 17000 11305
rect 19064 11296 19116 11348
rect 20168 11296 20220 11348
rect 15568 11228 15620 11280
rect 16028 11228 16080 11280
rect 12164 11160 12216 11212
rect 1584 11135 1636 11144
rect 1584 11101 1593 11135
rect 1593 11101 1627 11135
rect 1627 11101 1636 11135
rect 1584 11092 1636 11101
rect 12716 11160 12768 11212
rect 15016 11203 15068 11212
rect 15016 11169 15025 11203
rect 15025 11169 15059 11203
rect 15059 11169 15068 11203
rect 15016 11160 15068 11169
rect 15108 11203 15160 11212
rect 15108 11169 15117 11203
rect 15117 11169 15151 11203
rect 15151 11169 15160 11203
rect 15108 11160 15160 11169
rect 16120 11160 16172 11212
rect 20076 11228 20128 11280
rect 23296 11339 23348 11348
rect 23296 11305 23305 11339
rect 23305 11305 23339 11339
rect 23339 11305 23348 11339
rect 23296 11296 23348 11305
rect 26608 11296 26660 11348
rect 27160 11296 27212 11348
rect 23572 11228 23624 11280
rect 29000 11339 29052 11348
rect 29000 11305 29009 11339
rect 29009 11305 29043 11339
rect 29043 11305 29052 11339
rect 29000 11296 29052 11305
rect 29368 11228 29420 11280
rect 18604 11203 18656 11212
rect 18604 11169 18613 11203
rect 18613 11169 18647 11203
rect 18647 11169 18656 11203
rect 18604 11160 18656 11169
rect 19708 11160 19760 11212
rect 20628 11160 20680 11212
rect 22468 11160 22520 11212
rect 24032 11160 24084 11212
rect 24492 11160 24544 11212
rect 27528 11160 27580 11212
rect 29184 11160 29236 11212
rect 29644 11160 29696 11212
rect 18512 11135 18564 11144
rect 18512 11101 18521 11135
rect 18521 11101 18555 11135
rect 18555 11101 18564 11135
rect 18512 11092 18564 11101
rect 18972 11092 19024 11144
rect 24308 11092 24360 11144
rect 25964 11092 26016 11144
rect 26700 11092 26752 11144
rect 10600 11067 10652 11076
rect 10600 11033 10609 11067
rect 10609 11033 10643 11067
rect 10643 11033 10652 11067
rect 10600 11024 10652 11033
rect 11428 10956 11480 11008
rect 11704 10956 11756 11008
rect 11888 11024 11940 11076
rect 13360 10956 13412 11008
rect 15108 11024 15160 11076
rect 16120 11067 16172 11076
rect 16120 11033 16129 11067
rect 16129 11033 16163 11067
rect 16163 11033 16172 11067
rect 16120 11024 16172 11033
rect 15016 10956 15068 11008
rect 15752 10999 15804 11008
rect 15752 10965 15761 10999
rect 15761 10965 15795 10999
rect 15795 10965 15804 10999
rect 15752 10956 15804 10965
rect 17500 10956 17552 11008
rect 18236 10956 18288 11008
rect 20904 11024 20956 11076
rect 21088 11024 21140 11076
rect 23756 11067 23808 11076
rect 23756 11033 23765 11067
rect 23765 11033 23799 11067
rect 23799 11033 23808 11067
rect 23756 11024 23808 11033
rect 24860 11067 24912 11076
rect 24860 11033 24869 11067
rect 24869 11033 24903 11067
rect 24903 11033 24912 11067
rect 24860 11024 24912 11033
rect 26884 11135 26936 11144
rect 26884 11101 26893 11135
rect 26893 11101 26927 11135
rect 26927 11101 26936 11135
rect 26884 11092 26936 11101
rect 31392 11296 31444 11348
rect 34612 11296 34664 11348
rect 35072 11296 35124 11348
rect 31760 11160 31812 11212
rect 32680 11160 32732 11212
rect 32864 11203 32916 11212
rect 32864 11169 32873 11203
rect 32873 11169 32907 11203
rect 32907 11169 32916 11203
rect 32864 11160 32916 11169
rect 33600 11160 33652 11212
rect 34244 11160 34296 11212
rect 37372 11228 37424 11280
rect 39120 11160 39172 11212
rect 20812 10956 20864 11008
rect 21640 10956 21692 11008
rect 24676 10956 24728 11008
rect 29368 11024 29420 11076
rect 29736 11067 29788 11076
rect 29736 11033 29745 11067
rect 29745 11033 29779 11067
rect 29779 11033 29788 11067
rect 29736 11024 29788 11033
rect 30380 11024 30432 11076
rect 33784 11092 33836 11144
rect 34152 11092 34204 11144
rect 35624 11092 35676 11144
rect 37280 11092 37332 11144
rect 39212 11092 39264 11144
rect 47124 11296 47176 11348
rect 44180 11228 44232 11280
rect 40040 11092 40092 11144
rect 49148 11203 49200 11212
rect 49148 11169 49157 11203
rect 49157 11169 49191 11203
rect 49191 11169 49200 11203
rect 49148 11160 49200 11169
rect 28724 10956 28776 11008
rect 29460 10956 29512 11008
rect 30288 10956 30340 11008
rect 32312 10956 32364 11008
rect 33876 11067 33928 11076
rect 33876 11033 33885 11067
rect 33885 11033 33919 11067
rect 33919 11033 33928 11067
rect 35256 11067 35308 11076
rect 33876 11024 33928 11033
rect 35256 11033 35265 11067
rect 35265 11033 35299 11067
rect 35299 11033 35308 11067
rect 35256 11024 35308 11033
rect 35992 11067 36044 11076
rect 35992 11033 36001 11067
rect 36001 11033 36035 11067
rect 36035 11033 36044 11067
rect 35992 11024 36044 11033
rect 36728 11024 36780 11076
rect 37740 11067 37792 11076
rect 37740 11033 37749 11067
rect 37749 11033 37783 11067
rect 37783 11033 37792 11067
rect 37740 11024 37792 11033
rect 40132 11067 40184 11076
rect 40132 11033 40141 11067
rect 40141 11033 40175 11067
rect 40175 11033 40184 11067
rect 40132 11024 40184 11033
rect 40776 11024 40828 11076
rect 44180 11024 44232 11076
rect 46940 11024 46992 11076
rect 33324 10956 33376 11008
rect 35164 10999 35216 11008
rect 35164 10965 35173 10999
rect 35173 10965 35207 10999
rect 35207 10965 35216 10999
rect 35164 10956 35216 10965
rect 39304 10999 39356 11008
rect 39304 10965 39313 10999
rect 39313 10965 39347 10999
rect 39347 10965 39356 10999
rect 39304 10956 39356 10965
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 1860 10752 1912 10804
rect 11428 10752 11480 10804
rect 11704 10752 11756 10804
rect 12532 10752 12584 10804
rect 15200 10752 15252 10804
rect 1216 10684 1268 10736
rect 1308 10616 1360 10668
rect 14924 10684 14976 10736
rect 10324 10616 10376 10668
rect 12256 10616 12308 10668
rect 13820 10591 13872 10600
rect 13820 10557 13829 10591
rect 13829 10557 13863 10591
rect 13863 10557 13872 10591
rect 13820 10548 13872 10557
rect 17776 10684 17828 10736
rect 16488 10616 16540 10668
rect 16580 10616 16632 10668
rect 18328 10752 18380 10804
rect 18788 10795 18840 10804
rect 18788 10761 18797 10795
rect 18797 10761 18831 10795
rect 18831 10761 18840 10795
rect 18788 10752 18840 10761
rect 19616 10752 19668 10804
rect 20720 10795 20772 10804
rect 20720 10761 20729 10795
rect 20729 10761 20763 10795
rect 20763 10761 20772 10795
rect 20720 10752 20772 10761
rect 20904 10752 20956 10804
rect 22652 10752 22704 10804
rect 23572 10752 23624 10804
rect 24400 10752 24452 10804
rect 24492 10752 24544 10804
rect 25320 10795 25372 10804
rect 25320 10761 25329 10795
rect 25329 10761 25363 10795
rect 25363 10761 25372 10795
rect 25320 10752 25372 10761
rect 25964 10752 26016 10804
rect 31484 10752 31536 10804
rect 33324 10795 33376 10804
rect 33324 10761 33333 10795
rect 33333 10761 33367 10795
rect 33367 10761 33376 10795
rect 33324 10752 33376 10761
rect 18604 10684 18656 10736
rect 21456 10684 21508 10736
rect 12808 10480 12860 10532
rect 14832 10480 14884 10532
rect 2504 10455 2556 10464
rect 2504 10421 2513 10455
rect 2513 10421 2547 10455
rect 2547 10421 2556 10455
rect 2504 10412 2556 10421
rect 11244 10455 11296 10464
rect 11244 10421 11253 10455
rect 11253 10421 11287 10455
rect 11287 10421 11296 10455
rect 11244 10412 11296 10421
rect 12716 10412 12768 10464
rect 14372 10455 14424 10464
rect 14372 10421 14381 10455
rect 14381 10421 14415 10455
rect 14415 10421 14424 10455
rect 14372 10412 14424 10421
rect 15384 10548 15436 10600
rect 16212 10591 16264 10600
rect 16212 10557 16221 10591
rect 16221 10557 16255 10591
rect 16255 10557 16264 10591
rect 16212 10548 16264 10557
rect 16396 10548 16448 10600
rect 18696 10659 18748 10668
rect 18696 10625 18705 10659
rect 18705 10625 18739 10659
rect 18739 10625 18748 10659
rect 18696 10616 18748 10625
rect 19892 10659 19944 10668
rect 19892 10625 19901 10659
rect 19901 10625 19935 10659
rect 19935 10625 19944 10659
rect 19892 10616 19944 10625
rect 20536 10616 20588 10668
rect 20996 10616 21048 10668
rect 21088 10616 21140 10668
rect 24032 10684 24084 10736
rect 24676 10727 24728 10736
rect 24676 10693 24685 10727
rect 24685 10693 24719 10727
rect 24719 10693 24728 10727
rect 24676 10684 24728 10693
rect 27620 10684 27672 10736
rect 29276 10684 29328 10736
rect 24584 10659 24636 10668
rect 24584 10625 24593 10659
rect 24593 10625 24627 10659
rect 24627 10625 24636 10659
rect 24584 10616 24636 10625
rect 18788 10548 18840 10600
rect 18880 10591 18932 10600
rect 18880 10557 18889 10591
rect 18889 10557 18923 10591
rect 18923 10557 18932 10591
rect 18880 10548 18932 10557
rect 21180 10548 21232 10600
rect 16672 10480 16724 10532
rect 16764 10480 16816 10532
rect 22008 10591 22060 10600
rect 22008 10557 22017 10591
rect 22017 10557 22051 10591
rect 22051 10557 22060 10591
rect 22008 10548 22060 10557
rect 22284 10591 22336 10600
rect 22284 10557 22293 10591
rect 22293 10557 22327 10591
rect 22327 10557 22336 10591
rect 22284 10548 22336 10557
rect 22376 10548 22428 10600
rect 26608 10616 26660 10668
rect 27068 10616 27120 10668
rect 29644 10616 29696 10668
rect 29920 10684 29972 10736
rect 40132 10752 40184 10804
rect 40776 10752 40828 10804
rect 35532 10684 35584 10736
rect 49240 10684 49292 10736
rect 31300 10659 31352 10668
rect 31300 10625 31309 10659
rect 31309 10625 31343 10659
rect 31343 10625 31352 10659
rect 31300 10616 31352 10625
rect 35164 10616 35216 10668
rect 35716 10616 35768 10668
rect 36452 10659 36504 10668
rect 36452 10625 36461 10659
rect 36461 10625 36495 10659
rect 36495 10625 36504 10659
rect 36452 10616 36504 10625
rect 27252 10548 27304 10600
rect 17592 10412 17644 10464
rect 18328 10455 18380 10464
rect 18328 10421 18337 10455
rect 18337 10421 18371 10455
rect 18371 10421 18380 10455
rect 18328 10412 18380 10421
rect 28816 10548 28868 10600
rect 29000 10548 29052 10600
rect 31576 10591 31628 10600
rect 31576 10557 31585 10591
rect 31585 10557 31619 10591
rect 31619 10557 31628 10591
rect 31576 10548 31628 10557
rect 22744 10412 22796 10464
rect 26608 10455 26660 10464
rect 26608 10421 26617 10455
rect 26617 10421 26651 10455
rect 26651 10421 26660 10455
rect 26608 10412 26660 10421
rect 29276 10412 29328 10464
rect 30932 10523 30984 10532
rect 30932 10489 30941 10523
rect 30941 10489 30975 10523
rect 30975 10489 30984 10523
rect 30932 10480 30984 10489
rect 33784 10591 33836 10600
rect 33784 10557 33793 10591
rect 33793 10557 33827 10591
rect 33827 10557 33836 10591
rect 33784 10548 33836 10557
rect 35808 10548 35860 10600
rect 37280 10616 37332 10668
rect 36636 10548 36688 10600
rect 39488 10616 39540 10668
rect 46940 10616 46992 10668
rect 47032 10548 47084 10600
rect 31392 10412 31444 10464
rect 31484 10412 31536 10464
rect 33416 10412 33468 10464
rect 35900 10480 35952 10532
rect 40040 10480 40092 10532
rect 36544 10412 36596 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 12624 10208 12676 10260
rect 12808 10208 12860 10260
rect 13268 10208 13320 10260
rect 16488 10208 16540 10260
rect 16672 10208 16724 10260
rect 17224 10208 17276 10260
rect 18972 10208 19024 10260
rect 19432 10208 19484 10260
rect 22560 10208 22612 10260
rect 26608 10208 26660 10260
rect 26700 10251 26752 10260
rect 26700 10217 26709 10251
rect 26709 10217 26743 10251
rect 26743 10217 26752 10251
rect 26700 10208 26752 10217
rect 27252 10208 27304 10260
rect 19800 10140 19852 10192
rect 21732 10140 21784 10192
rect 1860 10115 1912 10124
rect 1860 10081 1869 10115
rect 1869 10081 1903 10115
rect 1903 10081 1912 10115
rect 1860 10072 1912 10081
rect 10416 10072 10468 10124
rect 12532 10072 12584 10124
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 13544 10072 13596 10081
rect 14280 10115 14332 10124
rect 14280 10081 14289 10115
rect 14289 10081 14323 10115
rect 14323 10081 14332 10115
rect 14280 10072 14332 10081
rect 16304 10072 16356 10124
rect 18512 10072 18564 10124
rect 18880 10072 18932 10124
rect 19524 10072 19576 10124
rect 20628 10072 20680 10124
rect 22008 10072 22060 10124
rect 23296 10115 23348 10124
rect 23296 10081 23305 10115
rect 23305 10081 23339 10115
rect 23339 10081 23348 10115
rect 23296 10072 23348 10081
rect 27620 10072 27672 10124
rect 29368 10251 29420 10260
rect 29368 10217 29377 10251
rect 29377 10217 29411 10251
rect 29411 10217 29420 10251
rect 29368 10208 29420 10217
rect 31760 10208 31812 10260
rect 32496 10208 32548 10260
rect 36544 10208 36596 10260
rect 36636 10251 36688 10260
rect 36636 10217 36645 10251
rect 36645 10217 36679 10251
rect 36679 10217 36688 10251
rect 36636 10208 36688 10217
rect 28816 10140 28868 10192
rect 29828 10140 29880 10192
rect 30196 10140 30248 10192
rect 34796 10140 34848 10192
rect 46940 10140 46992 10192
rect 1308 10004 1360 10056
rect 13360 10004 13412 10056
rect 16764 10047 16816 10056
rect 16764 10013 16773 10047
rect 16773 10013 16807 10047
rect 16807 10013 16816 10047
rect 16764 10004 16816 10013
rect 18604 10004 18656 10056
rect 11428 9936 11480 9988
rect 14096 9936 14148 9988
rect 15292 9936 15344 9988
rect 16396 9936 16448 9988
rect 16488 9936 16540 9988
rect 17500 9936 17552 9988
rect 11244 9868 11296 9920
rect 13268 9868 13320 9920
rect 19340 9868 19392 9920
rect 21088 9936 21140 9988
rect 21364 9868 21416 9920
rect 21456 9868 21508 9920
rect 22836 10004 22888 10056
rect 25964 10004 26016 10056
rect 26976 10047 27028 10056
rect 26976 10013 26985 10047
rect 26985 10013 27019 10047
rect 27019 10013 27028 10047
rect 26976 10004 27028 10013
rect 28540 10004 28592 10056
rect 29368 10004 29420 10056
rect 22560 9979 22612 9988
rect 22560 9945 22569 9979
rect 22569 9945 22603 9979
rect 22603 9945 22612 9979
rect 22560 9936 22612 9945
rect 24124 9936 24176 9988
rect 31300 10072 31352 10124
rect 31392 10072 31444 10124
rect 33416 10072 33468 10124
rect 34336 10072 34388 10124
rect 34428 10115 34480 10124
rect 34428 10081 34437 10115
rect 34437 10081 34471 10115
rect 34471 10081 34480 10115
rect 34428 10072 34480 10081
rect 39488 10115 39540 10124
rect 39488 10081 39497 10115
rect 39497 10081 39531 10115
rect 39531 10081 39540 10115
rect 39488 10072 39540 10081
rect 45836 10072 45888 10124
rect 49148 10115 49200 10124
rect 49148 10081 49157 10115
rect 49157 10081 49191 10115
rect 49191 10081 49200 10115
rect 49148 10072 49200 10081
rect 30380 10047 30432 10056
rect 30380 10013 30389 10047
rect 30389 10013 30423 10047
rect 30423 10013 30432 10047
rect 30380 10004 30432 10013
rect 33324 10004 33376 10056
rect 33692 10047 33744 10056
rect 22008 9868 22060 9920
rect 24032 9911 24084 9920
rect 24032 9877 24041 9911
rect 24041 9877 24075 9911
rect 24075 9877 24084 9911
rect 24032 9868 24084 9877
rect 24952 9868 25004 9920
rect 26424 9868 26476 9920
rect 30564 9936 30616 9988
rect 30656 9979 30708 9988
rect 30656 9945 30665 9979
rect 30665 9945 30699 9979
rect 30699 9945 30708 9979
rect 30656 9936 30708 9945
rect 32312 9936 32364 9988
rect 33692 10013 33701 10047
rect 33701 10013 33735 10047
rect 33735 10013 33744 10047
rect 33692 10004 33744 10013
rect 33784 10004 33836 10056
rect 34888 10047 34940 10056
rect 34888 10013 34897 10047
rect 34897 10013 34931 10047
rect 34931 10013 34940 10047
rect 34888 10004 34940 10013
rect 33508 9936 33560 9988
rect 36544 9936 36596 9988
rect 34244 9868 34296 9920
rect 35440 9868 35492 9920
rect 39304 10004 39356 10056
rect 38292 9979 38344 9988
rect 38292 9945 38301 9979
rect 38301 9945 38335 9979
rect 38335 9945 38344 9979
rect 38292 9936 38344 9945
rect 40316 9936 40368 9988
rect 44180 10004 44232 10056
rect 46664 10004 46716 10056
rect 46756 9936 46808 9988
rect 47308 9979 47360 9988
rect 47308 9945 47317 9979
rect 47317 9945 47351 9979
rect 47351 9945 47360 9979
rect 47308 9936 47360 9945
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 1308 9664 1360 9716
rect 13820 9664 13872 9716
rect 16212 9664 16264 9716
rect 19064 9664 19116 9716
rect 20444 9664 20496 9716
rect 21088 9664 21140 9716
rect 12716 9596 12768 9648
rect 1308 9528 1360 9580
rect 12532 9528 12584 9580
rect 1860 9503 1912 9512
rect 1860 9469 1869 9503
rect 1869 9469 1903 9503
rect 1903 9469 1912 9503
rect 1860 9460 1912 9469
rect 13360 9460 13412 9512
rect 14004 9596 14056 9648
rect 15200 9596 15252 9648
rect 15844 9639 15896 9648
rect 15844 9605 15853 9639
rect 15853 9605 15887 9639
rect 15887 9605 15896 9639
rect 15844 9596 15896 9605
rect 16580 9596 16632 9648
rect 17592 9596 17644 9648
rect 20352 9596 20404 9648
rect 21088 9528 21140 9580
rect 21824 9528 21876 9580
rect 21916 9528 21968 9580
rect 23388 9664 23440 9716
rect 26424 9664 26476 9716
rect 26976 9664 27028 9716
rect 23112 9639 23164 9648
rect 23112 9605 23121 9639
rect 23121 9605 23155 9639
rect 23155 9605 23164 9639
rect 23112 9596 23164 9605
rect 23756 9596 23808 9648
rect 26056 9596 26108 9648
rect 22376 9571 22428 9580
rect 22376 9537 22385 9571
rect 22385 9537 22419 9571
rect 22419 9537 22428 9571
rect 22376 9528 22428 9537
rect 23296 9528 23348 9580
rect 26148 9571 26200 9580
rect 26148 9537 26157 9571
rect 26157 9537 26191 9571
rect 26191 9537 26200 9571
rect 26148 9528 26200 9537
rect 11244 9324 11296 9376
rect 13912 9503 13964 9512
rect 13912 9469 13921 9503
rect 13921 9469 13955 9503
rect 13955 9469 13964 9503
rect 13912 9460 13964 9469
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 17132 9503 17184 9512
rect 17132 9469 17141 9503
rect 17141 9469 17175 9503
rect 17175 9469 17184 9503
rect 17132 9460 17184 9469
rect 17684 9460 17736 9512
rect 14280 9324 14332 9376
rect 16856 9324 16908 9376
rect 17868 9324 17920 9376
rect 19616 9503 19668 9512
rect 19616 9469 19625 9503
rect 19625 9469 19659 9503
rect 19659 9469 19668 9503
rect 19616 9460 19668 9469
rect 19708 9460 19760 9512
rect 22192 9460 22244 9512
rect 22468 9503 22520 9512
rect 22468 9469 22477 9503
rect 22477 9469 22511 9503
rect 22511 9469 22520 9503
rect 22468 9460 22520 9469
rect 23480 9460 23532 9512
rect 25504 9460 25556 9512
rect 26424 9503 26476 9512
rect 26424 9469 26433 9503
rect 26433 9469 26467 9503
rect 26467 9469 26476 9503
rect 26424 9460 26476 9469
rect 29276 9664 29328 9716
rect 29276 9528 29328 9580
rect 21180 9324 21232 9376
rect 21272 9324 21324 9376
rect 21824 9324 21876 9376
rect 27436 9392 27488 9444
rect 22560 9324 22612 9376
rect 23848 9324 23900 9376
rect 27068 9367 27120 9376
rect 27068 9333 27077 9367
rect 27077 9333 27111 9367
rect 27111 9333 27120 9367
rect 27068 9324 27120 9333
rect 27252 9367 27304 9376
rect 27252 9333 27261 9367
rect 27261 9333 27295 9367
rect 27295 9333 27304 9367
rect 27252 9324 27304 9333
rect 29092 9460 29144 9512
rect 30288 9596 30340 9648
rect 34336 9664 34388 9716
rect 34980 9664 35032 9716
rect 35440 9664 35492 9716
rect 37280 9707 37332 9716
rect 37280 9673 37289 9707
rect 37289 9673 37323 9707
rect 37323 9673 37332 9707
rect 37280 9664 37332 9673
rect 32312 9571 32364 9580
rect 32312 9537 32321 9571
rect 32321 9537 32355 9571
rect 32355 9537 32364 9571
rect 32312 9528 32364 9537
rect 32404 9528 32456 9580
rect 30012 9503 30064 9512
rect 30012 9469 30021 9503
rect 30021 9469 30055 9503
rect 30055 9469 30064 9503
rect 30012 9460 30064 9469
rect 32220 9460 32272 9512
rect 29552 9392 29604 9444
rect 31668 9392 31720 9444
rect 35716 9596 35768 9648
rect 36544 9596 36596 9648
rect 49332 9596 49384 9648
rect 35532 9528 35584 9580
rect 47216 9528 47268 9580
rect 33876 9503 33928 9512
rect 33876 9469 33885 9503
rect 33885 9469 33919 9503
rect 33919 9469 33928 9503
rect 33876 9460 33928 9469
rect 34520 9460 34572 9512
rect 38384 9460 38436 9512
rect 29092 9324 29144 9376
rect 29184 9324 29236 9376
rect 31484 9367 31536 9376
rect 31484 9333 31493 9367
rect 31493 9333 31527 9367
rect 31527 9333 31536 9367
rect 31484 9324 31536 9333
rect 35532 9324 35584 9376
rect 36728 9367 36780 9376
rect 36728 9333 36737 9367
rect 36737 9333 36771 9367
rect 36771 9333 36780 9367
rect 36728 9324 36780 9333
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 12348 9120 12400 9172
rect 2412 8984 2464 9036
rect 11152 8984 11204 9036
rect 13728 9120 13780 9172
rect 18788 9120 18840 9172
rect 19708 9120 19760 9172
rect 19892 9120 19944 9172
rect 20812 9120 20864 9172
rect 22652 9120 22704 9172
rect 23572 9120 23624 9172
rect 24492 9120 24544 9172
rect 24860 9120 24912 9172
rect 27804 9120 27856 9172
rect 29920 9120 29972 9172
rect 21824 9052 21876 9104
rect 13636 9027 13688 9036
rect 13636 8993 13645 9027
rect 13645 8993 13679 9027
rect 13679 8993 13688 9027
rect 13636 8984 13688 8993
rect 14188 8984 14240 9036
rect 22376 9052 22428 9104
rect 30472 9120 30524 9172
rect 34520 9120 34572 9172
rect 36452 9120 36504 9172
rect 1216 8916 1268 8968
rect 14280 8959 14332 8968
rect 14280 8925 14289 8959
rect 14289 8925 14323 8959
rect 14323 8925 14332 8959
rect 14280 8916 14332 8925
rect 1308 8848 1360 8900
rect 12440 8848 12492 8900
rect 14556 8891 14608 8900
rect 14556 8857 14565 8891
rect 14565 8857 14599 8891
rect 14599 8857 14608 8891
rect 14556 8848 14608 8857
rect 15200 8848 15252 8900
rect 1768 8823 1820 8832
rect 1768 8789 1777 8823
rect 1777 8789 1811 8823
rect 1811 8789 1820 8823
rect 1768 8780 1820 8789
rect 2504 8823 2556 8832
rect 2504 8789 2513 8823
rect 2513 8789 2547 8823
rect 2547 8789 2556 8823
rect 2504 8780 2556 8789
rect 11980 8780 12032 8832
rect 16856 8916 16908 8968
rect 19432 8959 19484 8968
rect 19432 8925 19441 8959
rect 19441 8925 19475 8959
rect 19475 8925 19484 8959
rect 19432 8916 19484 8925
rect 17408 8891 17460 8900
rect 17408 8857 17417 8891
rect 17417 8857 17451 8891
rect 17451 8857 17460 8891
rect 17408 8848 17460 8857
rect 19708 8891 19760 8900
rect 19708 8857 19717 8891
rect 19717 8857 19751 8891
rect 19751 8857 19760 8891
rect 19708 8848 19760 8857
rect 20444 8848 20496 8900
rect 21548 8916 21600 8968
rect 22376 8916 22428 8968
rect 23480 8959 23532 8968
rect 23480 8925 23489 8959
rect 23489 8925 23523 8959
rect 23523 8925 23532 8959
rect 23480 8916 23532 8925
rect 23572 8959 23624 8968
rect 23572 8925 23581 8959
rect 23581 8925 23615 8959
rect 23615 8925 23624 8959
rect 23572 8916 23624 8925
rect 23848 8984 23900 9036
rect 24124 9027 24176 9036
rect 24124 8993 24133 9027
rect 24133 8993 24167 9027
rect 24167 8993 24176 9027
rect 24124 8984 24176 8993
rect 24584 8984 24636 9036
rect 32036 9052 32088 9104
rect 36820 9120 36872 9172
rect 40040 9052 40092 9104
rect 29000 8984 29052 9036
rect 30104 8984 30156 9036
rect 32864 8984 32916 9036
rect 33600 9027 33652 9036
rect 33600 8993 33609 9027
rect 33609 8993 33643 9027
rect 33643 8993 33652 9027
rect 33600 8984 33652 8993
rect 34612 8984 34664 9036
rect 34796 8984 34848 9036
rect 35440 9027 35492 9036
rect 35440 8993 35449 9027
rect 35449 8993 35483 9027
rect 35483 8993 35492 9027
rect 35440 8984 35492 8993
rect 35532 8984 35584 9036
rect 22560 8848 22612 8900
rect 23664 8848 23716 8900
rect 25596 8916 25648 8968
rect 27160 8916 27212 8968
rect 27252 8848 27304 8900
rect 16028 8823 16080 8832
rect 16028 8789 16037 8823
rect 16037 8789 16071 8823
rect 16071 8789 16080 8823
rect 16028 8780 16080 8789
rect 16488 8823 16540 8832
rect 16488 8789 16497 8823
rect 16497 8789 16531 8823
rect 16531 8789 16540 8823
rect 16488 8780 16540 8789
rect 17592 8780 17644 8832
rect 19064 8780 19116 8832
rect 19892 8780 19944 8832
rect 20076 8780 20128 8832
rect 20996 8780 21048 8832
rect 21272 8780 21324 8832
rect 29000 8848 29052 8900
rect 30748 8959 30800 8968
rect 30748 8925 30757 8959
rect 30757 8925 30791 8959
rect 30791 8925 30800 8959
rect 30748 8916 30800 8925
rect 33324 8959 33376 8968
rect 33324 8925 33333 8959
rect 33333 8925 33367 8959
rect 33367 8925 33376 8959
rect 33324 8916 33376 8925
rect 33416 8959 33468 8968
rect 33416 8925 33425 8959
rect 33425 8925 33459 8959
rect 33459 8925 33468 8959
rect 33416 8916 33468 8925
rect 33968 8916 34020 8968
rect 31300 8848 31352 8900
rect 32312 8848 32364 8900
rect 27804 8780 27856 8832
rect 29276 8823 29328 8832
rect 29276 8789 29285 8823
rect 29285 8789 29319 8823
rect 29319 8789 29328 8823
rect 29276 8780 29328 8789
rect 30380 8780 30432 8832
rect 31024 8780 31076 8832
rect 34152 8780 34204 8832
rect 34520 8823 34572 8832
rect 34520 8789 34529 8823
rect 34529 8789 34563 8823
rect 34563 8789 34572 8823
rect 34520 8780 34572 8789
rect 34612 8780 34664 8832
rect 36544 8848 36596 8900
rect 36820 8959 36872 8968
rect 36820 8925 36829 8959
rect 36829 8925 36863 8959
rect 36863 8925 36872 8959
rect 36820 8916 36872 8925
rect 49240 8984 49292 9036
rect 37280 8848 37332 8900
rect 47124 8916 47176 8968
rect 36268 8780 36320 8832
rect 42708 8848 42760 8900
rect 39580 8780 39632 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 13728 8619 13780 8628
rect 13728 8585 13737 8619
rect 13737 8585 13771 8619
rect 13771 8585 13780 8619
rect 13728 8576 13780 8585
rect 14556 8576 14608 8628
rect 15108 8619 15160 8628
rect 15108 8585 15117 8619
rect 15117 8585 15151 8619
rect 15151 8585 15160 8619
rect 15108 8576 15160 8585
rect 15752 8619 15804 8628
rect 15752 8585 15761 8619
rect 15761 8585 15795 8619
rect 15795 8585 15804 8619
rect 15752 8576 15804 8585
rect 15936 8576 15988 8628
rect 16396 8576 16448 8628
rect 1768 8508 1820 8560
rect 14188 8508 14240 8560
rect 14280 8508 14332 8560
rect 4068 8440 4120 8492
rect 13820 8440 13872 8492
rect 17224 8508 17276 8560
rect 18696 8576 18748 8628
rect 19432 8576 19484 8628
rect 17592 8508 17644 8560
rect 16856 8483 16908 8492
rect 1400 8372 1452 8424
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 20628 8576 20680 8628
rect 20996 8576 21048 8628
rect 22376 8576 22428 8628
rect 22744 8576 22796 8628
rect 24492 8619 24544 8628
rect 24492 8585 24501 8619
rect 24501 8585 24535 8619
rect 24535 8585 24544 8619
rect 24492 8576 24544 8585
rect 25504 8619 25556 8628
rect 25504 8585 25513 8619
rect 25513 8585 25547 8619
rect 25547 8585 25556 8619
rect 25504 8576 25556 8585
rect 26056 8576 26108 8628
rect 27620 8576 27672 8628
rect 20444 8508 20496 8560
rect 23664 8508 23716 8560
rect 25044 8440 25096 8492
rect 26424 8440 26476 8492
rect 29460 8576 29512 8628
rect 31024 8619 31076 8628
rect 31024 8585 31033 8619
rect 31033 8585 31067 8619
rect 31067 8585 31076 8619
rect 31024 8576 31076 8585
rect 31300 8576 31352 8628
rect 29092 8508 29144 8560
rect 30380 8508 30432 8560
rect 30748 8508 30800 8560
rect 33876 8576 33928 8628
rect 34244 8576 34296 8628
rect 34612 8619 34664 8628
rect 34612 8585 34621 8619
rect 34621 8585 34655 8619
rect 34655 8585 34664 8619
rect 34612 8576 34664 8585
rect 35348 8619 35400 8628
rect 35348 8585 35357 8619
rect 35357 8585 35391 8619
rect 35391 8585 35400 8619
rect 35348 8576 35400 8585
rect 44824 8576 44876 8628
rect 31392 8483 31444 8492
rect 31392 8449 31401 8483
rect 31401 8449 31435 8483
rect 31435 8449 31444 8483
rect 31392 8440 31444 8449
rect 35256 8483 35308 8492
rect 35256 8449 35265 8483
rect 35265 8449 35299 8483
rect 35299 8449 35308 8483
rect 35256 8440 35308 8449
rect 16120 8372 16172 8424
rect 18880 8372 18932 8424
rect 21456 8372 21508 8424
rect 21548 8372 21600 8424
rect 22100 8372 22152 8424
rect 25228 8372 25280 8424
rect 30380 8372 30432 8424
rect 30748 8372 30800 8424
rect 31668 8415 31720 8424
rect 31668 8381 31677 8415
rect 31677 8381 31711 8415
rect 31711 8381 31720 8415
rect 31668 8372 31720 8381
rect 36728 8440 36780 8492
rect 39580 8508 39632 8560
rect 47676 8508 47728 8560
rect 49148 8551 49200 8560
rect 49148 8517 49157 8551
rect 49157 8517 49191 8551
rect 49191 8517 49200 8551
rect 49148 8508 49200 8517
rect 18604 8347 18656 8356
rect 18604 8313 18613 8347
rect 18613 8313 18647 8347
rect 18647 8313 18656 8347
rect 18604 8304 18656 8313
rect 26056 8347 26108 8356
rect 26056 8313 26065 8347
rect 26065 8313 26099 8347
rect 26099 8313 26108 8347
rect 26056 8304 26108 8313
rect 32220 8304 32272 8356
rect 34060 8347 34112 8356
rect 34060 8313 34069 8347
rect 34069 8313 34103 8347
rect 34103 8313 34112 8347
rect 35808 8372 35860 8424
rect 41328 8440 41380 8492
rect 45836 8483 45888 8492
rect 45836 8449 45845 8483
rect 45845 8449 45879 8483
rect 45879 8449 45888 8483
rect 45836 8440 45888 8449
rect 46756 8440 46808 8492
rect 34060 8304 34112 8313
rect 41420 8304 41472 8356
rect 46848 8415 46900 8424
rect 46848 8381 46857 8415
rect 46857 8381 46891 8415
rect 46891 8381 46900 8415
rect 46848 8372 46900 8381
rect 47584 8304 47636 8356
rect 15384 8279 15436 8288
rect 15384 8245 15393 8279
rect 15393 8245 15427 8279
rect 15427 8245 15436 8279
rect 15384 8236 15436 8245
rect 16396 8279 16448 8288
rect 16396 8245 16405 8279
rect 16405 8245 16439 8279
rect 16439 8245 16448 8279
rect 16396 8236 16448 8245
rect 27804 8236 27856 8288
rect 32772 8236 32824 8288
rect 34428 8236 34480 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 1400 8032 1452 8084
rect 16580 8075 16632 8084
rect 16580 8041 16589 8075
rect 16589 8041 16623 8075
rect 16623 8041 16632 8075
rect 16580 8032 16632 8041
rect 17132 8032 17184 8084
rect 18696 8032 18748 8084
rect 20352 8032 20404 8084
rect 17868 7964 17920 8016
rect 20812 8032 20864 8084
rect 21824 8032 21876 8084
rect 25228 8075 25280 8084
rect 25228 8041 25237 8075
rect 25237 8041 25271 8075
rect 25271 8041 25280 8075
rect 25228 8032 25280 8041
rect 30380 8075 30432 8084
rect 30380 8041 30389 8075
rect 30389 8041 30423 8075
rect 30423 8041 30432 8075
rect 30380 8032 30432 8041
rect 35256 8032 35308 8084
rect 14832 7896 14884 7948
rect 16028 7939 16080 7948
rect 16028 7905 16037 7939
rect 16037 7905 16071 7939
rect 16071 7905 16080 7939
rect 16028 7896 16080 7905
rect 1308 7828 1360 7880
rect 15384 7828 15436 7880
rect 10692 7760 10744 7812
rect 14372 7760 14424 7812
rect 18420 7939 18472 7948
rect 18420 7905 18429 7939
rect 18429 7905 18463 7939
rect 18463 7905 18472 7939
rect 18420 7896 18472 7905
rect 18512 7939 18564 7948
rect 18512 7905 18521 7939
rect 18521 7905 18555 7939
rect 18555 7905 18564 7939
rect 18512 7896 18564 7905
rect 30656 7964 30708 8016
rect 18604 7828 18656 7880
rect 20720 7896 20772 7948
rect 22008 7896 22060 7948
rect 29000 7939 29052 7948
rect 29000 7905 29009 7939
rect 29009 7905 29043 7939
rect 29043 7905 29052 7939
rect 29000 7896 29052 7905
rect 31116 7896 31168 7948
rect 32680 7896 32732 7948
rect 49240 7896 49292 7948
rect 23848 7828 23900 7880
rect 29828 7828 29880 7880
rect 32220 7871 32272 7880
rect 32220 7837 32229 7871
rect 32229 7837 32263 7871
rect 32263 7837 32272 7871
rect 32220 7828 32272 7837
rect 34428 7828 34480 7880
rect 47032 7828 47084 7880
rect 15108 7735 15160 7744
rect 15108 7701 15117 7735
rect 15117 7701 15151 7735
rect 15151 7701 15160 7735
rect 15108 7692 15160 7701
rect 17776 7692 17828 7744
rect 21272 7760 21324 7812
rect 18604 7692 18656 7744
rect 19432 7735 19484 7744
rect 19432 7701 19441 7735
rect 19441 7701 19475 7735
rect 19475 7701 19484 7735
rect 19432 7692 19484 7701
rect 19800 7735 19852 7744
rect 19800 7701 19809 7735
rect 19809 7701 19843 7735
rect 19843 7701 19852 7735
rect 19800 7692 19852 7701
rect 20904 7692 20956 7744
rect 23296 7692 23348 7744
rect 28356 7760 28408 7812
rect 23664 7735 23716 7744
rect 23664 7701 23673 7735
rect 23673 7701 23707 7735
rect 23707 7701 23716 7735
rect 23664 7692 23716 7701
rect 27804 7692 27856 7744
rect 30748 7735 30800 7744
rect 30748 7701 30757 7735
rect 30757 7701 30791 7735
rect 30791 7701 30800 7735
rect 30748 7692 30800 7701
rect 40592 7760 40644 7812
rect 38660 7692 38712 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 16304 7488 16356 7540
rect 16028 7420 16080 7472
rect 18328 7488 18380 7540
rect 18696 7531 18748 7540
rect 18696 7497 18705 7531
rect 18705 7497 18739 7531
rect 18739 7497 18748 7531
rect 18696 7488 18748 7497
rect 19248 7488 19300 7540
rect 20352 7531 20404 7540
rect 20352 7497 20361 7531
rect 20361 7497 20395 7531
rect 20395 7497 20404 7531
rect 20352 7488 20404 7497
rect 21456 7531 21508 7540
rect 21456 7497 21465 7531
rect 21465 7497 21499 7531
rect 21499 7497 21508 7531
rect 21456 7488 21508 7497
rect 22284 7488 22336 7540
rect 23296 7488 23348 7540
rect 29644 7531 29696 7540
rect 29644 7497 29653 7531
rect 29653 7497 29687 7531
rect 29687 7497 29696 7531
rect 29644 7488 29696 7497
rect 31392 7531 31444 7540
rect 31392 7497 31401 7531
rect 31401 7497 31435 7531
rect 31435 7497 31444 7531
rect 31392 7488 31444 7497
rect 32864 7488 32916 7540
rect 37372 7531 37424 7540
rect 37372 7497 37381 7531
rect 37381 7497 37415 7531
rect 37415 7497 37424 7531
rect 37372 7488 37424 7497
rect 1308 7352 1360 7404
rect 14096 7352 14148 7404
rect 19800 7420 19852 7472
rect 20904 7420 20956 7472
rect 22468 7420 22520 7472
rect 29552 7420 29604 7472
rect 44824 7463 44876 7472
rect 44824 7429 44833 7463
rect 44833 7429 44867 7463
rect 44867 7429 44876 7463
rect 44824 7420 44876 7429
rect 49332 7420 49384 7472
rect 17316 7284 17368 7336
rect 18972 7284 19024 7336
rect 20812 7395 20864 7404
rect 20812 7361 20821 7395
rect 20821 7361 20855 7395
rect 20855 7361 20864 7395
rect 20812 7352 20864 7361
rect 21732 7352 21784 7404
rect 22744 7352 22796 7404
rect 31484 7352 31536 7404
rect 34060 7352 34112 7404
rect 21640 7284 21692 7336
rect 29736 7284 29788 7336
rect 46940 7352 46992 7404
rect 38660 7284 38712 7336
rect 47032 7284 47084 7336
rect 19524 7216 19576 7268
rect 15108 7148 15160 7200
rect 16396 7148 16448 7200
rect 18696 7148 18748 7200
rect 37924 7191 37976 7200
rect 37924 7157 37933 7191
rect 37933 7157 37967 7191
rect 37967 7157 37976 7191
rect 37924 7148 37976 7157
rect 47216 7216 47268 7268
rect 45744 7148 45796 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 18696 6944 18748 6996
rect 20352 6944 20404 6996
rect 31116 6944 31168 6996
rect 37924 6876 37976 6928
rect 47124 6876 47176 6928
rect 17408 6808 17460 6860
rect 19708 6808 19760 6860
rect 21364 6808 21416 6860
rect 30012 6808 30064 6860
rect 49148 6851 49200 6860
rect 49148 6817 49157 6851
rect 49157 6817 49191 6851
rect 49191 6817 49200 6851
rect 49148 6808 49200 6817
rect 1308 6740 1360 6792
rect 1216 6672 1268 6724
rect 19064 6740 19116 6792
rect 20076 6740 20128 6792
rect 21180 6740 21232 6792
rect 30472 6740 30524 6792
rect 40592 6740 40644 6792
rect 47676 6740 47728 6792
rect 27804 6672 27856 6724
rect 48872 6672 48924 6724
rect 2412 6604 2464 6656
rect 16396 6647 16448 6656
rect 16396 6613 16405 6647
rect 16405 6613 16439 6647
rect 16439 6613 16448 6647
rect 16396 6604 16448 6613
rect 17776 6647 17828 6656
rect 17776 6613 17785 6647
rect 17785 6613 17819 6647
rect 17819 6613 17828 6647
rect 17776 6604 17828 6613
rect 18880 6604 18932 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 1216 6400 1268 6452
rect 18696 6443 18748 6452
rect 18696 6409 18705 6443
rect 18705 6409 18739 6443
rect 18739 6409 18748 6443
rect 18696 6400 18748 6409
rect 19616 6400 19668 6452
rect 34152 6332 34204 6384
rect 41420 6332 41472 6384
rect 49332 6332 49384 6384
rect 1308 6264 1360 6316
rect 17868 6264 17920 6316
rect 18788 6264 18840 6316
rect 19432 6264 19484 6316
rect 42708 6264 42760 6316
rect 28448 6196 28500 6248
rect 36912 6196 36964 6248
rect 10048 6128 10100 6180
rect 21180 6128 21232 6180
rect 26056 6128 26108 6180
rect 35808 6128 35860 6180
rect 46940 6128 46992 6180
rect 22744 6060 22796 6112
rect 37648 6103 37700 6112
rect 37648 6069 37657 6103
rect 37657 6069 37691 6103
rect 37691 6069 37700 6103
rect 37648 6060 37700 6069
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 37648 5856 37700 5908
rect 47308 5856 47360 5908
rect 13452 5788 13504 5840
rect 1308 5652 1360 5704
rect 49240 5720 49292 5772
rect 2780 5652 2832 5704
rect 40040 5652 40092 5704
rect 47584 5652 47636 5704
rect 15476 5584 15528 5636
rect 45836 5584 45888 5636
rect 19340 5516 19392 5568
rect 24032 5516 24084 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 37280 5312 37332 5364
rect 31300 5244 31352 5296
rect 49148 5287 49200 5296
rect 49148 5253 49157 5287
rect 49157 5253 49191 5287
rect 49191 5253 49200 5287
rect 49148 5244 49200 5253
rect 37280 5176 37332 5228
rect 45744 5176 45796 5228
rect 47216 5176 47268 5228
rect 1308 5108 1360 5160
rect 10784 5108 10836 5160
rect 48320 5108 48372 5160
rect 40040 5040 40092 5092
rect 37924 5015 37976 5024
rect 37924 4981 37933 5015
rect 37933 4981 37967 5015
rect 37967 4981 37976 5015
rect 37924 4972 37976 4981
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 1308 4768 1360 4820
rect 5540 4768 5592 4820
rect 22376 4768 22428 4820
rect 36912 4811 36964 4820
rect 36912 4777 36921 4811
rect 36921 4777 36955 4811
rect 36955 4777 36964 4811
rect 36912 4768 36964 4777
rect 37924 4768 37976 4820
rect 47216 4768 47268 4820
rect 31668 4700 31720 4752
rect 26240 4675 26292 4684
rect 26240 4641 26249 4675
rect 26249 4641 26283 4675
rect 26283 4641 26292 4675
rect 26240 4632 26292 4641
rect 49424 4632 49476 4684
rect 1308 4564 1360 4616
rect 22468 4564 22520 4616
rect 22652 4564 22704 4616
rect 23296 4564 23348 4616
rect 27068 4564 27120 4616
rect 47032 4564 47084 4616
rect 23572 4496 23624 4548
rect 36912 4496 36964 4548
rect 19340 4428 19392 4480
rect 24032 4428 24084 4480
rect 24768 4428 24820 4480
rect 39396 4428 39448 4480
rect 44456 4428 44508 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 1400 4156 1452 4208
rect 23664 4224 23716 4276
rect 24768 4224 24820 4276
rect 1308 4088 1360 4140
rect 24032 4156 24084 4208
rect 27344 4199 27396 4208
rect 27344 4165 27353 4199
rect 27353 4165 27387 4199
rect 27387 4165 27396 4199
rect 27344 4156 27396 4165
rect 16488 4088 16540 4140
rect 27160 4131 27212 4140
rect 27160 4097 27169 4131
rect 27169 4097 27203 4131
rect 27203 4097 27212 4131
rect 27160 4088 27212 4097
rect 34244 4088 34296 4140
rect 39212 4088 39264 4140
rect 39304 4088 39356 4140
rect 47124 4088 47176 4140
rect 49332 4088 49384 4140
rect 17776 4020 17828 4072
rect 16488 3952 16540 4004
rect 20168 4063 20220 4072
rect 20168 4029 20177 4063
rect 20177 4029 20211 4063
rect 20211 4029 20220 4063
rect 20168 4020 20220 4029
rect 22008 4063 22060 4072
rect 22008 4029 22017 4063
rect 22017 4029 22051 4063
rect 22051 4029 22060 4063
rect 22008 4020 22060 4029
rect 22284 4063 22336 4072
rect 22284 4029 22293 4063
rect 22293 4029 22327 4063
rect 22327 4029 22336 4063
rect 22284 4020 22336 4029
rect 5540 3884 5592 3936
rect 7472 3884 7524 3936
rect 20720 3884 20772 3936
rect 22468 3884 22520 3936
rect 23664 3884 23716 3936
rect 24492 4020 24544 4072
rect 25688 4063 25740 4072
rect 25688 4029 25697 4063
rect 25697 4029 25731 4063
rect 25731 4029 25740 4063
rect 25688 4020 25740 4029
rect 24400 3952 24452 4004
rect 46664 4063 46716 4072
rect 46664 4029 46673 4063
rect 46673 4029 46707 4063
rect 46707 4029 46716 4063
rect 46664 4020 46716 4029
rect 27160 3952 27212 4004
rect 33600 3952 33652 4004
rect 30656 3884 30708 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 5356 3680 5408 3732
rect 15384 3612 15436 3664
rect 1124 3544 1176 3596
rect 17224 3544 17276 3596
rect 1308 3476 1360 3528
rect 7564 3476 7616 3528
rect 16488 3519 16540 3528
rect 16488 3485 16497 3519
rect 16497 3485 16531 3519
rect 16531 3485 16540 3519
rect 16488 3476 16540 3485
rect 22284 3680 22336 3732
rect 27344 3680 27396 3732
rect 39304 3680 39356 3732
rect 20720 3612 20772 3664
rect 21916 3612 21968 3664
rect 19800 3544 19852 3596
rect 21180 3587 21232 3596
rect 21180 3553 21189 3587
rect 21189 3553 21223 3587
rect 21223 3553 21232 3587
rect 21180 3544 21232 3553
rect 22100 3544 22152 3596
rect 23296 3544 23348 3596
rect 23572 3544 23624 3596
rect 37004 3612 37056 3664
rect 45560 3612 45612 3664
rect 34520 3544 34572 3596
rect 47676 3544 47728 3596
rect 49148 3587 49200 3596
rect 49148 3553 49157 3587
rect 49157 3553 49191 3587
rect 49191 3553 49200 3587
rect 49148 3544 49200 3553
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 22928 3476 22980 3528
rect 12532 3340 12584 3392
rect 24400 3408 24452 3460
rect 24492 3340 24544 3392
rect 35808 3476 35860 3528
rect 40040 3476 40092 3528
rect 46940 3476 46992 3528
rect 40868 3408 40920 3460
rect 43444 3408 43496 3460
rect 48688 3408 48740 3460
rect 25872 3340 25924 3392
rect 40960 3340 41012 3392
rect 49792 3340 49844 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 1308 3136 1360 3188
rect 17224 3136 17276 3188
rect 24216 3136 24268 3188
rect 16120 3068 16172 3120
rect 1308 3000 1360 3052
rect 14280 3000 14332 3052
rect 16396 3000 16448 3052
rect 11060 2932 11112 2984
rect 11244 2864 11296 2916
rect 22100 3068 22152 3120
rect 22928 3111 22980 3120
rect 22928 3077 22937 3111
rect 22937 3077 22971 3111
rect 22971 3077 22980 3111
rect 22928 3068 22980 3077
rect 23664 3068 23716 3120
rect 19524 3000 19576 3052
rect 22744 3043 22796 3052
rect 22744 3009 22753 3043
rect 22753 3009 22787 3043
rect 22787 3009 22796 3043
rect 22744 3000 22796 3009
rect 27712 3068 27764 3120
rect 30748 3136 30800 3188
rect 49240 3068 49292 3120
rect 27620 3000 27672 3052
rect 29092 3043 29144 3052
rect 29092 3009 29101 3043
rect 29101 3009 29135 3043
rect 29135 3009 29144 3043
rect 29092 3000 29144 3009
rect 39396 3000 39448 3052
rect 45836 3043 45888 3052
rect 45836 3009 45845 3043
rect 45845 3009 45879 3043
rect 45879 3009 45888 3043
rect 45836 3000 45888 3009
rect 47308 3000 47360 3052
rect 19800 2975 19852 2984
rect 19800 2941 19809 2975
rect 19809 2941 19843 2975
rect 19843 2941 19852 2975
rect 19800 2932 19852 2941
rect 22284 2932 22336 2984
rect 26516 2932 26568 2984
rect 46756 2932 46808 2984
rect 46848 2975 46900 2984
rect 46848 2941 46857 2975
rect 46857 2941 46891 2975
rect 46891 2941 46900 2975
rect 46848 2932 46900 2941
rect 22652 2864 22704 2916
rect 23388 2864 23440 2916
rect 2320 2839 2372 2848
rect 2320 2805 2329 2839
rect 2329 2805 2363 2839
rect 2363 2805 2372 2839
rect 2320 2796 2372 2805
rect 2780 2839 2832 2848
rect 2780 2805 2789 2839
rect 2789 2805 2823 2839
rect 2823 2805 2832 2839
rect 2780 2796 2832 2805
rect 3332 2796 3384 2848
rect 8852 2796 8904 2848
rect 19432 2796 19484 2848
rect 20996 2796 21048 2848
rect 24860 2796 24912 2848
rect 30840 2839 30892 2848
rect 30840 2805 30849 2839
rect 30849 2805 30883 2839
rect 30883 2805 30892 2839
rect 30840 2796 30892 2805
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 9496 2592 9548 2644
rect 11060 2592 11112 2644
rect 16396 2635 16448 2644
rect 16396 2601 16405 2635
rect 16405 2601 16439 2635
rect 16439 2601 16448 2635
rect 16396 2592 16448 2601
rect 20996 2635 21048 2644
rect 20996 2601 21005 2635
rect 21005 2601 21039 2635
rect 21039 2601 21048 2635
rect 20996 2592 21048 2601
rect 23664 2592 23716 2644
rect 27620 2592 27672 2644
rect 1308 2388 1360 2440
rect 2780 2456 2832 2508
rect 20904 2524 20956 2576
rect 11704 2456 11756 2508
rect 13820 2456 13872 2508
rect 22836 2524 22888 2576
rect 23296 2524 23348 2576
rect 23388 2524 23440 2576
rect 25872 2524 25924 2576
rect 27436 2524 27488 2576
rect 2320 2431 2372 2440
rect 1216 2320 1268 2372
rect 2320 2397 2329 2431
rect 2329 2397 2363 2431
rect 2363 2397 2372 2431
rect 2320 2388 2372 2397
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 9680 2388 9732 2440
rect 12532 2388 12584 2440
rect 15384 2388 15436 2440
rect 22008 2456 22060 2508
rect 24860 2499 24912 2508
rect 24860 2465 24869 2499
rect 24869 2465 24903 2499
rect 24903 2465 24912 2499
rect 24860 2456 24912 2465
rect 24952 2456 25004 2508
rect 27712 2524 27764 2576
rect 31668 2592 31720 2644
rect 33600 2592 33652 2644
rect 30840 2524 30892 2576
rect 10600 2320 10652 2372
rect 9496 2252 9548 2304
rect 12348 2252 12400 2304
rect 18328 2320 18380 2372
rect 24860 2320 24912 2372
rect 28632 2388 28684 2440
rect 30748 2388 30800 2440
rect 33140 2431 33192 2440
rect 33140 2397 33149 2431
rect 33149 2397 33183 2431
rect 33183 2397 33192 2431
rect 33140 2388 33192 2397
rect 34980 2388 35032 2440
rect 41328 2456 41380 2508
rect 49148 2499 49200 2508
rect 49148 2465 49157 2499
rect 49157 2465 49191 2499
rect 49191 2465 49200 2499
rect 49148 2456 49200 2465
rect 27436 2320 27488 2372
rect 27160 2252 27212 2304
rect 44456 2388 44508 2440
rect 47216 2388 47268 2440
rect 48504 2320 48556 2372
rect 30656 2252 30708 2304
rect 37096 2295 37148 2304
rect 37096 2261 37105 2295
rect 37105 2261 37139 2295
rect 37139 2261 37148 2295
rect 37096 2252 37148 2261
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
rect 1308 2048 1360 2100
rect 3240 2048 3292 2100
rect 22468 2048 22520 2100
rect 27160 2048 27212 2100
<< metal2 >>
rect 1582 26200 1638 27000
rect 2226 26200 2282 27000
rect 2870 26200 2926 27000
rect 3514 26200 3570 27000
rect 4158 26200 4214 27000
rect 4802 26330 4858 27000
rect 4802 26302 5120 26330
rect 4802 26200 4858 26302
rect 1596 22234 1624 26200
rect 2136 24608 2188 24614
rect 2136 24550 2188 24556
rect 1860 23860 1912 23866
rect 1860 23802 1912 23808
rect 1872 22642 1900 23802
rect 2148 23798 2176 24550
rect 2136 23792 2188 23798
rect 2136 23734 2188 23740
rect 1860 22636 1912 22642
rect 1860 22578 1912 22584
rect 1584 22228 1636 22234
rect 1584 22170 1636 22176
rect 2240 22166 2268 26200
rect 2778 24440 2834 24449
rect 2778 24375 2780 24384
rect 2832 24375 2834 24384
rect 2780 24346 2832 24352
rect 2320 24200 2372 24206
rect 2320 24142 2372 24148
rect 2228 22160 2280 22166
rect 2228 22102 2280 22108
rect 1308 22092 1360 22098
rect 1308 22034 1360 22040
rect 1320 20777 1348 22034
rect 1768 22024 1820 22030
rect 1768 21966 1820 21972
rect 1780 21622 1808 21966
rect 1768 21616 1820 21622
rect 1768 21558 1820 21564
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1306 20768 1362 20777
rect 1306 20703 1362 20712
rect 1412 19961 1440 21422
rect 1860 20460 1912 20466
rect 1860 20402 1912 20408
rect 1398 19952 1454 19961
rect 1398 19887 1454 19896
rect 1766 19952 1822 19961
rect 1766 19887 1822 19896
rect 1780 19854 1808 19887
rect 1768 19848 1820 19854
rect 1872 19825 1900 20402
rect 1768 19790 1820 19796
rect 1858 19816 1914 19825
rect 1858 19751 1914 19760
rect 2332 19174 2360 24142
rect 2780 23044 2832 23050
rect 2780 22986 2832 22992
rect 2792 22250 2820 22986
rect 2884 22710 2912 26200
rect 3054 25664 3110 25673
rect 3054 25599 3110 25608
rect 3068 24886 3096 25599
rect 3056 24880 3108 24886
rect 3056 24822 3108 24828
rect 3422 24848 3478 24857
rect 3422 24783 3424 24792
rect 3476 24783 3478 24792
rect 3424 24754 3476 24760
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 3528 24274 3556 26200
rect 3606 25256 3662 25265
rect 3606 25191 3662 25200
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3514 24032 3570 24041
rect 3514 23967 3570 23976
rect 3332 23724 3384 23730
rect 3332 23666 3384 23672
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 3146 22808 3202 22817
rect 3146 22743 3148 22752
rect 3200 22743 3202 22752
rect 3148 22714 3200 22720
rect 2872 22704 2924 22710
rect 2872 22646 2924 22652
rect 2872 22568 2924 22574
rect 2872 22510 2924 22516
rect 2700 22222 2820 22250
rect 2700 21593 2728 22222
rect 2686 21584 2742 21593
rect 2686 21519 2742 21528
rect 2778 21176 2834 21185
rect 2884 21162 2912 22510
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2834 21134 2912 21162
rect 2778 21111 2834 21120
rect 2780 20868 2832 20874
rect 2780 20810 2832 20816
rect 2792 19938 2820 20810
rect 2872 20392 2924 20398
rect 2872 20334 2924 20340
rect 2700 19910 2820 19938
rect 2700 19553 2728 19910
rect 2780 19780 2832 19786
rect 2780 19722 2832 19728
rect 2686 19544 2742 19553
rect 2686 19479 2742 19488
rect 2320 19168 2372 19174
rect 2320 19110 2372 19116
rect 2792 18873 2820 19722
rect 2884 19530 2912 20334
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2884 19502 3004 19530
rect 2872 19372 2924 19378
rect 2872 19314 2924 19320
rect 2778 18864 2834 18873
rect 2778 18799 2834 18808
rect 2780 18692 2832 18698
rect 2780 18634 2832 18640
rect 2792 18306 2820 18634
rect 2884 18329 2912 19314
rect 2976 19281 3004 19502
rect 2962 19272 3018 19281
rect 2962 19207 3018 19216
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 2700 18278 2820 18306
rect 2870 18320 2926 18329
rect 1780 17814 1808 18226
rect 2700 17921 2728 18278
rect 2870 18255 2926 18264
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 2686 17912 2742 17921
rect 2686 17847 2742 17856
rect 1768 17808 1820 17814
rect 1768 17750 1820 17756
rect 1216 17740 1268 17746
rect 1216 17682 1268 17688
rect 1228 17105 1256 17682
rect 2792 17513 2820 18158
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 3344 17746 3372 23666
rect 3422 23624 3478 23633
rect 3422 23559 3478 23568
rect 3436 23526 3464 23559
rect 3424 23520 3476 23526
rect 3424 23462 3476 23468
rect 3422 23216 3478 23225
rect 3422 23151 3478 23160
rect 3436 22506 3464 23151
rect 3424 22500 3476 22506
rect 3424 22442 3476 22448
rect 3424 21548 3476 21554
rect 3424 21490 3476 21496
rect 3436 21146 3464 21490
rect 3424 21140 3476 21146
rect 3424 21082 3476 21088
rect 3528 18834 3556 23967
rect 3620 21350 3648 25191
rect 3882 24848 3938 24857
rect 3882 24783 3938 24792
rect 3896 22642 3924 24783
rect 3976 24064 4028 24070
rect 3976 24006 4028 24012
rect 3988 23798 4016 24006
rect 3976 23792 4028 23798
rect 3976 23734 4028 23740
rect 4172 23662 4200 26200
rect 4896 24200 4948 24206
rect 4896 24142 4948 24148
rect 4804 23724 4856 23730
rect 4804 23666 4856 23672
rect 4160 23656 4212 23662
rect 4160 23598 4212 23604
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 4436 23112 4488 23118
rect 4436 23054 4488 23060
rect 3884 22636 3936 22642
rect 3884 22578 3936 22584
rect 3988 22273 4016 23054
rect 4344 23044 4396 23050
rect 4344 22986 4396 22992
rect 4252 22704 4304 22710
rect 4252 22646 4304 22652
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 3974 22264 4030 22273
rect 3974 22199 4030 22208
rect 3792 22092 3844 22098
rect 3792 22034 3844 22040
rect 3804 22001 3832 22034
rect 3790 21992 3846 22001
rect 3790 21927 3846 21936
rect 3976 21616 4028 21622
rect 3976 21558 4028 21564
rect 3608 21344 3660 21350
rect 3608 21286 3660 21292
rect 3988 21078 4016 21558
rect 3976 21072 4028 21078
rect 3976 21014 4028 21020
rect 3608 20460 3660 20466
rect 3608 20402 3660 20408
rect 3620 20058 3648 20402
rect 3884 20392 3936 20398
rect 3882 20360 3884 20369
rect 3936 20360 3938 20369
rect 3882 20295 3938 20304
rect 3608 20052 3660 20058
rect 3608 19994 3660 20000
rect 3516 18828 3568 18834
rect 3516 18770 3568 18776
rect 4080 18358 4108 22578
rect 4160 22568 4212 22574
rect 4158 22536 4160 22545
rect 4212 22536 4214 22545
rect 4158 22471 4214 22480
rect 4158 22128 4214 22137
rect 4158 22063 4214 22072
rect 4172 21010 4200 22063
rect 4264 21622 4292 22646
rect 4252 21616 4304 21622
rect 4252 21558 4304 21564
rect 4356 21486 4384 22986
rect 4344 21480 4396 21486
rect 4344 21422 4396 21428
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 4252 19780 4304 19786
rect 4252 19722 4304 19728
rect 4264 18766 4292 19722
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 4068 18352 4120 18358
rect 4068 18294 4120 18300
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 3332 17740 3384 17746
rect 3332 17682 3384 17688
rect 2778 17504 2834 17513
rect 2778 17439 2834 17448
rect 1308 17128 1360 17134
rect 1214 17096 1270 17105
rect 1308 17070 1360 17076
rect 1214 17031 1270 17040
rect 1320 16697 1348 17070
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 1306 16688 1362 16697
rect 1306 16623 1362 16632
rect 1308 16516 1360 16522
rect 1308 16458 1360 16464
rect 1320 16289 1348 16458
rect 1306 16280 1362 16289
rect 1306 16215 1362 16224
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 1320 15881 1348 15982
rect 1306 15872 1362 15881
rect 1306 15807 1362 15816
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 3528 15706 3556 18226
rect 4344 17672 4396 17678
rect 4344 17614 4396 17620
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4172 16590 4200 16934
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 3976 16448 4028 16454
rect 3976 16390 4028 16396
rect 3988 16250 4016 16390
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 4080 16182 4108 16526
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 4356 16046 4384 17614
rect 4448 17338 4476 23054
rect 4620 22228 4672 22234
rect 4620 22170 4672 22176
rect 4528 22160 4580 22166
rect 4528 22102 4580 22108
rect 4540 19922 4568 22102
rect 4528 19916 4580 19922
rect 4528 19858 4580 19864
rect 4632 19446 4660 22170
rect 4620 19440 4672 19446
rect 4620 19382 4672 19388
rect 4710 18320 4766 18329
rect 4710 18255 4712 18264
rect 4764 18255 4766 18264
rect 4712 18226 4764 18232
rect 4816 17338 4844 23666
rect 4908 17678 4936 24142
rect 5092 22574 5120 26302
rect 5446 26200 5502 27000
rect 6090 26200 6146 27000
rect 6734 26330 6790 27000
rect 6472 26302 6790 26330
rect 5264 24200 5316 24206
rect 5264 24142 5316 24148
rect 5276 23186 5304 24142
rect 5460 23662 5488 26200
rect 5908 24132 5960 24138
rect 5908 24074 5960 24080
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5264 23180 5316 23186
rect 5264 23122 5316 23128
rect 5816 22636 5868 22642
rect 5816 22578 5868 22584
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 5632 22500 5684 22506
rect 5632 22442 5684 22448
rect 5356 21616 5408 21622
rect 5356 21558 5408 21564
rect 5080 21548 5132 21554
rect 5080 21490 5132 21496
rect 5172 21548 5224 21554
rect 5172 21490 5224 21496
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 4436 17332 4488 17338
rect 4436 17274 4488 17280
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 5000 17202 5028 17478
rect 5092 17338 5120 21490
rect 5184 18154 5212 21490
rect 5264 19984 5316 19990
rect 5264 19926 5316 19932
rect 5276 19378 5304 19926
rect 5264 19372 5316 19378
rect 5264 19314 5316 19320
rect 5264 19236 5316 19242
rect 5264 19178 5316 19184
rect 5276 18630 5304 19178
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5172 18148 5224 18154
rect 5172 18090 5224 18096
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 4804 16584 4856 16590
rect 4802 16552 4804 16561
rect 4856 16552 4858 16561
rect 4802 16487 4858 16496
rect 4344 16040 4396 16046
rect 4344 15982 4396 15988
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 1308 15564 1360 15570
rect 1308 15506 1360 15512
rect 1320 15473 1348 15506
rect 1306 15464 1362 15473
rect 1306 15399 1362 15408
rect 1306 15056 1362 15065
rect 1306 14991 1362 15000
rect 1320 14958 1348 14991
rect 1308 14952 1360 14958
rect 1308 14894 1360 14900
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 1306 14648 1362 14657
rect 2950 14651 3258 14660
rect 1306 14583 1362 14592
rect 1320 14482 1348 14583
rect 1308 14476 1360 14482
rect 1308 14418 1360 14424
rect 938 14240 994 14249
rect 938 14175 994 14184
rect 952 13870 980 14175
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 940 13864 992 13870
rect 940 13806 992 13812
rect 2778 13832 2834 13841
rect 2778 13767 2834 13776
rect 1766 13424 1822 13433
rect 2792 13394 2820 13767
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 1766 13359 1822 13368
rect 2780 13388 2832 13394
rect 1780 13326 1808 13359
rect 2780 13330 2832 13336
rect 1768 13320 1820 13326
rect 3528 13297 3556 13874
rect 1768 13262 1820 13268
rect 3514 13288 3570 13297
rect 3514 13223 3570 13232
rect 1214 13016 1270 13025
rect 1214 12951 1270 12960
rect 1228 12782 1256 12951
rect 1308 12844 1360 12850
rect 1308 12786 1360 12792
rect 1216 12776 1268 12782
rect 1216 12718 1268 12724
rect 1320 12617 1348 12786
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 1306 12608 1362 12617
rect 1306 12543 1362 12552
rect 2792 12442 2820 12650
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 1308 12232 1360 12238
rect 1214 12200 1270 12209
rect 1308 12174 1360 12180
rect 1214 12135 1270 12144
rect 1228 11762 1256 12135
rect 1320 11801 1348 12174
rect 1306 11792 1362 11801
rect 1216 11756 1268 11762
rect 1306 11727 1362 11736
rect 1216 11698 1268 11704
rect 1228 11354 1256 11698
rect 1308 11688 1360 11694
rect 1308 11630 1360 11636
rect 1320 11393 1348 11630
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 1306 11384 1362 11393
rect 2950 11387 3258 11396
rect 1216 11348 1268 11354
rect 1306 11319 1362 11328
rect 1216 11290 1268 11296
rect 1768 11280 1820 11286
rect 1768 11222 1820 11228
rect 1584 11144 1636 11150
rect 1780 11121 1808 11222
rect 1584 11086 1636 11092
rect 1766 11112 1822 11121
rect 1596 10985 1624 11086
rect 1766 11047 1822 11056
rect 1582 10976 1638 10985
rect 1582 10911 1638 10920
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 1216 10736 1268 10742
rect 1216 10678 1268 10684
rect 1228 10169 1256 10678
rect 1308 10668 1360 10674
rect 1308 10610 1360 10616
rect 1320 10577 1348 10610
rect 1306 10568 1362 10577
rect 1306 10503 1362 10512
rect 1214 10160 1270 10169
rect 1872 10130 1900 10746
rect 2502 10568 2558 10577
rect 2502 10503 2558 10512
rect 2516 10470 2544 10503
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 1214 10095 1270 10104
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1308 10056 1360 10062
rect 1308 9998 1360 10004
rect 1320 9761 1348 9998
rect 1306 9752 1362 9761
rect 1306 9687 1308 9696
rect 1360 9687 1362 9696
rect 1308 9658 1360 9664
rect 1308 9580 1360 9586
rect 1308 9522 1360 9528
rect 1320 9353 1348 9522
rect 1860 9512 1912 9518
rect 1858 9480 1860 9489
rect 1912 9480 1914 9489
rect 1858 9415 1914 9424
rect 1306 9344 1362 9353
rect 1306 9279 1362 9288
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 1216 8968 1268 8974
rect 1216 8910 1268 8916
rect 1306 8936 1362 8945
rect 1228 8537 1256 8910
rect 1306 8871 1308 8880
rect 1360 8871 1362 8880
rect 1308 8842 1360 8848
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1780 8566 1808 8774
rect 1768 8560 1820 8566
rect 1214 8528 1270 8537
rect 1768 8502 1820 8508
rect 1214 8463 1270 8472
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 8129 1440 8366
rect 1398 8120 1454 8129
rect 1398 8055 1400 8064
rect 1452 8055 1454 8064
rect 1400 8026 1452 8032
rect 1308 7880 1360 7886
rect 1308 7822 1360 7828
rect 1320 7721 1348 7822
rect 1306 7712 1362 7721
rect 1306 7647 1362 7656
rect 1308 7404 1360 7410
rect 1308 7346 1360 7352
rect 1320 7313 1348 7346
rect 1306 7304 1362 7313
rect 1306 7239 1362 7248
rect 1214 6896 1270 6905
rect 1214 6831 1270 6840
rect 1228 6730 1256 6831
rect 1308 6792 1360 6798
rect 1308 6734 1360 6740
rect 1216 6724 1268 6730
rect 1216 6666 1268 6672
rect 1228 6458 1256 6666
rect 1320 6497 1348 6734
rect 2424 6662 2452 8978
rect 2502 8936 2558 8945
rect 2502 8871 2558 8880
rect 2516 8838 2544 8871
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 4080 8498 4108 13874
rect 4356 11898 4384 15982
rect 5276 12306 5304 18566
rect 5368 16454 5396 21558
rect 5446 21448 5502 21457
rect 5446 21383 5448 21392
rect 5500 21383 5502 21392
rect 5448 21354 5500 21360
rect 5644 21010 5672 22442
rect 5724 22432 5776 22438
rect 5724 22374 5776 22380
rect 5632 21004 5684 21010
rect 5632 20946 5684 20952
rect 5736 19854 5764 22374
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5644 16726 5672 17138
rect 5828 16794 5856 22578
rect 5920 22094 5948 24074
rect 6104 23186 6132 26200
rect 6184 24404 6236 24410
rect 6184 24346 6236 24352
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 5920 22066 6132 22094
rect 5908 20460 5960 20466
rect 5908 20402 5960 20408
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5460 14550 5488 16050
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 5644 12986 5672 16662
rect 5920 16250 5948 20402
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 6012 18970 6040 19790
rect 6104 19446 6132 22066
rect 6196 19922 6224 24346
rect 6472 24274 6500 26302
rect 6734 26200 6790 26302
rect 7378 26330 7434 27000
rect 7378 26302 7696 26330
rect 7378 26200 7434 26302
rect 7196 24812 7248 24818
rect 7196 24754 7248 24760
rect 6460 24268 6512 24274
rect 6460 24210 6512 24216
rect 6828 23724 6880 23730
rect 6828 23666 6880 23672
rect 6644 23520 6696 23526
rect 6644 23462 6696 23468
rect 6656 21486 6684 23462
rect 6840 23322 6868 23666
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 6840 22778 6868 23258
rect 7104 23112 7156 23118
rect 7104 23054 7156 23060
rect 6736 22772 6788 22778
rect 6736 22714 6788 22720
rect 6828 22772 6880 22778
rect 6828 22714 6880 22720
rect 6748 22098 6776 22714
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 6736 22092 6788 22098
rect 6736 22034 6788 22040
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6460 21140 6512 21146
rect 6460 21082 6512 21088
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6276 19508 6328 19514
rect 6276 19450 6328 19456
rect 6092 19440 6144 19446
rect 6092 19382 6144 19388
rect 6184 19168 6236 19174
rect 6184 19110 6236 19116
rect 6000 18964 6052 18970
rect 6000 18906 6052 18912
rect 6090 18864 6146 18873
rect 6196 18834 6224 19110
rect 6090 18799 6146 18808
rect 6184 18828 6236 18834
rect 6104 18154 6132 18799
rect 6184 18770 6236 18776
rect 6092 18148 6144 18154
rect 6092 18090 6144 18096
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 6288 15910 6316 19450
rect 6380 18358 6408 19858
rect 6472 18358 6500 21082
rect 6826 19408 6882 19417
rect 6826 19343 6882 19352
rect 6840 19310 6868 19343
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6552 19168 6604 19174
rect 6644 19168 6696 19174
rect 6552 19110 6604 19116
rect 6642 19136 6644 19145
rect 6696 19136 6698 19145
rect 6564 19009 6592 19110
rect 6642 19071 6698 19080
rect 6550 19000 6606 19009
rect 6550 18935 6606 18944
rect 6644 18896 6696 18902
rect 6644 18838 6696 18844
rect 6552 18624 6604 18630
rect 6552 18566 6604 18572
rect 6368 18352 6420 18358
rect 6368 18294 6420 18300
rect 6460 18352 6512 18358
rect 6460 18294 6512 18300
rect 6460 18080 6512 18086
rect 6460 18022 6512 18028
rect 6472 16590 6500 18022
rect 6564 17202 6592 18566
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6656 17134 6684 18838
rect 6644 17128 6696 17134
rect 6644 17070 6696 17076
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 6380 16250 6408 16526
rect 6932 16454 6960 22578
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 7024 19310 7052 20878
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 7024 17746 7052 18022
rect 7012 17740 7064 17746
rect 7012 17682 7064 17688
rect 7116 17202 7144 23054
rect 7208 20398 7236 24754
rect 7378 24304 7434 24313
rect 7378 24239 7434 24248
rect 7392 24206 7420 24239
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 7668 22574 7696 26302
rect 8022 26200 8078 27000
rect 8666 26200 8722 27000
rect 9310 26200 9366 27000
rect 9954 26200 10010 27000
rect 10598 26330 10654 27000
rect 10598 26302 10732 26330
rect 10598 26200 10654 26302
rect 8036 24698 8064 26200
rect 7852 24670 8064 24698
rect 7852 23186 7880 24670
rect 8680 24274 8708 26200
rect 8668 24268 8720 24274
rect 8668 24210 8720 24216
rect 8852 24064 8904 24070
rect 8852 24006 8904 24012
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8576 23248 8628 23254
rect 8576 23190 8628 23196
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 8588 22098 8616 23190
rect 8576 22092 8628 22098
rect 8576 22034 8628 22040
rect 7656 22024 7708 22030
rect 7932 22024 7984 22030
rect 7656 21966 7708 21972
rect 7930 21992 7932 22001
rect 7984 21992 7986 22001
rect 7288 21548 7340 21554
rect 7288 21490 7340 21496
rect 7300 20602 7328 21490
rect 7668 21146 7696 21966
rect 7930 21927 7986 21936
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 7748 21616 7800 21622
rect 7748 21558 7800 21564
rect 7656 21140 7708 21146
rect 7656 21082 7708 21088
rect 7288 20596 7340 20602
rect 7288 20538 7340 20544
rect 7196 20392 7248 20398
rect 7196 20334 7248 20340
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 7208 18290 7236 18906
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7288 18420 7340 18426
rect 7288 18362 7340 18368
rect 7300 18329 7328 18362
rect 7286 18320 7342 18329
rect 7196 18284 7248 18290
rect 7286 18255 7342 18264
rect 7196 18226 7248 18232
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6656 15026 6684 15302
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6932 13326 6960 15370
rect 7392 13870 7420 18702
rect 7668 15434 7696 19654
rect 7760 19378 7788 21558
rect 7840 21480 7892 21486
rect 7838 21448 7840 21457
rect 7892 21448 7894 21457
rect 7838 21383 7894 21392
rect 7852 20942 7880 21383
rect 8024 21072 8076 21078
rect 8024 21014 8076 21020
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 8036 20806 8064 21014
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8024 20800 8076 20806
rect 8024 20742 8076 20748
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 7838 20496 7894 20505
rect 7838 20431 7894 20440
rect 7852 19854 7880 20431
rect 8312 20398 8340 20946
rect 8864 20466 8892 24006
rect 9324 23798 9352 26200
rect 9864 24880 9916 24886
rect 9864 24822 9916 24828
rect 9680 24200 9732 24206
rect 9680 24142 9732 24148
rect 9312 23792 9364 23798
rect 9312 23734 9364 23740
rect 9128 23656 9180 23662
rect 9128 23598 9180 23604
rect 9140 22030 9168 23598
rect 9692 23594 9720 24142
rect 9680 23588 9732 23594
rect 9680 23530 9732 23536
rect 9402 23216 9458 23225
rect 9402 23151 9404 23160
rect 9456 23151 9458 23160
rect 9404 23122 9456 23128
rect 9220 23112 9272 23118
rect 9218 23080 9220 23089
rect 9272 23080 9274 23089
rect 9218 23015 9274 23024
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 9232 21690 9260 23015
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9680 22568 9732 22574
rect 9680 22510 9732 22516
rect 9404 22432 9456 22438
rect 9404 22374 9456 22380
rect 9416 22094 9444 22374
rect 9416 22066 9628 22094
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 9220 21684 9272 21690
rect 9220 21626 9272 21632
rect 9034 21584 9090 21593
rect 9034 21519 9090 21528
rect 9048 21078 9076 21519
rect 9036 21072 9088 21078
rect 9036 21014 9088 21020
rect 8852 20460 8904 20466
rect 8852 20402 8904 20408
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 7932 19848 7984 19854
rect 7932 19790 7984 19796
rect 7944 19700 7972 19790
rect 7852 19672 7972 19700
rect 7748 19372 7800 19378
rect 7748 19314 7800 19320
rect 7852 19242 7880 19672
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 7944 19378 7972 19450
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 8760 19372 8812 19378
rect 8760 19314 8812 19320
rect 7944 19242 7972 19314
rect 7840 19236 7892 19242
rect 7840 19178 7892 19184
rect 7932 19236 7984 19242
rect 7932 19178 7984 19184
rect 7748 18896 7800 18902
rect 7748 18838 7800 18844
rect 7760 18358 7788 18838
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 8484 18692 8536 18698
rect 8484 18634 8536 18640
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 7748 18352 7800 18358
rect 7748 18294 7800 18300
rect 8312 18170 8340 18634
rect 8496 18306 8524 18634
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 8680 18358 8708 18566
rect 8668 18352 8720 18358
rect 8496 18278 8616 18306
rect 8668 18294 8720 18300
rect 8312 18142 8432 18170
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8312 17338 8340 18022
rect 8404 17882 8432 18142
rect 8588 18086 8616 18278
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8484 17808 8536 17814
rect 8484 17750 8536 17756
rect 8574 17776 8630 17785
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8024 16992 8076 16998
rect 8024 16934 8076 16940
rect 8036 16590 8064 16934
rect 8496 16726 8524 17750
rect 8574 17711 8630 17720
rect 8588 17678 8616 17711
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8588 16794 8616 17614
rect 8680 16794 8708 18294
rect 8772 17338 8800 19314
rect 8864 17814 8892 20402
rect 8944 19236 8996 19242
rect 8944 19178 8996 19184
rect 8852 17808 8904 17814
rect 8852 17750 8904 17756
rect 8760 17332 8812 17338
rect 8760 17274 8812 17280
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8484 16720 8536 16726
rect 8484 16662 8536 16668
rect 8956 16658 8984 19178
rect 9140 18850 9168 20402
rect 9416 20398 9444 21830
rect 9600 21350 9628 22066
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9600 21078 9628 21286
rect 9692 21146 9720 22510
rect 9784 21486 9812 22578
rect 9876 22098 9904 24822
rect 9968 22574 9996 26200
rect 10704 23798 10732 26302
rect 11242 26200 11298 27000
rect 11886 26200 11942 27000
rect 12530 26200 12586 27000
rect 13174 26330 13230 27000
rect 13174 26302 13400 26330
rect 13174 26200 13230 26302
rect 10968 24608 11020 24614
rect 10968 24550 11020 24556
rect 10784 24200 10836 24206
rect 10784 24142 10836 24148
rect 10796 23798 10824 24142
rect 10692 23792 10744 23798
rect 10692 23734 10744 23740
rect 10784 23792 10836 23798
rect 10784 23734 10836 23740
rect 10048 23724 10100 23730
rect 10048 23666 10100 23672
rect 9956 22568 10008 22574
rect 9956 22510 10008 22516
rect 10060 22098 10088 23666
rect 10416 22500 10468 22506
rect 10416 22442 10468 22448
rect 9864 22092 9916 22098
rect 9864 22034 9916 22040
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 10322 21856 10378 21865
rect 10322 21791 10378 21800
rect 10336 21622 10364 21791
rect 10324 21616 10376 21622
rect 10324 21558 10376 21564
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 10324 21480 10376 21486
rect 10324 21422 10376 21428
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9588 21072 9640 21078
rect 9640 21020 10180 21026
rect 9588 21014 10180 21020
rect 9600 20998 10180 21014
rect 9496 20936 9548 20942
rect 9496 20878 9548 20884
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9220 19712 9272 19718
rect 9220 19654 9272 19660
rect 9048 18834 9168 18850
rect 9036 18828 9168 18834
rect 9088 18822 9168 18828
rect 9036 18770 9088 18776
rect 9140 18193 9168 18822
rect 9232 18737 9260 19654
rect 9312 19372 9364 19378
rect 9312 19314 9364 19320
rect 9218 18728 9274 18737
rect 9218 18663 9274 18672
rect 9126 18184 9182 18193
rect 9126 18119 9182 18128
rect 9324 17320 9352 19314
rect 9508 19310 9536 20878
rect 9956 20868 10008 20874
rect 9956 20810 10008 20816
rect 9968 20210 9996 20810
rect 9876 20182 9996 20210
rect 9876 19514 9904 20182
rect 9956 19916 10008 19922
rect 9956 19858 10008 19864
rect 9968 19514 9996 19858
rect 10152 19786 10180 20998
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10140 19780 10192 19786
rect 10060 19740 10140 19768
rect 9864 19508 9916 19514
rect 9864 19450 9916 19456
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 10060 19394 10088 19740
rect 10140 19722 10192 19728
rect 9968 19366 10088 19394
rect 10140 19372 10192 19378
rect 9496 19304 9548 19310
rect 9496 19246 9548 19252
rect 9678 18864 9734 18873
rect 9678 18799 9680 18808
rect 9732 18799 9734 18808
rect 9680 18770 9732 18776
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 9232 17292 9352 17320
rect 9128 17060 9180 17066
rect 9128 17002 9180 17008
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8312 16114 8340 16594
rect 8852 16448 8904 16454
rect 8852 16390 8904 16396
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 7656 15428 7708 15434
rect 7656 15370 7708 15376
rect 8680 15366 8708 15982
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 8864 15094 8892 16390
rect 8956 16182 8984 16390
rect 9140 16250 9168 17002
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 8944 16176 8996 16182
rect 8944 16118 8996 16124
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 8852 15088 8904 15094
rect 8852 15030 8904 15036
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 9048 13530 9076 15302
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 9232 12753 9260 17292
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9324 16425 9352 17138
rect 9416 17105 9444 17614
rect 9402 17096 9458 17105
rect 9402 17031 9458 17040
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9310 16416 9366 16425
rect 9310 16351 9366 16360
rect 9416 15473 9444 16458
rect 9508 15910 9536 18634
rect 9864 18624 9916 18630
rect 9968 18612 9996 19366
rect 10140 19314 10192 19320
rect 10046 19272 10102 19281
rect 10046 19207 10102 19216
rect 10060 18766 10088 19207
rect 10152 19145 10180 19314
rect 10138 19136 10194 19145
rect 10138 19071 10194 19080
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 9916 18584 9996 18612
rect 9864 18566 9916 18572
rect 9968 18290 9996 18584
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9600 16522 9628 18158
rect 9956 17808 10008 17814
rect 9956 17750 10008 17756
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9588 16516 9640 16522
rect 9588 16458 9640 16464
rect 9692 16046 9720 17478
rect 9876 17270 9904 17478
rect 9968 17338 9996 17750
rect 10152 17649 10180 19071
rect 10138 17640 10194 17649
rect 10138 17575 10194 17584
rect 10244 17513 10272 20402
rect 10336 19446 10364 21422
rect 10428 21146 10456 22442
rect 10690 21720 10746 21729
rect 10690 21655 10746 21664
rect 10416 21140 10468 21146
rect 10416 21082 10468 21088
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 10416 19984 10468 19990
rect 10416 19926 10468 19932
rect 10324 19440 10376 19446
rect 10324 19382 10376 19388
rect 10324 18896 10376 18902
rect 10324 18838 10376 18844
rect 10336 18426 10364 18838
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10428 18154 10456 19926
rect 10520 19174 10548 20402
rect 10600 19712 10652 19718
rect 10600 19654 10652 19660
rect 10508 19168 10560 19174
rect 10508 19110 10560 19116
rect 10416 18148 10468 18154
rect 10416 18090 10468 18096
rect 10324 17536 10376 17542
rect 10230 17504 10286 17513
rect 10324 17478 10376 17484
rect 10230 17439 10286 17448
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 9864 17264 9916 17270
rect 9864 17206 9916 17212
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9862 16280 9918 16289
rect 9862 16215 9918 16224
rect 9876 16182 9904 16215
rect 9864 16176 9916 16182
rect 9864 16118 9916 16124
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9864 15972 9916 15978
rect 9864 15914 9916 15920
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9772 15632 9824 15638
rect 9772 15574 9824 15580
rect 9680 15496 9732 15502
rect 9402 15464 9458 15473
rect 9680 15438 9732 15444
rect 9402 15399 9404 15408
rect 9456 15399 9458 15408
rect 9404 15370 9456 15376
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9508 12782 9536 15302
rect 9692 14618 9720 15438
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9600 13870 9628 14282
rect 9784 14074 9812 15574
rect 9876 15162 9904 15914
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9862 14104 9918 14113
rect 9772 14068 9824 14074
rect 9862 14039 9864 14048
rect 9772 14010 9824 14016
rect 9916 14039 9918 14048
rect 9864 14010 9916 14016
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9968 13705 9996 17138
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 10138 16688 10194 16697
rect 10138 16623 10140 16632
rect 10192 16623 10194 16632
rect 10140 16594 10192 16600
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 10060 16046 10088 16526
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 10152 15638 10180 16186
rect 10140 15632 10192 15638
rect 10140 15574 10192 15580
rect 10244 15366 10272 16730
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10336 15162 10364 17478
rect 10428 16658 10456 18090
rect 10520 17746 10548 19110
rect 10612 19009 10640 19654
rect 10598 19000 10654 19009
rect 10598 18935 10654 18944
rect 10508 17740 10560 17746
rect 10508 17682 10560 17688
rect 10612 17626 10640 18935
rect 10520 17598 10640 17626
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10324 14340 10376 14346
rect 10324 14282 10376 14288
rect 10336 13977 10364 14282
rect 10322 13968 10378 13977
rect 10232 13932 10284 13938
rect 10322 13903 10378 13912
rect 10232 13874 10284 13880
rect 10244 13841 10272 13874
rect 10324 13864 10376 13870
rect 10230 13832 10286 13841
rect 10324 13806 10376 13812
rect 10230 13767 10286 13776
rect 9954 13696 10010 13705
rect 9954 13631 10010 13640
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9876 12986 9904 13330
rect 9954 13288 10010 13297
rect 9954 13223 9956 13232
rect 10008 13223 10010 13232
rect 9956 13194 10008 13200
rect 10336 13161 10364 13806
rect 10322 13152 10378 13161
rect 10322 13087 10378 13096
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9496 12776 9548 12782
rect 9218 12744 9274 12753
rect 9496 12718 9548 12724
rect 9218 12679 9274 12688
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 1306 6488 1362 6497
rect 1216 6452 1268 6458
rect 1306 6423 1362 6432
rect 1216 6394 1268 6400
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 1320 6089 1348 6258
rect 1306 6080 1362 6089
rect 1306 6015 1362 6024
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 1308 5704 1360 5710
rect 1306 5672 1308 5681
rect 2780 5704 2832 5710
rect 1360 5672 1362 5681
rect 2780 5646 2832 5652
rect 1306 5607 1362 5616
rect 2792 5273 2820 5646
rect 2778 5264 2834 5273
rect 2778 5199 2834 5208
rect 1308 5160 1360 5166
rect 1308 5102 1360 5108
rect 1320 4865 1348 5102
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 1306 4856 1362 4865
rect 2950 4859 3258 4868
rect 1306 4791 1308 4800
rect 1360 4791 1362 4800
rect 5540 4820 5592 4826
rect 1308 4762 1360 4768
rect 5540 4762 5592 4768
rect 1308 4616 1360 4622
rect 1308 4558 1360 4564
rect 1320 4457 1348 4558
rect 1306 4448 1362 4457
rect 1306 4383 1362 4392
rect 1400 4208 1452 4214
rect 1400 4150 1452 4156
rect 1308 4140 1360 4146
rect 1308 4082 1360 4088
rect 1320 3641 1348 4082
rect 1412 4049 1440 4150
rect 1398 4040 1454 4049
rect 1398 3975 1454 3984
rect 5552 3942 5580 4762
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 1306 3632 1362 3641
rect 1124 3596 1176 3602
rect 1306 3567 1362 3576
rect 1124 3538 1176 3544
rect 1136 800 1164 3538
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1320 3233 1348 3470
rect 1306 3224 1362 3233
rect 1306 3159 1308 3168
rect 1360 3159 1362 3168
rect 1308 3130 1360 3136
rect 1308 3052 1360 3058
rect 1308 2994 1360 3000
rect 1320 2825 1348 2994
rect 2320 2848 2372 2854
rect 1306 2816 1362 2825
rect 2320 2790 2372 2796
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 3332 2848 3384 2854
rect 3332 2790 3384 2796
rect 1306 2751 1362 2760
rect 2332 2446 2360 2790
rect 2792 2514 2820 2790
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 1308 2440 1360 2446
rect 1306 2408 1308 2417
rect 2320 2440 2372 2446
rect 1360 2408 1362 2417
rect 1216 2372 1268 2378
rect 2320 2382 2372 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 1306 2343 1362 2352
rect 1216 2314 1268 2320
rect 1228 2009 1256 2314
rect 3252 2106 3280 2382
rect 1308 2100 1360 2106
rect 1308 2042 1360 2048
rect 3240 2100 3292 2106
rect 3240 2042 3292 2048
rect 1214 2000 1270 2009
rect 1214 1935 1270 1944
rect 1320 1601 1348 2042
rect 1306 1592 1362 1601
rect 1306 1527 1362 1536
rect 3344 1442 3372 2790
rect 3252 1414 3372 1442
rect 3252 800 3280 1414
rect 5368 800 5396 3674
rect 7484 800 7512 3878
rect 7576 3534 7604 12038
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 9876 11898 9904 12922
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9876 11354 9904 11834
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 10060 6186 10088 12650
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 10244 11286 10272 12038
rect 10232 11280 10284 11286
rect 10232 11222 10284 11228
rect 10336 10674 10364 13087
rect 10428 12986 10456 14758
rect 10520 14618 10548 17598
rect 10598 17368 10654 17377
rect 10598 17303 10654 17312
rect 10612 17134 10640 17303
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10598 16280 10654 16289
rect 10598 16215 10654 16224
rect 10612 16182 10640 16215
rect 10600 16176 10652 16182
rect 10600 16118 10652 16124
rect 10598 15872 10654 15881
rect 10598 15807 10654 15816
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10416 12640 10468 12646
rect 10416 12582 10468 12588
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10428 10130 10456 12582
rect 10612 11830 10640 15807
rect 10704 15502 10732 21655
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 10796 18698 10824 19654
rect 10784 18692 10836 18698
rect 10784 18634 10836 18640
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10796 17678 10824 18022
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10796 15570 10824 17614
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10888 16794 10916 17070
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10980 16182 11008 24550
rect 11256 23186 11284 26200
rect 11796 24676 11848 24682
rect 11796 24618 11848 24624
rect 11612 24200 11664 24206
rect 11612 24142 11664 24148
rect 11244 23180 11296 23186
rect 11244 23122 11296 23128
rect 11518 22808 11574 22817
rect 11518 22743 11574 22752
rect 11532 22273 11560 22743
rect 11624 22574 11652 24142
rect 11808 23730 11836 24618
rect 11796 23724 11848 23730
rect 11796 23666 11848 23672
rect 11702 22672 11758 22681
rect 11702 22607 11758 22616
rect 11612 22568 11664 22574
rect 11612 22510 11664 22516
rect 11518 22264 11574 22273
rect 11518 22199 11574 22208
rect 11060 21956 11112 21962
rect 11060 21898 11112 21904
rect 11072 18170 11100 21898
rect 11152 21480 11204 21486
rect 11150 21448 11152 21457
rect 11204 21448 11206 21457
rect 11150 21383 11206 21392
rect 11624 20398 11652 22510
rect 11716 22098 11744 22607
rect 11796 22568 11848 22574
rect 11794 22536 11796 22545
rect 11848 22536 11850 22545
rect 11794 22471 11850 22480
rect 11808 22166 11836 22471
rect 11900 22166 11928 26200
rect 11978 24712 12034 24721
rect 11978 24647 12034 24656
rect 11992 22574 12020 24647
rect 12544 24138 12572 26200
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12532 24132 12584 24138
rect 12532 24074 12584 24080
rect 12440 24064 12492 24070
rect 12440 24006 12492 24012
rect 12070 23760 12126 23769
rect 12070 23695 12072 23704
rect 12124 23695 12126 23704
rect 12072 23666 12124 23672
rect 12452 23118 12480 24006
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13268 23316 13320 23322
rect 13268 23258 13320 23264
rect 12440 23112 12492 23118
rect 12440 23054 12492 23060
rect 11980 22568 12032 22574
rect 11980 22510 12032 22516
rect 13280 22438 13308 23258
rect 13372 23186 13400 26302
rect 13818 26200 13874 27000
rect 14462 26200 14518 27000
rect 15106 26330 15162 27000
rect 14752 26302 15162 26330
rect 13452 24404 13504 24410
rect 13452 24346 13504 24352
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 13268 22432 13320 22438
rect 13268 22374 13320 22380
rect 13360 22432 13412 22438
rect 13360 22374 13412 22380
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 11796 22160 11848 22166
rect 11796 22102 11848 22108
rect 11888 22160 11940 22166
rect 11888 22102 11940 22108
rect 11704 22092 11756 22098
rect 11704 22034 11756 22040
rect 11796 22024 11848 22030
rect 11796 21966 11848 21972
rect 11808 21690 11836 21966
rect 13372 21690 13400 22374
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 13360 21684 13412 21690
rect 13360 21626 13412 21632
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11704 20528 11756 20534
rect 11702 20496 11704 20505
rect 11756 20496 11758 20505
rect 11702 20431 11758 20440
rect 11612 20392 11664 20398
rect 11612 20334 11664 20340
rect 11520 20324 11572 20330
rect 11520 20266 11572 20272
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 11164 20058 11192 20198
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 11336 19440 11388 19446
rect 11336 19382 11388 19388
rect 11152 19236 11204 19242
rect 11152 19178 11204 19184
rect 11164 18290 11192 19178
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 11072 18142 11192 18170
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 10968 16176 11020 16182
rect 11072 16153 11100 18022
rect 11164 17882 11192 18142
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11256 17490 11284 18022
rect 11348 17610 11376 19382
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11336 17604 11388 17610
rect 11336 17546 11388 17552
rect 11164 17462 11284 17490
rect 10968 16118 11020 16124
rect 11058 16144 11114 16153
rect 11058 16079 11114 16088
rect 11164 15910 11192 17462
rect 11440 17320 11468 17818
rect 11532 17542 11560 20266
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11716 17542 11744 19790
rect 11794 19408 11850 19417
rect 11794 19343 11796 19352
rect 11848 19343 11850 19352
rect 11796 19314 11848 19320
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11808 18902 11836 19110
rect 11796 18896 11848 18902
rect 11796 18838 11848 18844
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11256 17292 11468 17320
rect 11256 16590 11284 17292
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 11348 16402 11376 16526
rect 11256 16374 11376 16402
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10692 15496 10744 15502
rect 10692 15438 10744 15444
rect 11164 15434 11192 15846
rect 11256 15706 11284 16374
rect 11440 16250 11468 17138
rect 11520 16448 11572 16454
rect 11520 16390 11572 16396
rect 11612 16448 11664 16454
rect 11612 16390 11664 16396
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 11532 15706 11560 16390
rect 11624 16250 11652 16390
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 11152 15428 11204 15434
rect 11152 15370 11204 15376
rect 11520 15428 11572 15434
rect 11520 15370 11572 15376
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 10980 14929 11008 14962
rect 10966 14920 11022 14929
rect 10966 14855 11022 14864
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 10704 14249 10732 14758
rect 11072 14550 11100 14758
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 10690 14240 10746 14249
rect 10690 14175 10746 14184
rect 10600 11824 10652 11830
rect 10600 11766 10652 11772
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 8850 5128 8906 5137
rect 8850 5063 8906 5072
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 8864 2854 8892 5063
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9508 2310 9536 2586
rect 9680 2440 9732 2446
rect 9600 2388 9680 2394
rect 9600 2382 9732 2388
rect 9600 2366 9720 2382
rect 10612 2378 10640 11018
rect 10704 7818 10732 14175
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10888 12170 10916 13262
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 11072 12986 11100 13194
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10980 12186 11008 12718
rect 10876 12164 10928 12170
rect 10980 12158 11100 12186
rect 10876 12106 10928 12112
rect 10888 11898 10916 12106
rect 11072 12102 11100 12158
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10796 5166 10824 11290
rect 10888 11218 10916 11834
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 11164 9042 11192 14962
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11256 14006 11284 14214
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11348 12850 11376 14214
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11440 12730 11468 14350
rect 11532 14074 11560 15370
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11532 13394 11560 14010
rect 11520 13388 11572 13394
rect 11572 13348 11652 13376
rect 11520 13330 11572 13336
rect 11624 13258 11652 13348
rect 11612 13252 11664 13258
rect 11612 13194 11664 13200
rect 11348 12702 11468 12730
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11256 9926 11284 10406
rect 11348 10033 11376 12702
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11440 11014 11468 12582
rect 11624 12170 11652 13194
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11624 11098 11652 12106
rect 11808 11665 11836 18226
rect 11888 16516 11940 16522
rect 11888 16458 11940 16464
rect 11900 13002 11928 16458
rect 11992 16454 12020 21490
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12912 21100 13308 21128
rect 12912 21010 12940 21100
rect 13280 21010 13308 21100
rect 12900 21004 12952 21010
rect 13268 21004 13320 21010
rect 12900 20946 12952 20952
rect 13004 20964 13216 20992
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12256 20800 12308 20806
rect 12256 20742 12308 20748
rect 12268 20534 12296 20742
rect 12256 20528 12308 20534
rect 12256 20470 12308 20476
rect 12072 20460 12124 20466
rect 12072 20402 12124 20408
rect 12084 20369 12112 20402
rect 12348 20392 12400 20398
rect 12070 20360 12126 20369
rect 12348 20334 12400 20340
rect 12070 20295 12126 20304
rect 12360 20058 12388 20334
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12452 20058 12480 20198
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12072 19440 12124 19446
rect 12072 19382 12124 19388
rect 12084 18154 12112 19382
rect 12360 18222 12388 19858
rect 12544 19718 12572 20878
rect 12808 20868 12860 20874
rect 13004 20856 13032 20964
rect 13188 20874 13216 20964
rect 13268 20946 13320 20952
rect 13464 20942 13492 24346
rect 13832 22574 13860 26200
rect 14280 24336 14332 24342
rect 14280 24278 14332 24284
rect 14292 23186 14320 24278
rect 14476 24274 14504 26200
rect 14464 24268 14516 24274
rect 14464 24210 14516 24216
rect 14752 23798 14780 26302
rect 15106 26200 15162 26302
rect 15750 26330 15806 27000
rect 15750 26302 15884 26330
rect 15750 26200 15806 26302
rect 15016 24064 15068 24070
rect 15016 24006 15068 24012
rect 14740 23792 14792 23798
rect 14740 23734 14792 23740
rect 14740 23656 14792 23662
rect 14740 23598 14792 23604
rect 14280 23180 14332 23186
rect 14280 23122 14332 23128
rect 14556 23180 14608 23186
rect 14556 23122 14608 23128
rect 14096 23044 14148 23050
rect 14096 22986 14148 22992
rect 13820 22568 13872 22574
rect 13820 22510 13872 22516
rect 13912 22228 13964 22234
rect 13912 22170 13964 22176
rect 13636 22160 13688 22166
rect 13636 22102 13688 22108
rect 13648 21554 13676 22102
rect 13636 21548 13688 21554
rect 13636 21490 13688 21496
rect 13452 20936 13504 20942
rect 13452 20878 13504 20884
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 12860 20828 13032 20856
rect 13084 20868 13136 20874
rect 12808 20810 12860 20816
rect 13084 20810 13136 20816
rect 13176 20868 13228 20874
rect 13176 20810 13228 20816
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12714 20768 12770 20777
rect 12636 20398 12664 20742
rect 12714 20703 12770 20712
rect 12728 20466 12756 20703
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 13096 20330 13124 20810
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 13084 20324 13136 20330
rect 13084 20266 13136 20272
rect 13636 20256 13688 20262
rect 13636 20198 13688 20204
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12452 19530 12480 19654
rect 12636 19530 12664 19994
rect 13648 19854 13676 20198
rect 13636 19848 13688 19854
rect 13636 19790 13688 19796
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 12452 19502 12664 19530
rect 13360 19508 13412 19514
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12452 18970 12480 19110
rect 12544 18970 12572 19502
rect 13360 19450 13412 19456
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12348 18216 12400 18222
rect 12348 18158 12400 18164
rect 12072 18148 12124 18154
rect 12072 18090 12124 18096
rect 12360 17746 12388 18158
rect 12452 18086 12480 18702
rect 12544 18272 12572 18906
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 12544 18244 12664 18272
rect 12532 18148 12584 18154
rect 12532 18090 12584 18096
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 12452 17678 12480 18022
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12162 17232 12218 17241
rect 12162 17167 12164 17176
rect 12216 17167 12218 17176
rect 12164 17138 12216 17144
rect 12164 17060 12216 17066
rect 12164 17002 12216 17008
rect 12072 16516 12124 16522
rect 12072 16458 12124 16464
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 12084 16182 12112 16458
rect 12072 16176 12124 16182
rect 12072 16118 12124 16124
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 11992 15201 12020 16050
rect 12072 15904 12124 15910
rect 12070 15872 12072 15881
rect 12124 15872 12126 15881
rect 12070 15807 12126 15816
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 11978 15192 12034 15201
rect 12084 15162 12112 15302
rect 11978 15127 12034 15136
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 11980 15088 12032 15094
rect 12084 15065 12112 15098
rect 11980 15030 12032 15036
rect 12070 15056 12126 15065
rect 11992 14414 12020 15030
rect 12070 14991 12126 15000
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 12176 14328 12204 17002
rect 12268 14958 12296 17478
rect 12452 17270 12480 17614
rect 12544 17338 12572 18090
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12440 17264 12492 17270
rect 12440 17206 12492 17212
rect 12636 17202 12664 18244
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 12452 16590 12480 17002
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12348 16108 12400 16114
rect 12348 16050 12400 16056
rect 12360 15638 12388 16050
rect 12348 15632 12400 15638
rect 12348 15574 12400 15580
rect 12544 15094 12572 16934
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12636 15570 12664 15982
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 12728 15026 12756 17682
rect 12820 15162 12848 18362
rect 13372 18222 13400 19450
rect 13452 19304 13504 19310
rect 13452 19246 13504 19252
rect 13464 18222 13492 19246
rect 13648 19145 13676 19654
rect 13634 19136 13690 19145
rect 13634 19071 13690 19080
rect 13740 19009 13768 20742
rect 13832 20398 13860 20878
rect 13924 20602 13952 22170
rect 14108 21162 14136 22986
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 14292 22098 14320 22918
rect 14464 22704 14516 22710
rect 14464 22646 14516 22652
rect 14280 22092 14332 22098
rect 14280 22034 14332 22040
rect 14372 21956 14424 21962
rect 14372 21898 14424 21904
rect 14188 21888 14240 21894
rect 14188 21830 14240 21836
rect 14200 21321 14228 21830
rect 14186 21312 14242 21321
rect 14186 21247 14242 21256
rect 14016 21134 14136 21162
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 13820 20392 13872 20398
rect 13820 20334 13872 20340
rect 13832 19922 13860 20334
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 13726 19000 13782 19009
rect 13726 18935 13782 18944
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13556 18329 13584 18838
rect 13832 18834 13860 19858
rect 14016 19310 14044 21134
rect 14384 21010 14412 21898
rect 14188 21004 14240 21010
rect 14188 20946 14240 20952
rect 14372 21004 14424 21010
rect 14372 20946 14424 20952
rect 14200 20398 14228 20946
rect 14188 20392 14240 20398
rect 14188 20334 14240 20340
rect 14384 19990 14412 20946
rect 14476 20806 14504 22646
rect 14464 20800 14516 20806
rect 14464 20742 14516 20748
rect 14372 19984 14424 19990
rect 14372 19926 14424 19932
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13542 18320 13598 18329
rect 13542 18255 13598 18264
rect 14004 18284 14056 18290
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13358 17912 13414 17921
rect 13358 17847 13414 17856
rect 13372 17814 13400 17847
rect 13360 17808 13412 17814
rect 13360 17750 13412 17756
rect 13556 17678 13584 18255
rect 14004 18226 14056 18232
rect 14016 18154 14044 18226
rect 14108 18170 14136 19790
rect 14568 19530 14596 23122
rect 14648 23044 14700 23050
rect 14648 22986 14700 22992
rect 14660 19825 14688 22986
rect 14752 22098 14780 23598
rect 14740 22092 14792 22098
rect 15028 22094 15056 24006
rect 15568 23860 15620 23866
rect 15568 23802 15620 23808
rect 15292 23792 15344 23798
rect 15292 23734 15344 23740
rect 15304 23594 15332 23734
rect 15292 23588 15344 23594
rect 15292 23530 15344 23536
rect 15028 22066 15148 22094
rect 14740 22034 14792 22040
rect 14832 21956 14884 21962
rect 14832 21898 14884 21904
rect 14738 21720 14794 21729
rect 14738 21655 14740 21664
rect 14792 21655 14794 21664
rect 14740 21626 14792 21632
rect 14646 19816 14702 19825
rect 14646 19751 14702 19760
rect 14476 19502 14596 19530
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14200 18290 14228 18702
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14004 18148 14056 18154
rect 14108 18142 14228 18170
rect 14004 18090 14056 18096
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13464 16998 13492 17478
rect 14016 17338 14044 18090
rect 14004 17332 14056 17338
rect 13924 17292 14004 17320
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13464 16658 13492 16934
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 12992 16448 13044 16454
rect 12992 16390 13044 16396
rect 13004 16182 13032 16390
rect 12992 16176 13044 16182
rect 12992 16118 13044 16124
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12348 14544 12400 14550
rect 12400 14504 12480 14532
rect 12348 14486 12400 14492
rect 12256 14340 12308 14346
rect 12176 14300 12256 14328
rect 12256 14282 12308 14288
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 11900 12974 12020 13002
rect 12084 12986 12112 13126
rect 12268 12986 12296 13670
rect 11794 11656 11850 11665
rect 11794 11591 11850 11600
rect 11624 11082 11928 11098
rect 11624 11076 11940 11082
rect 11624 11070 11888 11076
rect 11888 11018 11940 11024
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11716 10810 11744 10950
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11334 10024 11390 10033
rect 11440 9994 11468 10746
rect 11334 9959 11390 9968
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11256 9382 11284 9862
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11072 2650 11100 2926
rect 11256 2922 11284 9318
rect 11992 8838 12020 12974
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 12268 12306 12296 12786
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12072 11552 12124 11558
rect 12070 11520 12072 11529
rect 12124 11520 12126 11529
rect 12070 11455 12126 11464
rect 12176 11218 12204 11630
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12268 10674 12296 12038
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12360 9178 12388 13738
rect 12452 13546 12480 14504
rect 12544 14006 12572 14894
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13360 14476 13412 14482
rect 13464 14464 13492 14758
rect 13544 14476 13596 14482
rect 13464 14436 13544 14464
rect 13360 14418 13412 14424
rect 13544 14418 13596 14424
rect 13372 14006 13400 14418
rect 13450 14376 13506 14385
rect 13450 14311 13506 14320
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 13360 14000 13412 14006
rect 13360 13942 13412 13948
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12624 13864 12676 13870
rect 12622 13832 12624 13841
rect 12676 13832 12678 13841
rect 12622 13767 12678 13776
rect 12452 13518 12664 13546
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 12452 11529 12480 13398
rect 12532 13388 12584 13394
rect 12532 13330 12584 13336
rect 12544 12850 12572 13330
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12636 11778 12664 13518
rect 12544 11750 12664 11778
rect 12438 11520 12494 11529
rect 12438 11455 12494 11464
rect 12544 10810 12572 11750
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12636 10266 12664 11630
rect 12728 11218 12756 13874
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12808 13456 12860 13462
rect 12808 13398 12860 13404
rect 12820 12782 12848 13398
rect 13372 13326 13400 13806
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13372 12918 13400 13262
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12820 12434 12848 12582
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13084 12436 13136 12442
rect 12820 12406 12940 12434
rect 12912 11801 12940 12406
rect 13084 12378 13136 12384
rect 13096 12170 13124 12378
rect 13084 12164 13136 12170
rect 13084 12106 13136 12112
rect 13372 11898 13400 12854
rect 13464 12170 13492 14311
rect 13556 13394 13584 14418
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 12898 11792 12954 11801
rect 12898 11727 12954 11736
rect 13450 11792 13506 11801
rect 13450 11727 13506 11736
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12544 9586 12572 10066
rect 12728 9654 12756 10406
rect 12820 10266 12848 10474
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13280 9926 13308 10202
rect 13372 10062 13400 10950
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 13372 9518 13400 9998
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12440 8900 12492 8906
rect 12440 8842 12492 8848
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 12452 6914 12480 8842
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12360 6886 12480 6914
rect 11244 2916 11296 2922
rect 11244 2858 11296 2864
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 10600 2372 10652 2378
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 9600 800 9628 2366
rect 10600 2314 10652 2320
rect 11716 800 11744 2450
rect 12360 2310 12388 6886
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 13464 5846 13492 11727
rect 13556 10130 13584 13330
rect 13648 11642 13676 16526
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13740 15502 13768 15982
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13924 15094 13952 17292
rect 14004 17274 14056 17280
rect 14004 16652 14056 16658
rect 14004 16594 14056 16600
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 14016 16046 14044 16594
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 13912 15088 13964 15094
rect 13912 15030 13964 15036
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13832 13530 13860 14418
rect 13924 14278 13952 15030
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13740 12238 13768 13262
rect 13924 12306 13952 13942
rect 14016 13734 14044 15982
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13728 12232 13780 12238
rect 13924 12209 13952 12242
rect 13910 12200 13966 12209
rect 13728 12174 13780 12180
rect 13832 12158 13910 12186
rect 13648 11614 13768 11642
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13648 9042 13676 11494
rect 13740 10713 13768 11614
rect 13832 11132 13860 12158
rect 13910 12135 13966 12144
rect 13910 12064 13966 12073
rect 13910 11999 13966 12008
rect 13924 11286 13952 11999
rect 14016 11762 14044 13670
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 13912 11280 13964 11286
rect 13912 11222 13964 11228
rect 13832 11104 13952 11132
rect 13726 10704 13782 10713
rect 13726 10639 13782 10648
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13832 9722 13860 10542
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13740 8634 13768 9114
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13832 8498 13860 9658
rect 13924 9518 13952 11104
rect 14108 9994 14136 16594
rect 14200 15609 14228 18142
rect 14292 18086 14320 18702
rect 14384 18193 14412 19110
rect 14370 18184 14426 18193
rect 14370 18119 14426 18128
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 14292 17746 14320 18022
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14384 16658 14412 17478
rect 14476 16794 14504 19502
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14568 18970 14596 19314
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14844 18204 14872 21898
rect 15120 21690 15148 22066
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15108 21684 15160 21690
rect 15108 21626 15160 21632
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 14936 19174 14964 21490
rect 15016 21480 15068 21486
rect 15016 21422 15068 21428
rect 15028 21010 15056 21422
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 15106 20904 15162 20913
rect 15106 20839 15162 20848
rect 15120 20602 15148 20839
rect 15212 20618 15240 21966
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 15304 21486 15332 21830
rect 15580 21690 15608 23802
rect 15856 22710 15884 26302
rect 16394 26200 16450 27000
rect 17038 26200 17094 27000
rect 17682 26330 17738 27000
rect 17682 26302 17908 26330
rect 17682 26200 17738 26302
rect 16408 23186 16436 26200
rect 17052 23798 17080 26200
rect 17132 24200 17184 24206
rect 17776 24200 17828 24206
rect 17132 24142 17184 24148
rect 17774 24168 17776 24177
rect 17828 24168 17830 24177
rect 17040 23792 17092 23798
rect 17040 23734 17092 23740
rect 16764 23656 16816 23662
rect 16764 23598 16816 23604
rect 16396 23180 16448 23186
rect 16396 23122 16448 23128
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 16486 22808 16542 22817
rect 16684 22778 16712 23054
rect 16486 22743 16542 22752
rect 16580 22772 16632 22778
rect 15844 22704 15896 22710
rect 15844 22646 15896 22652
rect 16026 22128 16082 22137
rect 16026 22063 16082 22072
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 15304 21146 15332 21422
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15108 20596 15160 20602
rect 15212 20590 15332 20618
rect 15108 20538 15160 20544
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15212 19990 15240 20402
rect 15200 19984 15252 19990
rect 15200 19926 15252 19932
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 14924 19168 14976 19174
rect 14924 19110 14976 19116
rect 15120 18714 15148 19654
rect 15304 18834 15332 20590
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15396 20058 15424 20538
rect 15476 20324 15528 20330
rect 15476 20266 15528 20272
rect 15488 20058 15516 20266
rect 15764 20097 15792 21286
rect 15936 20936 15988 20942
rect 15856 20896 15936 20924
rect 15750 20088 15806 20097
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15476 20052 15528 20058
rect 15750 20023 15806 20032
rect 15476 19994 15528 20000
rect 15856 19990 15884 20896
rect 15936 20878 15988 20884
rect 15936 20528 15988 20534
rect 15936 20470 15988 20476
rect 15844 19984 15896 19990
rect 15844 19926 15896 19932
rect 15568 19440 15620 19446
rect 15568 19382 15620 19388
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 15120 18686 15332 18714
rect 15304 18630 15332 18686
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 15292 18624 15344 18630
rect 15292 18566 15344 18572
rect 15212 18426 15240 18566
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 14844 18176 14964 18204
rect 14936 17882 14964 18176
rect 15488 17921 15516 18226
rect 15474 17912 15530 17921
rect 14924 17876 14976 17882
rect 15474 17847 15530 17856
rect 14924 17818 14976 17824
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 14922 17640 14978 17649
rect 14556 17604 14608 17610
rect 14922 17575 14978 17584
rect 14556 17546 14608 17552
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14476 16250 14504 16390
rect 14464 16244 14516 16250
rect 14464 16186 14516 16192
rect 14568 15706 14596 17546
rect 14646 17096 14702 17105
rect 14646 17031 14702 17040
rect 14832 17060 14884 17066
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14186 15600 14242 15609
rect 14186 15535 14242 15544
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14292 14890 14320 15438
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14280 14884 14332 14890
rect 14280 14826 14332 14832
rect 14278 14512 14334 14521
rect 14278 14447 14334 14456
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14200 14006 14228 14214
rect 14188 14000 14240 14006
rect 14188 13942 14240 13948
rect 14200 13462 14228 13942
rect 14188 13456 14240 13462
rect 14188 13398 14240 13404
rect 14200 12900 14228 13398
rect 14292 13258 14320 14447
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14476 13433 14504 13466
rect 14462 13424 14518 13433
rect 14462 13359 14518 13368
rect 14370 13288 14426 13297
rect 14280 13252 14332 13258
rect 14370 13223 14372 13232
rect 14280 13194 14332 13200
rect 14424 13223 14426 13232
rect 14372 13194 14424 13200
rect 14372 12912 14424 12918
rect 14200 12872 14372 12900
rect 14200 11830 14228 12872
rect 14372 12854 14424 12860
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14292 11830 14320 12174
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14280 11824 14332 11830
rect 14280 11766 14332 11772
rect 14292 10130 14320 11766
rect 14568 11354 14596 15302
rect 14660 14929 14688 17031
rect 14832 17002 14884 17008
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14752 16794 14780 16934
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14844 16590 14872 17002
rect 14832 16584 14884 16590
rect 14832 16526 14884 16532
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14844 15910 14872 16050
rect 14936 15994 14964 17575
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 15028 16182 15056 16934
rect 15120 16658 15148 17682
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 15212 16561 15240 17682
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15396 17202 15424 17274
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15198 16552 15254 16561
rect 15198 16487 15254 16496
rect 15016 16176 15068 16182
rect 15016 16118 15068 16124
rect 14936 15966 15056 15994
rect 14832 15904 14884 15910
rect 14884 15864 14964 15892
rect 14832 15846 14884 15852
rect 14936 15162 14964 15864
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 14646 14920 14702 14929
rect 14646 14855 14702 14864
rect 14844 14346 14872 15098
rect 14832 14340 14884 14346
rect 14832 14282 14884 14288
rect 14924 14272 14976 14278
rect 14922 14240 14924 14249
rect 14976 14240 14978 14249
rect 14922 14175 14978 14184
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14660 11121 14688 13738
rect 15028 13433 15056 15966
rect 15108 15564 15160 15570
rect 15108 15506 15160 15512
rect 15120 14074 15148 15506
rect 15292 15088 15344 15094
rect 15292 15030 15344 15036
rect 15304 14822 15332 15030
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15304 14385 15332 14758
rect 15290 14376 15346 14385
rect 15290 14311 15346 14320
rect 15108 14068 15160 14074
rect 15108 14010 15160 14016
rect 15120 13569 15148 14010
rect 15106 13560 15162 13569
rect 15106 13495 15162 13504
rect 15200 13524 15252 13530
rect 15014 13424 15070 13433
rect 15014 13359 15070 13368
rect 14832 13184 14884 13190
rect 14830 13152 14832 13161
rect 14924 13184 14976 13190
rect 14884 13152 14886 13161
rect 14924 13126 14976 13132
rect 14830 13087 14886 13096
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14752 11626 14780 11698
rect 14740 11620 14792 11626
rect 14740 11562 14792 11568
rect 14832 11552 14884 11558
rect 14830 11520 14832 11529
rect 14884 11520 14886 11529
rect 14830 11455 14886 11464
rect 14646 11112 14702 11121
rect 14646 11047 14702 11056
rect 14936 10742 14964 13126
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 15028 11218 15056 11494
rect 15120 11218 15148 13495
rect 15200 13466 15252 13472
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15106 11112 15162 11121
rect 15106 11047 15108 11056
rect 15160 11047 15162 11056
rect 15108 11018 15160 11024
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 14924 10736 14976 10742
rect 14924 10678 14976 10684
rect 14832 10532 14884 10538
rect 14832 10474 14884 10480
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 14004 9648 14056 9654
rect 14056 9596 14136 9602
rect 14004 9590 14136 9596
rect 14016 9574 14136 9590
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 14108 7410 14136 9574
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14200 8566 14228 8978
rect 14292 8974 14320 9318
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14292 8566 14320 8910
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 14280 8560 14332 8566
rect 14280 8502 14332 8508
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 13452 5840 13504 5846
rect 13452 5782 13504 5788
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12544 2446 12572 3334
rect 14292 3058 14320 8502
rect 14384 7818 14412 10406
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14568 8634 14596 8842
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14844 7954 14872 10474
rect 15028 10305 15056 10950
rect 15212 10810 15240 13466
rect 15384 13252 15436 13258
rect 15384 13194 15436 13200
rect 15396 13161 15424 13194
rect 15382 13152 15438 13161
rect 15382 13087 15438 13096
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15304 12170 15332 12718
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15014 10296 15070 10305
rect 15014 10231 15070 10240
rect 15304 9994 15332 12106
rect 15396 10606 15424 13087
rect 15488 11898 15516 17070
rect 15580 17066 15608 19382
rect 15856 18698 15884 19926
rect 15948 19854 15976 20470
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 16040 19310 16068 22063
rect 16118 21584 16174 21593
rect 16118 21519 16120 21528
rect 16172 21519 16174 21528
rect 16120 21490 16172 21496
rect 16396 20800 16448 20806
rect 16394 20768 16396 20777
rect 16448 20768 16450 20777
rect 16394 20703 16450 20712
rect 16118 20496 16174 20505
rect 16118 20431 16120 20440
rect 16172 20431 16174 20440
rect 16120 20402 16172 20408
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 16224 19961 16252 20198
rect 16210 19952 16266 19961
rect 16210 19887 16266 19896
rect 16304 19780 16356 19786
rect 16304 19722 16356 19728
rect 16210 19680 16266 19689
rect 16210 19615 16266 19624
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 15844 18692 15896 18698
rect 15844 18634 15896 18640
rect 15856 18086 15884 18634
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15856 17678 15884 18022
rect 16040 17882 16068 18158
rect 16028 17876 16080 17882
rect 16028 17818 16080 17824
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15936 17536 15988 17542
rect 15934 17504 15936 17513
rect 15988 17504 15990 17513
rect 15934 17439 15990 17448
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 15580 13530 15608 15370
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15672 13394 15700 16186
rect 15764 15706 15792 16526
rect 15948 16114 15976 17439
rect 16132 17134 16160 18906
rect 16224 18426 16252 19615
rect 16316 19514 16344 19722
rect 16304 19508 16356 19514
rect 16304 19450 16356 19456
rect 16302 19000 16358 19009
rect 16302 18935 16304 18944
rect 16356 18935 16358 18944
rect 16304 18906 16356 18912
rect 16408 18902 16436 20703
rect 16500 19360 16528 22743
rect 16580 22714 16632 22720
rect 16672 22772 16724 22778
rect 16672 22714 16724 22720
rect 16592 22137 16620 22714
rect 16578 22128 16634 22137
rect 16776 22094 16804 23598
rect 17144 23361 17172 24142
rect 17774 24103 17830 24112
rect 17408 24064 17460 24070
rect 17408 24006 17460 24012
rect 17224 23724 17276 23730
rect 17224 23666 17276 23672
rect 17236 23526 17264 23666
rect 17224 23520 17276 23526
rect 17224 23462 17276 23468
rect 17130 23352 17186 23361
rect 17130 23287 17132 23296
rect 17184 23287 17186 23296
rect 17132 23258 17184 23264
rect 17132 23112 17184 23118
rect 17132 23054 17184 23060
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 16868 22438 16896 22578
rect 17144 22438 17172 23054
rect 16856 22432 16908 22438
rect 16856 22374 16908 22380
rect 17132 22432 17184 22438
rect 17132 22374 17184 22380
rect 16856 22228 16908 22234
rect 16856 22170 16908 22176
rect 16578 22063 16634 22072
rect 16684 22066 16804 22094
rect 16684 19514 16712 22066
rect 16868 21962 16896 22170
rect 17132 22160 17184 22166
rect 17132 22102 17184 22108
rect 16856 21956 16908 21962
rect 16776 21916 16856 21944
rect 16776 20942 16804 21916
rect 16856 21898 16908 21904
rect 17040 21888 17092 21894
rect 16946 21856 17002 21865
rect 17040 21830 17092 21836
rect 16946 21791 17002 21800
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16868 21049 16896 21286
rect 16960 21146 16988 21791
rect 17052 21622 17080 21830
rect 17144 21622 17172 22102
rect 17040 21616 17092 21622
rect 17040 21558 17092 21564
rect 17132 21616 17184 21622
rect 17132 21558 17184 21564
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 16854 21040 16910 21049
rect 16854 20975 16910 20984
rect 16764 20936 16816 20942
rect 16764 20878 16816 20884
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16776 20262 16804 20402
rect 17052 20398 17080 21558
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 17130 21176 17186 21185
rect 17236 21146 17264 21490
rect 17130 21111 17186 21120
rect 17224 21140 17276 21146
rect 17144 20641 17172 21111
rect 17224 21082 17276 21088
rect 17316 20800 17368 20806
rect 17316 20742 17368 20748
rect 17130 20632 17186 20641
rect 17130 20567 17186 20576
rect 17040 20392 17092 20398
rect 17040 20334 17092 20340
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16856 20256 16908 20262
rect 16856 20198 16908 20204
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16500 19332 16620 19360
rect 16592 19009 16620 19332
rect 16578 19000 16634 19009
rect 16578 18935 16634 18944
rect 16396 18896 16448 18902
rect 16776 18873 16804 20198
rect 16396 18838 16448 18844
rect 16762 18864 16818 18873
rect 16762 18799 16818 18808
rect 16488 18692 16540 18698
rect 16488 18634 16540 18640
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 16212 18420 16264 18426
rect 16212 18362 16264 18368
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 16316 16980 16344 18566
rect 16500 18154 16528 18634
rect 16868 18442 16896 20198
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 16960 19854 16988 19994
rect 16948 19848 17000 19854
rect 16948 19790 17000 19796
rect 16960 19310 16988 19790
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 17038 19136 17094 19145
rect 17038 19071 17094 19080
rect 17052 18834 17080 19071
rect 17040 18828 17092 18834
rect 17040 18770 17092 18776
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16684 18414 16896 18442
rect 16488 18148 16540 18154
rect 16488 18090 16540 18096
rect 16394 17096 16450 17105
rect 16394 17031 16450 17040
rect 16132 16952 16344 16980
rect 16028 16720 16080 16726
rect 16028 16662 16080 16668
rect 16040 16250 16068 16662
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 15948 16017 15976 16050
rect 15934 16008 15990 16017
rect 15934 15943 15990 15952
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15856 15570 15884 15846
rect 15844 15564 15896 15570
rect 15844 15506 15896 15512
rect 15934 15192 15990 15201
rect 15934 15127 15990 15136
rect 15948 13870 15976 15127
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 16040 14278 16068 14554
rect 16132 14278 16160 16952
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16224 14482 16252 16730
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16316 15745 16344 15982
rect 16302 15736 16358 15745
rect 16302 15671 16358 15680
rect 16408 14618 16436 17031
rect 16500 16726 16528 18090
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16592 17542 16620 18022
rect 16684 17746 16712 18414
rect 16764 18216 16816 18222
rect 16960 18193 16988 18566
rect 17144 18426 17172 18702
rect 17132 18420 17184 18426
rect 17132 18362 17184 18368
rect 16764 18158 16816 18164
rect 16946 18184 17002 18193
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16592 17202 16620 17478
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16488 16720 16540 16726
rect 16488 16662 16540 16668
rect 16672 16516 16724 16522
rect 16672 16458 16724 16464
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 16224 14385 16252 14418
rect 16210 14376 16266 14385
rect 16210 14311 16266 14320
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 16132 14074 16160 14214
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16118 13968 16174 13977
rect 16118 13903 16174 13912
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15658 13152 15714 13161
rect 15658 13087 15714 13096
rect 15476 11892 15528 11898
rect 15528 11852 15608 11880
rect 15476 11834 15528 11840
rect 15474 11792 15530 11801
rect 15474 11727 15476 11736
rect 15528 11727 15530 11736
rect 15476 11698 15528 11704
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15304 9738 15332 9930
rect 15212 9710 15332 9738
rect 15212 9654 15240 9710
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15106 9344 15162 9353
rect 15106 9279 15162 9288
rect 15120 8634 15148 9279
rect 15212 8906 15240 9590
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15212 8514 15240 8842
rect 15120 8486 15240 8514
rect 14832 7948 14884 7954
rect 14832 7890 14884 7896
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 15120 7750 15148 8486
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15396 7886 15424 8230
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15108 7744 15160 7750
rect 15108 7686 15160 7692
rect 15120 7206 15148 7686
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15488 5642 15516 11494
rect 15580 11286 15608 11852
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15672 10577 15700 13087
rect 15948 12986 15976 13806
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 16026 12880 16082 12889
rect 16026 12815 16028 12824
rect 16080 12815 16082 12824
rect 16028 12786 16080 12792
rect 16132 12617 16160 13903
rect 16224 13326 16252 14214
rect 16394 13968 16450 13977
rect 16394 13903 16450 13912
rect 16408 13802 16436 13903
rect 16500 13802 16528 14758
rect 16684 14482 16712 16458
rect 16776 15162 16804 18158
rect 16946 18119 17002 18128
rect 17040 18148 17092 18154
rect 17040 18090 17092 18096
rect 17052 17066 17080 18090
rect 17040 17060 17092 17066
rect 17040 17002 17092 17008
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16960 16794 16988 16934
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 17130 16688 17186 16697
rect 17130 16623 17186 16632
rect 17144 15502 17172 16623
rect 17236 16250 17264 19314
rect 17328 18970 17356 20742
rect 17420 20466 17448 24006
rect 17592 23316 17644 23322
rect 17592 23258 17644 23264
rect 17500 23044 17552 23050
rect 17500 22986 17552 22992
rect 17512 22030 17540 22986
rect 17604 22982 17632 23258
rect 17592 22976 17644 22982
rect 17592 22918 17644 22924
rect 17776 22976 17828 22982
rect 17776 22918 17828 22924
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17788 21894 17816 22918
rect 17880 22760 17908 26302
rect 18326 26200 18382 27000
rect 18970 26200 19026 27000
rect 19614 26200 19670 27000
rect 20258 26200 20314 27000
rect 20902 26200 20958 27000
rect 21546 26330 21602 27000
rect 21192 26302 21602 26330
rect 18340 24274 18368 26200
rect 18328 24268 18380 24274
rect 18328 24210 18380 24216
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18984 23798 19012 26200
rect 19628 24970 19656 26200
rect 19352 24942 19656 24970
rect 19352 24290 19380 24942
rect 19432 24812 19484 24818
rect 19432 24754 19484 24760
rect 19444 24342 19472 24754
rect 19616 24608 19668 24614
rect 19616 24550 19668 24556
rect 19260 24274 19380 24290
rect 19432 24336 19484 24342
rect 19432 24278 19484 24284
rect 19248 24268 19380 24274
rect 19300 24262 19380 24268
rect 19248 24210 19300 24216
rect 19628 24206 19656 24550
rect 19616 24200 19668 24206
rect 19616 24142 19668 24148
rect 19156 24064 19208 24070
rect 19156 24006 19208 24012
rect 18972 23792 19024 23798
rect 18972 23734 19024 23740
rect 18788 23724 18840 23730
rect 18788 23666 18840 23672
rect 18328 23656 18380 23662
rect 18328 23598 18380 23604
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17880 22732 18184 22760
rect 17868 22432 17920 22438
rect 17868 22374 17920 22380
rect 17880 21978 17908 22374
rect 18052 22024 18104 22030
rect 17880 21972 18052 21978
rect 17880 21966 18104 21972
rect 17880 21950 18092 21966
rect 18156 21962 18184 22732
rect 18144 21956 18196 21962
rect 17776 21888 17828 21894
rect 17776 21830 17828 21836
rect 17880 21434 17908 21950
rect 18144 21898 18196 21904
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17960 21480 18012 21486
rect 17788 21428 17960 21434
rect 17788 21422 18012 21428
rect 17788 21406 18000 21422
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 17512 21010 17540 21286
rect 17590 21040 17646 21049
rect 17500 21004 17552 21010
rect 17590 20975 17646 20984
rect 17500 20946 17552 20952
rect 17408 20460 17460 20466
rect 17408 20402 17460 20408
rect 17604 19802 17632 20975
rect 17788 20398 17816 21406
rect 18340 21078 18368 23598
rect 18604 23248 18656 23254
rect 18604 23190 18656 23196
rect 18420 23044 18472 23050
rect 18420 22986 18472 22992
rect 18432 22710 18460 22986
rect 18616 22778 18644 23190
rect 18800 23186 18828 23666
rect 19168 23662 19196 24006
rect 19156 23656 19208 23662
rect 19156 23598 19208 23604
rect 19062 23488 19118 23497
rect 19062 23423 19118 23432
rect 18788 23180 18840 23186
rect 18788 23122 18840 23128
rect 19076 22778 19104 23423
rect 19628 23322 19656 24142
rect 20272 24138 20300 26200
rect 20536 24744 20588 24750
rect 20536 24686 20588 24692
rect 20260 24132 20312 24138
rect 20260 24074 20312 24080
rect 20548 23882 20576 24686
rect 20916 24274 20944 26200
rect 21192 24857 21220 26302
rect 21546 26200 21602 26302
rect 22190 26200 22246 27000
rect 22834 26200 22890 27000
rect 23478 26200 23534 27000
rect 24122 26330 24178 27000
rect 23952 26302 24178 26330
rect 24676 26376 24728 26382
rect 24676 26318 24728 26324
rect 21270 25528 21326 25537
rect 21270 25463 21326 25472
rect 21178 24848 21234 24857
rect 21178 24783 21234 24792
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20272 23866 20576 23882
rect 19708 23860 19760 23866
rect 19708 23802 19760 23808
rect 20272 23860 20588 23866
rect 20272 23854 20536 23860
rect 19720 23322 19748 23802
rect 20166 23352 20222 23361
rect 19616 23316 19668 23322
rect 19616 23258 19668 23264
rect 19708 23316 19760 23322
rect 20166 23287 20222 23296
rect 19708 23258 19760 23264
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 18604 22772 18656 22778
rect 18604 22714 18656 22720
rect 19064 22772 19116 22778
rect 19064 22714 19116 22720
rect 18420 22704 18472 22710
rect 18420 22646 18472 22652
rect 18432 22234 18460 22646
rect 18420 22228 18472 22234
rect 18420 22170 18472 22176
rect 18328 21072 18380 21078
rect 18328 21014 18380 21020
rect 17958 20904 18014 20913
rect 17958 20839 17960 20848
rect 18012 20839 18014 20848
rect 17960 20810 18012 20816
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18432 20466 18460 22170
rect 18616 22001 18644 22714
rect 19524 22704 19576 22710
rect 19904 22681 19932 23054
rect 20180 22681 20208 23287
rect 19524 22646 19576 22652
rect 19890 22672 19946 22681
rect 19432 22568 19484 22574
rect 19432 22510 19484 22516
rect 18788 22500 18840 22506
rect 18788 22442 18840 22448
rect 18602 21992 18658 22001
rect 18602 21927 18658 21936
rect 18800 21010 18828 22442
rect 19444 22094 19472 22510
rect 19352 22066 19472 22094
rect 19352 22030 19380 22066
rect 19340 22024 19392 22030
rect 18878 21992 18934 22001
rect 19340 21966 19392 21972
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 18878 21927 18934 21936
rect 18892 21049 18920 21927
rect 19444 21894 19472 21966
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 18878 21040 18934 21049
rect 18788 21004 18840 21010
rect 18878 20975 18934 20984
rect 19338 21040 19394 21049
rect 19338 20975 19394 20984
rect 18788 20946 18840 20952
rect 18604 20800 18656 20806
rect 18604 20742 18656 20748
rect 18420 20460 18472 20466
rect 18420 20402 18472 20408
rect 17776 20392 17828 20398
rect 17776 20334 17828 20340
rect 17788 19922 17816 20334
rect 18328 20256 18380 20262
rect 18328 20198 18380 20204
rect 17776 19916 17828 19922
rect 17776 19858 17828 19864
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17512 19774 17632 19802
rect 17316 18964 17368 18970
rect 17316 18906 17368 18912
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17420 17377 17448 18022
rect 17406 17368 17462 17377
rect 17406 17303 17462 17312
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17420 16726 17448 17070
rect 17408 16720 17460 16726
rect 17408 16662 17460 16668
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17132 15496 17184 15502
rect 17132 15438 17184 15444
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16762 14920 16818 14929
rect 16762 14855 16818 14864
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16578 14104 16634 14113
rect 16578 14039 16634 14048
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16488 13796 16540 13802
rect 16488 13738 16540 13744
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 16118 12608 16174 12617
rect 16118 12543 16174 12552
rect 16026 12200 16082 12209
rect 16026 12135 16082 12144
rect 16040 12102 16068 12135
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15658 10568 15714 10577
rect 15658 10503 15714 10512
rect 15764 8634 15792 10950
rect 15842 10296 15898 10305
rect 15842 10231 15898 10240
rect 15856 9654 15884 10231
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 15948 8634 15976 12038
rect 16040 11286 16068 12038
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 16132 11218 16160 12543
rect 16316 12434 16344 13670
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16500 12782 16528 13262
rect 16592 13258 16620 14039
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16580 12912 16632 12918
rect 16580 12854 16632 12860
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16592 12714 16620 12854
rect 16580 12708 16632 12714
rect 16580 12650 16632 12656
rect 16316 12406 16436 12434
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16224 11354 16252 11494
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 16040 7954 16068 8774
rect 16132 8430 16160 11018
rect 16408 10606 16436 12406
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16500 11898 16528 12174
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16592 11778 16620 11834
rect 16500 11750 16620 11778
rect 16500 11354 16528 11750
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16396 10600 16448 10606
rect 16396 10542 16448 10548
rect 16224 9722 16252 10542
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 16040 7478 16068 7890
rect 16316 7546 16344 10066
rect 16408 9994 16436 10542
rect 16500 10266 16528 10610
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16500 10169 16528 10202
rect 16486 10160 16542 10169
rect 16486 10095 16542 10104
rect 16396 9988 16448 9994
rect 16396 9930 16448 9936
rect 16488 9988 16540 9994
rect 16488 9930 16540 9936
rect 16500 9674 16528 9930
rect 16408 9646 16528 9674
rect 16592 9654 16620 10610
rect 16776 10538 16804 14855
rect 16868 14822 16896 15302
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 17144 14958 17172 15098
rect 17132 14952 17184 14958
rect 17132 14894 17184 14900
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16960 14414 16988 14554
rect 17040 14476 17092 14482
rect 17040 14418 17092 14424
rect 16948 14408 17000 14414
rect 16854 14376 16910 14385
rect 16948 14350 17000 14356
rect 16854 14311 16910 14320
rect 16868 13546 16896 14311
rect 16960 13734 16988 14350
rect 16948 13728 17000 13734
rect 16948 13670 17000 13676
rect 16868 13518 16988 13546
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16868 12850 16896 12922
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16868 11762 16896 12786
rect 16960 12306 16988 13518
rect 17052 12918 17080 14418
rect 17144 14278 17172 14894
rect 17236 14414 17264 15846
rect 17512 15688 17540 19774
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17604 19310 17632 19654
rect 17788 19378 17816 19858
rect 17880 19446 17908 19858
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17868 19440 17920 19446
rect 17868 19382 17920 19388
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17592 19304 17644 19310
rect 18340 19281 18368 20198
rect 18432 19854 18460 20402
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 17592 19246 17644 19252
rect 18326 19272 18382 19281
rect 18326 19207 18382 19216
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 17696 18902 17724 19110
rect 17684 18896 17736 18902
rect 17684 18838 17736 18844
rect 17868 18692 17920 18698
rect 17868 18634 17920 18640
rect 17880 18426 17908 18634
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17868 18420 17920 18426
rect 18432 18408 18460 19790
rect 18616 19786 18644 20742
rect 19352 20618 19380 20975
rect 19076 20602 19380 20618
rect 19064 20596 19380 20602
rect 19116 20590 19380 20596
rect 19064 20538 19116 20544
rect 19536 20058 19564 22646
rect 19890 22607 19946 22616
rect 20166 22672 20222 22681
rect 20166 22607 20222 22616
rect 20272 22094 20300 23854
rect 20536 23802 20588 23808
rect 21284 23798 21312 25463
rect 21732 24404 21784 24410
rect 21732 24346 21784 24352
rect 20352 23792 20404 23798
rect 20352 23734 20404 23740
rect 20996 23792 21048 23798
rect 20996 23734 21048 23740
rect 21272 23792 21324 23798
rect 21272 23734 21324 23740
rect 21640 23792 21692 23798
rect 21640 23734 21692 23740
rect 20364 22930 20392 23734
rect 20628 23520 20680 23526
rect 20628 23462 20680 23468
rect 20640 23050 20668 23462
rect 20628 23044 20680 23050
rect 20628 22986 20680 22992
rect 20720 23044 20772 23050
rect 20720 22986 20772 22992
rect 20732 22930 20760 22986
rect 20364 22902 20760 22930
rect 20364 22710 20392 22902
rect 20352 22704 20404 22710
rect 20352 22646 20404 22652
rect 20352 22094 20404 22098
rect 20272 22092 20404 22094
rect 20272 22066 20352 22092
rect 20352 22034 20404 22040
rect 20444 22092 20496 22098
rect 20444 22034 20496 22040
rect 20628 22092 20680 22098
rect 20628 22034 20680 22040
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 19996 21185 20024 21830
rect 20088 21622 20116 21966
rect 20168 21956 20220 21962
rect 20168 21898 20220 21904
rect 20076 21616 20128 21622
rect 20076 21558 20128 21564
rect 20088 21418 20116 21558
rect 20180 21486 20208 21898
rect 20456 21622 20484 22034
rect 20640 21690 20668 22034
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 20628 21684 20680 21690
rect 20628 21626 20680 21632
rect 20444 21616 20496 21622
rect 20444 21558 20496 21564
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 20076 21412 20128 21418
rect 20076 21354 20128 21360
rect 19982 21176 20038 21185
rect 19982 21111 20038 21120
rect 19614 20768 19670 20777
rect 19614 20703 19670 20712
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 18604 19780 18656 19786
rect 18604 19722 18656 19728
rect 18604 19440 18656 19446
rect 18604 19382 18656 19388
rect 18694 19408 18750 19417
rect 17868 18362 17920 18368
rect 18340 18380 18460 18408
rect 18510 18456 18566 18465
rect 18510 18391 18566 18400
rect 17684 18216 17736 18222
rect 17684 18158 17736 18164
rect 17696 17338 17724 18158
rect 18340 17746 18368 18380
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 18328 17740 18380 17746
rect 18328 17682 18380 17688
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17684 17332 17736 17338
rect 17684 17274 17736 17280
rect 17774 17232 17830 17241
rect 17774 17167 17830 17176
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17420 15660 17540 15688
rect 17316 15088 17368 15094
rect 17420 15076 17448 15660
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 17368 15048 17448 15076
rect 17316 15030 17368 15036
rect 17328 14822 17356 15030
rect 17512 14822 17540 15506
rect 17604 15366 17632 16730
rect 17682 16144 17738 16153
rect 17682 16079 17684 16088
rect 17736 16079 17738 16088
rect 17684 16050 17736 16056
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17500 14816 17552 14822
rect 17500 14758 17552 14764
rect 17408 14476 17460 14482
rect 17512 14464 17540 14758
rect 17460 14436 17540 14464
rect 17408 14418 17460 14424
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 17222 14240 17278 14249
rect 17222 14175 17278 14184
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17144 13161 17172 13874
rect 17130 13152 17186 13161
rect 17130 13087 17186 13096
rect 17236 13002 17264 14175
rect 17328 13938 17356 14350
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17420 14074 17448 14214
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17604 13977 17632 15302
rect 17696 14521 17724 15438
rect 17682 14512 17738 14521
rect 17682 14447 17738 14456
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17696 14006 17724 14350
rect 17788 14249 17816 17167
rect 17880 17134 17908 17614
rect 18328 17604 18380 17610
rect 18328 17546 18380 17552
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 18340 16522 18368 17546
rect 18328 16516 18380 16522
rect 18328 16458 18380 16464
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17880 14958 17908 15846
rect 17972 15638 18000 15846
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17868 14340 17920 14346
rect 17868 14282 17920 14288
rect 17774 14240 17830 14249
rect 17774 14175 17830 14184
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17684 14000 17736 14006
rect 17590 13968 17646 13977
rect 17316 13932 17368 13938
rect 17684 13942 17736 13948
rect 17590 13903 17646 13912
rect 17316 13874 17368 13880
rect 17406 13832 17462 13841
rect 17406 13767 17462 13776
rect 17314 13560 17370 13569
rect 17314 13495 17370 13504
rect 17328 13394 17356 13495
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17144 12974 17264 13002
rect 17040 12912 17092 12918
rect 17040 12854 17092 12860
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 17144 12102 17172 12974
rect 17420 12434 17448 13767
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17328 12406 17448 12434
rect 17222 12200 17278 12209
rect 17222 12135 17278 12144
rect 17236 12102 17264 12135
rect 17132 12096 17184 12102
rect 17130 12064 17132 12073
rect 17224 12096 17276 12102
rect 17184 12064 17186 12073
rect 17224 12038 17276 12044
rect 17130 11999 17186 12008
rect 17236 11937 17264 12038
rect 17222 11928 17278 11937
rect 17222 11863 17278 11872
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16946 11656 17002 11665
rect 16946 11591 17002 11600
rect 16960 11354 16988 11591
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16672 10532 16724 10538
rect 16672 10474 16724 10480
rect 16764 10532 16816 10538
rect 16764 10474 16816 10480
rect 16684 10266 16712 10474
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16776 9674 16804 9998
rect 16580 9648 16632 9654
rect 16408 8634 16436 9646
rect 16776 9646 16896 9674
rect 16580 9590 16632 9596
rect 16868 9518 16896 9646
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 16868 9382 16896 9454
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16868 8974 16896 9318
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16408 8294 16436 8570
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16028 7472 16080 7478
rect 16028 7414 16080 7420
rect 16408 7206 16436 8230
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16408 6662 16436 7142
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 15476 5636 15528 5642
rect 15476 5578 15528 5584
rect 15384 3664 15436 3670
rect 15384 3606 15436 3612
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 13832 800 13860 2450
rect 15396 2446 15424 3606
rect 16120 3120 16172 3126
rect 16120 3062 16172 3068
rect 16132 2774 16160 3062
rect 16408 3058 16436 6598
rect 16500 4146 16528 8774
rect 16868 8498 16896 8910
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16578 8256 16634 8265
rect 16578 8191 16634 8200
rect 16592 8090 16620 8191
rect 17144 8090 17172 9454
rect 17236 8566 17264 10202
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17328 7342 17356 12406
rect 17512 12170 17540 13330
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17500 12164 17552 12170
rect 17500 12106 17552 12112
rect 17500 11008 17552 11014
rect 17500 10950 17552 10956
rect 17512 9994 17540 10950
rect 17604 10470 17632 13126
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 17500 9988 17552 9994
rect 17552 9948 17632 9976
rect 17500 9930 17552 9936
rect 17604 9654 17632 9948
rect 17592 9648 17644 9654
rect 17592 9590 17644 9596
rect 17696 9518 17724 12242
rect 17788 10742 17816 14010
rect 17880 13988 17908 14282
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17880 13960 18000 13988
rect 17972 13326 18000 13960
rect 18144 13864 18196 13870
rect 18144 13806 18196 13812
rect 18156 13462 18184 13806
rect 18144 13456 18196 13462
rect 18144 13398 18196 13404
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17776 10736 17828 10742
rect 17776 10678 17828 10684
rect 17684 9512 17736 9518
rect 17684 9454 17736 9460
rect 17880 9382 17908 12106
rect 18248 12084 18276 12786
rect 18340 12238 18368 16458
rect 18432 15706 18460 18226
rect 18524 18057 18552 18391
rect 18616 18222 18644 19382
rect 18694 19343 18750 19352
rect 19432 19372 19484 19378
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18510 18048 18566 18057
rect 18510 17983 18566 17992
rect 18616 17746 18644 18158
rect 18512 17740 18564 17746
rect 18512 17682 18564 17688
rect 18604 17740 18656 17746
rect 18604 17682 18656 17688
rect 18524 17202 18552 17682
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 18616 16998 18644 17682
rect 18604 16992 18656 16998
rect 18604 16934 18656 16940
rect 18616 16114 18644 16934
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18604 15972 18656 15978
rect 18604 15914 18656 15920
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 18420 15428 18472 15434
rect 18420 15370 18472 15376
rect 18432 14890 18460 15370
rect 18420 14884 18472 14890
rect 18420 14826 18472 14832
rect 18420 14544 18472 14550
rect 18420 14486 18472 14492
rect 18432 13326 18460 14486
rect 18524 14006 18552 15846
rect 18616 15706 18644 15914
rect 18604 15700 18656 15706
rect 18604 15642 18656 15648
rect 18708 15162 18736 19343
rect 19432 19314 19484 19320
rect 19444 18766 19472 19314
rect 19628 18850 19656 20703
rect 20088 20534 20116 21354
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20260 20868 20312 20874
rect 20260 20810 20312 20816
rect 20076 20528 20128 20534
rect 20076 20470 20128 20476
rect 19800 20392 19852 20398
rect 19800 20334 19852 20340
rect 19706 20088 19762 20097
rect 19706 20023 19762 20032
rect 19536 18822 19656 18850
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19260 18630 19288 18702
rect 19248 18624 19300 18630
rect 19248 18566 19300 18572
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19260 18290 19288 18566
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19154 18048 19210 18057
rect 19154 17983 19210 17992
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18984 17338 19012 17478
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 18878 15736 18934 15745
rect 18878 15671 18934 15680
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18892 14958 18920 15671
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18602 14512 18658 14521
rect 18708 14482 18736 14554
rect 18602 14447 18604 14456
rect 18656 14447 18658 14456
rect 18696 14476 18748 14482
rect 18604 14418 18656 14424
rect 18696 14418 18748 14424
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18800 13841 18828 14894
rect 18878 14784 18934 14793
rect 18878 14719 18934 14728
rect 18892 14113 18920 14719
rect 18878 14104 18934 14113
rect 18878 14039 18934 14048
rect 18786 13832 18842 13841
rect 18786 13767 18842 13776
rect 18604 13456 18656 13462
rect 18604 13398 18656 13404
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18616 12782 18644 13398
rect 18892 12866 18920 14039
rect 18800 12838 18920 12866
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 18248 12056 18368 12084
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18236 11756 18288 11762
rect 18340 11744 18368 12056
rect 18288 11716 18368 11744
rect 18236 11698 18288 11704
rect 18248 11014 18276 11698
rect 18328 11620 18380 11626
rect 18328 11562 18380 11568
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18340 10810 18368 11562
rect 18328 10804 18380 10810
rect 18328 10746 18380 10752
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17408 8900 17460 8906
rect 17408 8842 17460 8848
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17420 6866 17448 8842
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17604 8566 17632 8774
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17776 7744 17828 7750
rect 17776 7686 17828 7692
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17788 6662 17816 7686
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 17788 4078 17816 6598
rect 17880 6322 17908 7958
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18340 7546 18368 10406
rect 18432 7954 18460 12582
rect 18604 12436 18656 12442
rect 18604 12378 18656 12384
rect 18616 11529 18644 12378
rect 18602 11520 18658 11529
rect 18602 11455 18658 11464
rect 18616 11218 18644 11455
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18512 11144 18564 11150
rect 18510 11112 18512 11121
rect 18564 11112 18566 11121
rect 18510 11047 18566 11056
rect 18800 10810 18828 12838
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18604 10736 18656 10742
rect 18604 10678 18656 10684
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18524 7954 18552 10066
rect 18616 10062 18644 10678
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18604 10056 18656 10062
rect 18602 10024 18604 10033
rect 18656 10024 18658 10033
rect 18602 9959 18658 9968
rect 18708 8634 18736 10610
rect 18892 10606 18920 12718
rect 18984 11150 19012 15438
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 19076 14385 19104 14418
rect 19062 14376 19118 14385
rect 19062 14311 19118 14320
rect 19168 14278 19196 17983
rect 19352 17898 19380 18566
rect 19260 17870 19380 17898
rect 19260 16794 19288 17870
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19352 17202 19380 17682
rect 19536 17678 19564 18822
rect 19616 18760 19668 18766
rect 19614 18728 19616 18737
rect 19668 18728 19670 18737
rect 19614 18663 19670 18672
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19260 16522 19288 16730
rect 19430 16552 19486 16561
rect 19248 16516 19300 16522
rect 19430 16487 19486 16496
rect 19248 16458 19300 16464
rect 19444 16454 19472 16487
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19260 15434 19288 16186
rect 19352 16046 19380 16390
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19338 15736 19394 15745
rect 19338 15671 19394 15680
rect 19352 15570 19380 15671
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 19168 13784 19196 14214
rect 19076 13756 19196 13784
rect 19076 13462 19104 13756
rect 19154 13696 19210 13705
rect 19154 13631 19210 13640
rect 19064 13456 19116 13462
rect 19064 13398 19116 13404
rect 19064 13252 19116 13258
rect 19064 13194 19116 13200
rect 19076 11354 19104 13194
rect 19168 12714 19196 13631
rect 19260 13530 19288 15370
rect 19522 15192 19578 15201
rect 19522 15127 19578 15136
rect 19536 13938 19564 15127
rect 19720 14278 19748 20023
rect 19812 19990 19840 20334
rect 19800 19984 19852 19990
rect 19800 19926 19852 19932
rect 19812 17241 19840 19926
rect 19892 19780 19944 19786
rect 19892 19722 19944 19728
rect 19904 18902 19932 19722
rect 20088 19310 20116 20470
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19892 18896 19944 18902
rect 19892 18838 19944 18844
rect 19904 18737 19932 18838
rect 19890 18728 19946 18737
rect 19890 18663 19946 18672
rect 19996 18358 20024 18906
rect 19984 18352 20036 18358
rect 20088 18340 20116 19246
rect 20168 18352 20220 18358
rect 20088 18312 20168 18340
rect 19984 18294 20036 18300
rect 20168 18294 20220 18300
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 19904 17882 19932 18158
rect 19892 17876 19944 17882
rect 19892 17818 19944 17824
rect 20180 17649 20208 18294
rect 20272 17882 20300 20810
rect 20364 20777 20392 21286
rect 20350 20768 20406 20777
rect 20350 20703 20406 20712
rect 20456 20602 20484 21558
rect 20628 21480 20680 21486
rect 20628 21422 20680 21428
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 20548 21146 20576 21286
rect 20640 21146 20668 21422
rect 20536 21140 20588 21146
rect 20536 21082 20588 21088
rect 20628 21140 20680 21146
rect 20628 21082 20680 21088
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 20352 20528 20404 20534
rect 20352 20470 20404 20476
rect 20364 20262 20392 20470
rect 20352 20256 20404 20262
rect 20352 20198 20404 20204
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20166 17640 20222 17649
rect 20364 17610 20392 20198
rect 20444 19848 20496 19854
rect 20444 19790 20496 19796
rect 20456 17746 20484 19790
rect 20536 19440 20588 19446
rect 20536 19382 20588 19388
rect 20444 17740 20496 17746
rect 20444 17682 20496 17688
rect 20166 17575 20222 17584
rect 20352 17604 20404 17610
rect 20180 17270 20208 17575
rect 20352 17546 20404 17552
rect 20168 17264 20220 17270
rect 19798 17232 19854 17241
rect 20168 17206 20220 17212
rect 19798 17167 19854 17176
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 19800 16448 19852 16454
rect 19800 16390 19852 16396
rect 19812 15162 19840 16390
rect 20088 16250 20116 17070
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20180 16726 20208 16934
rect 20168 16720 20220 16726
rect 20168 16662 20220 16668
rect 20076 16244 20128 16250
rect 20076 16186 20128 16192
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19800 15156 19852 15162
rect 19800 15098 19852 15104
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19812 14550 19840 14962
rect 19800 14544 19852 14550
rect 19800 14486 19852 14492
rect 19708 14272 19760 14278
rect 19708 14214 19760 14220
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 19616 13864 19668 13870
rect 19616 13806 19668 13812
rect 19708 13864 19760 13870
rect 19708 13806 19760 13812
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19628 13326 19656 13806
rect 19616 13320 19668 13326
rect 19616 13262 19668 13268
rect 19720 12986 19748 13806
rect 19812 13394 19840 14486
rect 19904 13530 19932 15302
rect 20088 14958 20116 16186
rect 20352 15564 20404 15570
rect 20352 15506 20404 15512
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 19996 13530 20024 14894
rect 20364 14414 20392 15506
rect 20548 15366 20576 19382
rect 20640 18834 20668 21082
rect 20732 20602 20760 21898
rect 21008 21321 21036 23734
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 21088 23044 21140 23050
rect 21088 22986 21140 22992
rect 21100 22710 21128 22986
rect 21088 22704 21140 22710
rect 21088 22646 21140 22652
rect 21192 22642 21220 23122
rect 21180 22636 21232 22642
rect 21180 22578 21232 22584
rect 21192 22030 21220 22578
rect 21652 22234 21680 23734
rect 21640 22228 21692 22234
rect 21640 22170 21692 22176
rect 21180 22024 21232 22030
rect 21180 21966 21232 21972
rect 20994 21312 21050 21321
rect 20994 21247 21050 21256
rect 21192 21010 21220 21966
rect 21744 21865 21772 24346
rect 22008 23112 22060 23118
rect 22008 23054 22060 23060
rect 21824 22704 21876 22710
rect 21824 22646 21876 22652
rect 21836 22234 21864 22646
rect 22020 22642 22048 23054
rect 22100 22976 22152 22982
rect 22098 22944 22100 22953
rect 22152 22944 22154 22953
rect 22098 22879 22154 22888
rect 22008 22636 22060 22642
rect 22008 22578 22060 22584
rect 21824 22228 21876 22234
rect 21824 22170 21876 22176
rect 21836 22094 21864 22170
rect 21836 22066 21956 22094
rect 21730 21856 21786 21865
rect 21730 21791 21786 21800
rect 21270 21720 21326 21729
rect 21270 21655 21326 21664
rect 21284 21554 21312 21655
rect 21928 21554 21956 22066
rect 22020 21554 22048 22578
rect 22112 22438 22140 22879
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 21272 21548 21324 21554
rect 21272 21490 21324 21496
rect 21548 21548 21600 21554
rect 21548 21490 21600 21496
rect 21916 21548 21968 21554
rect 21916 21490 21968 21496
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 21560 21146 21588 21490
rect 21928 21350 21956 21490
rect 22098 21448 22154 21457
rect 22098 21383 22154 21392
rect 22112 21350 22140 21383
rect 21916 21344 21968 21350
rect 21916 21286 21968 21292
rect 22100 21344 22152 21350
rect 22100 21286 22152 21292
rect 21548 21140 21600 21146
rect 21548 21082 21600 21088
rect 21454 21040 21510 21049
rect 21180 21004 21232 21010
rect 21928 21010 21956 21286
rect 22112 21185 22140 21286
rect 22098 21176 22154 21185
rect 22098 21111 22154 21120
rect 21454 20975 21510 20984
rect 21732 21004 21784 21010
rect 21180 20946 21232 20952
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 21100 20262 21128 20402
rect 21180 20392 21232 20398
rect 21468 20369 21496 20975
rect 21732 20946 21784 20952
rect 21916 21004 21968 21010
rect 21916 20946 21968 20952
rect 21180 20334 21232 20340
rect 21454 20360 21510 20369
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 20996 19780 21048 19786
rect 20996 19722 21048 19728
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20732 16522 20760 19314
rect 21008 19310 21036 19722
rect 20996 19304 21048 19310
rect 20996 19246 21048 19252
rect 20812 18624 20864 18630
rect 20812 18566 20864 18572
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20824 15706 20852 18566
rect 20902 17640 20958 17649
rect 20902 17575 20904 17584
rect 20956 17575 20958 17584
rect 20904 17546 20956 17552
rect 20916 17270 20944 17546
rect 20904 17264 20956 17270
rect 20904 17206 20956 17212
rect 20916 16726 20944 17206
rect 20904 16720 20956 16726
rect 20904 16662 20956 16668
rect 20916 16522 20944 16662
rect 20904 16516 20956 16522
rect 20904 16458 20956 16464
rect 20916 16182 20944 16458
rect 20904 16176 20956 16182
rect 20904 16118 20956 16124
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20916 15570 20944 16118
rect 21008 15910 21036 19246
rect 21088 17740 21140 17746
rect 21088 17682 21140 17688
rect 21100 16658 21128 17682
rect 21192 17241 21220 20334
rect 21510 20318 21588 20346
rect 21454 20295 21510 20304
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 21284 19514 21312 19994
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 21284 18358 21312 18702
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 21468 18426 21496 18566
rect 21456 18420 21508 18426
rect 21456 18362 21508 18368
rect 21272 18352 21324 18358
rect 21272 18294 21324 18300
rect 21364 17536 21416 17542
rect 21364 17478 21416 17484
rect 21178 17232 21234 17241
rect 21178 17167 21234 17176
rect 21088 16652 21140 16658
rect 21088 16594 21140 16600
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20536 15360 20588 15366
rect 20456 15320 20536 15348
rect 20456 14822 20484 15320
rect 20536 15302 20588 15308
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 20088 13734 20116 14214
rect 20076 13728 20128 13734
rect 20076 13670 20128 13676
rect 19892 13524 19944 13530
rect 19892 13466 19944 13472
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 19800 13388 19852 13394
rect 19800 13330 19852 13336
rect 20088 13190 20116 13670
rect 20076 13184 20128 13190
rect 20076 13126 20128 13132
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 19708 12980 19760 12986
rect 19708 12922 19760 12928
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19156 12708 19208 12714
rect 19156 12650 19208 12656
rect 19432 12164 19484 12170
rect 19432 12106 19484 12112
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18800 9178 18828 10542
rect 18892 10130 18920 10542
rect 18972 10260 19024 10266
rect 18972 10202 19024 10208
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 18512 7948 18564 7954
rect 18512 7890 18564 7896
rect 18616 7886 18644 8298
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18616 7426 18644 7686
rect 18708 7546 18736 8026
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18616 7398 18736 7426
rect 18708 7206 18736 7398
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18708 7002 18736 7142
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 18708 6458 18736 6938
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18800 6322 18828 9114
rect 18880 8424 18932 8430
rect 18880 8366 18932 8372
rect 18892 6662 18920 8366
rect 18984 7342 19012 10202
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 19076 8838 19104 9658
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 19076 6798 19104 8774
rect 19260 7546 19288 11630
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19352 9926 19380 11494
rect 19444 10266 19472 12106
rect 19432 10260 19484 10266
rect 19432 10202 19484 10208
rect 19536 10130 19564 12786
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19628 10810 19656 12718
rect 19720 12306 19748 12922
rect 20272 12646 20300 13126
rect 20260 12640 20312 12646
rect 20258 12608 20260 12617
rect 20312 12608 20314 12617
rect 20258 12543 20314 12552
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 19890 11928 19946 11937
rect 20548 11898 20576 14962
rect 20732 14074 20760 15098
rect 20904 14952 20956 14958
rect 20904 14894 20956 14900
rect 20916 14278 20944 14894
rect 21100 14482 21128 16594
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 21088 14476 21140 14482
rect 21088 14418 21140 14424
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20626 12744 20682 12753
rect 20626 12679 20628 12688
rect 20680 12679 20682 12688
rect 20628 12650 20680 12656
rect 20916 12434 20944 14214
rect 21008 14074 21036 14350
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 20916 12406 21036 12434
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 19890 11863 19946 11872
rect 20076 11892 20128 11898
rect 19904 11694 19932 11863
rect 20076 11834 20128 11840
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 19892 11688 19944 11694
rect 19812 11648 19892 11676
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19720 11218 19748 11494
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19616 10804 19668 10810
rect 19616 10746 19668 10752
rect 19812 10198 19840 11648
rect 19892 11630 19944 11636
rect 20088 11626 20116 11834
rect 20824 11830 20852 12242
rect 20812 11824 20864 11830
rect 20812 11766 20864 11772
rect 20168 11688 20220 11694
rect 21008 11665 21036 12406
rect 20168 11630 20220 11636
rect 20994 11656 21050 11665
rect 20076 11620 20128 11626
rect 20076 11562 20128 11568
rect 20180 11354 20208 11630
rect 20994 11591 21050 11600
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20076 11280 20128 11286
rect 20076 11222 20128 11228
rect 19890 10840 19946 10849
rect 19890 10775 19946 10784
rect 19904 10674 19932 10775
rect 19892 10668 19944 10674
rect 19892 10610 19944 10616
rect 19904 10305 19932 10610
rect 19890 10296 19946 10305
rect 19890 10231 19946 10240
rect 19800 10192 19852 10198
rect 19800 10134 19852 10140
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19616 9512 19668 9518
rect 19616 9454 19668 9460
rect 19708 9512 19760 9518
rect 19708 9454 19760 9460
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 19444 8634 19472 8910
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 18880 6656 18932 6662
rect 18880 6598 18932 6604
rect 19444 6322 19472 7686
rect 19524 7268 19576 7274
rect 19524 7210 19576 7216
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 19352 4486 19380 5510
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 16488 4004 16540 4010
rect 16488 3946 16540 3952
rect 16500 3534 16528 3946
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 17236 3194 17264 3538
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 15948 2746 16160 2774
rect 15384 2440 15436 2446
rect 15384 2382 15436 2388
rect 15948 800 15976 2746
rect 16408 2650 16436 2994
rect 19444 2854 19472 3470
rect 19536 3058 19564 7210
rect 19628 6458 19656 9454
rect 19720 9178 19748 9454
rect 19708 9172 19760 9178
rect 19708 9114 19760 9120
rect 19892 9172 19944 9178
rect 19892 9114 19944 9120
rect 19708 8900 19760 8906
rect 19708 8842 19760 8848
rect 19720 6866 19748 8842
rect 19904 8838 19932 9114
rect 20088 8838 20116 11222
rect 20628 11212 20680 11218
rect 20628 11154 20680 11160
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20364 9722 20484 9738
rect 20364 9716 20496 9722
rect 20364 9710 20444 9716
rect 20364 9654 20392 9710
rect 20444 9658 20496 9664
rect 20352 9648 20404 9654
rect 20404 9596 20484 9602
rect 20352 9590 20484 9596
rect 20364 9574 20484 9590
rect 20456 8906 20484 9574
rect 20548 8945 20576 10610
rect 20640 10130 20668 11154
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 20812 11008 20864 11014
rect 20812 10950 20864 10956
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20732 10713 20760 10746
rect 20718 10704 20774 10713
rect 20718 10639 20774 10648
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 20534 8936 20590 8945
rect 20444 8900 20496 8906
rect 20534 8871 20590 8880
rect 20444 8842 20496 8848
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 20076 8832 20128 8838
rect 20076 8774 20128 8780
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19812 7478 19840 7686
rect 19800 7472 19852 7478
rect 19800 7414 19852 7420
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 20088 6798 20116 8774
rect 20456 8566 20484 8842
rect 20640 8634 20668 10066
rect 20824 9178 20852 10950
rect 20916 10810 20944 11018
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 21008 10674 21036 11591
rect 21100 11082 21128 13874
rect 21192 12918 21220 15098
rect 21284 14958 21312 15302
rect 21272 14952 21324 14958
rect 21272 14894 21324 14900
rect 21376 13530 21404 17478
rect 21560 16182 21588 20318
rect 21744 19854 21772 20946
rect 22006 20632 22062 20641
rect 22006 20567 22008 20576
rect 22060 20567 22062 20576
rect 22008 20538 22060 20544
rect 21824 19984 21876 19990
rect 21824 19926 21876 19932
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21732 19712 21784 19718
rect 21732 19654 21784 19660
rect 21744 19514 21772 19654
rect 21732 19508 21784 19514
rect 21732 19450 21784 19456
rect 21836 19378 21864 19926
rect 22100 19780 22152 19786
rect 22100 19722 22152 19728
rect 22008 19712 22060 19718
rect 22008 19654 22060 19660
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 22020 19310 22048 19654
rect 22112 19378 22140 19722
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22008 19304 22060 19310
rect 22008 19246 22060 19252
rect 22006 19000 22062 19009
rect 22006 18935 22062 18944
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 21732 18624 21784 18630
rect 21732 18566 21784 18572
rect 21744 18086 21772 18566
rect 21732 18080 21784 18086
rect 21732 18022 21784 18028
rect 21548 16176 21600 16182
rect 21548 16118 21600 16124
rect 21560 15450 21588 16118
rect 21744 15570 21772 18022
rect 21928 17542 21956 18770
rect 22020 18086 22048 18935
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 21916 17536 21968 17542
rect 21916 17478 21968 17484
rect 21928 15638 21956 17478
rect 22020 17066 22048 17614
rect 22008 17060 22060 17066
rect 22008 17002 22060 17008
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 22020 15638 22048 16050
rect 21916 15632 21968 15638
rect 21916 15574 21968 15580
rect 22008 15632 22060 15638
rect 22008 15574 22060 15580
rect 21732 15564 21784 15570
rect 21732 15506 21784 15512
rect 21468 15422 21588 15450
rect 21468 15026 21496 15422
rect 21548 15360 21600 15366
rect 21548 15302 21600 15308
rect 21640 15360 21692 15366
rect 21640 15302 21692 15308
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21364 13524 21416 13530
rect 21364 13466 21416 13472
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21284 13161 21312 13262
rect 21270 13152 21326 13161
rect 21270 13087 21326 13096
rect 21180 12912 21232 12918
rect 21180 12854 21232 12860
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 21192 12170 21220 12718
rect 21272 12708 21324 12714
rect 21272 12650 21324 12656
rect 21284 12238 21312 12650
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21180 12164 21232 12170
rect 21180 12106 21232 12112
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 21284 11694 21312 12038
rect 21376 11694 21404 13330
rect 21468 12102 21496 14758
rect 21560 12918 21588 15302
rect 21652 15162 21680 15302
rect 21640 15156 21692 15162
rect 21640 15098 21692 15104
rect 21652 14929 21680 15098
rect 21732 15088 21784 15094
rect 21732 15030 21784 15036
rect 21638 14920 21694 14929
rect 21638 14855 21694 14864
rect 21744 14618 21772 15030
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 21732 14476 21784 14482
rect 21732 14418 21784 14424
rect 21744 14278 21772 14418
rect 21916 14340 21968 14346
rect 21916 14282 21968 14288
rect 21732 14272 21784 14278
rect 21732 14214 21784 14220
rect 21928 13870 21956 14282
rect 21916 13864 21968 13870
rect 21916 13806 21968 13812
rect 22112 13326 22140 19314
rect 22204 17202 22232 26200
rect 22468 25356 22520 25362
rect 22468 25298 22520 25304
rect 22284 24404 22336 24410
rect 22284 24346 22336 24352
rect 22296 23866 22324 24346
rect 22376 24336 22428 24342
rect 22376 24278 22428 24284
rect 22388 23866 22416 24278
rect 22480 23866 22508 25298
rect 22560 24200 22612 24206
rect 22612 24148 22784 24154
rect 22560 24142 22784 24148
rect 22572 24138 22784 24142
rect 22572 24132 22796 24138
rect 22572 24126 22744 24132
rect 22744 24074 22796 24080
rect 22284 23860 22336 23866
rect 22284 23802 22336 23808
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22468 23860 22520 23866
rect 22468 23802 22520 23808
rect 22480 23497 22508 23802
rect 22742 23760 22798 23769
rect 22742 23695 22798 23704
rect 22560 23656 22612 23662
rect 22560 23598 22612 23604
rect 22466 23488 22522 23497
rect 22466 23423 22522 23432
rect 22572 23322 22600 23598
rect 22560 23316 22612 23322
rect 22560 23258 22612 23264
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 22480 22098 22508 22918
rect 22652 22568 22704 22574
rect 22652 22510 22704 22516
rect 22664 22166 22692 22510
rect 22756 22438 22784 23695
rect 22848 23089 22876 26200
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23388 24268 23440 24274
rect 23388 24210 23440 24216
rect 23296 23520 23348 23526
rect 23296 23462 23348 23468
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23112 23180 23164 23186
rect 23112 23122 23164 23128
rect 22834 23080 22890 23089
rect 22834 23015 22890 23024
rect 23124 22953 23152 23122
rect 23110 22944 23166 22953
rect 23110 22879 23166 22888
rect 23308 22710 23336 23462
rect 23400 23254 23428 24210
rect 23388 23248 23440 23254
rect 23388 23190 23440 23196
rect 23296 22704 23348 22710
rect 23492 22692 23520 26200
rect 23572 23860 23624 23866
rect 23572 23802 23624 23808
rect 23584 23225 23612 23802
rect 23664 23656 23716 23662
rect 23716 23604 23888 23610
rect 23664 23598 23888 23604
rect 23676 23582 23888 23598
rect 23570 23216 23626 23225
rect 23570 23151 23626 23160
rect 23664 23180 23716 23186
rect 23664 23122 23716 23128
rect 23572 22704 23624 22710
rect 23492 22664 23572 22692
rect 23296 22646 23348 22652
rect 23572 22646 23624 22652
rect 22744 22432 22796 22438
rect 22744 22374 22796 22380
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 22652 22160 22704 22166
rect 22652 22102 22704 22108
rect 22834 22128 22890 22137
rect 22468 22092 22520 22098
rect 22468 22034 22520 22040
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 22296 21146 22324 21626
rect 22376 21412 22428 21418
rect 22376 21354 22428 21360
rect 22388 21321 22416 21354
rect 22374 21312 22430 21321
rect 22374 21247 22430 21256
rect 22284 21140 22336 21146
rect 22284 21082 22336 21088
rect 22560 20800 22612 20806
rect 22560 20742 22612 20748
rect 22468 20528 22520 20534
rect 22468 20470 22520 20476
rect 22480 19854 22508 20470
rect 22468 19848 22520 19854
rect 22468 19790 22520 19796
rect 22468 19712 22520 19718
rect 22468 19654 22520 19660
rect 22480 19378 22508 19654
rect 22468 19372 22520 19378
rect 22468 19314 22520 19320
rect 22376 19236 22428 19242
rect 22376 19178 22428 19184
rect 22388 18970 22416 19178
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 22296 17746 22324 18702
rect 22284 17740 22336 17746
rect 22284 17682 22336 17688
rect 22296 17202 22324 17682
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 22376 17128 22428 17134
rect 22376 17070 22428 17076
rect 22388 16454 22416 17070
rect 22376 16448 22428 16454
rect 22376 16390 22428 16396
rect 22284 15904 22336 15910
rect 22284 15846 22336 15852
rect 22296 14006 22324 15846
rect 22376 15632 22428 15638
rect 22374 15600 22376 15609
rect 22428 15600 22430 15609
rect 22374 15535 22430 15544
rect 22480 15484 22508 19314
rect 22572 18630 22600 20742
rect 22664 19310 22692 22102
rect 22744 22092 22796 22098
rect 23308 22094 23336 22646
rect 22834 22063 22890 22072
rect 23216 22066 23428 22094
rect 22744 22034 22796 22040
rect 22756 21010 22784 22034
rect 22848 21078 22876 22063
rect 23216 22030 23244 22066
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 23296 22024 23348 22030
rect 23296 21966 23348 21972
rect 23020 21888 23072 21894
rect 23020 21830 23072 21836
rect 23032 21622 23060 21830
rect 23020 21616 23072 21622
rect 23020 21558 23072 21564
rect 23308 21486 23336 21966
rect 23400 21622 23428 22066
rect 23388 21616 23440 21622
rect 23388 21558 23440 21564
rect 23296 21480 23348 21486
rect 23296 21422 23348 21428
rect 23400 21434 23428 21558
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22836 21072 22888 21078
rect 22836 21014 22888 21020
rect 22744 21004 22796 21010
rect 22744 20946 22796 20952
rect 22836 20936 22888 20942
rect 22834 20904 22836 20913
rect 22888 20904 22890 20913
rect 22744 20868 22796 20874
rect 22834 20839 22890 20848
rect 22744 20810 22796 20816
rect 22756 20602 22784 20810
rect 23308 20806 23336 21422
rect 23400 21406 23520 21434
rect 23296 20800 23348 20806
rect 23296 20742 23348 20748
rect 22744 20596 22796 20602
rect 22744 20538 22796 20544
rect 23492 20466 23520 21406
rect 23676 20890 23704 23122
rect 23860 23118 23888 23582
rect 23848 23112 23900 23118
rect 23846 23080 23848 23089
rect 23900 23080 23902 23089
rect 23846 23015 23902 23024
rect 23756 22976 23808 22982
rect 23756 22918 23808 22924
rect 23768 22234 23796 22918
rect 23952 22545 23980 26302
rect 24122 26200 24178 26302
rect 24688 26160 24716 26318
rect 24766 26200 24822 27000
rect 25410 26200 25466 27000
rect 26054 26330 26110 27000
rect 25792 26302 26110 26330
rect 24780 26160 24808 26200
rect 24688 26132 24808 26160
rect 25228 25764 25280 25770
rect 25228 25706 25280 25712
rect 24032 25560 24084 25566
rect 24032 25502 24084 25508
rect 24044 24206 24072 25502
rect 24860 24404 24912 24410
rect 24860 24346 24912 24352
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 24872 24313 24900 24346
rect 24858 24304 24914 24313
rect 24858 24239 24914 24248
rect 24032 24200 24084 24206
rect 24032 24142 24084 24148
rect 24044 23050 24072 24142
rect 24676 23860 24728 23866
rect 24676 23802 24728 23808
rect 24124 23724 24176 23730
rect 24124 23666 24176 23672
rect 24136 23497 24164 23666
rect 24122 23488 24178 23497
rect 24122 23423 24178 23432
rect 24032 23044 24084 23050
rect 24032 22986 24084 22992
rect 24216 23044 24268 23050
rect 24216 22986 24268 22992
rect 24124 22568 24176 22574
rect 23938 22536 23994 22545
rect 24124 22510 24176 22516
rect 23938 22471 23994 22480
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23754 21176 23810 21185
rect 23754 21111 23810 21120
rect 23768 21010 23796 21111
rect 23756 21004 23808 21010
rect 23756 20946 23808 20952
rect 23848 21004 23900 21010
rect 23848 20946 23900 20952
rect 23676 20862 23796 20890
rect 23664 20800 23716 20806
rect 23662 20768 23664 20777
rect 23716 20768 23718 20777
rect 23662 20703 23718 20712
rect 22836 20460 22888 20466
rect 22836 20402 22888 20408
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 22652 19304 22704 19310
rect 22652 19246 22704 19252
rect 22742 19272 22798 19281
rect 22742 19207 22798 19216
rect 22560 18624 22612 18630
rect 22560 18566 22612 18572
rect 22756 16658 22784 19207
rect 22848 17814 22876 20402
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23296 19780 23348 19786
rect 23296 19722 23348 19728
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23204 18352 23256 18358
rect 23204 18294 23256 18300
rect 23216 18086 23244 18294
rect 23308 18290 23336 19722
rect 23400 19378 23428 20334
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23492 19334 23520 20402
rect 23768 20398 23796 20862
rect 23860 20641 23888 20946
rect 23846 20632 23902 20641
rect 23846 20567 23902 20576
rect 24136 20398 24164 22510
rect 24228 22098 24256 22986
rect 24400 22704 24452 22710
rect 24452 22664 24624 22692
rect 24400 22646 24452 22652
rect 24596 22574 24624 22664
rect 24308 22568 24360 22574
rect 24308 22510 24360 22516
rect 24584 22568 24636 22574
rect 24584 22510 24636 22516
rect 24216 22092 24268 22098
rect 24216 22034 24268 22040
rect 24320 21894 24348 22510
rect 24584 22432 24636 22438
rect 24584 22374 24636 22380
rect 24596 22137 24624 22374
rect 24582 22128 24638 22137
rect 24582 22063 24638 22072
rect 24688 22094 24716 23802
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 24872 22642 24900 23598
rect 25148 22778 25176 24346
rect 25136 22772 25188 22778
rect 25136 22714 25188 22720
rect 24860 22636 24912 22642
rect 24860 22578 24912 22584
rect 24872 22216 24900 22578
rect 25136 22228 25188 22234
rect 24872 22188 25136 22216
rect 25136 22170 25188 22176
rect 25134 22128 25190 22137
rect 24688 22066 25084 22094
rect 24308 21888 24360 21894
rect 24308 21830 24360 21836
rect 23756 20392 23808 20398
rect 23756 20334 23808 20340
rect 24124 20392 24176 20398
rect 24124 20334 24176 20340
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 23756 19916 23808 19922
rect 23756 19858 23808 19864
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23584 19514 23612 19654
rect 23572 19508 23624 19514
rect 23572 19450 23624 19456
rect 23400 18630 23428 19314
rect 23492 19306 23612 19334
rect 23480 19168 23532 19174
rect 23478 19136 23480 19145
rect 23532 19136 23534 19145
rect 23478 19071 23534 19080
rect 23584 18766 23612 19306
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 23400 18358 23428 18566
rect 23388 18352 23440 18358
rect 23388 18294 23440 18300
rect 23296 18284 23348 18290
rect 23296 18226 23348 18232
rect 23204 18080 23256 18086
rect 23204 18022 23256 18028
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22836 17808 22888 17814
rect 22836 17750 22888 17756
rect 23308 17610 23336 18226
rect 23296 17604 23348 17610
rect 23296 17546 23348 17552
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23308 16794 23336 17546
rect 23296 16788 23348 16794
rect 23296 16730 23348 16736
rect 22744 16652 22796 16658
rect 22744 16594 22796 16600
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22652 15904 22704 15910
rect 22652 15846 22704 15852
rect 22572 15638 22600 15846
rect 22664 15706 22692 15846
rect 22652 15700 22704 15706
rect 22652 15642 22704 15648
rect 22560 15632 22612 15638
rect 22560 15574 22612 15580
rect 22388 15456 22508 15484
rect 22560 15496 22612 15502
rect 22388 14226 22416 15456
rect 22560 15438 22612 15444
rect 22466 14240 22522 14249
rect 22388 14198 22466 14226
rect 22466 14175 22522 14184
rect 22284 14000 22336 14006
rect 22204 13948 22284 13954
rect 22204 13942 22336 13948
rect 22204 13926 22324 13942
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 21640 13184 21692 13190
rect 21638 13152 21640 13161
rect 21692 13152 21694 13161
rect 21638 13087 21694 13096
rect 21548 12912 21600 12918
rect 21600 12860 21680 12866
rect 21548 12854 21680 12860
rect 21560 12838 21680 12854
rect 21546 12608 21602 12617
rect 21546 12543 21602 12552
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21088 11076 21140 11082
rect 21088 11018 21140 11024
rect 21100 10674 21128 11018
rect 20996 10668 21048 10674
rect 20996 10610 21048 10616
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 21100 9994 21128 10610
rect 21180 10600 21232 10606
rect 21180 10542 21232 10548
rect 21088 9988 21140 9994
rect 21088 9930 21140 9936
rect 21100 9722 21128 9930
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21100 9586 21128 9658
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 21192 9382 21220 10542
rect 21284 9382 21312 11630
rect 21456 10736 21508 10742
rect 21456 10678 21508 10684
rect 21468 9926 21496 10678
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21456 9920 21508 9926
rect 21456 9862 21508 9868
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 20812 9172 20864 9178
rect 20812 9114 20864 9120
rect 20996 8832 21048 8838
rect 20996 8774 21048 8780
rect 21008 8634 21036 8774
rect 20628 8628 20680 8634
rect 20996 8628 21048 8634
rect 20680 8588 20760 8616
rect 20628 8570 20680 8576
rect 20444 8560 20496 8566
rect 20444 8502 20496 8508
rect 20456 8242 20484 8502
rect 20364 8214 20484 8242
rect 20364 8090 20392 8214
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 20364 7546 20392 8026
rect 20732 7954 20760 8588
rect 20996 8570 21048 8576
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20364 7002 20392 7482
rect 20824 7410 20852 8026
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 20916 7478 20944 7686
rect 20904 7472 20956 7478
rect 20904 7414 20956 7420
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20352 6996 20404 7002
rect 20352 6938 20404 6944
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 19800 3596 19852 3602
rect 19800 3538 19852 3544
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 19812 2990 19840 3538
rect 19800 2984 19852 2990
rect 19800 2926 19852 2932
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 18328 2372 18380 2378
rect 18328 2314 18380 2320
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 1122 0 1178 800
rect 3238 0 3294 800
rect 5354 0 5410 800
rect 7470 0 7526 800
rect 9586 0 9642 800
rect 11702 0 11758 800
rect 13818 0 13874 800
rect 15934 0 15990 800
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18340 762 18368 2314
rect 20180 800 20208 4014
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20732 3670 20760 3878
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 20916 2582 20944 7414
rect 21192 6798 21220 9318
rect 21272 8832 21324 8838
rect 21272 8774 21324 8780
rect 21284 7818 21312 8774
rect 21272 7812 21324 7818
rect 21272 7754 21324 7760
rect 21376 6866 21404 9862
rect 21560 8974 21588 12543
rect 21652 12442 21680 12838
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 21640 12164 21692 12170
rect 21640 12106 21692 12112
rect 21652 11014 21680 12106
rect 21640 11008 21692 11014
rect 21640 10950 21692 10956
rect 21548 8968 21600 8974
rect 21548 8910 21600 8916
rect 21560 8430 21588 8910
rect 21456 8424 21508 8430
rect 21548 8424 21600 8430
rect 21456 8366 21508 8372
rect 21546 8392 21548 8401
rect 21600 8392 21602 8401
rect 21468 7546 21496 8366
rect 21546 8327 21602 8336
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21652 7342 21680 10950
rect 21836 10282 21864 12582
rect 21744 10254 21864 10282
rect 21744 10198 21772 10254
rect 21732 10192 21784 10198
rect 21732 10134 21784 10140
rect 21744 7410 21772 10134
rect 21928 9586 21956 12786
rect 22008 12776 22060 12782
rect 22008 12718 22060 12724
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 22020 11898 22048 12718
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 22112 11830 22140 12718
rect 22100 11824 22152 11830
rect 22100 11766 22152 11772
rect 22100 11552 22152 11558
rect 22204 11540 22232 13926
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 22152 11512 22232 11540
rect 22100 11494 22152 11500
rect 22190 10704 22246 10713
rect 22296 10690 22324 13126
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22388 11937 22416 12786
rect 22480 12646 22508 14175
rect 22468 12640 22520 12646
rect 22468 12582 22520 12588
rect 22572 12442 22600 15438
rect 22652 14544 22704 14550
rect 22652 14486 22704 14492
rect 22664 12986 22692 14486
rect 22756 14482 22784 16594
rect 23768 16522 23796 19858
rect 23860 18358 23888 20198
rect 24136 19990 24164 20334
rect 23940 19984 23992 19990
rect 23940 19926 23992 19932
rect 24124 19984 24176 19990
rect 24124 19926 24176 19932
rect 23952 18850 23980 19926
rect 24032 19440 24084 19446
rect 24032 19382 24084 19388
rect 24044 18970 24072 19382
rect 24032 18964 24084 18970
rect 24032 18906 24084 18912
rect 23952 18822 24072 18850
rect 24044 18766 24072 18822
rect 23940 18760 23992 18766
rect 23940 18702 23992 18708
rect 24032 18760 24084 18766
rect 24032 18702 24084 18708
rect 23848 18352 23900 18358
rect 23848 18294 23900 18300
rect 23952 17184 23980 18702
rect 24044 18630 24072 18702
rect 24032 18624 24084 18630
rect 24032 18566 24084 18572
rect 24032 17196 24084 17202
rect 23952 17156 24032 17184
rect 24032 17138 24084 17144
rect 23938 16960 23994 16969
rect 23938 16895 23994 16904
rect 23952 16726 23980 16895
rect 24044 16726 24072 17138
rect 23940 16720 23992 16726
rect 23846 16688 23902 16697
rect 23940 16662 23992 16668
rect 24032 16720 24084 16726
rect 24032 16662 24084 16668
rect 23846 16623 23902 16632
rect 23756 16516 23808 16522
rect 23756 16458 23808 16464
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23480 16448 23532 16454
rect 23480 16390 23532 16396
rect 22848 16250 22876 16390
rect 22836 16244 22888 16250
rect 22836 16186 22888 16192
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22834 15464 22890 15473
rect 22834 15399 22890 15408
rect 22744 14476 22796 14482
rect 22744 14418 22796 14424
rect 22756 13258 22784 14418
rect 22744 13252 22796 13258
rect 22744 13194 22796 13200
rect 22652 12980 22704 12986
rect 22652 12922 22704 12928
rect 22848 12850 22876 15399
rect 23308 15201 23336 16390
rect 23388 15564 23440 15570
rect 23388 15506 23440 15512
rect 23294 15192 23350 15201
rect 23294 15127 23350 15136
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 23020 14340 23072 14346
rect 23020 14282 23072 14288
rect 23032 13870 23060 14282
rect 23296 14272 23348 14278
rect 23400 14260 23428 15506
rect 23492 15162 23520 16390
rect 23664 16176 23716 16182
rect 23664 16118 23716 16124
rect 23572 16040 23624 16046
rect 23572 15982 23624 15988
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23480 14612 23532 14618
rect 23480 14554 23532 14560
rect 23492 14346 23520 14554
rect 23480 14340 23532 14346
rect 23480 14282 23532 14288
rect 23348 14232 23428 14260
rect 23296 14214 23348 14220
rect 23400 14090 23428 14232
rect 23296 14068 23348 14074
rect 23400 14062 23520 14090
rect 23296 14010 23348 14016
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23112 13456 23164 13462
rect 23110 13424 23112 13433
rect 23164 13424 23166 13433
rect 23110 13359 23166 13368
rect 23204 13184 23256 13190
rect 23204 13126 23256 13132
rect 23308 13138 23336 14010
rect 23492 13870 23520 14062
rect 23480 13864 23532 13870
rect 23480 13806 23532 13812
rect 22836 12844 22888 12850
rect 23216 12832 23244 13126
rect 23308 13110 23428 13138
rect 23400 12832 23428 13110
rect 23584 12986 23612 15982
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23480 12844 23532 12850
rect 23216 12804 23336 12832
rect 22836 12786 22888 12792
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 22744 12300 22796 12306
rect 22744 12242 22796 12248
rect 22468 12096 22520 12102
rect 22468 12038 22520 12044
rect 22560 12096 22612 12102
rect 22560 12038 22612 12044
rect 22374 11928 22430 11937
rect 22374 11863 22376 11872
rect 22428 11863 22430 11872
rect 22376 11834 22428 11840
rect 22480 11218 22508 12038
rect 22572 11626 22600 12038
rect 22652 11756 22704 11762
rect 22652 11698 22704 11704
rect 22560 11620 22612 11626
rect 22560 11562 22612 11568
rect 22664 11506 22692 11698
rect 22756 11694 22784 12242
rect 22744 11688 22796 11694
rect 22744 11630 22796 11636
rect 22572 11478 22692 11506
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 22296 10662 22416 10690
rect 22190 10639 22246 10648
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 22020 10130 22048 10542
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 21824 9580 21876 9586
rect 21824 9522 21876 9528
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21836 9466 21864 9522
rect 22020 9466 22048 9862
rect 22204 9518 22232 10639
rect 22388 10606 22416 10662
rect 22284 10600 22336 10606
rect 22284 10542 22336 10548
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 21836 9438 22048 9466
rect 22192 9512 22244 9518
rect 22192 9454 22244 9460
rect 21824 9376 21876 9382
rect 21824 9318 21876 9324
rect 21836 9194 21864 9318
rect 21836 9166 21956 9194
rect 21824 9104 21876 9110
rect 21824 9046 21876 9052
rect 21836 8090 21864 9046
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21732 7404 21784 7410
rect 21732 7346 21784 7352
rect 21640 7336 21692 7342
rect 21640 7278 21692 7284
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 21180 6180 21232 6186
rect 21180 6122 21232 6128
rect 21192 3602 21220 6122
rect 21928 3670 21956 9166
rect 22100 8424 22152 8430
rect 22020 8372 22100 8378
rect 22020 8366 22152 8372
rect 22020 8350 22140 8366
rect 22020 7954 22048 8350
rect 22008 7948 22060 7954
rect 22008 7890 22060 7896
rect 22020 4078 22048 7890
rect 22296 7546 22324 10542
rect 22572 10266 22600 11478
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22572 9994 22600 10202
rect 22560 9988 22612 9994
rect 22560 9930 22612 9936
rect 22376 9580 22428 9586
rect 22376 9522 22428 9528
rect 22388 9110 22416 9522
rect 22468 9512 22520 9518
rect 22468 9454 22520 9460
rect 22376 9104 22428 9110
rect 22480 9081 22508 9454
rect 22560 9376 22612 9382
rect 22560 9318 22612 9324
rect 22376 9046 22428 9052
rect 22466 9072 22522 9081
rect 22466 9007 22522 9016
rect 22376 8968 22428 8974
rect 22376 8910 22428 8916
rect 22388 8634 22416 8910
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 22388 4826 22416 8570
rect 22480 7478 22508 9007
rect 22572 8906 22600 9318
rect 22664 9178 22692 10746
rect 22744 10464 22796 10470
rect 22744 10406 22796 10412
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 22560 8900 22612 8906
rect 22560 8842 22612 8848
rect 22756 8634 22784 10406
rect 22848 10062 22876 12582
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23308 11354 23336 12804
rect 23400 12804 23480 12832
rect 23400 11830 23428 12804
rect 23480 12786 23532 12792
rect 23676 12374 23704 16118
rect 23860 15502 23888 16623
rect 23940 15904 23992 15910
rect 24044 15892 24072 16662
rect 23992 15864 24072 15892
rect 23940 15846 23992 15852
rect 23848 15496 23900 15502
rect 23848 15438 23900 15444
rect 23756 14816 23808 14822
rect 23756 14758 23808 14764
rect 23768 14618 23796 14758
rect 23756 14612 23808 14618
rect 23756 14554 23808 14560
rect 23952 14414 23980 15846
rect 24136 14890 24164 19926
rect 24214 17368 24270 17377
rect 24214 17303 24216 17312
rect 24268 17303 24270 17312
rect 24216 17274 24268 17280
rect 24320 17105 24348 21830
rect 24596 21049 24624 22063
rect 25056 22030 25084 22066
rect 25240 22094 25268 25706
rect 25424 24682 25452 26200
rect 25504 24812 25556 24818
rect 25504 24754 25556 24760
rect 25412 24676 25464 24682
rect 25412 24618 25464 24624
rect 25320 22976 25372 22982
rect 25320 22918 25372 22924
rect 25190 22072 25268 22094
rect 25134 22066 25268 22072
rect 25134 22063 25190 22066
rect 25044 22024 25096 22030
rect 25044 21966 25096 21972
rect 25148 21690 25176 22063
rect 25136 21684 25188 21690
rect 25136 21626 25188 21632
rect 25228 21480 25280 21486
rect 25228 21422 25280 21428
rect 24768 21344 24820 21350
rect 24768 21286 24820 21292
rect 24780 21146 24808 21286
rect 24768 21140 24820 21146
rect 24768 21082 24820 21088
rect 24582 21040 24638 21049
rect 24582 20975 24638 20984
rect 24768 20936 24820 20942
rect 25240 20890 25268 21422
rect 24768 20878 24820 20884
rect 24400 20528 24452 20534
rect 24400 20470 24452 20476
rect 24584 20528 24636 20534
rect 24584 20470 24636 20476
rect 24412 19446 24440 20470
rect 24596 20398 24624 20470
rect 24584 20392 24636 20398
rect 24584 20334 24636 20340
rect 24674 20088 24730 20097
rect 24674 20023 24730 20032
rect 24688 19854 24716 20023
rect 24676 19848 24728 19854
rect 24676 19790 24728 19796
rect 24492 19712 24544 19718
rect 24490 19680 24492 19689
rect 24544 19680 24546 19689
rect 24490 19615 24546 19624
rect 24400 19440 24452 19446
rect 24400 19382 24452 19388
rect 24676 18624 24728 18630
rect 24676 18566 24728 18572
rect 24584 18148 24636 18154
rect 24584 18090 24636 18096
rect 24596 17882 24624 18090
rect 24492 17876 24544 17882
rect 24492 17818 24544 17824
rect 24584 17876 24636 17882
rect 24584 17818 24636 17824
rect 24306 17096 24362 17105
rect 24504 17066 24532 17818
rect 24306 17031 24362 17040
rect 24492 17060 24544 17066
rect 24492 17002 24544 17008
rect 24308 16448 24360 16454
rect 24308 16390 24360 16396
rect 24124 14884 24176 14890
rect 24124 14826 24176 14832
rect 23940 14408 23992 14414
rect 23940 14350 23992 14356
rect 24032 14408 24084 14414
rect 24032 14350 24084 14356
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23860 13530 23888 14214
rect 24044 14074 24072 14350
rect 24216 14272 24268 14278
rect 24216 14214 24268 14220
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 23848 13524 23900 13530
rect 23848 13466 23900 13472
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23768 12986 23796 13330
rect 23756 12980 23808 12986
rect 23756 12922 23808 12928
rect 23860 12918 23888 13466
rect 23848 12912 23900 12918
rect 23848 12854 23900 12860
rect 23664 12368 23716 12374
rect 23664 12310 23716 12316
rect 23754 12200 23810 12209
rect 23754 12135 23810 12144
rect 23388 11824 23440 11830
rect 23388 11766 23440 11772
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23572 11280 23624 11286
rect 23572 11222 23624 11228
rect 23294 11112 23350 11121
rect 23294 11047 23350 11056
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23308 10248 23336 11047
rect 23584 10810 23612 11222
rect 23768 11121 23796 12135
rect 24044 11218 24072 14010
rect 24228 12918 24256 14214
rect 24124 12912 24176 12918
rect 24124 12854 24176 12860
rect 24216 12912 24268 12918
rect 24216 12854 24268 12860
rect 24136 12434 24164 12854
rect 24136 12406 24256 12434
rect 24032 11212 24084 11218
rect 24032 11154 24084 11160
rect 23754 11112 23810 11121
rect 23754 11047 23756 11056
rect 23808 11047 23810 11056
rect 23756 11018 23808 11024
rect 23572 10804 23624 10810
rect 23572 10746 23624 10752
rect 23124 10220 23336 10248
rect 22836 10056 22888 10062
rect 22836 9998 22888 10004
rect 23124 9654 23152 10220
rect 23296 10124 23348 10130
rect 23296 10066 23348 10072
rect 23112 9648 23164 9654
rect 23112 9590 23164 9596
rect 23308 9586 23336 10066
rect 23388 9716 23440 9722
rect 23388 9658 23440 9664
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 23400 9489 23428 9658
rect 23480 9512 23532 9518
rect 23386 9480 23442 9489
rect 23584 9466 23612 10746
rect 24032 10736 24084 10742
rect 24032 10678 24084 10684
rect 24044 9926 24072 10678
rect 24124 9988 24176 9994
rect 24124 9930 24176 9936
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 23756 9648 23808 9654
rect 23756 9590 23808 9596
rect 23768 9466 23796 9590
rect 23532 9460 23612 9466
rect 23480 9454 23612 9460
rect 23492 9438 23612 9454
rect 23676 9438 23796 9466
rect 23386 9415 23442 9424
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 23572 9172 23624 9178
rect 23572 9114 23624 9120
rect 23584 8974 23612 9114
rect 23480 8968 23532 8974
rect 23478 8936 23480 8945
rect 23572 8968 23624 8974
rect 23532 8936 23534 8945
rect 23572 8910 23624 8916
rect 23676 8906 23704 9438
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 23860 9042 23888 9318
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23478 8871 23534 8880
rect 23664 8900 23716 8906
rect 23664 8842 23716 8848
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 22468 7472 22520 7478
rect 22468 7414 22520 7420
rect 22756 7410 22784 8570
rect 23676 8566 23704 8842
rect 23664 8560 23716 8566
rect 23664 8502 23716 8508
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23676 7750 23704 8502
rect 23860 7886 23888 8978
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 23664 7744 23716 7750
rect 23664 7686 23716 7692
rect 23308 7546 23336 7686
rect 23296 7540 23348 7546
rect 23296 7482 23348 7488
rect 22744 7404 22796 7410
rect 22744 7346 22796 7352
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22744 6112 22796 6118
rect 22744 6054 22796 6060
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 22468 4616 22520 4622
rect 22468 4558 22520 4564
rect 22652 4616 22704 4622
rect 22652 4558 22704 4564
rect 22008 4072 22060 4078
rect 22008 4014 22060 4020
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 21916 3664 21968 3670
rect 21916 3606 21968 3612
rect 21180 3596 21232 3602
rect 21180 3538 21232 3544
rect 20996 2848 21048 2854
rect 20996 2790 21048 2796
rect 21008 2650 21036 2790
rect 20996 2644 21048 2650
rect 20996 2586 21048 2592
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 22020 2514 22048 4014
rect 22296 3738 22324 4014
rect 22480 3942 22508 4558
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 22284 3732 22336 3738
rect 22284 3674 22336 3680
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 22112 3126 22140 3538
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 22284 2984 22336 2990
rect 22284 2926 22336 2932
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 22296 800 22324 2926
rect 22480 2106 22508 3878
rect 22664 2922 22692 4558
rect 22756 3058 22784 6054
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 23296 4616 23348 4622
rect 23296 4558 23348 4564
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 23308 3602 23336 4558
rect 23572 4548 23624 4554
rect 23572 4490 23624 4496
rect 23584 3602 23612 4490
rect 23676 4282 23704 7686
rect 24044 5574 24072 9862
rect 24136 9042 24164 9930
rect 24124 9036 24176 9042
rect 24124 8978 24176 8984
rect 24032 5568 24084 5574
rect 24032 5510 24084 5516
rect 24032 4480 24084 4486
rect 24032 4422 24084 4428
rect 23664 4276 23716 4282
rect 23664 4218 23716 4224
rect 24044 4214 24072 4422
rect 24032 4208 24084 4214
rect 24032 4150 24084 4156
rect 24228 4026 24256 12406
rect 24320 11150 24348 16390
rect 24688 16017 24716 18566
rect 24780 17814 24808 20878
rect 24872 20862 25268 20890
rect 24872 19530 24900 20862
rect 25136 20800 25188 20806
rect 25136 20742 25188 20748
rect 24950 19816 25006 19825
rect 24950 19751 25006 19760
rect 24964 19718 24992 19751
rect 24952 19712 25004 19718
rect 24952 19654 25004 19660
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 24872 19502 24992 19530
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 24768 17808 24820 17814
rect 24768 17750 24820 17756
rect 24780 17338 24808 17750
rect 24872 17338 24900 18226
rect 24964 17678 24992 19502
rect 25056 18834 25084 19654
rect 25148 18970 25176 20742
rect 25228 19916 25280 19922
rect 25228 19858 25280 19864
rect 25136 18964 25188 18970
rect 25136 18906 25188 18912
rect 25044 18828 25096 18834
rect 25044 18770 25096 18776
rect 25134 18456 25190 18465
rect 25134 18391 25136 18400
rect 25188 18391 25190 18400
rect 25136 18362 25188 18368
rect 25042 18320 25098 18329
rect 25042 18255 25044 18264
rect 25096 18255 25098 18264
rect 25044 18226 25096 18232
rect 25240 18222 25268 19858
rect 25332 19310 25360 22918
rect 25412 22092 25464 22098
rect 25412 22034 25464 22040
rect 25424 21894 25452 22034
rect 25412 21888 25464 21894
rect 25412 21830 25464 21836
rect 25424 20398 25452 21830
rect 25516 20534 25544 24754
rect 25792 24614 25820 26302
rect 26054 26200 26110 26302
rect 26698 26200 26754 27000
rect 27342 26330 27398 27000
rect 27986 26330 28042 27000
rect 28630 26330 28686 27000
rect 29274 26330 29330 27000
rect 29918 26330 29974 27000
rect 30562 26330 30618 27000
rect 31206 26330 31262 27000
rect 31482 26344 31538 26353
rect 27342 26302 27568 26330
rect 27342 26200 27398 26302
rect 27540 26246 27568 26302
rect 27986 26302 28488 26330
rect 27528 26240 27580 26246
rect 25872 25628 25924 25634
rect 25872 25570 25924 25576
rect 25780 24608 25832 24614
rect 25780 24550 25832 24556
rect 25778 23488 25834 23497
rect 25778 23423 25834 23432
rect 25596 23112 25648 23118
rect 25596 23054 25648 23060
rect 25608 21049 25636 23054
rect 25792 22166 25820 23423
rect 25780 22160 25832 22166
rect 25780 22102 25832 22108
rect 25594 21040 25650 21049
rect 25594 20975 25650 20984
rect 25504 20528 25556 20534
rect 25504 20470 25556 20476
rect 25608 20398 25636 20975
rect 25412 20392 25464 20398
rect 25412 20334 25464 20340
rect 25596 20392 25648 20398
rect 25596 20334 25648 20340
rect 25410 20088 25466 20097
rect 25410 20023 25466 20032
rect 25320 19304 25372 19310
rect 25320 19246 25372 19252
rect 25424 18630 25452 20023
rect 25504 19236 25556 19242
rect 25504 19178 25556 19184
rect 25412 18624 25464 18630
rect 25412 18566 25464 18572
rect 25516 18426 25544 19178
rect 25504 18420 25556 18426
rect 25504 18362 25556 18368
rect 25228 18216 25280 18222
rect 25228 18158 25280 18164
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 25056 17746 25084 18022
rect 25608 17746 25636 20334
rect 25792 20262 25820 22102
rect 25780 20256 25832 20262
rect 25780 20198 25832 20204
rect 25780 19712 25832 19718
rect 25780 19654 25832 19660
rect 25792 19446 25820 19654
rect 25780 19440 25832 19446
rect 25780 19382 25832 19388
rect 25688 19304 25740 19310
rect 25686 19272 25688 19281
rect 25740 19272 25742 19281
rect 25884 19242 25912 25570
rect 26608 24200 26660 24206
rect 26608 24142 26660 24148
rect 25964 24064 26016 24070
rect 25964 24006 26016 24012
rect 26516 24064 26568 24070
rect 26516 24006 26568 24012
rect 25976 23186 26004 24006
rect 26528 23798 26556 24006
rect 26516 23792 26568 23798
rect 26516 23734 26568 23740
rect 25964 23180 26016 23186
rect 25964 23122 26016 23128
rect 26424 22772 26476 22778
rect 26424 22714 26476 22720
rect 26148 22500 26200 22506
rect 26148 22442 26200 22448
rect 26160 22098 26188 22442
rect 26240 22432 26292 22438
rect 26240 22374 26292 22380
rect 26148 22092 26200 22098
rect 26148 22034 26200 22040
rect 26054 21584 26110 21593
rect 25964 21548 26016 21554
rect 26054 21519 26110 21528
rect 25964 21490 26016 21496
rect 25976 20602 26004 21490
rect 26068 20602 26096 21519
rect 26148 21412 26200 21418
rect 26148 21354 26200 21360
rect 26160 20806 26188 21354
rect 26252 21146 26280 22374
rect 26332 21888 26384 21894
rect 26436 21876 26464 22714
rect 26528 22710 26556 23734
rect 26620 23526 26648 24142
rect 26608 23520 26660 23526
rect 26608 23462 26660 23468
rect 26516 22704 26568 22710
rect 26712 22681 26740 26200
rect 27986 26200 28042 26302
rect 27528 26182 27580 26188
rect 28356 24744 28408 24750
rect 28356 24686 28408 24692
rect 27620 24336 27672 24342
rect 27620 24278 27672 24284
rect 27344 24200 27396 24206
rect 27344 24142 27396 24148
rect 26884 24132 26936 24138
rect 26884 24074 26936 24080
rect 26792 24064 26844 24070
rect 26792 24006 26844 24012
rect 26804 23866 26832 24006
rect 26792 23860 26844 23866
rect 26792 23802 26844 23808
rect 26896 22778 26924 24074
rect 26976 23112 27028 23118
rect 26976 23054 27028 23060
rect 26884 22772 26936 22778
rect 26884 22714 26936 22720
rect 26988 22710 27016 23054
rect 26976 22704 27028 22710
rect 26516 22646 26568 22652
rect 26698 22672 26754 22681
rect 26528 22506 26556 22646
rect 26976 22646 27028 22652
rect 26698 22607 26754 22616
rect 26516 22500 26568 22506
rect 26516 22442 26568 22448
rect 27252 22500 27304 22506
rect 27252 22442 27304 22448
rect 26608 22432 26660 22438
rect 26608 22374 26660 22380
rect 26620 22166 26648 22374
rect 27264 22234 27292 22442
rect 27356 22234 27384 24142
rect 27436 23724 27488 23730
rect 27436 23666 27488 23672
rect 27448 22982 27476 23666
rect 27528 23520 27580 23526
rect 27528 23462 27580 23468
rect 27436 22976 27488 22982
rect 27436 22918 27488 22924
rect 27448 22778 27476 22918
rect 27436 22772 27488 22778
rect 27436 22714 27488 22720
rect 27436 22636 27488 22642
rect 27436 22578 27488 22584
rect 27252 22228 27304 22234
rect 27252 22170 27304 22176
rect 27344 22228 27396 22234
rect 27344 22170 27396 22176
rect 26608 22160 26660 22166
rect 26608 22102 26660 22108
rect 26700 22160 26752 22166
rect 26700 22102 26752 22108
rect 26712 21978 26740 22102
rect 26384 21848 26464 21876
rect 26332 21830 26384 21836
rect 26240 21140 26292 21146
rect 26240 21082 26292 21088
rect 26148 20800 26200 20806
rect 26148 20742 26200 20748
rect 25964 20596 26016 20602
rect 25964 20538 26016 20544
rect 26056 20596 26108 20602
rect 26108 20556 26188 20584
rect 26056 20538 26108 20544
rect 25976 19378 26004 20538
rect 26056 20460 26108 20466
rect 26056 20402 26108 20408
rect 25964 19372 26016 19378
rect 26068 19360 26096 20402
rect 26160 19514 26188 20556
rect 26252 20466 26280 21082
rect 26330 21040 26386 21049
rect 26330 20975 26332 20984
rect 26384 20975 26386 20984
rect 26332 20946 26384 20952
rect 26332 20800 26384 20806
rect 26332 20742 26384 20748
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 26240 19712 26292 19718
rect 26238 19680 26240 19689
rect 26292 19680 26294 19689
rect 26238 19615 26294 19624
rect 26148 19508 26200 19514
rect 26200 19468 26280 19496
rect 26148 19450 26200 19456
rect 26068 19332 26188 19360
rect 25964 19314 26016 19320
rect 25686 19207 25742 19216
rect 25872 19236 25924 19242
rect 25872 19178 25924 19184
rect 25962 19000 26018 19009
rect 25962 18935 26018 18944
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 25596 17740 25648 17746
rect 25596 17682 25648 17688
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 25228 17672 25280 17678
rect 25228 17614 25280 17620
rect 25780 17672 25832 17678
rect 25780 17614 25832 17620
rect 25044 17536 25096 17542
rect 25044 17478 25096 17484
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 24860 17332 24912 17338
rect 24860 17274 24912 17280
rect 24952 17196 25004 17202
rect 24952 17138 25004 17144
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 24768 16176 24820 16182
rect 24872 16130 24900 16594
rect 24820 16124 24900 16130
rect 24768 16118 24900 16124
rect 24780 16102 24900 16118
rect 24674 16008 24730 16017
rect 24674 15943 24730 15952
rect 24400 15904 24452 15910
rect 24400 15846 24452 15852
rect 24412 14482 24440 15846
rect 24584 15632 24636 15638
rect 24490 15600 24546 15609
rect 24768 15632 24820 15638
rect 24636 15592 24768 15620
rect 24584 15574 24636 15580
rect 24768 15574 24820 15580
rect 24490 15535 24546 15544
rect 24504 15026 24532 15535
rect 24492 15020 24544 15026
rect 24492 14962 24544 14968
rect 24584 14952 24636 14958
rect 24768 14952 24820 14958
rect 24636 14900 24768 14906
rect 24584 14894 24820 14900
rect 24596 14878 24808 14894
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24400 14476 24452 14482
rect 24400 14418 24452 14424
rect 24504 13274 24532 14758
rect 24596 14618 24624 14878
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 24596 13297 24624 14554
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24412 13246 24532 13274
rect 24582 13288 24638 13297
rect 24308 11144 24360 11150
rect 24308 11086 24360 11092
rect 24412 10810 24440 13246
rect 24582 13223 24638 13232
rect 24492 13184 24544 13190
rect 24492 13126 24544 13132
rect 24504 12889 24532 13126
rect 24490 12880 24546 12889
rect 24490 12815 24546 12824
rect 24492 12232 24544 12238
rect 24492 12174 24544 12180
rect 24504 11830 24532 12174
rect 24688 12102 24716 14418
rect 24872 13938 24900 14418
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 24964 13530 24992 17138
rect 25056 16250 25084 17478
rect 25044 16244 25096 16250
rect 25044 16186 25096 16192
rect 25134 16144 25190 16153
rect 25134 16079 25190 16088
rect 25148 15745 25176 16079
rect 25134 15736 25190 15745
rect 25134 15671 25190 15680
rect 25148 15570 25176 15671
rect 25136 15564 25188 15570
rect 25136 15506 25188 15512
rect 25148 14822 25176 15506
rect 25136 14816 25188 14822
rect 25240 14793 25268 17614
rect 25504 17128 25556 17134
rect 25318 17096 25374 17105
rect 25504 17070 25556 17076
rect 25318 17031 25374 17040
rect 25136 14758 25188 14764
rect 25226 14784 25282 14793
rect 25226 14719 25282 14728
rect 25228 14000 25280 14006
rect 25228 13942 25280 13948
rect 25136 13864 25188 13870
rect 25136 13806 25188 13812
rect 25148 13530 25176 13806
rect 24952 13524 25004 13530
rect 24952 13466 25004 13472
rect 25136 13524 25188 13530
rect 25136 13466 25188 13472
rect 25240 13326 25268 13942
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 25228 13320 25280 13326
rect 25228 13262 25280 13268
rect 24676 12096 24728 12102
rect 24676 12038 24728 12044
rect 24492 11824 24544 11830
rect 24492 11766 24544 11772
rect 24504 11218 24532 11766
rect 24492 11212 24544 11218
rect 24492 11154 24544 11160
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 24400 10804 24452 10810
rect 24400 10746 24452 10752
rect 24492 10804 24544 10810
rect 24492 10746 24544 10752
rect 24504 9178 24532 10746
rect 24688 10742 24716 10950
rect 24676 10736 24728 10742
rect 24676 10678 24728 10684
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24492 9172 24544 9178
rect 24492 9114 24544 9120
rect 24504 8634 24532 9114
rect 24596 9042 24624 10610
rect 24872 9178 24900 11018
rect 24964 9926 24992 13262
rect 25332 13172 25360 17031
rect 25410 15464 25466 15473
rect 25410 15399 25466 15408
rect 25424 15366 25452 15399
rect 25412 15360 25464 15366
rect 25412 15302 25464 15308
rect 25424 14822 25452 15302
rect 25412 14816 25464 14822
rect 25412 14758 25464 14764
rect 25424 14113 25452 14758
rect 25516 14278 25544 17070
rect 25792 16522 25820 17614
rect 25780 16516 25832 16522
rect 25780 16458 25832 16464
rect 25792 15094 25820 16458
rect 25872 16244 25924 16250
rect 25976 16232 26004 18935
rect 26160 18698 26188 19332
rect 26252 19281 26280 19468
rect 26238 19272 26294 19281
rect 26238 19207 26294 19216
rect 26148 18692 26200 18698
rect 26148 18634 26200 18640
rect 26344 18034 26372 20742
rect 26436 18630 26464 21848
rect 26528 21950 26740 21978
rect 26884 22024 26936 22030
rect 26884 21966 26936 21972
rect 26528 18970 26556 21950
rect 26700 21888 26752 21894
rect 26700 21830 26752 21836
rect 26608 21548 26660 21554
rect 26608 21490 26660 21496
rect 26516 18964 26568 18970
rect 26516 18906 26568 18912
rect 26620 18834 26648 21490
rect 26712 20058 26740 21830
rect 26792 20868 26844 20874
rect 26792 20810 26844 20816
rect 26804 20058 26832 20810
rect 26700 20052 26752 20058
rect 26700 19994 26752 20000
rect 26792 20052 26844 20058
rect 26792 19994 26844 20000
rect 26700 19372 26752 19378
rect 26700 19314 26752 19320
rect 26712 19145 26740 19314
rect 26698 19136 26754 19145
rect 26698 19071 26754 19080
rect 26896 18873 26924 21966
rect 27158 21720 27214 21729
rect 27158 21655 27160 21664
rect 27212 21655 27214 21664
rect 27160 21626 27212 21632
rect 27264 20466 27292 22170
rect 27344 21888 27396 21894
rect 27342 21856 27344 21865
rect 27396 21856 27398 21865
rect 27342 21791 27398 21800
rect 27356 20602 27384 21791
rect 27344 20596 27396 20602
rect 27344 20538 27396 20544
rect 27252 20460 27304 20466
rect 27252 20402 27304 20408
rect 27342 20360 27398 20369
rect 27252 20324 27304 20330
rect 27342 20295 27398 20304
rect 27252 20266 27304 20272
rect 27068 20256 27120 20262
rect 27068 20198 27120 20204
rect 27080 19718 27108 20198
rect 27264 19718 27292 20266
rect 27068 19712 27120 19718
rect 27068 19654 27120 19660
rect 27252 19712 27304 19718
rect 27252 19654 27304 19660
rect 27080 19417 27108 19654
rect 27264 19417 27292 19654
rect 27066 19408 27122 19417
rect 27066 19343 27122 19352
rect 27250 19408 27306 19417
rect 27250 19343 27306 19352
rect 27160 19168 27212 19174
rect 27160 19110 27212 19116
rect 27252 19168 27304 19174
rect 27252 19110 27304 19116
rect 26882 18864 26938 18873
rect 26608 18828 26660 18834
rect 27172 18834 27200 19110
rect 26882 18799 26938 18808
rect 27160 18828 27212 18834
rect 26608 18770 26660 18776
rect 27160 18770 27212 18776
rect 26608 18692 26660 18698
rect 26608 18634 26660 18640
rect 26424 18624 26476 18630
rect 26424 18566 26476 18572
rect 26516 18284 26568 18290
rect 26516 18226 26568 18232
rect 26424 18216 26476 18222
rect 26424 18158 26476 18164
rect 26160 18006 26372 18034
rect 26160 17785 26188 18006
rect 26146 17776 26202 17785
rect 26146 17711 26202 17720
rect 26056 17536 26108 17542
rect 26056 17478 26108 17484
rect 25924 16204 26004 16232
rect 25872 16186 25924 16192
rect 25872 15360 25924 15366
rect 25976 15337 26004 16204
rect 25872 15302 25924 15308
rect 25962 15328 26018 15337
rect 25780 15088 25832 15094
rect 25780 15030 25832 15036
rect 25688 15020 25740 15026
rect 25688 14962 25740 14968
rect 25596 14816 25648 14822
rect 25596 14758 25648 14764
rect 25608 14550 25636 14758
rect 25596 14544 25648 14550
rect 25596 14486 25648 14492
rect 25504 14272 25556 14278
rect 25504 14214 25556 14220
rect 25410 14104 25466 14113
rect 25410 14039 25466 14048
rect 25240 13144 25360 13172
rect 25240 12714 25268 13144
rect 25424 13002 25452 14039
rect 25516 13326 25544 14214
rect 25504 13320 25556 13326
rect 25504 13262 25556 13268
rect 25332 12974 25452 13002
rect 25228 12708 25280 12714
rect 25228 12650 25280 12656
rect 25332 10810 25360 12974
rect 25412 12708 25464 12714
rect 25412 12650 25464 12656
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 25424 10577 25452 12650
rect 25596 12436 25648 12442
rect 25596 12378 25648 12384
rect 25608 11898 25636 12378
rect 25596 11892 25648 11898
rect 25596 11834 25648 11840
rect 25410 10568 25466 10577
rect 25410 10503 25466 10512
rect 24952 9920 25004 9926
rect 25004 9880 25084 9908
rect 24952 9862 25004 9868
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 24584 9036 24636 9042
rect 24584 8978 24636 8984
rect 24492 8628 24544 8634
rect 24492 8570 24544 8576
rect 25056 8498 25084 9880
rect 25504 9512 25556 9518
rect 25504 9454 25556 9460
rect 25516 8634 25544 9454
rect 25608 8974 25636 11834
rect 25596 8968 25648 8974
rect 25596 8910 25648 8916
rect 25504 8628 25556 8634
rect 25504 8570 25556 8576
rect 25044 8492 25096 8498
rect 25044 8434 25096 8440
rect 25228 8424 25280 8430
rect 25228 8366 25280 8372
rect 25240 8090 25268 8366
rect 25228 8084 25280 8090
rect 25228 8026 25280 8032
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24780 4282 24808 4422
rect 24768 4276 24820 4282
rect 24768 4218 24820 4224
rect 24492 4072 24544 4078
rect 24228 4010 24440 4026
rect 24492 4014 24544 4020
rect 24228 4004 24452 4010
rect 24228 3998 24400 4004
rect 23664 3936 23716 3942
rect 23664 3878 23716 3884
rect 23296 3596 23348 3602
rect 23296 3538 23348 3544
rect 23572 3596 23624 3602
rect 23572 3538 23624 3544
rect 22928 3528 22980 3534
rect 22928 3470 22980 3476
rect 22940 3126 22968 3470
rect 22928 3120 22980 3126
rect 22848 3068 22928 3074
rect 22848 3062 22980 3068
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 22848 3046 22968 3062
rect 22652 2916 22704 2922
rect 22652 2858 22704 2864
rect 22848 2582 22876 3046
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 23308 2582 23336 3538
rect 23676 3126 23704 3878
rect 24228 3194 24256 3998
rect 24400 3946 24452 3952
rect 24400 3460 24452 3466
rect 24400 3402 24452 3408
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 23664 3120 23716 3126
rect 23664 3062 23716 3068
rect 23388 2916 23440 2922
rect 23388 2858 23440 2864
rect 23400 2582 23428 2858
rect 23676 2650 23704 3062
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 22836 2576 22888 2582
rect 22836 2518 22888 2524
rect 23296 2576 23348 2582
rect 23296 2518 23348 2524
rect 23388 2576 23440 2582
rect 23388 2518 23440 2524
rect 22468 2100 22520 2106
rect 22468 2042 22520 2048
rect 24412 800 24440 3402
rect 24504 3398 24532 4014
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 24780 2394 24808 4218
rect 25700 4078 25728 14962
rect 25884 13258 25912 15302
rect 25962 15263 26018 15272
rect 25872 13252 25924 13258
rect 25872 13194 25924 13200
rect 25976 12782 26004 15263
rect 26068 15162 26096 17478
rect 26436 16250 26464 18158
rect 26528 17270 26556 18226
rect 26620 17746 26648 18634
rect 27264 18426 27292 19110
rect 27252 18420 27304 18426
rect 27252 18362 27304 18368
rect 27356 18306 27384 20295
rect 27264 18278 27384 18306
rect 26792 18216 26844 18222
rect 26792 18158 26844 18164
rect 26608 17740 26660 17746
rect 26608 17682 26660 17688
rect 26516 17264 26568 17270
rect 26516 17206 26568 17212
rect 26424 16244 26476 16250
rect 26424 16186 26476 16192
rect 26436 16046 26464 16186
rect 26424 16040 26476 16046
rect 26424 15982 26476 15988
rect 26148 15700 26200 15706
rect 26528 15688 26556 17206
rect 26620 16998 26648 17682
rect 26608 16992 26660 16998
rect 26608 16934 26660 16940
rect 26620 16522 26648 16934
rect 26608 16516 26660 16522
rect 26608 16458 26660 16464
rect 26620 16250 26648 16458
rect 26608 16244 26660 16250
rect 26608 16186 26660 16192
rect 26804 15706 26832 18158
rect 27160 18080 27212 18086
rect 27160 18022 27212 18028
rect 27068 17264 27120 17270
rect 27068 17206 27120 17212
rect 27080 17105 27108 17206
rect 27066 17096 27122 17105
rect 27066 17031 27122 17040
rect 27172 16697 27200 18022
rect 27158 16688 27214 16697
rect 27158 16623 27214 16632
rect 27160 16176 27212 16182
rect 27066 16144 27122 16153
rect 27160 16118 27212 16124
rect 27066 16079 27122 16088
rect 26792 15700 26844 15706
rect 26528 15660 26740 15688
rect 26148 15642 26200 15648
rect 26056 15156 26108 15162
rect 26056 15098 26108 15104
rect 26056 13184 26108 13190
rect 26056 13126 26108 13132
rect 25964 12776 26016 12782
rect 25964 12718 26016 12724
rect 26068 12442 26096 13126
rect 26160 12889 26188 15642
rect 26238 15600 26294 15609
rect 26238 15535 26294 15544
rect 26424 15564 26476 15570
rect 26252 15366 26280 15535
rect 26424 15506 26476 15512
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26240 15360 26292 15366
rect 26240 15302 26292 15308
rect 26240 14816 26292 14822
rect 26240 14758 26292 14764
rect 26252 14346 26280 14758
rect 26240 14340 26292 14346
rect 26240 14282 26292 14288
rect 26436 14074 26464 15506
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 26146 12880 26202 12889
rect 26146 12815 26202 12824
rect 26056 12436 26108 12442
rect 26056 12378 26108 12384
rect 26332 12368 26384 12374
rect 26238 12336 26294 12345
rect 26332 12310 26384 12316
rect 26238 12271 26294 12280
rect 25964 12232 26016 12238
rect 25964 12174 26016 12180
rect 25976 11898 26004 12174
rect 26252 12102 26280 12271
rect 26240 12096 26292 12102
rect 26240 12038 26292 12044
rect 25964 11892 26016 11898
rect 25964 11834 26016 11840
rect 25976 11150 26004 11834
rect 26344 11694 26372 12310
rect 26332 11688 26384 11694
rect 26332 11630 26384 11636
rect 26620 11354 26648 15506
rect 26712 15434 26740 15660
rect 26792 15642 26844 15648
rect 26976 15700 27028 15706
rect 26976 15642 27028 15648
rect 26988 15609 27016 15642
rect 27080 15638 27108 16079
rect 27068 15632 27120 15638
rect 26974 15600 27030 15609
rect 27068 15574 27120 15580
rect 26974 15535 27030 15544
rect 26700 15428 26752 15434
rect 26700 15370 26752 15376
rect 26792 15360 26844 15366
rect 26976 15360 27028 15366
rect 26792 15302 26844 15308
rect 26974 15328 26976 15337
rect 27028 15328 27030 15337
rect 26804 14822 26832 15302
rect 26974 15263 27030 15272
rect 27080 15162 27108 15574
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 27080 15065 27108 15098
rect 27066 15056 27122 15065
rect 27066 14991 27122 15000
rect 27172 14890 27200 16118
rect 27264 15162 27292 18278
rect 27342 18184 27398 18193
rect 27342 18119 27398 18128
rect 27356 16250 27384 18119
rect 27448 16454 27476 22578
rect 27540 21010 27568 23462
rect 27632 23186 27660 24278
rect 28368 24206 28396 24686
rect 28356 24200 28408 24206
rect 28356 24142 28408 24148
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 28172 23724 28224 23730
rect 28172 23666 28224 23672
rect 27804 23520 27856 23526
rect 27804 23462 27856 23468
rect 27620 23180 27672 23186
rect 27620 23122 27672 23128
rect 27712 22704 27764 22710
rect 27712 22646 27764 22652
rect 27620 22160 27672 22166
rect 27620 22102 27672 22108
rect 27528 21004 27580 21010
rect 27528 20946 27580 20952
rect 27632 20874 27660 22102
rect 27620 20868 27672 20874
rect 27620 20810 27672 20816
rect 27620 20528 27672 20534
rect 27620 20470 27672 20476
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 27540 18902 27568 19790
rect 27632 19310 27660 20470
rect 27724 20262 27752 22646
rect 27816 22574 27844 23462
rect 28184 23050 28212 23666
rect 28460 23225 28488 26302
rect 28630 26314 28948 26330
rect 28630 26308 28960 26314
rect 28630 26302 28908 26308
rect 28630 26200 28686 26302
rect 28908 26250 28960 26256
rect 29274 26302 29592 26330
rect 29274 26200 29330 26302
rect 29564 25809 29592 26302
rect 29918 26302 30420 26330
rect 29918 26200 29974 26302
rect 30102 26208 30158 26217
rect 30102 26143 30158 26152
rect 29550 25800 29606 25809
rect 29550 25735 29606 25744
rect 29828 25492 29880 25498
rect 29828 25434 29880 25440
rect 28632 25288 28684 25294
rect 28632 25230 28684 25236
rect 28540 23792 28592 23798
rect 28540 23734 28592 23740
rect 28446 23216 28502 23225
rect 28356 23180 28408 23186
rect 28446 23151 28502 23160
rect 28356 23122 28408 23128
rect 28172 23044 28224 23050
rect 28172 22986 28224 22992
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 27804 22568 27856 22574
rect 27804 22510 27856 22516
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 28172 21616 28224 21622
rect 28368 21593 28396 23122
rect 28552 22094 28580 23734
rect 28644 22710 28672 25230
rect 29644 24336 29696 24342
rect 29644 24278 29696 24284
rect 29368 24132 29420 24138
rect 29368 24074 29420 24080
rect 29380 23866 29408 24074
rect 29656 24070 29684 24278
rect 29644 24064 29696 24070
rect 29644 24006 29696 24012
rect 29368 23860 29420 23866
rect 29368 23802 29420 23808
rect 29000 23588 29052 23594
rect 29000 23530 29052 23536
rect 28724 23044 28776 23050
rect 28724 22986 28776 22992
rect 28632 22704 28684 22710
rect 28632 22646 28684 22652
rect 28460 22066 28580 22094
rect 28172 21558 28224 21564
rect 28354 21584 28410 21593
rect 28184 21486 28212 21558
rect 28354 21519 28410 21528
rect 28172 21480 28224 21486
rect 28172 21422 28224 21428
rect 28262 21176 28318 21185
rect 28262 21111 28318 21120
rect 27804 20868 27856 20874
rect 27804 20810 27856 20816
rect 27816 20641 27844 20810
rect 28276 20788 28304 21111
rect 28276 20777 28396 20788
rect 28276 20768 28410 20777
rect 28276 20760 28354 20768
rect 27950 20700 28258 20709
rect 28354 20703 28410 20712
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27802 20632 27858 20641
rect 27950 20635 28258 20644
rect 27802 20567 27858 20576
rect 27712 20256 27764 20262
rect 27712 20198 27764 20204
rect 27712 20052 27764 20058
rect 27712 19994 27764 20000
rect 27620 19304 27672 19310
rect 27620 19246 27672 19252
rect 27724 19009 27752 19994
rect 27816 19292 27844 20567
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 28368 19514 28396 20703
rect 28356 19508 28408 19514
rect 28356 19450 28408 19456
rect 27896 19304 27948 19310
rect 27816 19264 27896 19292
rect 27896 19246 27948 19252
rect 28080 19236 28132 19242
rect 28080 19178 28132 19184
rect 28092 19009 28120 19178
rect 27710 19000 27766 19009
rect 27710 18935 27766 18944
rect 28078 19000 28134 19009
rect 28078 18935 28134 18944
rect 27528 18896 27580 18902
rect 27528 18838 27580 18844
rect 27528 18760 27580 18766
rect 27528 18702 27580 18708
rect 27540 16522 27568 18702
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 27712 18420 27764 18426
rect 27712 18362 27764 18368
rect 27620 18080 27672 18086
rect 27620 18022 27672 18028
rect 27632 16969 27660 18022
rect 27618 16960 27674 16969
rect 27618 16895 27674 16904
rect 27528 16516 27580 16522
rect 27528 16458 27580 16464
rect 27436 16448 27488 16454
rect 27436 16390 27488 16396
rect 27344 16244 27396 16250
rect 27344 16186 27396 16192
rect 27528 16244 27580 16250
rect 27528 16186 27580 16192
rect 27436 16108 27488 16114
rect 27436 16050 27488 16056
rect 27448 16017 27476 16050
rect 27434 16008 27490 16017
rect 27344 15972 27396 15978
rect 27434 15943 27490 15952
rect 27344 15914 27396 15920
rect 27252 15156 27304 15162
rect 27252 15098 27304 15104
rect 27250 15056 27306 15065
rect 27250 14991 27252 15000
rect 27304 14991 27306 15000
rect 27252 14962 27304 14968
rect 27160 14884 27212 14890
rect 27080 14844 27160 14872
rect 26792 14816 26844 14822
rect 26792 14758 26844 14764
rect 27080 14414 27108 14844
rect 27160 14826 27212 14832
rect 27160 14476 27212 14482
rect 27160 14418 27212 14424
rect 27068 14408 27120 14414
rect 27068 14350 27120 14356
rect 27080 14006 27108 14350
rect 26792 14000 26844 14006
rect 26792 13942 26844 13948
rect 27068 14000 27120 14006
rect 27068 13942 27120 13948
rect 26804 12918 26832 13942
rect 27068 13320 27120 13326
rect 27068 13262 27120 13268
rect 26976 13184 27028 13190
rect 26976 13126 27028 13132
rect 26792 12912 26844 12918
rect 26792 12854 26844 12860
rect 26804 12238 26832 12854
rect 26988 12306 27016 13126
rect 27080 12986 27108 13262
rect 27172 12986 27200 14418
rect 27068 12980 27120 12986
rect 27068 12922 27120 12928
rect 27160 12980 27212 12986
rect 27160 12922 27212 12928
rect 27356 12374 27384 15914
rect 27448 15638 27476 15943
rect 27540 15706 27568 16186
rect 27528 15700 27580 15706
rect 27528 15642 27580 15648
rect 27436 15632 27488 15638
rect 27436 15574 27488 15580
rect 27724 15502 27752 18362
rect 28356 17740 28408 17746
rect 28356 17682 28408 17688
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27802 17368 27858 17377
rect 27950 17371 28258 17380
rect 27802 17303 27804 17312
rect 27856 17303 27858 17312
rect 27804 17274 27856 17280
rect 27988 17264 28040 17270
rect 27802 17232 27858 17241
rect 27988 17206 28040 17212
rect 28078 17232 28134 17241
rect 27802 17167 27804 17176
rect 27856 17167 27858 17176
rect 27804 17138 27856 17144
rect 28000 17105 28028 17206
rect 28078 17167 28134 17176
rect 28092 17134 28120 17167
rect 28080 17128 28132 17134
rect 27986 17096 28042 17105
rect 27896 17060 27948 17066
rect 27816 17020 27896 17048
rect 27712 15496 27764 15502
rect 27712 15438 27764 15444
rect 27436 15360 27488 15366
rect 27436 15302 27488 15308
rect 27448 13462 27476 15302
rect 27436 13456 27488 13462
rect 27436 13398 27488 13404
rect 27620 13456 27672 13462
rect 27620 13398 27672 13404
rect 27632 13161 27660 13398
rect 27816 13394 27844 17020
rect 28080 17070 28132 17076
rect 27986 17031 28042 17040
rect 27896 17002 27948 17008
rect 28368 16658 28396 17682
rect 28356 16652 28408 16658
rect 28356 16594 28408 16600
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 28368 16114 28396 16594
rect 28460 16590 28488 22066
rect 28632 21888 28684 21894
rect 28630 21856 28632 21865
rect 28684 21856 28686 21865
rect 28630 21791 28686 21800
rect 28736 21690 28764 22986
rect 28908 22092 28960 22098
rect 28908 22034 28960 22040
rect 28816 22024 28868 22030
rect 28816 21966 28868 21972
rect 28828 21729 28856 21966
rect 28814 21720 28870 21729
rect 28540 21684 28592 21690
rect 28540 21626 28592 21632
rect 28724 21684 28776 21690
rect 28814 21655 28870 21664
rect 28724 21626 28776 21632
rect 28552 20942 28580 21626
rect 28632 21616 28684 21622
rect 28632 21558 28684 21564
rect 28644 21486 28672 21558
rect 28920 21486 28948 22034
rect 28632 21480 28684 21486
rect 28816 21480 28868 21486
rect 28632 21422 28684 21428
rect 28814 21448 28816 21457
rect 28908 21480 28960 21486
rect 28868 21448 28870 21457
rect 28908 21422 28960 21428
rect 28814 21383 28870 21392
rect 28540 20936 28592 20942
rect 28540 20878 28592 20884
rect 28724 20800 28776 20806
rect 28724 20742 28776 20748
rect 28540 20392 28592 20398
rect 28540 20334 28592 20340
rect 28552 18970 28580 20334
rect 28632 19916 28684 19922
rect 28632 19858 28684 19864
rect 28644 19378 28672 19858
rect 28736 19514 28764 20742
rect 28828 20505 28856 21383
rect 29012 21010 29040 23530
rect 29092 22976 29144 22982
rect 29090 22944 29092 22953
rect 29276 22976 29328 22982
rect 29144 22944 29146 22953
rect 29276 22918 29328 22924
rect 29368 22976 29420 22982
rect 29368 22918 29420 22924
rect 29090 22879 29146 22888
rect 29104 21554 29132 22879
rect 29288 21622 29316 22918
rect 29380 22522 29408 22918
rect 29380 22494 29500 22522
rect 29368 22228 29420 22234
rect 29368 22170 29420 22176
rect 29380 21962 29408 22170
rect 29368 21956 29420 21962
rect 29368 21898 29420 21904
rect 29276 21616 29328 21622
rect 29472 21570 29500 22494
rect 29656 22094 29684 24006
rect 29736 23656 29788 23662
rect 29736 23598 29788 23604
rect 29748 22438 29776 23598
rect 29840 23322 29868 25434
rect 29918 24168 29974 24177
rect 29918 24103 29974 24112
rect 29932 24070 29960 24103
rect 29920 24064 29972 24070
rect 29920 24006 29972 24012
rect 29828 23316 29880 23322
rect 29828 23258 29880 23264
rect 30012 23248 30064 23254
rect 30012 23190 30064 23196
rect 30024 22710 30052 23190
rect 30116 23066 30144 26143
rect 30392 25401 30420 26302
rect 30562 26302 30788 26330
rect 30562 26200 30618 26302
rect 30378 25392 30434 25401
rect 30378 25327 30434 25336
rect 30288 24608 30340 24614
rect 30288 24550 30340 24556
rect 30196 24404 30248 24410
rect 30196 24346 30248 24352
rect 30208 23186 30236 24346
rect 30300 24342 30328 24550
rect 30288 24336 30340 24342
rect 30288 24278 30340 24284
rect 30288 24200 30340 24206
rect 30288 24142 30340 24148
rect 30300 23526 30328 24142
rect 30564 23792 30616 23798
rect 30564 23734 30616 23740
rect 30288 23520 30340 23526
rect 30288 23462 30340 23468
rect 30300 23186 30328 23462
rect 30196 23180 30248 23186
rect 30196 23122 30248 23128
rect 30288 23180 30340 23186
rect 30288 23122 30340 23128
rect 30116 23038 30236 23066
rect 30104 22976 30156 22982
rect 30104 22918 30156 22924
rect 30012 22704 30064 22710
rect 30012 22646 30064 22652
rect 29736 22432 29788 22438
rect 29736 22374 29788 22380
rect 29920 22432 29972 22438
rect 29920 22374 29972 22380
rect 29932 22166 29960 22374
rect 29920 22160 29972 22166
rect 29920 22102 29972 22108
rect 29656 22066 29868 22094
rect 29644 22024 29696 22030
rect 29644 21966 29696 21972
rect 29276 21558 29328 21564
rect 29092 21548 29144 21554
rect 29092 21490 29144 21496
rect 29000 21004 29052 21010
rect 29000 20946 29052 20952
rect 28908 20800 28960 20806
rect 28908 20742 28960 20748
rect 28814 20496 28870 20505
rect 28814 20431 28870 20440
rect 28920 20346 28948 20742
rect 29288 20618 29316 21558
rect 29380 21542 29500 21570
rect 29552 21548 29604 21554
rect 29380 21350 29408 21542
rect 29552 21490 29604 21496
rect 29460 21480 29512 21486
rect 29460 21422 29512 21428
rect 29368 21344 29420 21350
rect 29368 21286 29420 21292
rect 29288 20590 29408 20618
rect 29276 20528 29328 20534
rect 28998 20496 29054 20505
rect 29276 20470 29328 20476
rect 28998 20431 29054 20440
rect 28828 20318 28948 20346
rect 28828 20058 28856 20318
rect 28816 20052 28868 20058
rect 28816 19994 28868 20000
rect 28908 19984 28960 19990
rect 28908 19926 28960 19932
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 28828 19553 28856 19790
rect 28814 19544 28870 19553
rect 28724 19508 28776 19514
rect 28814 19479 28870 19488
rect 28724 19450 28776 19456
rect 28632 19372 28684 19378
rect 28632 19314 28684 19320
rect 28724 19372 28776 19378
rect 28724 19314 28776 19320
rect 28540 18964 28592 18970
rect 28540 18906 28592 18912
rect 28632 18760 28684 18766
rect 28632 18702 28684 18708
rect 28540 18624 28592 18630
rect 28540 18566 28592 18572
rect 28552 17513 28580 18566
rect 28644 18290 28672 18702
rect 28632 18284 28684 18290
rect 28632 18226 28684 18232
rect 28632 18080 28684 18086
rect 28632 18022 28684 18028
rect 28538 17504 28594 17513
rect 28538 17439 28594 17448
rect 28448 16584 28500 16590
rect 28448 16526 28500 16532
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 28368 15094 28396 16050
rect 28644 15638 28672 18022
rect 28736 16130 28764 19314
rect 28920 18306 28948 19926
rect 28828 18278 28948 18306
rect 28828 18222 28856 18278
rect 28816 18216 28868 18222
rect 28816 18158 28868 18164
rect 28908 18216 28960 18222
rect 28908 18158 28960 18164
rect 28816 17808 28868 17814
rect 28816 17750 28868 17756
rect 28828 17678 28856 17750
rect 28816 17672 28868 17678
rect 28814 17640 28816 17649
rect 28868 17640 28870 17649
rect 28814 17575 28870 17584
rect 28920 17542 28948 18158
rect 29012 17814 29040 20431
rect 29288 20398 29316 20470
rect 29276 20392 29328 20398
rect 29276 20334 29328 20340
rect 29184 20256 29236 20262
rect 29184 20198 29236 20204
rect 29196 19700 29224 20198
rect 29288 20058 29316 20334
rect 29380 20058 29408 20590
rect 29276 20052 29328 20058
rect 29276 19994 29328 20000
rect 29368 20052 29420 20058
rect 29368 19994 29420 20000
rect 29276 19712 29328 19718
rect 29196 19672 29276 19700
rect 29276 19654 29328 19660
rect 29288 19446 29316 19654
rect 29276 19440 29328 19446
rect 29276 19382 29328 19388
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 29092 18624 29144 18630
rect 29092 18566 29144 18572
rect 29104 18086 29132 18566
rect 29092 18080 29144 18086
rect 29092 18022 29144 18028
rect 29000 17808 29052 17814
rect 29000 17750 29052 17756
rect 29104 17649 29132 18022
rect 29090 17640 29146 17649
rect 29090 17575 29146 17584
rect 28908 17536 28960 17542
rect 28908 17478 28960 17484
rect 29090 17368 29146 17377
rect 29090 17303 29092 17312
rect 29144 17303 29146 17312
rect 29092 17274 29144 17280
rect 29092 17128 29144 17134
rect 29090 17096 29092 17105
rect 29144 17096 29146 17105
rect 29090 17031 29146 17040
rect 29000 16992 29052 16998
rect 29052 16952 29132 16980
rect 29000 16934 29052 16940
rect 29000 16720 29052 16726
rect 29000 16662 29052 16668
rect 28908 16584 28960 16590
rect 28908 16526 28960 16532
rect 28920 16182 28948 16526
rect 28908 16176 28960 16182
rect 28736 16102 28856 16130
rect 28908 16118 28960 16124
rect 28724 16040 28776 16046
rect 28724 15982 28776 15988
rect 28632 15632 28684 15638
rect 28632 15574 28684 15580
rect 28540 15564 28592 15570
rect 28540 15506 28592 15512
rect 28356 15088 28408 15094
rect 28356 15030 28408 15036
rect 28448 15088 28500 15094
rect 28448 15030 28500 15036
rect 28080 14884 28132 14890
rect 28460 14872 28488 15030
rect 28132 14844 28488 14872
rect 28080 14826 28132 14832
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 28460 14074 28488 14844
rect 28552 14482 28580 15506
rect 28736 15502 28764 15982
rect 28724 15496 28776 15502
rect 28724 15438 28776 15444
rect 28724 15156 28776 15162
rect 28724 15098 28776 15104
rect 28736 14906 28764 15098
rect 28828 14906 28856 16102
rect 28920 15638 28948 16118
rect 28908 15632 28960 15638
rect 28908 15574 28960 15580
rect 28736 14878 28856 14906
rect 28908 14952 28960 14958
rect 28908 14894 28960 14900
rect 28736 14550 28764 14878
rect 28816 14816 28868 14822
rect 28816 14758 28868 14764
rect 28724 14544 28776 14550
rect 28724 14486 28776 14492
rect 28540 14476 28592 14482
rect 28540 14418 28592 14424
rect 28632 14272 28684 14278
rect 28632 14214 28684 14220
rect 28448 14068 28500 14074
rect 28448 14010 28500 14016
rect 27804 13388 27856 13394
rect 27804 13330 27856 13336
rect 27618 13152 27674 13161
rect 27618 13087 27674 13096
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 27712 12912 27764 12918
rect 27712 12854 27764 12860
rect 28172 12912 28224 12918
rect 28460 12900 28488 14010
rect 28540 13728 28592 13734
rect 28540 13670 28592 13676
rect 28224 12872 28488 12900
rect 28172 12854 28224 12860
rect 27620 12436 27672 12442
rect 27724 12434 27752 12854
rect 27724 12406 27844 12434
rect 27620 12378 27672 12384
rect 27344 12368 27396 12374
rect 27344 12310 27396 12316
rect 26976 12300 27028 12306
rect 26976 12242 27028 12248
rect 27528 12300 27580 12306
rect 27528 12242 27580 12248
rect 26792 12232 26844 12238
rect 26792 12174 26844 12180
rect 27160 12232 27212 12238
rect 27160 12174 27212 12180
rect 27172 11626 27200 12174
rect 27344 12096 27396 12102
rect 27344 12038 27396 12044
rect 27356 11898 27384 12038
rect 27344 11892 27396 11898
rect 27344 11834 27396 11840
rect 27344 11756 27396 11762
rect 27344 11698 27396 11704
rect 27160 11620 27212 11626
rect 27160 11562 27212 11568
rect 26608 11348 26660 11354
rect 26608 11290 26660 11296
rect 27160 11348 27212 11354
rect 27160 11290 27212 11296
rect 25964 11144 26016 11150
rect 25964 11086 26016 11092
rect 25976 10810 26004 11086
rect 25964 10804 26016 10810
rect 25964 10746 26016 10752
rect 25976 10062 26004 10746
rect 26620 10674 26648 11290
rect 26700 11144 26752 11150
rect 26700 11086 26752 11092
rect 26884 11144 26936 11150
rect 26936 11104 27016 11132
rect 26884 11086 26936 11092
rect 26608 10668 26660 10674
rect 26608 10610 26660 10616
rect 26608 10464 26660 10470
rect 26608 10406 26660 10412
rect 26620 10266 26648 10406
rect 26712 10266 26740 11086
rect 26608 10260 26660 10266
rect 26608 10202 26660 10208
rect 26700 10260 26752 10266
rect 26700 10202 26752 10208
rect 26988 10062 27016 11104
rect 27068 10668 27120 10674
rect 27068 10610 27120 10616
rect 27080 10169 27108 10610
rect 27066 10160 27122 10169
rect 27066 10095 27122 10104
rect 25964 10056 26016 10062
rect 25964 9998 26016 10004
rect 26976 10056 27028 10062
rect 26976 9998 27028 10004
rect 26424 9920 26476 9926
rect 26424 9862 26476 9868
rect 26436 9722 26464 9862
rect 26988 9722 27016 9998
rect 26424 9716 26476 9722
rect 26424 9658 26476 9664
rect 26976 9716 27028 9722
rect 26976 9658 27028 9664
rect 26056 9648 26108 9654
rect 26054 9616 26056 9625
rect 26108 9616 26110 9625
rect 26054 9551 26110 9560
rect 26148 9580 26200 9586
rect 26068 8634 26096 9551
rect 26148 9522 26200 9528
rect 26160 9081 26188 9522
rect 26424 9512 26476 9518
rect 26424 9454 26476 9460
rect 26146 9072 26202 9081
rect 26146 9007 26202 9016
rect 26056 8628 26108 8634
rect 26056 8570 26108 8576
rect 26160 8378 26188 9007
rect 26436 8498 26464 9454
rect 27080 9382 27108 10095
rect 27068 9376 27120 9382
rect 27068 9318 27120 9324
rect 26424 8492 26476 8498
rect 26424 8434 26476 8440
rect 26068 8362 26188 8378
rect 26056 8356 26188 8362
rect 26108 8350 26188 8356
rect 26056 8298 26108 8304
rect 26068 6186 26096 8298
rect 26056 6180 26108 6186
rect 26056 6122 26108 6128
rect 26238 5128 26294 5137
rect 26238 5063 26294 5072
rect 26252 4690 26280 5063
rect 26240 4684 26292 4690
rect 26240 4626 26292 4632
rect 27080 4622 27108 9318
rect 27172 8974 27200 11290
rect 27356 10849 27384 11698
rect 27436 11688 27488 11694
rect 27434 11656 27436 11665
rect 27488 11656 27490 11665
rect 27434 11591 27490 11600
rect 27540 11218 27568 12242
rect 27632 12102 27660 12378
rect 27620 12096 27672 12102
rect 27620 12038 27672 12044
rect 27528 11212 27580 11218
rect 27528 11154 27580 11160
rect 27342 10840 27398 10849
rect 27342 10775 27398 10784
rect 27620 10736 27672 10742
rect 27620 10678 27672 10684
rect 27252 10600 27304 10606
rect 27252 10542 27304 10548
rect 27264 10266 27292 10542
rect 27252 10260 27304 10266
rect 27632 10248 27660 10678
rect 27252 10202 27304 10208
rect 27448 10220 27660 10248
rect 27264 9382 27292 10202
rect 27448 9450 27476 10220
rect 27620 10124 27672 10130
rect 27620 10066 27672 10072
rect 27436 9444 27488 9450
rect 27436 9386 27488 9392
rect 27252 9376 27304 9382
rect 27252 9318 27304 9324
rect 27160 8968 27212 8974
rect 27160 8910 27212 8916
rect 27264 8906 27292 9318
rect 27252 8900 27304 8906
rect 27252 8842 27304 8848
rect 27632 8634 27660 10066
rect 27816 9178 27844 12406
rect 28460 12186 28488 12872
rect 28552 12714 28580 13670
rect 28540 12708 28592 12714
rect 28540 12650 28592 12656
rect 28460 12158 28580 12186
rect 28356 12096 28408 12102
rect 28356 12038 28408 12044
rect 28448 12096 28500 12102
rect 28448 12038 28500 12044
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 27804 9172 27856 9178
rect 27804 9114 27856 9120
rect 27804 8832 27856 8838
rect 27804 8774 27856 8780
rect 27620 8628 27672 8634
rect 27620 8570 27672 8576
rect 27816 8294 27844 8774
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 27804 8288 27856 8294
rect 27804 8230 27856 8236
rect 27816 7750 27844 8230
rect 28368 7818 28396 12038
rect 28460 11898 28488 12038
rect 28448 11892 28500 11898
rect 28448 11834 28500 11840
rect 28448 11756 28500 11762
rect 28448 11698 28500 11704
rect 28356 7812 28408 7818
rect 28356 7754 28408 7760
rect 27804 7744 27856 7750
rect 27804 7686 27856 7692
rect 27816 6730 27844 7686
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27804 6724 27856 6730
rect 27804 6666 27856 6672
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 28460 6254 28488 11698
rect 28552 10996 28580 12158
rect 28644 11121 28672 14214
rect 28736 13705 28764 14486
rect 28722 13696 28778 13705
rect 28722 13631 28778 13640
rect 28828 12306 28856 14758
rect 28816 12300 28868 12306
rect 28816 12242 28868 12248
rect 28814 11792 28870 11801
rect 28814 11727 28870 11736
rect 28828 11694 28856 11727
rect 28816 11688 28868 11694
rect 28816 11630 28868 11636
rect 28630 11112 28686 11121
rect 28630 11047 28686 11056
rect 28724 11008 28776 11014
rect 28552 10968 28724 10996
rect 28552 10062 28580 10968
rect 28724 10950 28776 10956
rect 28816 10600 28868 10606
rect 28920 10588 28948 14894
rect 29012 13938 29040 16662
rect 29104 15162 29132 16952
rect 29196 16658 29224 18702
rect 29288 18612 29316 19382
rect 29380 18766 29408 19994
rect 29472 19922 29500 21422
rect 29460 19916 29512 19922
rect 29460 19858 29512 19864
rect 29460 19712 29512 19718
rect 29460 19654 29512 19660
rect 29368 18760 29420 18766
rect 29368 18702 29420 18708
rect 29472 18698 29500 19654
rect 29564 18970 29592 21490
rect 29656 20602 29684 21966
rect 29840 21865 29868 22066
rect 29826 21856 29882 21865
rect 29826 21791 29882 21800
rect 29736 21072 29788 21078
rect 29736 21014 29788 21020
rect 29748 20913 29776 21014
rect 29734 20904 29790 20913
rect 29734 20839 29790 20848
rect 29840 20602 29868 21791
rect 29920 20936 29972 20942
rect 29920 20878 29972 20884
rect 29644 20596 29696 20602
rect 29644 20538 29696 20544
rect 29828 20596 29880 20602
rect 29828 20538 29880 20544
rect 29736 20392 29788 20398
rect 29736 20334 29788 20340
rect 29644 19916 29696 19922
rect 29644 19858 29696 19864
rect 29656 19378 29684 19858
rect 29644 19372 29696 19378
rect 29644 19314 29696 19320
rect 29552 18964 29604 18970
rect 29552 18906 29604 18912
rect 29656 18834 29684 19314
rect 29644 18828 29696 18834
rect 29644 18770 29696 18776
rect 29460 18692 29512 18698
rect 29460 18634 29512 18640
rect 29288 18584 29408 18612
rect 29276 17536 29328 17542
rect 29276 17478 29328 17484
rect 29184 16652 29236 16658
rect 29184 16594 29236 16600
rect 29184 16448 29236 16454
rect 29184 16390 29236 16396
rect 29196 15570 29224 16390
rect 29288 16250 29316 17478
rect 29380 17202 29408 18584
rect 29552 18216 29604 18222
rect 29552 18158 29604 18164
rect 29368 17196 29420 17202
rect 29368 17138 29420 17144
rect 29380 16794 29408 17138
rect 29458 17096 29514 17105
rect 29458 17031 29514 17040
rect 29472 16998 29500 17031
rect 29460 16992 29512 16998
rect 29460 16934 29512 16940
rect 29368 16788 29420 16794
rect 29368 16730 29420 16736
rect 29276 16244 29328 16250
rect 29276 16186 29328 16192
rect 29184 15564 29236 15570
rect 29184 15506 29236 15512
rect 29092 15156 29144 15162
rect 29092 15098 29144 15104
rect 29092 14612 29144 14618
rect 29092 14554 29144 14560
rect 29000 13932 29052 13938
rect 29000 13874 29052 13880
rect 29012 12918 29040 13874
rect 29104 13530 29132 14554
rect 29276 14272 29328 14278
rect 29274 14240 29276 14249
rect 29460 14272 29512 14278
rect 29328 14240 29330 14249
rect 29460 14214 29512 14220
rect 29274 14175 29330 14184
rect 29288 14006 29316 14175
rect 29276 14000 29328 14006
rect 29276 13942 29328 13948
rect 29368 13728 29420 13734
rect 29368 13670 29420 13676
rect 29092 13524 29144 13530
rect 29092 13466 29144 13472
rect 29380 12986 29408 13670
rect 29472 13530 29500 14214
rect 29460 13524 29512 13530
rect 29460 13466 29512 13472
rect 29368 12980 29420 12986
rect 29368 12922 29420 12928
rect 29000 12912 29052 12918
rect 29000 12854 29052 12860
rect 29276 12844 29328 12850
rect 29276 12786 29328 12792
rect 29092 12232 29144 12238
rect 29092 12174 29144 12180
rect 29104 11830 29132 12174
rect 29182 11928 29238 11937
rect 29182 11863 29238 11872
rect 29092 11824 29144 11830
rect 29092 11766 29144 11772
rect 28998 11656 29054 11665
rect 28998 11591 29054 11600
rect 29012 11354 29040 11591
rect 29196 11370 29224 11863
rect 29288 11558 29316 12786
rect 29380 12238 29408 12922
rect 29472 12646 29500 13466
rect 29564 12850 29592 18158
rect 29644 17128 29696 17134
rect 29644 17070 29696 17076
rect 29552 12844 29604 12850
rect 29552 12786 29604 12792
rect 29460 12640 29512 12646
rect 29460 12582 29512 12588
rect 29472 12345 29500 12582
rect 29458 12336 29514 12345
rect 29458 12271 29514 12280
rect 29368 12232 29420 12238
rect 29368 12174 29420 12180
rect 29460 11824 29512 11830
rect 29460 11766 29512 11772
rect 29368 11688 29420 11694
rect 29368 11630 29420 11636
rect 29276 11552 29328 11558
rect 29276 11494 29328 11500
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 29104 11342 29224 11370
rect 29012 11257 29040 11290
rect 28998 11248 29054 11257
rect 28998 11183 29054 11192
rect 29000 10600 29052 10606
rect 28920 10560 29000 10588
rect 28816 10542 28868 10548
rect 29000 10542 29052 10548
rect 28828 10198 28856 10542
rect 28816 10192 28868 10198
rect 28816 10134 28868 10140
rect 28540 10056 28592 10062
rect 28540 9998 28592 10004
rect 29104 9602 29132 11342
rect 29184 11212 29236 11218
rect 29184 11154 29236 11160
rect 29012 9574 29132 9602
rect 29012 9042 29040 9574
rect 29092 9512 29144 9518
rect 29092 9454 29144 9460
rect 29104 9382 29132 9454
rect 29196 9382 29224 11154
rect 29288 10742 29316 11494
rect 29380 11286 29408 11630
rect 29368 11280 29420 11286
rect 29368 11222 29420 11228
rect 29368 11076 29420 11082
rect 29368 11018 29420 11024
rect 29276 10736 29328 10742
rect 29276 10678 29328 10684
rect 29276 10464 29328 10470
rect 29276 10406 29328 10412
rect 29288 9722 29316 10406
rect 29380 10266 29408 11018
rect 29472 11014 29500 11766
rect 29552 11552 29604 11558
rect 29552 11494 29604 11500
rect 29460 11008 29512 11014
rect 29460 10950 29512 10956
rect 29368 10260 29420 10266
rect 29368 10202 29420 10208
rect 29368 10056 29420 10062
rect 29368 9998 29420 10004
rect 29276 9716 29328 9722
rect 29276 9658 29328 9664
rect 29276 9580 29328 9586
rect 29380 9568 29408 9998
rect 29564 9568 29592 11494
rect 29656 11218 29684 17070
rect 29748 16590 29776 20334
rect 29828 18828 29880 18834
rect 29828 18770 29880 18776
rect 29736 16584 29788 16590
rect 29736 16526 29788 16532
rect 29736 16448 29788 16454
rect 29736 16390 29788 16396
rect 29748 16289 29776 16390
rect 29734 16280 29790 16289
rect 29734 16215 29790 16224
rect 29840 15094 29868 18770
rect 29932 18465 29960 20878
rect 30024 20534 30052 22646
rect 30116 21146 30144 22918
rect 30208 22094 30236 23038
rect 30380 22568 30432 22574
rect 30380 22510 30432 22516
rect 30288 22432 30340 22438
rect 30288 22374 30340 22380
rect 30300 22234 30328 22374
rect 30392 22234 30420 22510
rect 30288 22228 30340 22234
rect 30288 22170 30340 22176
rect 30380 22228 30432 22234
rect 30380 22170 30432 22176
rect 30208 22066 30328 22094
rect 30194 21856 30250 21865
rect 30194 21791 30250 21800
rect 30208 21622 30236 21791
rect 30196 21616 30248 21622
rect 30196 21558 30248 21564
rect 30196 21344 30248 21350
rect 30196 21286 30248 21292
rect 30104 21140 30156 21146
rect 30104 21082 30156 21088
rect 30104 21004 30156 21010
rect 30104 20946 30156 20952
rect 30116 20806 30144 20946
rect 30104 20800 30156 20806
rect 30104 20742 30156 20748
rect 30104 20596 30156 20602
rect 30104 20538 30156 20544
rect 30012 20528 30064 20534
rect 30012 20470 30064 20476
rect 30116 19718 30144 20538
rect 30208 20398 30236 21286
rect 30196 20392 30248 20398
rect 30196 20334 30248 20340
rect 30300 20262 30328 22066
rect 30378 21584 30434 21593
rect 30378 21519 30434 21528
rect 30392 20534 30420 21519
rect 30472 21344 30524 21350
rect 30472 21286 30524 21292
rect 30380 20528 30432 20534
rect 30380 20470 30432 20476
rect 30380 20324 30432 20330
rect 30380 20266 30432 20272
rect 30288 20256 30340 20262
rect 30288 20198 30340 20204
rect 30194 19952 30250 19961
rect 30194 19887 30250 19896
rect 30208 19854 30236 19887
rect 30392 19854 30420 20266
rect 30196 19848 30248 19854
rect 30380 19848 30432 19854
rect 30196 19790 30248 19796
rect 30286 19816 30342 19825
rect 30104 19712 30156 19718
rect 30208 19689 30236 19790
rect 30380 19790 30432 19796
rect 30286 19751 30342 19760
rect 30104 19654 30156 19660
rect 30194 19680 30250 19689
rect 30194 19615 30250 19624
rect 30300 19496 30328 19751
rect 30208 19468 30328 19496
rect 30104 18964 30156 18970
rect 30104 18906 30156 18912
rect 30116 18630 30144 18906
rect 30012 18624 30064 18630
rect 30012 18566 30064 18572
rect 30104 18624 30156 18630
rect 30104 18566 30156 18572
rect 29918 18456 29974 18465
rect 29918 18391 29974 18400
rect 29920 17332 29972 17338
rect 29920 17274 29972 17280
rect 29932 17241 29960 17274
rect 29918 17232 29974 17241
rect 29918 17167 29974 17176
rect 29920 16652 29972 16658
rect 29920 16594 29972 16600
rect 29828 15088 29880 15094
rect 29828 15030 29880 15036
rect 29736 12912 29788 12918
rect 29736 12854 29788 12860
rect 29748 12442 29776 12854
rect 29736 12436 29788 12442
rect 29736 12378 29788 12384
rect 29644 11212 29696 11218
rect 29644 11154 29696 11160
rect 29748 11082 29776 12378
rect 29840 11626 29868 15030
rect 29932 11937 29960 16594
rect 30024 13190 30052 18566
rect 30104 18420 30156 18426
rect 30208 18408 30236 19468
rect 30288 19372 30340 19378
rect 30288 19314 30340 19320
rect 30156 18380 30236 18408
rect 30104 18362 30156 18368
rect 30104 18284 30156 18290
rect 30104 18226 30156 18232
rect 30116 17270 30144 18226
rect 30104 17264 30156 17270
rect 30104 17206 30156 17212
rect 30208 16454 30236 18380
rect 30300 17882 30328 19314
rect 30378 18864 30434 18873
rect 30378 18799 30434 18808
rect 30392 18426 30420 18799
rect 30380 18420 30432 18426
rect 30380 18362 30432 18368
rect 30484 18154 30512 21286
rect 30576 21146 30604 23734
rect 30656 22976 30708 22982
rect 30656 22918 30708 22924
rect 30564 21140 30616 21146
rect 30564 21082 30616 21088
rect 30564 20868 30616 20874
rect 30564 20810 30616 20816
rect 30576 20777 30604 20810
rect 30562 20768 30618 20777
rect 30562 20703 30618 20712
rect 30668 20584 30696 22918
rect 30760 22817 30788 26302
rect 31206 26302 31482 26330
rect 31206 26200 31262 26302
rect 31482 26279 31538 26288
rect 31850 26330 31906 27000
rect 31850 26302 32168 26330
rect 31850 26200 31906 26302
rect 31942 25936 31998 25945
rect 31942 25871 31998 25880
rect 31852 25696 31904 25702
rect 31852 25638 31904 25644
rect 31576 25424 31628 25430
rect 31576 25366 31628 25372
rect 31484 24200 31536 24206
rect 31484 24142 31536 24148
rect 31116 24132 31168 24138
rect 31116 24074 31168 24080
rect 31300 24132 31352 24138
rect 31300 24074 31352 24080
rect 30932 23792 30984 23798
rect 30932 23734 30984 23740
rect 30944 23254 30972 23734
rect 30932 23248 30984 23254
rect 30932 23190 30984 23196
rect 30944 23050 30972 23190
rect 31024 23112 31076 23118
rect 31024 23054 31076 23060
rect 30840 23044 30892 23050
rect 30840 22986 30892 22992
rect 30932 23044 30984 23050
rect 30932 22986 30984 22992
rect 30746 22808 30802 22817
rect 30852 22778 30880 22986
rect 30746 22743 30802 22752
rect 30840 22772 30892 22778
rect 30840 22714 30892 22720
rect 30748 21480 30800 21486
rect 30748 21422 30800 21428
rect 30760 21010 30788 21422
rect 30840 21412 30892 21418
rect 30840 21354 30892 21360
rect 30748 21004 30800 21010
rect 30748 20946 30800 20952
rect 30668 20556 30788 20584
rect 30656 20256 30708 20262
rect 30562 20224 30618 20233
rect 30656 20198 30708 20204
rect 30562 20159 30618 20168
rect 30576 18222 30604 20159
rect 30564 18216 30616 18222
rect 30564 18158 30616 18164
rect 30472 18148 30524 18154
rect 30472 18090 30524 18096
rect 30288 17876 30340 17882
rect 30288 17818 30340 17824
rect 30380 17876 30432 17882
rect 30380 17818 30432 17824
rect 30392 17678 30420 17818
rect 30380 17672 30432 17678
rect 30380 17614 30432 17620
rect 30392 16726 30420 17614
rect 30564 16992 30616 16998
rect 30564 16934 30616 16940
rect 30380 16720 30432 16726
rect 30380 16662 30432 16668
rect 30472 16720 30524 16726
rect 30472 16662 30524 16668
rect 30380 16516 30432 16522
rect 30380 16458 30432 16464
rect 30196 16448 30248 16454
rect 30196 16390 30248 16396
rect 30288 16448 30340 16454
rect 30288 16390 30340 16396
rect 30208 16114 30236 16390
rect 30300 16182 30328 16390
rect 30392 16250 30420 16458
rect 30380 16244 30432 16250
rect 30380 16186 30432 16192
rect 30288 16176 30340 16182
rect 30288 16118 30340 16124
rect 30196 16108 30248 16114
rect 30196 16050 30248 16056
rect 30380 15972 30432 15978
rect 30380 15914 30432 15920
rect 30102 15872 30158 15881
rect 30102 15807 30158 15816
rect 30116 14958 30144 15807
rect 30288 15496 30340 15502
rect 30288 15438 30340 15444
rect 30104 14952 30156 14958
rect 30104 14894 30156 14900
rect 30104 14816 30156 14822
rect 30104 14758 30156 14764
rect 30116 13326 30144 14758
rect 30196 14272 30248 14278
rect 30196 14214 30248 14220
rect 30208 13977 30236 14214
rect 30194 13968 30250 13977
rect 30194 13903 30250 13912
rect 30300 13734 30328 15438
rect 30392 14482 30420 15914
rect 30380 14476 30432 14482
rect 30380 14418 30432 14424
rect 30484 14278 30512 16662
rect 30472 14272 30524 14278
rect 30472 14214 30524 14220
rect 30380 14068 30432 14074
rect 30380 14010 30432 14016
rect 30288 13728 30340 13734
rect 30288 13670 30340 13676
rect 30196 13388 30248 13394
rect 30196 13330 30248 13336
rect 30104 13320 30156 13326
rect 30104 13262 30156 13268
rect 30012 13184 30064 13190
rect 30012 13126 30064 13132
rect 30010 12880 30066 12889
rect 30010 12815 30066 12824
rect 30024 12306 30052 12815
rect 30104 12640 30156 12646
rect 30104 12582 30156 12588
rect 30012 12300 30064 12306
rect 30012 12242 30064 12248
rect 29918 11928 29974 11937
rect 30116 11880 30144 12582
rect 29918 11863 29974 11872
rect 30024 11852 30144 11880
rect 29828 11620 29880 11626
rect 29828 11562 29880 11568
rect 29736 11076 29788 11082
rect 29736 11018 29788 11024
rect 30024 10962 30052 11852
rect 30104 11756 30156 11762
rect 30104 11698 30156 11704
rect 29748 10934 30052 10962
rect 29644 10668 29696 10674
rect 29644 10610 29696 10616
rect 29328 9540 29408 9568
rect 29472 9540 29592 9568
rect 29276 9522 29328 9528
rect 29092 9376 29144 9382
rect 29092 9318 29144 9324
rect 29184 9376 29236 9382
rect 29184 9318 29236 9324
rect 29000 9036 29052 9042
rect 29000 8978 29052 8984
rect 29000 8900 29052 8906
rect 29000 8842 29052 8848
rect 29012 7954 29040 8842
rect 29104 8566 29132 9318
rect 29288 8838 29316 9522
rect 29276 8832 29328 8838
rect 29276 8774 29328 8780
rect 29472 8634 29500 9540
rect 29552 9444 29604 9450
rect 29552 9386 29604 9392
rect 29460 8628 29512 8634
rect 29460 8570 29512 8576
rect 29092 8560 29144 8566
rect 29092 8502 29144 8508
rect 29000 7948 29052 7954
rect 29000 7890 29052 7896
rect 28448 6248 28500 6254
rect 28448 6190 28500 6196
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 27068 4616 27120 4622
rect 27068 4558 27120 4564
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 27344 4208 27396 4214
rect 27344 4150 27396 4156
rect 27160 4140 27212 4146
rect 27160 4082 27212 4088
rect 25688 4072 25740 4078
rect 25688 4014 25740 4020
rect 27172 4010 27200 4082
rect 27160 4004 27212 4010
rect 27160 3946 27212 3952
rect 27356 3738 27384 4150
rect 27344 3732 27396 3738
rect 27344 3674 27396 3680
rect 25872 3392 25924 3398
rect 25872 3334 25924 3340
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 24872 2514 24900 2790
rect 25884 2582 25912 3334
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 27712 3120 27764 3126
rect 27712 3062 27764 3068
rect 27620 3052 27672 3058
rect 27620 2994 27672 3000
rect 26516 2984 26568 2990
rect 26516 2926 26568 2932
rect 25872 2576 25924 2582
rect 25872 2518 25924 2524
rect 24860 2508 24912 2514
rect 24860 2450 24912 2456
rect 24952 2508 25004 2514
rect 24952 2450 25004 2456
rect 24964 2394 24992 2450
rect 24780 2372 24992 2394
rect 24780 2366 24860 2372
rect 24912 2366 24992 2372
rect 24860 2314 24912 2320
rect 26528 800 26556 2926
rect 27632 2650 27660 2994
rect 27620 2644 27672 2650
rect 27620 2586 27672 2592
rect 27724 2582 27752 3062
rect 29104 3058 29132 8502
rect 29564 7478 29592 9386
rect 29656 7546 29684 10610
rect 29644 7540 29696 7546
rect 29644 7482 29696 7488
rect 29552 7472 29604 7478
rect 29552 7414 29604 7420
rect 29748 7342 29776 10934
rect 29920 10736 29972 10742
rect 29920 10678 29972 10684
rect 29828 10192 29880 10198
rect 29828 10134 29880 10140
rect 29840 7886 29868 10134
rect 29932 9178 29960 10678
rect 30012 9512 30064 9518
rect 30012 9454 30064 9460
rect 29920 9172 29972 9178
rect 29920 9114 29972 9120
rect 29828 7880 29880 7886
rect 29828 7822 29880 7828
rect 29736 7336 29788 7342
rect 29736 7278 29788 7284
rect 30024 6866 30052 9454
rect 30116 9042 30144 11698
rect 30208 10198 30236 13330
rect 30300 12918 30328 13670
rect 30288 12912 30340 12918
rect 30288 12854 30340 12860
rect 30288 12164 30340 12170
rect 30288 12106 30340 12112
rect 30300 11898 30328 12106
rect 30392 12102 30420 14010
rect 30472 13184 30524 13190
rect 30472 13126 30524 13132
rect 30484 12170 30512 13126
rect 30472 12164 30524 12170
rect 30472 12106 30524 12112
rect 30380 12096 30432 12102
rect 30380 12038 30432 12044
rect 30288 11892 30340 11898
rect 30288 11834 30340 11840
rect 30484 11778 30512 12106
rect 30300 11750 30512 11778
rect 30300 11014 30328 11750
rect 30380 11076 30432 11082
rect 30380 11018 30432 11024
rect 30288 11008 30340 11014
rect 30288 10950 30340 10956
rect 30196 10192 30248 10198
rect 30196 10134 30248 10140
rect 30392 10062 30420 11018
rect 30576 10577 30604 16934
rect 30668 16250 30696 20198
rect 30760 19961 30788 20556
rect 30746 19952 30802 19961
rect 30746 19887 30802 19896
rect 30746 19544 30802 19553
rect 30746 19479 30802 19488
rect 30760 18970 30788 19479
rect 30852 19446 30880 21354
rect 31036 21332 31064 23054
rect 31128 21457 31156 24074
rect 31208 23112 31260 23118
rect 31208 23054 31260 23060
rect 31220 22506 31248 23054
rect 31208 22500 31260 22506
rect 31208 22442 31260 22448
rect 31220 22098 31248 22442
rect 31208 22092 31260 22098
rect 31208 22034 31260 22040
rect 31208 21956 31260 21962
rect 31208 21898 31260 21904
rect 31114 21448 31170 21457
rect 31114 21383 31170 21392
rect 31036 21304 31156 21332
rect 31128 20330 31156 21304
rect 31220 20924 31248 21898
rect 31312 21486 31340 24074
rect 31496 22982 31524 24142
rect 31484 22976 31536 22982
rect 31484 22918 31536 22924
rect 31390 22128 31446 22137
rect 31390 22063 31446 22072
rect 31404 21962 31432 22063
rect 31392 21956 31444 21962
rect 31392 21898 31444 21904
rect 31300 21480 31352 21486
rect 31300 21422 31352 21428
rect 31300 20936 31352 20942
rect 31220 20896 31300 20924
rect 31220 20534 31248 20896
rect 31300 20878 31352 20884
rect 31300 20800 31352 20806
rect 31300 20742 31352 20748
rect 31208 20528 31260 20534
rect 31208 20470 31260 20476
rect 31208 20392 31260 20398
rect 31208 20334 31260 20340
rect 31116 20324 31168 20330
rect 31116 20266 31168 20272
rect 30932 20256 30984 20262
rect 31220 20233 31248 20334
rect 30932 20198 30984 20204
rect 31206 20224 31262 20233
rect 30840 19440 30892 19446
rect 30840 19382 30892 19388
rect 30748 18964 30800 18970
rect 30748 18906 30800 18912
rect 30760 18834 30788 18906
rect 30748 18828 30800 18834
rect 30748 18770 30800 18776
rect 30852 17882 30880 19382
rect 30944 19378 30972 20198
rect 31206 20159 31262 20168
rect 31312 20074 31340 20742
rect 31390 20632 31446 20641
rect 31390 20567 31446 20576
rect 31404 20097 31432 20567
rect 31128 20046 31340 20074
rect 31390 20088 31446 20097
rect 31024 19848 31076 19854
rect 31024 19790 31076 19796
rect 30932 19372 30984 19378
rect 30932 19314 30984 19320
rect 30932 18080 30984 18086
rect 30932 18022 30984 18028
rect 30840 17876 30892 17882
rect 30840 17818 30892 17824
rect 30838 17776 30894 17785
rect 30838 17711 30894 17720
rect 30748 17264 30800 17270
rect 30748 17206 30800 17212
rect 30760 17134 30788 17206
rect 30748 17128 30800 17134
rect 30748 17070 30800 17076
rect 30656 16244 30708 16250
rect 30656 16186 30708 16192
rect 30760 16130 30788 17070
rect 30668 16102 30788 16130
rect 30562 10568 30618 10577
rect 30562 10503 30618 10512
rect 30668 10248 30696 16102
rect 30852 16046 30880 17711
rect 30944 16182 30972 18022
rect 31036 17678 31064 19790
rect 31128 18426 31156 20046
rect 31390 20023 31446 20032
rect 31298 19952 31354 19961
rect 31404 19922 31432 20023
rect 31496 19922 31524 22918
rect 31588 20874 31616 25366
rect 31668 24064 31720 24070
rect 31668 24006 31720 24012
rect 31680 23186 31708 24006
rect 31668 23180 31720 23186
rect 31668 23122 31720 23128
rect 31864 22953 31892 25638
rect 31850 22944 31906 22953
rect 31850 22879 31906 22888
rect 31760 22772 31812 22778
rect 31760 22714 31812 22720
rect 31668 22568 31720 22574
rect 31668 22510 31720 22516
rect 31680 22234 31708 22510
rect 31668 22228 31720 22234
rect 31668 22170 31720 22176
rect 31772 21894 31800 22714
rect 31760 21888 31812 21894
rect 31760 21830 31812 21836
rect 31760 21684 31812 21690
rect 31760 21626 31812 21632
rect 31666 21448 31722 21457
rect 31666 21383 31722 21392
rect 31576 20868 31628 20874
rect 31576 20810 31628 20816
rect 31298 19887 31354 19896
rect 31392 19916 31444 19922
rect 31312 19854 31340 19887
rect 31392 19858 31444 19864
rect 31484 19916 31536 19922
rect 31484 19858 31536 19864
rect 31300 19848 31352 19854
rect 31300 19790 31352 19796
rect 31208 19780 31260 19786
rect 31208 19722 31260 19728
rect 31220 19378 31248 19722
rect 31208 19372 31260 19378
rect 31208 19314 31260 19320
rect 31220 18766 31248 19314
rect 31576 19236 31628 19242
rect 31576 19178 31628 19184
rect 31482 19136 31538 19145
rect 31482 19071 31538 19080
rect 31208 18760 31260 18766
rect 31208 18702 31260 18708
rect 31392 18692 31444 18698
rect 31392 18634 31444 18640
rect 31300 18624 31352 18630
rect 31300 18566 31352 18572
rect 31116 18420 31168 18426
rect 31116 18362 31168 18368
rect 31024 17672 31076 17678
rect 31024 17614 31076 17620
rect 31022 17368 31078 17377
rect 31022 17303 31078 17312
rect 31036 16726 31064 17303
rect 31208 16992 31260 16998
rect 31208 16934 31260 16940
rect 31024 16720 31076 16726
rect 31024 16662 31076 16668
rect 30932 16176 30984 16182
rect 30932 16118 30984 16124
rect 30840 16040 30892 16046
rect 30840 15982 30892 15988
rect 31116 15972 31168 15978
rect 31116 15914 31168 15920
rect 31128 15881 31156 15914
rect 31114 15872 31170 15881
rect 31114 15807 31170 15816
rect 31024 15428 31076 15434
rect 31024 15370 31076 15376
rect 31036 15337 31064 15370
rect 31116 15360 31168 15366
rect 31022 15328 31078 15337
rect 31116 15302 31168 15308
rect 31022 15263 31078 15272
rect 30748 14952 30800 14958
rect 30748 14894 30800 14900
rect 31024 14952 31076 14958
rect 31024 14894 31076 14900
rect 30760 14793 30788 14894
rect 30932 14884 30984 14890
rect 30932 14826 30984 14832
rect 30746 14784 30802 14793
rect 30746 14719 30802 14728
rect 30840 14612 30892 14618
rect 30944 14600 30972 14826
rect 30892 14572 30972 14600
rect 30840 14554 30892 14560
rect 30748 14476 30800 14482
rect 30748 14418 30800 14424
rect 30760 11626 30788 14418
rect 31036 14414 31064 14894
rect 31128 14414 31156 15302
rect 31024 14408 31076 14414
rect 31024 14350 31076 14356
rect 31116 14408 31168 14414
rect 31116 14350 31168 14356
rect 30840 13864 30892 13870
rect 30840 13806 30892 13812
rect 31114 13832 31170 13841
rect 30852 13462 30880 13806
rect 31114 13767 31170 13776
rect 30840 13456 30892 13462
rect 30840 13398 30892 13404
rect 31024 12640 31076 12646
rect 31024 12582 31076 12588
rect 31036 12345 31064 12582
rect 31022 12336 31078 12345
rect 31022 12271 31078 12280
rect 30930 12064 30986 12073
rect 30930 11999 30986 12008
rect 30748 11620 30800 11626
rect 30748 11562 30800 11568
rect 30944 10538 30972 11999
rect 30932 10532 30984 10538
rect 30932 10474 30984 10480
rect 30576 10220 30696 10248
rect 30380 10056 30432 10062
rect 30576 10033 30604 10220
rect 30380 9998 30432 10004
rect 30562 10024 30618 10033
rect 30392 9908 30420 9998
rect 30562 9959 30564 9968
rect 30616 9959 30618 9968
rect 30656 9988 30708 9994
rect 30564 9930 30616 9936
rect 30656 9930 30708 9936
rect 30300 9880 30420 9908
rect 30300 9654 30328 9880
rect 30288 9648 30340 9654
rect 30288 9590 30340 9596
rect 30472 9172 30524 9178
rect 30472 9114 30524 9120
rect 30104 9036 30156 9042
rect 30104 8978 30156 8984
rect 30380 8832 30432 8838
rect 30380 8774 30432 8780
rect 30392 8566 30420 8774
rect 30380 8560 30432 8566
rect 30380 8502 30432 8508
rect 30380 8424 30432 8430
rect 30380 8366 30432 8372
rect 30392 8090 30420 8366
rect 30380 8084 30432 8090
rect 30380 8026 30432 8032
rect 30012 6860 30064 6866
rect 30012 6802 30064 6808
rect 30484 6798 30512 9114
rect 30668 8022 30696 9930
rect 30748 8968 30800 8974
rect 30748 8910 30800 8916
rect 30760 8566 30788 8910
rect 31024 8832 31076 8838
rect 31024 8774 31076 8780
rect 31036 8634 31064 8774
rect 31024 8628 31076 8634
rect 31024 8570 31076 8576
rect 30748 8560 30800 8566
rect 30748 8502 30800 8508
rect 30748 8424 30800 8430
rect 30748 8366 30800 8372
rect 30656 8016 30708 8022
rect 30656 7958 30708 7964
rect 30760 7750 30788 8366
rect 31128 7954 31156 13767
rect 31220 11880 31248 16934
rect 31312 13734 31340 18566
rect 31404 18222 31432 18634
rect 31392 18216 31444 18222
rect 31392 18158 31444 18164
rect 31392 16992 31444 16998
rect 31392 16934 31444 16940
rect 31404 16658 31432 16934
rect 31392 16652 31444 16658
rect 31392 16594 31444 16600
rect 31390 16280 31446 16289
rect 31390 16215 31446 16224
rect 31300 13728 31352 13734
rect 31300 13670 31352 13676
rect 31404 13138 31432 16215
rect 31496 14414 31524 19071
rect 31588 18222 31616 19178
rect 31680 18601 31708 21383
rect 31772 21350 31800 21626
rect 31760 21344 31812 21350
rect 31760 21286 31812 21292
rect 31760 21072 31812 21078
rect 31760 21014 31812 21020
rect 31772 19378 31800 21014
rect 31864 20942 31892 22879
rect 31852 20936 31904 20942
rect 31852 20878 31904 20884
rect 31852 20800 31904 20806
rect 31852 20742 31904 20748
rect 31864 19689 31892 20742
rect 31850 19680 31906 19689
rect 31850 19615 31906 19624
rect 31760 19372 31812 19378
rect 31760 19314 31812 19320
rect 31852 19372 31904 19378
rect 31852 19314 31904 19320
rect 31864 18850 31892 19314
rect 31772 18822 31892 18850
rect 31666 18592 31722 18601
rect 31666 18527 31722 18536
rect 31772 18358 31800 18822
rect 31956 18714 31984 25871
rect 32140 25129 32168 26302
rect 32494 26200 32550 27000
rect 33138 26330 33194 27000
rect 33138 26302 33456 26330
rect 32586 26208 32642 26217
rect 32508 26160 32536 26200
rect 32508 26152 32586 26160
rect 33138 26200 33194 26302
rect 33428 26178 33456 26302
rect 33782 26200 33838 27000
rect 34426 26200 34482 27000
rect 35070 26330 35126 27000
rect 35714 26330 35770 27000
rect 36358 26330 36414 27000
rect 35070 26302 35480 26330
rect 35070 26200 35126 26302
rect 32508 26143 32642 26152
rect 33416 26172 33468 26178
rect 32508 26132 32628 26143
rect 33416 26114 33468 26120
rect 33796 26042 33824 26200
rect 34440 26110 34468 26200
rect 34428 26104 34480 26110
rect 34428 26046 34480 26052
rect 33784 26036 33836 26042
rect 33784 25978 33836 25984
rect 32126 25120 32182 25129
rect 32126 25055 32182 25064
rect 33324 25016 33376 25022
rect 33324 24958 33376 24964
rect 32218 24712 32274 24721
rect 32218 24647 32274 24656
rect 32128 24064 32180 24070
rect 32128 24006 32180 24012
rect 32140 23905 32168 24006
rect 32126 23896 32182 23905
rect 32126 23831 32182 23840
rect 32140 23050 32168 23831
rect 32128 23044 32180 23050
rect 32128 22986 32180 22992
rect 32140 21962 32168 22986
rect 32128 21956 32180 21962
rect 32128 21898 32180 21904
rect 32140 21690 32168 21898
rect 32232 21865 32260 24647
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 32680 23724 32732 23730
rect 32680 23666 32732 23672
rect 32588 23656 32640 23662
rect 32588 23598 32640 23604
rect 32600 22953 32628 23598
rect 32586 22944 32642 22953
rect 32586 22879 32642 22888
rect 32496 22636 32548 22642
rect 32496 22578 32548 22584
rect 32508 22234 32536 22578
rect 32496 22228 32548 22234
rect 32496 22170 32548 22176
rect 32600 22166 32628 22879
rect 32588 22160 32640 22166
rect 32588 22102 32640 22108
rect 32312 22092 32364 22098
rect 32312 22034 32364 22040
rect 32218 21856 32274 21865
rect 32218 21791 32274 21800
rect 32128 21684 32180 21690
rect 32128 21626 32180 21632
rect 32036 21480 32088 21486
rect 32036 21422 32088 21428
rect 32048 19514 32076 21422
rect 32140 20913 32168 21626
rect 32126 20904 32182 20913
rect 32126 20839 32182 20848
rect 32232 19922 32260 21791
rect 32324 20942 32352 22034
rect 32692 21894 32720 23666
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 32864 23180 32916 23186
rect 32864 23122 32916 23128
rect 32772 22568 32824 22574
rect 32772 22510 32824 22516
rect 32680 21888 32732 21894
rect 32680 21830 32732 21836
rect 32404 21684 32456 21690
rect 32404 21626 32456 21632
rect 32416 21078 32444 21626
rect 32496 21480 32548 21486
rect 32496 21422 32548 21428
rect 32508 21350 32536 21422
rect 32496 21344 32548 21350
rect 32496 21286 32548 21292
rect 32588 21344 32640 21350
rect 32588 21286 32640 21292
rect 32404 21072 32456 21078
rect 32404 21014 32456 21020
rect 32312 20936 32364 20942
rect 32312 20878 32364 20884
rect 32324 20398 32352 20878
rect 32312 20392 32364 20398
rect 32312 20334 32364 20340
rect 32220 19916 32272 19922
rect 32220 19858 32272 19864
rect 32128 19712 32180 19718
rect 32128 19654 32180 19660
rect 32036 19508 32088 19514
rect 32036 19450 32088 19456
rect 32036 19168 32088 19174
rect 32036 19110 32088 19116
rect 32048 18902 32076 19110
rect 32036 18896 32088 18902
rect 32036 18838 32088 18844
rect 31864 18686 31984 18714
rect 31760 18352 31812 18358
rect 31760 18294 31812 18300
rect 31576 18216 31628 18222
rect 31576 18158 31628 18164
rect 31576 18080 31628 18086
rect 31576 18022 31628 18028
rect 31484 14408 31536 14414
rect 31484 14350 31536 14356
rect 31482 13288 31538 13297
rect 31482 13223 31484 13232
rect 31536 13223 31538 13232
rect 31484 13194 31536 13200
rect 31404 13110 31524 13138
rect 31392 12844 31444 12850
rect 31392 12786 31444 12792
rect 31404 12374 31432 12786
rect 31392 12368 31444 12374
rect 31392 12310 31444 12316
rect 31300 11892 31352 11898
rect 31220 11852 31300 11880
rect 31300 11834 31352 11840
rect 31404 11354 31432 12310
rect 31392 11348 31444 11354
rect 31392 11290 31444 11296
rect 31496 10810 31524 13110
rect 31588 12782 31616 18022
rect 31758 17912 31814 17921
rect 31758 17847 31814 17856
rect 31668 17740 31720 17746
rect 31668 17682 31720 17688
rect 31680 16522 31708 17682
rect 31772 16998 31800 17847
rect 31760 16992 31812 16998
rect 31760 16934 31812 16940
rect 31758 16552 31814 16561
rect 31668 16516 31720 16522
rect 31758 16487 31760 16496
rect 31668 16458 31720 16464
rect 31812 16487 31814 16496
rect 31760 16458 31812 16464
rect 31680 14482 31708 16458
rect 31864 15706 31892 18686
rect 32036 18624 32088 18630
rect 32036 18566 32088 18572
rect 31944 17876 31996 17882
rect 31944 17818 31996 17824
rect 31956 17678 31984 17818
rect 31944 17672 31996 17678
rect 31944 17614 31996 17620
rect 32048 17338 32076 18566
rect 32036 17332 32088 17338
rect 32036 17274 32088 17280
rect 31944 16992 31996 16998
rect 31944 16934 31996 16940
rect 31956 16250 31984 16934
rect 32140 16794 32168 19654
rect 32220 19508 32272 19514
rect 32220 19450 32272 19456
rect 32232 19378 32260 19450
rect 32324 19378 32352 20334
rect 32508 19854 32536 21286
rect 32496 19848 32548 19854
rect 32496 19790 32548 19796
rect 32404 19712 32456 19718
rect 32404 19654 32456 19660
rect 32220 19372 32272 19378
rect 32220 19314 32272 19320
rect 32312 19372 32364 19378
rect 32312 19314 32364 19320
rect 32220 18828 32272 18834
rect 32220 18770 32272 18776
rect 32128 16788 32180 16794
rect 32128 16730 32180 16736
rect 31944 16244 31996 16250
rect 31944 16186 31996 16192
rect 31852 15700 31904 15706
rect 31852 15642 31904 15648
rect 32036 15496 32088 15502
rect 32036 15438 32088 15444
rect 31758 15328 31814 15337
rect 31758 15263 31814 15272
rect 31668 14476 31720 14482
rect 31668 14418 31720 14424
rect 31666 14240 31722 14249
rect 31666 14175 31722 14184
rect 31576 12776 31628 12782
rect 31574 12744 31576 12753
rect 31628 12744 31630 12753
rect 31574 12679 31630 12688
rect 31680 11200 31708 14175
rect 31772 12209 31800 15263
rect 32048 14550 32076 15438
rect 32036 14544 32088 14550
rect 32036 14486 32088 14492
rect 32036 14272 32088 14278
rect 32232 14249 32260 18770
rect 32312 18216 32364 18222
rect 32312 18158 32364 18164
rect 32324 15638 32352 18158
rect 32416 16538 32444 19654
rect 32496 18148 32548 18154
rect 32496 18090 32548 18096
rect 32508 17610 32536 18090
rect 32600 17882 32628 21286
rect 32784 21049 32812 22510
rect 32770 21040 32826 21049
rect 32876 21010 32904 23122
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 33336 22098 33364 24958
rect 34244 24812 34296 24818
rect 34244 24754 34296 24760
rect 34060 24744 34112 24750
rect 34060 24686 34112 24692
rect 33414 24304 33470 24313
rect 34072 24274 34100 24686
rect 34256 24274 34284 24754
rect 35256 24336 35308 24342
rect 35256 24278 35308 24284
rect 33414 24239 33470 24248
rect 34060 24268 34112 24274
rect 33428 22778 33456 24239
rect 34060 24210 34112 24216
rect 34244 24268 34296 24274
rect 34244 24210 34296 24216
rect 35072 24200 35124 24206
rect 35072 24142 35124 24148
rect 33876 24132 33928 24138
rect 33876 24074 33928 24080
rect 33600 24064 33652 24070
rect 33600 24006 33652 24012
rect 33612 23769 33640 24006
rect 33784 23792 33836 23798
rect 33598 23760 33654 23769
rect 33784 23734 33836 23740
rect 33598 23695 33654 23704
rect 33508 23656 33560 23662
rect 33508 23598 33560 23604
rect 33520 22778 33548 23598
rect 33796 23322 33824 23734
rect 33784 23316 33836 23322
rect 33784 23258 33836 23264
rect 33416 22772 33468 22778
rect 33416 22714 33468 22720
rect 33508 22772 33560 22778
rect 33508 22714 33560 22720
rect 33324 22092 33376 22098
rect 33324 22034 33376 22040
rect 33140 21888 33192 21894
rect 33060 21836 33140 21842
rect 33060 21830 33192 21836
rect 33060 21814 33180 21830
rect 33060 21486 33088 21814
rect 33428 21729 33456 22714
rect 33600 22704 33652 22710
rect 33652 22652 33732 22658
rect 33600 22646 33732 22652
rect 33612 22630 33732 22646
rect 33704 22506 33732 22630
rect 33692 22500 33744 22506
rect 33692 22442 33744 22448
rect 33796 22166 33824 23258
rect 33888 22710 33916 24074
rect 34242 23896 34298 23905
rect 34242 23831 34298 23840
rect 34256 23798 34284 23831
rect 34244 23792 34296 23798
rect 34244 23734 34296 23740
rect 33968 23112 34020 23118
rect 33968 23054 34020 23060
rect 33876 22704 33928 22710
rect 33876 22646 33928 22652
rect 33784 22160 33836 22166
rect 33784 22102 33836 22108
rect 33508 22092 33560 22098
rect 33508 22034 33560 22040
rect 33876 22092 33928 22098
rect 33876 22034 33928 22040
rect 33414 21720 33470 21729
rect 33414 21655 33470 21664
rect 33048 21480 33100 21486
rect 33048 21422 33100 21428
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 32770 20975 32826 20984
rect 32864 21004 32916 21010
rect 32864 20946 32916 20952
rect 33140 21004 33192 21010
rect 33140 20946 33192 20952
rect 33046 20904 33102 20913
rect 33152 20890 33180 20946
rect 33102 20862 33180 20890
rect 33046 20839 33048 20848
rect 33100 20839 33102 20848
rect 33048 20810 33100 20816
rect 33060 20534 33088 20810
rect 33048 20528 33100 20534
rect 33048 20470 33100 20476
rect 32680 20392 32732 20398
rect 32680 20334 32732 20340
rect 32692 19825 32720 20334
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 32864 19916 32916 19922
rect 32864 19858 32916 19864
rect 32956 19916 33008 19922
rect 32956 19858 33008 19864
rect 32772 19848 32824 19854
rect 32678 19816 32734 19825
rect 32772 19790 32824 19796
rect 32678 19751 32734 19760
rect 32784 19514 32812 19790
rect 32772 19508 32824 19514
rect 32772 19450 32824 19456
rect 32678 19408 32734 19417
rect 32678 19343 32734 19352
rect 32588 17876 32640 17882
rect 32588 17818 32640 17824
rect 32496 17604 32548 17610
rect 32496 17546 32548 17552
rect 32508 17270 32536 17546
rect 32600 17270 32628 17818
rect 32496 17264 32548 17270
rect 32496 17206 32548 17212
rect 32588 17264 32640 17270
rect 32588 17206 32640 17212
rect 32508 16658 32536 17206
rect 32496 16652 32548 16658
rect 32496 16594 32548 16600
rect 32416 16510 32536 16538
rect 32508 15745 32536 16510
rect 32692 16250 32720 19343
rect 32876 19224 32904 19858
rect 32968 19378 32996 19858
rect 33048 19712 33100 19718
rect 33048 19654 33100 19660
rect 33060 19378 33088 19654
rect 33428 19530 33456 21655
rect 33520 20058 33548 22034
rect 33888 21729 33916 22034
rect 33874 21720 33930 21729
rect 33874 21655 33930 21664
rect 33600 21548 33652 21554
rect 33600 21490 33652 21496
rect 33612 21321 33640 21490
rect 33692 21480 33744 21486
rect 33690 21448 33692 21457
rect 33744 21448 33746 21457
rect 33690 21383 33746 21392
rect 33598 21312 33654 21321
rect 33598 21247 33654 21256
rect 33888 20913 33916 21655
rect 33874 20904 33930 20913
rect 33874 20839 33930 20848
rect 33784 20800 33836 20806
rect 33980 20754 34008 23054
rect 34256 22710 34284 23734
rect 34888 23180 34940 23186
rect 34888 23122 34940 23128
rect 34900 22778 34928 23122
rect 34888 22772 34940 22778
rect 34888 22714 34940 22720
rect 34244 22704 34296 22710
rect 34058 22672 34114 22681
rect 34244 22646 34296 22652
rect 34058 22607 34114 22616
rect 33836 20748 34008 20754
rect 33784 20742 34008 20748
rect 33796 20726 34008 20742
rect 33980 20602 34008 20726
rect 33968 20596 34020 20602
rect 33968 20538 34020 20544
rect 33692 20324 33744 20330
rect 33692 20266 33744 20272
rect 33508 20052 33560 20058
rect 33508 19994 33560 20000
rect 33336 19502 33456 19530
rect 32956 19372 33008 19378
rect 32956 19314 33008 19320
rect 33048 19372 33100 19378
rect 33048 19314 33100 19320
rect 33232 19304 33284 19310
rect 33230 19272 33232 19281
rect 33284 19272 33286 19281
rect 32956 19236 33008 19242
rect 32876 19196 32956 19224
rect 33230 19207 33286 19216
rect 32956 19178 33008 19184
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 33140 18964 33192 18970
rect 33140 18906 33192 18912
rect 33152 18329 33180 18906
rect 33138 18320 33194 18329
rect 33138 18255 33140 18264
rect 33192 18255 33194 18264
rect 33140 18226 33192 18232
rect 32864 18216 32916 18222
rect 32864 18158 32916 18164
rect 32876 17882 32904 18158
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 32864 17876 32916 17882
rect 32864 17818 32916 17824
rect 32772 17536 32824 17542
rect 32772 17478 32824 17484
rect 32784 17338 32812 17478
rect 32772 17332 32824 17338
rect 32772 17274 32824 17280
rect 32876 16726 32904 17818
rect 33336 17762 33364 19502
rect 33508 19304 33560 19310
rect 33508 19246 33560 19252
rect 33520 18834 33548 19246
rect 33508 18828 33560 18834
rect 33508 18770 33560 18776
rect 33600 18624 33652 18630
rect 33600 18566 33652 18572
rect 33612 18465 33640 18566
rect 33414 18456 33470 18465
rect 33414 18391 33416 18400
rect 33468 18391 33470 18400
rect 33598 18456 33654 18465
rect 33598 18391 33654 18400
rect 33416 18362 33468 18368
rect 33600 18352 33652 18358
rect 33600 18294 33652 18300
rect 33244 17746 33364 17762
rect 33232 17740 33364 17746
rect 33284 17734 33364 17740
rect 33232 17682 33284 17688
rect 33244 17134 33272 17682
rect 33232 17128 33284 17134
rect 33232 17070 33284 17076
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 33508 16788 33560 16794
rect 33508 16730 33560 16736
rect 32864 16720 32916 16726
rect 32864 16662 32916 16668
rect 32876 16266 32904 16662
rect 32956 16652 33008 16658
rect 32956 16594 33008 16600
rect 32680 16244 32732 16250
rect 32680 16186 32732 16192
rect 32784 16238 32904 16266
rect 32494 15736 32550 15745
rect 32494 15671 32550 15680
rect 32312 15632 32364 15638
rect 32312 15574 32364 15580
rect 32784 15502 32812 16238
rect 32862 16144 32918 16153
rect 32862 16079 32918 16088
rect 32876 15570 32904 16079
rect 32968 16046 32996 16594
rect 32956 16040 33008 16046
rect 32956 15982 33008 15988
rect 33520 15994 33548 16730
rect 33612 16590 33640 18294
rect 33704 17746 33732 20266
rect 34072 20262 34100 22607
rect 34428 22568 34480 22574
rect 34428 22510 34480 22516
rect 34612 22568 34664 22574
rect 34612 22510 34664 22516
rect 34440 22386 34468 22510
rect 34440 22358 34560 22386
rect 34244 22228 34296 22234
rect 34244 22170 34296 22176
rect 34256 21622 34284 22170
rect 34336 22160 34388 22166
rect 34336 22102 34388 22108
rect 34244 21616 34296 21622
rect 34244 21558 34296 21564
rect 34152 20800 34204 20806
rect 34152 20742 34204 20748
rect 34060 20256 34112 20262
rect 34060 20198 34112 20204
rect 33874 20088 33930 20097
rect 33874 20023 33930 20032
rect 33968 20052 34020 20058
rect 33888 19922 33916 20023
rect 33968 19994 34020 20000
rect 33876 19916 33928 19922
rect 33876 19858 33928 19864
rect 33980 19378 34008 19994
rect 34060 19916 34112 19922
rect 34060 19858 34112 19864
rect 33876 19372 33928 19378
rect 33876 19314 33928 19320
rect 33968 19372 34020 19378
rect 33968 19314 34020 19320
rect 33888 19281 33916 19314
rect 33874 19272 33930 19281
rect 33874 19207 33930 19216
rect 33968 19236 34020 19242
rect 33968 19178 34020 19184
rect 33980 18873 34008 19178
rect 33782 18864 33838 18873
rect 33966 18864 34022 18873
rect 33782 18799 33838 18808
rect 33876 18828 33928 18834
rect 33796 17882 33824 18799
rect 33966 18799 34022 18808
rect 33876 18770 33928 18776
rect 33888 18612 33916 18770
rect 33968 18624 34020 18630
rect 33888 18584 33968 18612
rect 33968 18566 34020 18572
rect 33876 18216 33928 18222
rect 33876 18158 33928 18164
rect 33784 17876 33836 17882
rect 33784 17818 33836 17824
rect 33692 17740 33744 17746
rect 33692 17682 33744 17688
rect 33784 17536 33836 17542
rect 33784 17478 33836 17484
rect 33692 17060 33744 17066
rect 33692 17002 33744 17008
rect 33600 16584 33652 16590
rect 33600 16526 33652 16532
rect 33520 15966 33640 15994
rect 33416 15904 33468 15910
rect 33416 15846 33468 15852
rect 33508 15904 33560 15910
rect 33508 15846 33560 15852
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 33048 15632 33100 15638
rect 33048 15574 33100 15580
rect 32864 15564 32916 15570
rect 32864 15506 32916 15512
rect 32772 15496 32824 15502
rect 32772 15438 32824 15444
rect 33060 15366 33088 15574
rect 32772 15360 32824 15366
rect 32772 15302 32824 15308
rect 33048 15360 33100 15366
rect 33048 15302 33100 15308
rect 32680 15020 32732 15026
rect 32680 14962 32732 14968
rect 32588 14952 32640 14958
rect 32588 14894 32640 14900
rect 32600 14278 32628 14894
rect 32588 14272 32640 14278
rect 32036 14214 32088 14220
rect 32218 14240 32274 14249
rect 31852 13796 31904 13802
rect 31852 13738 31904 13744
rect 31864 12889 31892 13738
rect 31944 13252 31996 13258
rect 31944 13194 31996 13200
rect 31850 12880 31906 12889
rect 31850 12815 31906 12824
rect 31758 12200 31814 12209
rect 31758 12135 31814 12144
rect 31956 11694 31984 13194
rect 31944 11688 31996 11694
rect 32048 11665 32076 14214
rect 32588 14214 32640 14220
rect 32218 14175 32274 14184
rect 32220 13864 32272 13870
rect 32220 13806 32272 13812
rect 32588 13864 32640 13870
rect 32588 13806 32640 13812
rect 32232 13394 32260 13806
rect 32600 13433 32628 13806
rect 32586 13424 32642 13433
rect 32220 13388 32272 13394
rect 32586 13359 32642 13368
rect 32220 13330 32272 13336
rect 32128 13184 32180 13190
rect 32128 13126 32180 13132
rect 32140 11778 32168 13126
rect 32232 12850 32260 13330
rect 32312 13184 32364 13190
rect 32312 13126 32364 13132
rect 32324 12986 32352 13126
rect 32312 12980 32364 12986
rect 32312 12922 32364 12928
rect 32496 12912 32548 12918
rect 32496 12854 32548 12860
rect 32220 12844 32272 12850
rect 32220 12786 32272 12792
rect 32232 12306 32260 12786
rect 32220 12300 32272 12306
rect 32220 12242 32272 12248
rect 32140 11750 32444 11778
rect 32312 11688 32364 11694
rect 31944 11630 31996 11636
rect 32034 11656 32090 11665
rect 32312 11630 32364 11636
rect 32034 11591 32090 11600
rect 32324 11558 32352 11630
rect 31760 11552 31812 11558
rect 32312 11552 32364 11558
rect 31812 11500 32076 11506
rect 31760 11494 32076 11500
rect 32312 11494 32364 11500
rect 31772 11478 32076 11494
rect 31760 11212 31812 11218
rect 31680 11172 31760 11200
rect 31760 11154 31812 11160
rect 31574 11112 31630 11121
rect 31574 11047 31630 11056
rect 31484 10804 31536 10810
rect 31484 10746 31536 10752
rect 31300 10668 31352 10674
rect 31300 10610 31352 10616
rect 31312 10130 31340 10610
rect 31588 10606 31616 11047
rect 31576 10600 31628 10606
rect 31576 10542 31628 10548
rect 31392 10464 31444 10470
rect 31392 10406 31444 10412
rect 31484 10464 31536 10470
rect 31484 10406 31536 10412
rect 31404 10130 31432 10406
rect 31300 10124 31352 10130
rect 31300 10066 31352 10072
rect 31392 10124 31444 10130
rect 31392 10066 31444 10072
rect 31496 9382 31524 10406
rect 31772 10266 31800 11154
rect 31760 10260 31812 10266
rect 31760 10202 31812 10208
rect 31668 9444 31720 9450
rect 31668 9386 31720 9392
rect 31484 9376 31536 9382
rect 31484 9318 31536 9324
rect 31300 8900 31352 8906
rect 31300 8842 31352 8848
rect 31312 8634 31340 8842
rect 31300 8628 31352 8634
rect 31300 8570 31352 8576
rect 31116 7948 31168 7954
rect 31116 7890 31168 7896
rect 30748 7744 30800 7750
rect 30748 7686 30800 7692
rect 30472 6792 30524 6798
rect 30472 6734 30524 6740
rect 30656 3936 30708 3942
rect 30656 3878 30708 3884
rect 29092 3052 29144 3058
rect 29092 2994 29144 3000
rect 27436 2576 27488 2582
rect 27436 2518 27488 2524
rect 27712 2576 27764 2582
rect 27712 2518 27764 2524
rect 27448 2378 27476 2518
rect 28632 2440 28684 2446
rect 28632 2382 28684 2388
rect 27436 2372 27488 2378
rect 27436 2314 27488 2320
rect 27160 2304 27212 2310
rect 27160 2246 27212 2252
rect 27172 2106 27200 2246
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 27160 2100 27212 2106
rect 27160 2042 27212 2048
rect 28644 800 28672 2382
rect 30668 2310 30696 3878
rect 30760 3194 30788 7686
rect 31128 7002 31156 7890
rect 31116 6996 31168 7002
rect 31116 6938 31168 6944
rect 31312 5302 31340 8570
rect 31392 8492 31444 8498
rect 31392 8434 31444 8440
rect 31404 7546 31432 8434
rect 31392 7540 31444 7546
rect 31392 7482 31444 7488
rect 31496 7410 31524 9318
rect 31680 8430 31708 9386
rect 32048 9110 32076 11478
rect 32324 11014 32352 11494
rect 32312 11008 32364 11014
rect 32312 10950 32364 10956
rect 32324 9994 32352 10950
rect 32312 9988 32364 9994
rect 32312 9930 32364 9936
rect 32324 9586 32352 9930
rect 32416 9586 32444 11750
rect 32508 10266 32536 12854
rect 32692 11898 32720 14962
rect 32784 14074 32812 15302
rect 33230 15192 33286 15201
rect 33230 15127 33286 15136
rect 33244 14822 33272 15127
rect 33324 14952 33376 14958
rect 33324 14894 33376 14900
rect 33232 14816 33284 14822
rect 33232 14758 33284 14764
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 32864 14544 32916 14550
rect 32864 14486 32916 14492
rect 33230 14512 33286 14521
rect 32772 14068 32824 14074
rect 32772 14010 32824 14016
rect 32876 13326 32904 14486
rect 32956 14476 33008 14482
rect 33230 14447 33286 14456
rect 32956 14418 33008 14424
rect 32968 14249 32996 14418
rect 33140 14340 33192 14346
rect 33140 14282 33192 14288
rect 32954 14240 33010 14249
rect 32954 14175 33010 14184
rect 33152 13870 33180 14282
rect 33140 13864 33192 13870
rect 33140 13806 33192 13812
rect 33244 13716 33272 14447
rect 33336 14249 33364 14894
rect 33428 14414 33456 15846
rect 33520 14521 33548 15846
rect 33506 14512 33562 14521
rect 33612 14482 33640 15966
rect 33704 14793 33732 17002
rect 33796 15978 33824 17478
rect 33888 16998 33916 18158
rect 33980 18057 34008 18566
rect 34072 18442 34100 19858
rect 34164 19310 34192 20742
rect 34348 20369 34376 22102
rect 34532 22094 34560 22358
rect 34440 22066 34560 22094
rect 34440 21554 34468 22066
rect 34520 21888 34572 21894
rect 34520 21830 34572 21836
rect 34532 21593 34560 21830
rect 34518 21584 34574 21593
rect 34428 21548 34480 21554
rect 34518 21519 34574 21528
rect 34428 21490 34480 21496
rect 34334 20360 34390 20369
rect 34334 20295 34390 20304
rect 34428 19984 34480 19990
rect 34428 19926 34480 19932
rect 34152 19304 34204 19310
rect 34152 19246 34204 19252
rect 34072 18414 34376 18442
rect 34152 18352 34204 18358
rect 34152 18294 34204 18300
rect 33966 18048 34022 18057
rect 33966 17983 34022 17992
rect 33968 17808 34020 17814
rect 33968 17750 34020 17756
rect 33876 16992 33928 16998
rect 33876 16934 33928 16940
rect 33980 16250 34008 17750
rect 34060 17740 34112 17746
rect 34060 17682 34112 17688
rect 33968 16244 34020 16250
rect 33968 16186 34020 16192
rect 33876 16108 33928 16114
rect 33876 16050 33928 16056
rect 33784 15972 33836 15978
rect 33784 15914 33836 15920
rect 33784 15156 33836 15162
rect 33784 15098 33836 15104
rect 33690 14784 33746 14793
rect 33690 14719 33746 14728
rect 33796 14498 33824 15098
rect 33888 14618 33916 16050
rect 34072 15314 34100 17682
rect 34164 17270 34192 18294
rect 34152 17264 34204 17270
rect 34152 17206 34204 17212
rect 34164 16794 34192 17206
rect 34244 17128 34296 17134
rect 34244 17070 34296 17076
rect 34256 16998 34284 17070
rect 34244 16992 34296 16998
rect 34244 16934 34296 16940
rect 34152 16788 34204 16794
rect 34152 16730 34204 16736
rect 34164 16674 34192 16730
rect 34164 16646 34284 16674
rect 34152 16516 34204 16522
rect 34152 16458 34204 16464
rect 34164 16046 34192 16458
rect 34256 16454 34284 16646
rect 34244 16448 34296 16454
rect 34244 16390 34296 16396
rect 34152 16040 34204 16046
rect 34152 15982 34204 15988
rect 34164 15706 34192 15982
rect 34256 15706 34284 16390
rect 34152 15700 34204 15706
rect 34152 15642 34204 15648
rect 34244 15700 34296 15706
rect 34244 15642 34296 15648
rect 34256 15434 34284 15642
rect 34348 15570 34376 18414
rect 34336 15564 34388 15570
rect 34336 15506 34388 15512
rect 34244 15428 34296 15434
rect 34244 15370 34296 15376
rect 34072 15286 34284 15314
rect 34058 15192 34114 15201
rect 34058 15127 34114 15136
rect 33876 14612 33928 14618
rect 33876 14554 33928 14560
rect 33968 14612 34020 14618
rect 33968 14554 34020 14560
rect 33980 14498 34008 14554
rect 33506 14447 33562 14456
rect 33600 14476 33652 14482
rect 33796 14470 34008 14498
rect 33600 14418 33652 14424
rect 33416 14408 33468 14414
rect 34072 14362 34100 15127
rect 34152 14952 34204 14958
rect 34152 14894 34204 14900
rect 34164 14793 34192 14894
rect 34150 14784 34206 14793
rect 34150 14719 34206 14728
rect 34152 14476 34204 14482
rect 34152 14418 34204 14424
rect 33416 14350 33468 14356
rect 33888 14334 34100 14362
rect 33322 14240 33378 14249
rect 33322 14175 33378 14184
rect 33692 13932 33744 13938
rect 33692 13874 33744 13880
rect 33600 13864 33652 13870
rect 33600 13806 33652 13812
rect 33244 13688 33364 13716
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 32956 13456 33008 13462
rect 32956 13398 33008 13404
rect 32864 13320 32916 13326
rect 32864 13262 32916 13268
rect 32968 12900 32996 13398
rect 33336 13258 33364 13688
rect 33612 13410 33640 13806
rect 33520 13382 33640 13410
rect 33324 13252 33376 13258
rect 33324 13194 33376 13200
rect 32876 12872 32996 12900
rect 32770 11928 32826 11937
rect 32680 11892 32732 11898
rect 32770 11863 32826 11872
rect 32680 11834 32732 11840
rect 32784 11694 32812 11863
rect 32772 11688 32824 11694
rect 32772 11630 32824 11636
rect 32680 11212 32732 11218
rect 32680 11154 32732 11160
rect 32496 10260 32548 10266
rect 32496 10202 32548 10208
rect 32312 9580 32364 9586
rect 32312 9522 32364 9528
rect 32404 9580 32456 9586
rect 32404 9522 32456 9528
rect 32220 9512 32272 9518
rect 32220 9454 32272 9460
rect 32036 9104 32088 9110
rect 32036 9046 32088 9052
rect 31668 8424 31720 8430
rect 31668 8366 31720 8372
rect 32232 8362 32260 9454
rect 32324 8906 32352 9522
rect 32692 9489 32720 11154
rect 32678 9480 32734 9489
rect 32678 9415 32734 9424
rect 32312 8900 32364 8906
rect 32312 8842 32364 8848
rect 32220 8356 32272 8362
rect 32220 8298 32272 8304
rect 32232 7886 32260 8298
rect 32692 7954 32720 9415
rect 32784 8294 32812 11630
rect 32876 11218 32904 12872
rect 33324 12776 33376 12782
rect 33324 12718 33376 12724
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 33336 12434 33364 12718
rect 33244 12406 33364 12434
rect 33244 12170 33272 12406
rect 33232 12164 33284 12170
rect 33232 12106 33284 12112
rect 33244 11676 33272 12106
rect 33244 11648 33364 11676
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 32864 11212 32916 11218
rect 32864 11154 32916 11160
rect 33336 11014 33364 11648
rect 33324 11008 33376 11014
rect 33324 10950 33376 10956
rect 33336 10810 33364 10950
rect 33324 10804 33376 10810
rect 33324 10746 33376 10752
rect 33416 10464 33468 10470
rect 33416 10406 33468 10412
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 33428 10130 33456 10406
rect 33416 10124 33468 10130
rect 33416 10066 33468 10072
rect 33324 10056 33376 10062
rect 33324 9998 33376 10004
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 32864 9036 32916 9042
rect 32864 8978 32916 8984
rect 32772 8288 32824 8294
rect 32772 8230 32824 8236
rect 32680 7948 32732 7954
rect 32680 7890 32732 7896
rect 32220 7880 32272 7886
rect 32220 7822 32272 7828
rect 32876 7546 32904 8978
rect 33336 8974 33364 9998
rect 33520 9994 33548 13382
rect 33600 13252 33652 13258
rect 33600 13194 33652 13200
rect 33612 11558 33640 13194
rect 33704 12850 33732 13874
rect 33692 12844 33744 12850
rect 33692 12786 33744 12792
rect 33888 12434 33916 14334
rect 34058 14240 34114 14249
rect 34058 14175 34114 14184
rect 34072 13870 34100 14175
rect 34060 13864 34112 13870
rect 34060 13806 34112 13812
rect 33968 13728 34020 13734
rect 33968 13670 34020 13676
rect 33980 13394 34008 13670
rect 34164 13394 34192 14418
rect 33968 13388 34020 13394
rect 33968 13330 34020 13336
rect 34152 13388 34204 13394
rect 34152 13330 34204 13336
rect 34164 12714 34192 13330
rect 33968 12708 34020 12714
rect 33968 12650 34020 12656
rect 34152 12708 34204 12714
rect 34152 12650 34204 12656
rect 33796 12406 33916 12434
rect 33600 11552 33652 11558
rect 33600 11494 33652 11500
rect 33600 11212 33652 11218
rect 33600 11154 33652 11160
rect 33508 9988 33560 9994
rect 33508 9930 33560 9936
rect 33612 9042 33640 11154
rect 33796 11150 33824 12406
rect 33876 11552 33928 11558
rect 33876 11494 33928 11500
rect 33784 11144 33836 11150
rect 33784 11086 33836 11092
rect 33888 11082 33916 11494
rect 33980 11121 34008 12650
rect 34150 12608 34206 12617
rect 34150 12543 34206 12552
rect 34060 12368 34112 12374
rect 34060 12310 34112 12316
rect 33966 11112 34022 11121
rect 33876 11076 33928 11082
rect 33966 11047 34022 11056
rect 33876 11018 33928 11024
rect 33784 10600 33836 10606
rect 33784 10542 33836 10548
rect 33690 10160 33746 10169
rect 33690 10095 33746 10104
rect 33704 10062 33732 10095
rect 33796 10062 33824 10542
rect 33692 10056 33744 10062
rect 33692 9998 33744 10004
rect 33784 10056 33836 10062
rect 33784 9998 33836 10004
rect 33796 9500 33824 9998
rect 33876 9512 33928 9518
rect 33796 9472 33876 9500
rect 33876 9454 33928 9460
rect 33600 9036 33652 9042
rect 33600 8978 33652 8984
rect 33324 8968 33376 8974
rect 33416 8968 33468 8974
rect 33324 8910 33376 8916
rect 33414 8936 33416 8945
rect 33468 8936 33470 8945
rect 33414 8871 33470 8880
rect 33888 8634 33916 9454
rect 33968 8968 34020 8974
rect 33966 8936 33968 8945
rect 34020 8936 34022 8945
rect 33966 8871 34022 8880
rect 33876 8628 33928 8634
rect 33876 8570 33928 8576
rect 34072 8480 34100 12310
rect 34164 12306 34192 12543
rect 34152 12300 34204 12306
rect 34152 12242 34204 12248
rect 34256 12238 34284 15286
rect 34244 12232 34296 12238
rect 34244 12174 34296 12180
rect 34256 11218 34284 12174
rect 34244 11212 34296 11218
rect 34244 11154 34296 11160
rect 34152 11144 34204 11150
rect 34152 11086 34204 11092
rect 34164 8838 34192 11086
rect 34348 10985 34376 15506
rect 34440 13938 34468 19926
rect 34624 19514 34652 22510
rect 34704 22432 34756 22438
rect 34704 22374 34756 22380
rect 34716 20466 34744 22374
rect 34796 21548 34848 21554
rect 34796 21490 34848 21496
rect 34808 21185 34836 21490
rect 34794 21176 34850 21185
rect 34794 21111 34850 21120
rect 34900 21010 34928 22714
rect 34980 21616 35032 21622
rect 34980 21558 35032 21564
rect 34888 21004 34940 21010
rect 34888 20946 34940 20952
rect 34704 20460 34756 20466
rect 34704 20402 34756 20408
rect 34704 20052 34756 20058
rect 34704 19994 34756 20000
rect 34716 19786 34744 19994
rect 34704 19780 34756 19786
rect 34704 19722 34756 19728
rect 34612 19508 34664 19514
rect 34612 19450 34664 19456
rect 34704 19508 34756 19514
rect 34704 19450 34756 19456
rect 34520 19372 34572 19378
rect 34520 19314 34572 19320
rect 34532 18086 34560 19314
rect 34520 18080 34572 18086
rect 34520 18022 34572 18028
rect 34716 17882 34744 19450
rect 34794 18864 34850 18873
rect 34794 18799 34850 18808
rect 34704 17876 34756 17882
rect 34704 17818 34756 17824
rect 34612 17740 34664 17746
rect 34612 17682 34664 17688
rect 34520 17604 34572 17610
rect 34520 17546 34572 17552
rect 34532 15162 34560 17546
rect 34624 17202 34652 17682
rect 34704 17536 34756 17542
rect 34704 17478 34756 17484
rect 34612 17196 34664 17202
rect 34612 17138 34664 17144
rect 34624 16726 34652 17138
rect 34612 16720 34664 16726
rect 34612 16662 34664 16668
rect 34520 15156 34572 15162
rect 34520 15098 34572 15104
rect 34428 13932 34480 13938
rect 34428 13874 34480 13880
rect 34520 13864 34572 13870
rect 34520 13806 34572 13812
rect 34532 13530 34560 13806
rect 34428 13524 34480 13530
rect 34428 13466 34480 13472
rect 34520 13524 34572 13530
rect 34520 13466 34572 13472
rect 34440 13433 34468 13466
rect 34426 13424 34482 13433
rect 34426 13359 34482 13368
rect 34624 13326 34652 16662
rect 34716 15162 34744 17478
rect 34808 16794 34836 18799
rect 34900 17746 34928 20946
rect 34992 20913 35020 21558
rect 34978 20904 35034 20913
rect 34978 20839 35034 20848
rect 35084 20505 35112 24142
rect 35164 24064 35216 24070
rect 35164 24006 35216 24012
rect 35176 23798 35204 24006
rect 35164 23792 35216 23798
rect 35164 23734 35216 23740
rect 35164 23656 35216 23662
rect 35164 23598 35216 23604
rect 35176 21894 35204 23598
rect 35268 23050 35296 24278
rect 35348 24268 35400 24274
rect 35348 24210 35400 24216
rect 35360 24177 35388 24210
rect 35346 24168 35402 24177
rect 35346 24103 35402 24112
rect 35348 24064 35400 24070
rect 35348 24006 35400 24012
rect 35360 23526 35388 24006
rect 35348 23520 35400 23526
rect 35348 23462 35400 23468
rect 35452 23361 35480 26302
rect 35714 26302 36032 26330
rect 35714 26200 35770 26302
rect 35714 25256 35770 25265
rect 35714 25191 35770 25200
rect 35532 24132 35584 24138
rect 35532 24074 35584 24080
rect 35544 23866 35572 24074
rect 35622 23896 35678 23905
rect 35532 23860 35584 23866
rect 35622 23831 35624 23840
rect 35532 23802 35584 23808
rect 35676 23831 35678 23840
rect 35624 23802 35676 23808
rect 35532 23724 35584 23730
rect 35532 23666 35584 23672
rect 35438 23352 35494 23361
rect 35348 23316 35400 23322
rect 35438 23287 35494 23296
rect 35348 23258 35400 23264
rect 35360 23202 35388 23258
rect 35544 23202 35572 23666
rect 35624 23520 35676 23526
rect 35624 23462 35676 23468
rect 35360 23174 35572 23202
rect 35256 23044 35308 23050
rect 35256 22986 35308 22992
rect 35346 22536 35402 22545
rect 35544 22506 35572 23174
rect 35636 22778 35664 23462
rect 35728 22794 35756 25191
rect 36004 25158 36032 26302
rect 36358 26302 36768 26330
rect 36358 26200 36414 26302
rect 35992 25152 36044 25158
rect 35992 25094 36044 25100
rect 35808 25084 35860 25090
rect 35808 25026 35860 25032
rect 35820 24614 35848 25026
rect 36740 24886 36768 26302
rect 37002 26200 37058 27000
rect 37646 26200 37702 27000
rect 38290 26330 38346 27000
rect 38934 26330 38990 27000
rect 38290 26302 38516 26330
rect 38290 26200 38346 26302
rect 37016 25974 37044 26200
rect 37004 25968 37056 25974
rect 37004 25910 37056 25916
rect 37186 24984 37242 24993
rect 37660 24954 37688 26200
rect 37740 25220 37792 25226
rect 37740 25162 37792 25168
rect 37186 24919 37242 24928
rect 37648 24948 37700 24954
rect 36728 24880 36780 24886
rect 36728 24822 36780 24828
rect 36544 24676 36596 24682
rect 36544 24618 36596 24624
rect 35808 24608 35860 24614
rect 35808 24550 35860 24556
rect 36268 24404 36320 24410
rect 36268 24346 36320 24352
rect 35808 24268 35860 24274
rect 35808 24210 35860 24216
rect 35820 23322 35848 24210
rect 36084 24064 36136 24070
rect 36084 24006 36136 24012
rect 36176 24064 36228 24070
rect 36176 24006 36228 24012
rect 35992 23860 36044 23866
rect 35992 23802 36044 23808
rect 35808 23316 35860 23322
rect 35808 23258 35860 23264
rect 35820 22964 35848 23258
rect 36004 23050 36032 23802
rect 36096 23497 36124 24006
rect 36082 23488 36138 23497
rect 36082 23423 36138 23432
rect 35992 23044 36044 23050
rect 35992 22986 36044 22992
rect 35900 22976 35952 22982
rect 35820 22936 35900 22964
rect 35900 22918 35952 22924
rect 35624 22772 35676 22778
rect 35728 22766 35848 22794
rect 35624 22714 35676 22720
rect 35346 22471 35402 22480
rect 35532 22500 35584 22506
rect 35254 21992 35310 22001
rect 35254 21927 35310 21936
rect 35268 21894 35296 21927
rect 35164 21888 35216 21894
rect 35164 21830 35216 21836
rect 35256 21888 35308 21894
rect 35256 21830 35308 21836
rect 35164 21412 35216 21418
rect 35164 21354 35216 21360
rect 35070 20496 35126 20505
rect 35070 20431 35126 20440
rect 35072 19712 35124 19718
rect 35072 19654 35124 19660
rect 35084 19394 35112 19654
rect 35176 19514 35204 21354
rect 35256 20460 35308 20466
rect 35256 20402 35308 20408
rect 35164 19508 35216 19514
rect 35164 19450 35216 19456
rect 35084 19378 35204 19394
rect 35084 19372 35216 19378
rect 35084 19366 35164 19372
rect 34980 19304 35032 19310
rect 34980 19246 35032 19252
rect 34888 17740 34940 17746
rect 34888 17682 34940 17688
rect 34992 17610 35020 19246
rect 34980 17604 35032 17610
rect 34980 17546 35032 17552
rect 34888 17128 34940 17134
rect 34888 17070 34940 17076
rect 34796 16788 34848 16794
rect 34796 16730 34848 16736
rect 34808 16658 34836 16730
rect 34796 16652 34848 16658
rect 34796 16594 34848 16600
rect 34796 16176 34848 16182
rect 34794 16144 34796 16153
rect 34848 16144 34850 16153
rect 34794 16079 34850 16088
rect 34900 16046 34928 17070
rect 34992 17066 35020 17546
rect 34980 17060 35032 17066
rect 34980 17002 35032 17008
rect 34980 16448 35032 16454
rect 34980 16390 35032 16396
rect 34992 16250 35020 16390
rect 35084 16289 35112 19366
rect 35164 19314 35216 19320
rect 35268 19145 35296 20402
rect 35360 20058 35388 22471
rect 35532 22442 35584 22448
rect 35820 21690 35848 22766
rect 35900 22432 35952 22438
rect 35900 22374 35952 22380
rect 35912 22137 35940 22374
rect 35898 22128 35954 22137
rect 35898 22063 35954 22072
rect 35912 22030 35940 22063
rect 35900 22024 35952 22030
rect 35900 21966 35952 21972
rect 35808 21684 35860 21690
rect 35808 21626 35860 21632
rect 35440 21344 35492 21350
rect 35440 21286 35492 21292
rect 35716 21344 35768 21350
rect 35716 21286 35768 21292
rect 35348 20052 35400 20058
rect 35348 19994 35400 20000
rect 35348 19712 35400 19718
rect 35346 19680 35348 19689
rect 35400 19680 35402 19689
rect 35346 19615 35402 19624
rect 35254 19136 35310 19145
rect 35254 19071 35310 19080
rect 35254 19000 35310 19009
rect 35254 18935 35310 18944
rect 35268 18834 35296 18935
rect 35348 18896 35400 18902
rect 35348 18838 35400 18844
rect 35256 18828 35308 18834
rect 35256 18770 35308 18776
rect 35360 18086 35388 18838
rect 35348 18080 35400 18086
rect 35348 18022 35400 18028
rect 35348 17536 35400 17542
rect 35348 17478 35400 17484
rect 35070 16280 35126 16289
rect 34980 16244 35032 16250
rect 35360 16250 35388 17478
rect 35452 17134 35480 21286
rect 35728 21146 35756 21286
rect 35716 21140 35768 21146
rect 35716 21082 35768 21088
rect 35622 21040 35678 21049
rect 35622 20975 35678 20984
rect 35636 20466 35664 20975
rect 35820 20602 35848 21626
rect 36004 21622 36032 22986
rect 36188 21894 36216 24006
rect 36280 23526 36308 24346
rect 36556 24274 36584 24618
rect 36728 24608 36780 24614
rect 36728 24550 36780 24556
rect 36740 24274 36768 24550
rect 36544 24268 36596 24274
rect 36544 24210 36596 24216
rect 36728 24268 36780 24274
rect 36728 24210 36780 24216
rect 36452 23656 36504 23662
rect 36452 23598 36504 23604
rect 36268 23520 36320 23526
rect 36268 23462 36320 23468
rect 36464 22953 36492 23598
rect 36912 23520 36964 23526
rect 36912 23462 36964 23468
rect 36728 22976 36780 22982
rect 36450 22944 36506 22953
rect 36728 22918 36780 22924
rect 36450 22879 36506 22888
rect 36740 22438 36768 22918
rect 36728 22432 36780 22438
rect 36728 22374 36780 22380
rect 36176 21888 36228 21894
rect 36176 21830 36228 21836
rect 36452 21888 36504 21894
rect 36452 21830 36504 21836
rect 36544 21888 36596 21894
rect 36544 21830 36596 21836
rect 35992 21616 36044 21622
rect 35992 21558 36044 21564
rect 36176 21480 36228 21486
rect 36176 21422 36228 21428
rect 36188 20602 36216 21422
rect 36360 21344 36412 21350
rect 36360 21286 36412 21292
rect 35808 20596 35860 20602
rect 35808 20538 35860 20544
rect 36176 20596 36228 20602
rect 36176 20538 36228 20544
rect 36268 20528 36320 20534
rect 36266 20496 36268 20505
rect 36320 20496 36322 20505
rect 35624 20460 35676 20466
rect 35624 20402 35676 20408
rect 35808 20460 35860 20466
rect 36266 20431 36322 20440
rect 35808 20402 35860 20408
rect 35716 20392 35768 20398
rect 35716 20334 35768 20340
rect 35532 20256 35584 20262
rect 35532 20198 35584 20204
rect 35440 17128 35492 17134
rect 35440 17070 35492 17076
rect 35070 16215 35126 16224
rect 35348 16244 35400 16250
rect 34980 16186 35032 16192
rect 35348 16186 35400 16192
rect 34888 16040 34940 16046
rect 34888 15982 34940 15988
rect 34900 15502 34928 15982
rect 34888 15496 34940 15502
rect 34888 15438 34940 15444
rect 34704 15156 34756 15162
rect 34704 15098 34756 15104
rect 34796 14544 34848 14550
rect 34796 14486 34848 14492
rect 34612 13320 34664 13326
rect 34612 13262 34664 13268
rect 34624 12918 34652 13262
rect 34808 12918 34836 14486
rect 34900 14482 34928 15438
rect 34992 15201 35020 16186
rect 35070 16144 35126 16153
rect 35360 16130 35388 16186
rect 35070 16079 35126 16088
rect 35268 16102 35388 16130
rect 34978 15192 35034 15201
rect 34978 15127 35034 15136
rect 35084 14822 35112 16079
rect 35162 15872 35218 15881
rect 35162 15807 35218 15816
rect 35176 15570 35204 15807
rect 35164 15564 35216 15570
rect 35164 15506 35216 15512
rect 35268 15366 35296 16102
rect 35348 16040 35400 16046
rect 35348 15982 35400 15988
rect 35440 16040 35492 16046
rect 35440 15982 35492 15988
rect 35360 15745 35388 15982
rect 35346 15736 35402 15745
rect 35346 15671 35402 15680
rect 35256 15360 35308 15366
rect 35256 15302 35308 15308
rect 35072 14816 35124 14822
rect 35072 14758 35124 14764
rect 34888 14476 34940 14482
rect 34888 14418 34940 14424
rect 35452 14346 35480 15982
rect 35544 14958 35572 20198
rect 35622 20088 35678 20097
rect 35622 20023 35678 20032
rect 35636 19990 35664 20023
rect 35624 19984 35676 19990
rect 35624 19926 35676 19932
rect 35624 19440 35676 19446
rect 35624 19382 35676 19388
rect 35636 18834 35664 19382
rect 35728 19378 35756 20334
rect 35820 19718 35848 20402
rect 36084 20256 36136 20262
rect 36084 20198 36136 20204
rect 35898 19952 35954 19961
rect 36096 19922 36124 20198
rect 35898 19887 35954 19896
rect 36084 19916 36136 19922
rect 35912 19854 35940 19887
rect 36084 19858 36136 19864
rect 35900 19848 35952 19854
rect 35900 19790 35952 19796
rect 35808 19712 35860 19718
rect 35808 19654 35860 19660
rect 35900 19712 35952 19718
rect 35900 19654 35952 19660
rect 35716 19372 35768 19378
rect 35716 19314 35768 19320
rect 35808 19304 35860 19310
rect 35808 19246 35860 19252
rect 35820 18873 35848 19246
rect 35806 18864 35862 18873
rect 35624 18828 35676 18834
rect 35806 18799 35862 18808
rect 35624 18770 35676 18776
rect 35912 18698 35940 19654
rect 35992 19372 36044 19378
rect 35992 19314 36044 19320
rect 35900 18692 35952 18698
rect 35900 18634 35952 18640
rect 35808 18624 35860 18630
rect 35808 18566 35860 18572
rect 35716 18148 35768 18154
rect 35716 18090 35768 18096
rect 35728 17746 35756 18090
rect 35716 17740 35768 17746
rect 35716 17682 35768 17688
rect 35624 17672 35676 17678
rect 35624 17614 35676 17620
rect 35636 15620 35664 17614
rect 35728 16658 35756 17682
rect 35820 17270 35848 18566
rect 35808 17264 35860 17270
rect 35808 17206 35860 17212
rect 35900 16788 35952 16794
rect 35900 16730 35952 16736
rect 35716 16652 35768 16658
rect 35716 16594 35768 16600
rect 35806 16416 35862 16425
rect 35806 16351 35862 16360
rect 35636 15592 35756 15620
rect 35532 14952 35584 14958
rect 35532 14894 35584 14900
rect 35164 14340 35216 14346
rect 35164 14282 35216 14288
rect 35440 14340 35492 14346
rect 35440 14282 35492 14288
rect 35072 14068 35124 14074
rect 35072 14010 35124 14016
rect 35084 13954 35112 14010
rect 34992 13926 35112 13954
rect 34992 13734 35020 13926
rect 34980 13728 35032 13734
rect 34980 13670 35032 13676
rect 35072 13728 35124 13734
rect 35072 13670 35124 13676
rect 34612 12912 34664 12918
rect 34612 12854 34664 12860
rect 34796 12912 34848 12918
rect 34796 12854 34848 12860
rect 34428 12844 34480 12850
rect 34428 12786 34480 12792
rect 34440 12073 34468 12786
rect 34520 12096 34572 12102
rect 34426 12064 34482 12073
rect 34520 12038 34572 12044
rect 34426 11999 34482 12008
rect 34532 11694 34560 12038
rect 34520 11688 34572 11694
rect 34520 11630 34572 11636
rect 34624 11354 34652 12854
rect 34888 12776 34940 12782
rect 34702 12744 34758 12753
rect 34888 12718 34940 12724
rect 34702 12679 34758 12688
rect 34716 12306 34744 12679
rect 34704 12300 34756 12306
rect 34704 12242 34756 12248
rect 34612 11348 34664 11354
rect 34612 11290 34664 11296
rect 34716 11257 34744 12242
rect 34794 11928 34850 11937
rect 34794 11863 34850 11872
rect 34808 11830 34836 11863
rect 34796 11824 34848 11830
rect 34796 11766 34848 11772
rect 34900 11694 34928 12718
rect 35084 12434 35112 13670
rect 35176 12646 35204 14282
rect 35728 14074 35756 15592
rect 35820 14890 35848 16351
rect 35808 14884 35860 14890
rect 35808 14826 35860 14832
rect 35624 14068 35676 14074
rect 35624 14010 35676 14016
rect 35716 14068 35768 14074
rect 35716 14010 35768 14016
rect 35348 13184 35400 13190
rect 35348 13126 35400 13132
rect 35164 12640 35216 12646
rect 35164 12582 35216 12588
rect 34992 12406 35112 12434
rect 34888 11688 34940 11694
rect 34888 11630 34940 11636
rect 34702 11248 34758 11257
rect 34702 11183 34758 11192
rect 34334 10976 34390 10985
rect 34334 10911 34390 10920
rect 34348 10130 34376 10911
rect 34796 10192 34848 10198
rect 34426 10160 34482 10169
rect 34336 10124 34388 10130
rect 34796 10134 34848 10140
rect 34426 10095 34428 10104
rect 34336 10066 34388 10072
rect 34480 10095 34482 10104
rect 34428 10066 34480 10072
rect 34244 9920 34296 9926
rect 34244 9862 34296 9868
rect 34152 8832 34204 8838
rect 34152 8774 34204 8780
rect 34256 8634 34284 9862
rect 34348 9722 34376 10066
rect 34336 9716 34388 9722
rect 34336 9658 34388 9664
rect 34520 9512 34572 9518
rect 34520 9454 34572 9460
rect 34532 9178 34560 9454
rect 34520 9172 34572 9178
rect 34520 9114 34572 9120
rect 34808 9042 34836 10134
rect 34900 10062 34928 11630
rect 34888 10056 34940 10062
rect 34888 9998 34940 10004
rect 34992 9722 35020 12406
rect 35072 11620 35124 11626
rect 35072 11562 35124 11568
rect 35084 11354 35112 11562
rect 35164 11552 35216 11558
rect 35164 11494 35216 11500
rect 35072 11348 35124 11354
rect 35072 11290 35124 11296
rect 35176 11014 35204 11494
rect 35254 11112 35310 11121
rect 35254 11047 35256 11056
rect 35308 11047 35310 11056
rect 35256 11018 35308 11024
rect 35164 11008 35216 11014
rect 35164 10950 35216 10956
rect 35176 10674 35204 10950
rect 35164 10668 35216 10674
rect 35164 10610 35216 10616
rect 34980 9716 35032 9722
rect 34980 9658 35032 9664
rect 34612 9036 34664 9042
rect 34612 8978 34664 8984
rect 34796 9036 34848 9042
rect 34796 8978 34848 8984
rect 34624 8838 34652 8978
rect 34520 8832 34572 8838
rect 34520 8774 34572 8780
rect 34612 8832 34664 8838
rect 34612 8774 34664 8780
rect 34244 8628 34296 8634
rect 34244 8570 34296 8576
rect 34072 8452 34192 8480
rect 34060 8356 34112 8362
rect 34060 8298 34112 8304
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 32864 7540 32916 7546
rect 32864 7482 32916 7488
rect 34072 7410 34100 8298
rect 31484 7404 31536 7410
rect 31484 7346 31536 7352
rect 34060 7404 34112 7410
rect 34060 7346 34112 7352
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 34164 6390 34192 8452
rect 34428 8288 34480 8294
rect 34428 8230 34480 8236
rect 34440 7886 34468 8230
rect 34428 7880 34480 7886
rect 34428 7822 34480 7828
rect 34152 6384 34204 6390
rect 34152 6326 34204 6332
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 34242 5672 34298 5681
rect 34242 5607 34298 5616
rect 31300 5296 31352 5302
rect 31300 5238 31352 5244
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 31668 4752 31720 4758
rect 31668 4694 31720 4700
rect 30748 3188 30800 3194
rect 30748 3130 30800 3136
rect 30840 2848 30892 2854
rect 30840 2790 30892 2796
rect 30852 2582 30880 2790
rect 31680 2650 31708 4694
rect 34256 4146 34284 5607
rect 34244 4140 34296 4146
rect 34244 4082 34296 4088
rect 33600 4004 33652 4010
rect 33600 3946 33652 3952
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 33612 2650 33640 3946
rect 34532 3602 34560 8774
rect 34624 8634 34652 8774
rect 35360 8634 35388 13126
rect 35440 12708 35492 12714
rect 35440 12650 35492 12656
rect 35452 12170 35480 12650
rect 35636 12434 35664 14010
rect 35716 13456 35768 13462
rect 35716 13398 35768 13404
rect 35728 13326 35756 13398
rect 35716 13320 35768 13326
rect 35716 13262 35768 13268
rect 35728 12986 35756 13262
rect 35808 13252 35860 13258
rect 35808 13194 35860 13200
rect 35820 12986 35848 13194
rect 35716 12980 35768 12986
rect 35716 12922 35768 12928
rect 35808 12980 35860 12986
rect 35808 12922 35860 12928
rect 35544 12406 35664 12434
rect 35440 12164 35492 12170
rect 35440 12106 35492 12112
rect 35544 10742 35572 12406
rect 35728 12306 35756 12922
rect 35716 12300 35768 12306
rect 35716 12242 35768 12248
rect 35624 11552 35676 11558
rect 35624 11494 35676 11500
rect 35636 11150 35664 11494
rect 35624 11144 35676 11150
rect 35624 11086 35676 11092
rect 35532 10736 35584 10742
rect 35532 10678 35584 10684
rect 35716 10668 35768 10674
rect 35716 10610 35768 10616
rect 35440 9920 35492 9926
rect 35440 9862 35492 9868
rect 35452 9722 35480 9862
rect 35440 9716 35492 9722
rect 35440 9658 35492 9664
rect 35452 9042 35480 9658
rect 35728 9654 35756 10610
rect 35808 10600 35860 10606
rect 35808 10542 35860 10548
rect 35716 9648 35768 9654
rect 35716 9590 35768 9596
rect 35532 9580 35584 9586
rect 35532 9522 35584 9528
rect 35544 9489 35572 9522
rect 35530 9480 35586 9489
rect 35530 9415 35586 9424
rect 35532 9376 35584 9382
rect 35532 9318 35584 9324
rect 35544 9042 35572 9318
rect 35440 9036 35492 9042
rect 35440 8978 35492 8984
rect 35532 9036 35584 9042
rect 35532 8978 35584 8984
rect 34612 8628 34664 8634
rect 34612 8570 34664 8576
rect 35348 8628 35400 8634
rect 35348 8570 35400 8576
rect 35256 8492 35308 8498
rect 35256 8434 35308 8440
rect 35268 8090 35296 8434
rect 35820 8430 35848 10542
rect 35912 10538 35940 16730
rect 36004 15026 36032 19314
rect 36096 17746 36124 19858
rect 36372 19394 36400 21286
rect 36464 20330 36492 21830
rect 36452 20324 36504 20330
rect 36452 20266 36504 20272
rect 36452 19712 36504 19718
rect 36452 19654 36504 19660
rect 36464 19514 36492 19654
rect 36452 19508 36504 19514
rect 36452 19450 36504 19456
rect 36372 19366 36492 19394
rect 36084 17740 36136 17746
rect 36084 17682 36136 17688
rect 36268 17332 36320 17338
rect 36268 17274 36320 17280
rect 36176 15496 36228 15502
rect 36176 15438 36228 15444
rect 36084 15360 36136 15366
rect 36084 15302 36136 15308
rect 35992 15020 36044 15026
rect 35992 14962 36044 14968
rect 36096 14278 36124 15302
rect 36188 14346 36216 15438
rect 36280 15162 36308 17274
rect 36360 17196 36412 17202
rect 36360 17138 36412 17144
rect 36372 16794 36400 17138
rect 36360 16788 36412 16794
rect 36360 16730 36412 16736
rect 36360 16108 36412 16114
rect 36464 16096 36492 19366
rect 36556 18970 36584 21830
rect 36636 21480 36688 21486
rect 36636 21422 36688 21428
rect 36648 20806 36676 21422
rect 36740 21010 36768 22374
rect 36924 21622 36952 23462
rect 37096 22636 37148 22642
rect 37096 22578 37148 22584
rect 36912 21616 36964 21622
rect 36912 21558 36964 21564
rect 36820 21344 36872 21350
rect 36820 21286 36872 21292
rect 36728 21004 36780 21010
rect 36728 20946 36780 20952
rect 36636 20800 36688 20806
rect 36636 20742 36688 20748
rect 36648 20233 36676 20742
rect 36740 20398 36768 20946
rect 36832 20466 36860 21286
rect 36924 21146 36952 21558
rect 36912 21140 36964 21146
rect 36912 21082 36964 21088
rect 36820 20460 36872 20466
rect 36820 20402 36872 20408
rect 36728 20392 36780 20398
rect 36728 20334 36780 20340
rect 36634 20224 36690 20233
rect 36634 20159 36690 20168
rect 36648 19174 36676 20159
rect 37004 19304 37056 19310
rect 36910 19272 36966 19281
rect 37004 19246 37056 19252
rect 36910 19207 36966 19216
rect 36924 19174 36952 19207
rect 36636 19168 36688 19174
rect 36636 19110 36688 19116
rect 36912 19168 36964 19174
rect 36912 19110 36964 19116
rect 36544 18964 36596 18970
rect 36544 18906 36596 18912
rect 36636 18692 36688 18698
rect 36636 18634 36688 18640
rect 36648 17746 36676 18634
rect 36912 18624 36964 18630
rect 36912 18566 36964 18572
rect 36924 18465 36952 18566
rect 36910 18456 36966 18465
rect 36910 18391 36966 18400
rect 36910 18320 36966 18329
rect 36910 18255 36966 18264
rect 36924 18222 36952 18255
rect 36820 18216 36872 18222
rect 36820 18158 36872 18164
rect 36912 18216 36964 18222
rect 36912 18158 36964 18164
rect 36636 17740 36688 17746
rect 36636 17682 36688 17688
rect 36726 17504 36782 17513
rect 36726 17439 36782 17448
rect 36544 17128 36596 17134
rect 36544 17070 36596 17076
rect 36412 16068 36492 16096
rect 36360 16050 36412 16056
rect 36360 15972 36412 15978
rect 36360 15914 36412 15920
rect 36268 15156 36320 15162
rect 36268 15098 36320 15104
rect 36268 14816 36320 14822
rect 36268 14758 36320 14764
rect 36176 14340 36228 14346
rect 36176 14282 36228 14288
rect 36084 14272 36136 14278
rect 36084 14214 36136 14220
rect 36096 13802 36124 14214
rect 36084 13796 36136 13802
rect 36084 13738 36136 13744
rect 36188 13734 36216 14282
rect 36176 13728 36228 13734
rect 36176 13670 36228 13676
rect 36188 13462 36216 13670
rect 36176 13456 36228 13462
rect 36176 13398 36228 13404
rect 36188 12306 36216 13398
rect 36176 12300 36228 12306
rect 36176 12242 36228 12248
rect 35992 11552 36044 11558
rect 35992 11494 36044 11500
rect 36004 11082 36032 11494
rect 35992 11076 36044 11082
rect 35992 11018 36044 11024
rect 35900 10532 35952 10538
rect 35900 10474 35952 10480
rect 36280 9625 36308 14758
rect 36372 14006 36400 15914
rect 36556 14550 36584 17070
rect 36634 16688 36690 16697
rect 36634 16623 36690 16632
rect 36648 16454 36676 16623
rect 36740 16590 36768 17439
rect 36728 16584 36780 16590
rect 36728 16526 36780 16532
rect 36636 16448 36688 16454
rect 36636 16390 36688 16396
rect 36740 16182 36768 16526
rect 36728 16176 36780 16182
rect 36728 16118 36780 16124
rect 36832 16017 36860 18158
rect 37016 16794 37044 19246
rect 37108 18193 37136 22578
rect 37200 22094 37228 24919
rect 37648 24890 37700 24896
rect 37752 23746 37780 25162
rect 37830 24440 37886 24449
rect 37830 24375 37886 24384
rect 37844 24206 37872 24375
rect 37924 24268 37976 24274
rect 37924 24210 37976 24216
rect 38384 24268 38436 24274
rect 38384 24210 38436 24216
rect 37832 24200 37884 24206
rect 37936 24177 37964 24210
rect 37832 24142 37884 24148
rect 37922 24168 37978 24177
rect 37922 24103 37978 24112
rect 38292 24132 38344 24138
rect 38292 24074 38344 24080
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 37660 23718 37780 23746
rect 37464 23180 37516 23186
rect 37464 23122 37516 23128
rect 37476 22642 37504 23122
rect 37464 22636 37516 22642
rect 37464 22578 37516 22584
rect 37200 22066 37320 22094
rect 37188 22024 37240 22030
rect 37188 21966 37240 21972
rect 37200 21146 37228 21966
rect 37292 21894 37320 22066
rect 37476 21962 37504 22578
rect 37464 21956 37516 21962
rect 37464 21898 37516 21904
rect 37556 21956 37608 21962
rect 37556 21898 37608 21904
rect 37280 21888 37332 21894
rect 37280 21830 37332 21836
rect 37188 21140 37240 21146
rect 37188 21082 37240 21088
rect 37292 21026 37320 21830
rect 37476 21468 37504 21898
rect 37568 21622 37596 21898
rect 37556 21616 37608 21622
rect 37556 21558 37608 21564
rect 37660 21570 37688 23718
rect 37738 23624 37794 23633
rect 37738 23559 37794 23568
rect 37752 21672 37780 23559
rect 38304 22982 38332 24074
rect 38292 22976 38344 22982
rect 38292 22918 38344 22924
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 38292 22092 38344 22098
rect 38292 22034 38344 22040
rect 38396 22094 38424 24210
rect 38488 22817 38516 26302
rect 38934 26302 39344 26330
rect 38934 26200 38990 26302
rect 38660 25764 38712 25770
rect 38660 25706 38712 25712
rect 38568 23792 38620 23798
rect 38568 23734 38620 23740
rect 38474 22808 38530 22817
rect 38474 22743 38530 22752
rect 38580 22234 38608 23734
rect 38568 22228 38620 22234
rect 38568 22170 38620 22176
rect 38396 22080 38516 22094
rect 38568 22092 38620 22098
rect 38396 22066 38568 22080
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 37752 21644 37872 21672
rect 37660 21542 37780 21570
rect 37648 21480 37700 21486
rect 37476 21440 37648 21468
rect 37648 21422 37700 21428
rect 37372 21344 37424 21350
rect 37372 21286 37424 21292
rect 37556 21344 37608 21350
rect 37556 21286 37608 21292
rect 37200 20998 37320 21026
rect 37200 20466 37228 20998
rect 37280 20800 37332 20806
rect 37384 20754 37412 21286
rect 37332 20748 37412 20754
rect 37280 20742 37412 20748
rect 37292 20726 37412 20742
rect 37292 20602 37320 20726
rect 37280 20596 37332 20602
rect 37280 20538 37332 20544
rect 37188 20460 37240 20466
rect 37188 20402 37240 20408
rect 37278 20360 37334 20369
rect 37278 20295 37334 20304
rect 37292 20058 37320 20295
rect 37188 20052 37240 20058
rect 37188 19994 37240 20000
rect 37280 20052 37332 20058
rect 37280 19994 37332 20000
rect 37200 19378 37228 19994
rect 37372 19916 37424 19922
rect 37372 19858 37424 19864
rect 37464 19916 37516 19922
rect 37464 19858 37516 19864
rect 37280 19780 37332 19786
rect 37280 19722 37332 19728
rect 37188 19372 37240 19378
rect 37188 19314 37240 19320
rect 37188 19236 37240 19242
rect 37188 19178 37240 19184
rect 37200 18766 37228 19178
rect 37188 18760 37240 18766
rect 37188 18702 37240 18708
rect 37292 18408 37320 19722
rect 37200 18380 37320 18408
rect 37094 18184 37150 18193
rect 37094 18119 37150 18128
rect 37200 18086 37228 18380
rect 37384 18358 37412 19858
rect 37476 18358 37504 19858
rect 37568 19009 37596 21286
rect 37660 20942 37688 21422
rect 37752 21418 37780 21542
rect 37740 21412 37792 21418
rect 37740 21354 37792 21360
rect 37648 20936 37700 20942
rect 37648 20878 37700 20884
rect 37660 20380 37688 20878
rect 37740 20392 37792 20398
rect 37660 20352 37740 20380
rect 37740 20334 37792 20340
rect 37648 19712 37700 19718
rect 37648 19654 37700 19660
rect 37554 19000 37610 19009
rect 37554 18935 37610 18944
rect 37556 18896 37608 18902
rect 37556 18838 37608 18844
rect 37372 18352 37424 18358
rect 37372 18294 37424 18300
rect 37464 18352 37516 18358
rect 37464 18294 37516 18300
rect 37280 18284 37332 18290
rect 37280 18226 37332 18232
rect 37188 18080 37240 18086
rect 37188 18022 37240 18028
rect 37188 17672 37240 17678
rect 37188 17614 37240 17620
rect 37096 16992 37148 16998
rect 37096 16934 37148 16940
rect 37004 16788 37056 16794
rect 37004 16730 37056 16736
rect 37004 16584 37056 16590
rect 37004 16526 37056 16532
rect 36912 16516 36964 16522
rect 36912 16458 36964 16464
rect 36924 16425 36952 16458
rect 36910 16416 36966 16425
rect 36910 16351 36966 16360
rect 36912 16244 36964 16250
rect 36912 16186 36964 16192
rect 36818 16008 36874 16017
rect 36818 15943 36874 15952
rect 36924 15366 36952 16186
rect 37016 16046 37044 16526
rect 37004 16040 37056 16046
rect 37004 15982 37056 15988
rect 36912 15360 36964 15366
rect 36912 15302 36964 15308
rect 36636 14952 36688 14958
rect 36636 14894 36688 14900
rect 36544 14544 36596 14550
rect 36544 14486 36596 14492
rect 36360 14000 36412 14006
rect 36360 13942 36412 13948
rect 36556 13938 36584 14486
rect 36544 13932 36596 13938
rect 36544 13874 36596 13880
rect 36452 13320 36504 13326
rect 36452 13262 36504 13268
rect 36464 12918 36492 13262
rect 36452 12912 36504 12918
rect 36452 12854 36504 12860
rect 36452 12776 36504 12782
rect 36452 12718 36504 12724
rect 36464 12481 36492 12718
rect 36450 12472 36506 12481
rect 36648 12442 36676 14894
rect 36728 14000 36780 14006
rect 36728 13942 36780 13948
rect 36740 13394 36768 13942
rect 36728 13388 36780 13394
rect 36728 13330 36780 13336
rect 36450 12407 36452 12416
rect 36504 12407 36506 12416
rect 36636 12436 36688 12442
rect 36452 12378 36504 12384
rect 36924 12434 36952 15302
rect 37108 14822 37136 16934
rect 37200 16590 37228 17614
rect 37188 16584 37240 16590
rect 37188 16526 37240 16532
rect 37200 16114 37228 16526
rect 37188 16108 37240 16114
rect 37188 16050 37240 16056
rect 37200 15638 37228 16050
rect 37188 15632 37240 15638
rect 37188 15574 37240 15580
rect 37096 14816 37148 14822
rect 37096 14758 37148 14764
rect 37292 14074 37320 18226
rect 37384 17814 37412 18294
rect 37464 18080 37516 18086
rect 37464 18022 37516 18028
rect 37372 17808 37424 17814
rect 37372 17750 37424 17756
rect 37476 17678 37504 18022
rect 37464 17672 37516 17678
rect 37464 17614 37516 17620
rect 37372 16992 37424 16998
rect 37372 16934 37424 16940
rect 37384 16726 37412 16934
rect 37372 16720 37424 16726
rect 37372 16662 37424 16668
rect 37384 16250 37412 16662
rect 37464 16584 37516 16590
rect 37464 16526 37516 16532
rect 37372 16244 37424 16250
rect 37372 16186 37424 16192
rect 37476 16046 37504 16526
rect 37464 16040 37516 16046
rect 37464 15982 37516 15988
rect 37476 15502 37504 15982
rect 37464 15496 37516 15502
rect 37464 15438 37516 15444
rect 37476 14958 37504 15438
rect 37464 14952 37516 14958
rect 37464 14894 37516 14900
rect 37372 14884 37424 14890
rect 37372 14826 37424 14832
rect 37188 14068 37240 14074
rect 37188 14010 37240 14016
rect 37280 14068 37332 14074
rect 37280 14010 37332 14016
rect 37200 13954 37228 14010
rect 37278 13968 37334 13977
rect 37200 13926 37278 13954
rect 37278 13903 37334 13912
rect 37096 13864 37148 13870
rect 37096 13806 37148 13812
rect 37108 12442 37136 13806
rect 37188 13728 37240 13734
rect 37188 13670 37240 13676
rect 37200 13258 37228 13670
rect 37188 13252 37240 13258
rect 37188 13194 37240 13200
rect 37096 12436 37148 12442
rect 36924 12406 37044 12434
rect 36636 12378 36688 12384
rect 36728 12300 36780 12306
rect 36728 12242 36780 12248
rect 36740 11830 36768 12242
rect 36728 11824 36780 11830
rect 36728 11766 36780 11772
rect 36740 11082 36768 11766
rect 36728 11076 36780 11082
rect 36728 11018 36780 11024
rect 36452 10668 36504 10674
rect 36452 10610 36504 10616
rect 36266 9616 36322 9625
rect 36266 9551 36322 9560
rect 36280 8838 36308 9551
rect 36464 9178 36492 10610
rect 36636 10600 36688 10606
rect 36636 10542 36688 10548
rect 36544 10464 36596 10470
rect 36544 10406 36596 10412
rect 36556 10266 36584 10406
rect 36648 10266 36676 10542
rect 36544 10260 36596 10266
rect 36544 10202 36596 10208
rect 36636 10260 36688 10266
rect 36636 10202 36688 10208
rect 36740 10146 36768 11018
rect 36556 10118 36768 10146
rect 36556 9994 36584 10118
rect 36544 9988 36596 9994
rect 36544 9930 36596 9936
rect 36556 9654 36584 9930
rect 36544 9648 36596 9654
rect 36544 9590 36596 9596
rect 36452 9172 36504 9178
rect 36452 9114 36504 9120
rect 36556 8906 36584 9590
rect 36728 9376 36780 9382
rect 36728 9318 36780 9324
rect 36544 8900 36596 8906
rect 36544 8842 36596 8848
rect 36268 8832 36320 8838
rect 36268 8774 36320 8780
rect 36740 8498 36768 9318
rect 36820 9172 36872 9178
rect 36820 9114 36872 9120
rect 36832 8974 36860 9114
rect 36820 8968 36872 8974
rect 36820 8910 36872 8916
rect 36728 8492 36780 8498
rect 36728 8434 36780 8440
rect 35808 8424 35860 8430
rect 35808 8366 35860 8372
rect 35256 8084 35308 8090
rect 35256 8026 35308 8032
rect 36912 6248 36964 6254
rect 36912 6190 36964 6196
rect 35808 6180 35860 6186
rect 35808 6122 35860 6128
rect 34520 3596 34572 3602
rect 34520 3538 34572 3544
rect 35820 3534 35848 6122
rect 36924 4826 36952 6190
rect 36912 4820 36964 4826
rect 36912 4762 36964 4768
rect 36924 4554 36952 4762
rect 36912 4548 36964 4554
rect 36912 4490 36964 4496
rect 37016 3670 37044 12406
rect 37096 12378 37148 12384
rect 37188 12368 37240 12374
rect 37188 12310 37240 12316
rect 37280 12368 37332 12374
rect 37280 12310 37332 12316
rect 37200 11234 37228 12310
rect 37292 11898 37320 12310
rect 37280 11892 37332 11898
rect 37280 11834 37332 11840
rect 37384 11830 37412 14826
rect 37476 14482 37504 14894
rect 37568 14793 37596 18838
rect 37660 17338 37688 19654
rect 37752 19378 37780 20334
rect 37740 19372 37792 19378
rect 37740 19314 37792 19320
rect 37844 19310 37872 21644
rect 38304 21350 38332 22034
rect 38396 21486 38424 22066
rect 38488 22052 38568 22066
rect 38568 22034 38620 22040
rect 38568 21616 38620 21622
rect 38474 21584 38530 21593
rect 38568 21558 38620 21564
rect 38474 21519 38530 21528
rect 38384 21480 38436 21486
rect 38384 21422 38436 21428
rect 38292 21344 38344 21350
rect 38292 21286 38344 21292
rect 38488 21185 38516 21519
rect 38474 21176 38530 21185
rect 38474 21111 38530 21120
rect 38580 20874 38608 21558
rect 38568 20868 38620 20874
rect 38568 20810 38620 20816
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 37924 20596 37976 20602
rect 37924 20538 37976 20544
rect 37936 19922 37964 20538
rect 37924 19916 37976 19922
rect 37924 19858 37976 19864
rect 38672 19718 38700 25706
rect 38936 25696 38988 25702
rect 38936 25638 38988 25644
rect 38948 25294 38976 25638
rect 38844 25288 38896 25294
rect 38844 25230 38896 25236
rect 38936 25288 38988 25294
rect 38936 25230 38988 25236
rect 38752 24812 38804 24818
rect 38752 24754 38804 24760
rect 38764 23322 38792 24754
rect 38752 23316 38804 23322
rect 38752 23258 38804 23264
rect 38752 22432 38804 22438
rect 38752 22374 38804 22380
rect 38764 22166 38792 22374
rect 38856 22234 38884 25230
rect 39212 24608 39264 24614
rect 39212 24550 39264 24556
rect 39120 24200 39172 24206
rect 39120 24142 39172 24148
rect 39026 23896 39082 23905
rect 38936 23860 38988 23866
rect 39026 23831 39082 23840
rect 38936 23802 38988 23808
rect 38948 23769 38976 23802
rect 38934 23760 38990 23769
rect 38934 23695 38990 23704
rect 39040 23186 39068 23831
rect 39028 23180 39080 23186
rect 39028 23122 39080 23128
rect 38844 22228 38896 22234
rect 38844 22170 38896 22176
rect 38752 22160 38804 22166
rect 39132 22137 39160 24142
rect 38752 22102 38804 22108
rect 39118 22128 39174 22137
rect 39118 22063 39174 22072
rect 38752 21616 38804 21622
rect 38752 21558 38804 21564
rect 38764 20534 38792 21558
rect 39028 21480 39080 21486
rect 39028 21422 39080 21428
rect 39224 21468 39252 24550
rect 39316 23186 39344 26302
rect 39578 26200 39634 27000
rect 39854 26616 39910 26625
rect 39854 26551 39910 26560
rect 39486 25936 39542 25945
rect 39486 25871 39542 25880
rect 39394 24440 39450 24449
rect 39394 24375 39396 24384
rect 39448 24375 39450 24384
rect 39396 24346 39448 24352
rect 39500 24274 39528 25871
rect 39488 24268 39540 24274
rect 39488 24210 39540 24216
rect 39396 24200 39448 24206
rect 39396 24142 39448 24148
rect 39408 23662 39436 24142
rect 39500 23730 39528 24210
rect 39488 23724 39540 23730
rect 39488 23666 39540 23672
rect 39396 23656 39448 23662
rect 39396 23598 39448 23604
rect 39396 23248 39448 23254
rect 39394 23216 39396 23225
rect 39488 23248 39540 23254
rect 39448 23216 39450 23225
rect 39304 23180 39356 23186
rect 39488 23190 39540 23196
rect 39394 23151 39450 23160
rect 39304 23122 39356 23128
rect 39500 23050 39528 23190
rect 39488 23044 39540 23050
rect 39488 22986 39540 22992
rect 39304 22976 39356 22982
rect 39304 22918 39356 22924
rect 39316 21570 39344 22918
rect 39500 22710 39528 22986
rect 39592 22710 39620 26200
rect 39868 25945 39896 26551
rect 40040 26240 40092 26246
rect 40222 26200 40278 27000
rect 41418 26480 41474 26489
rect 41418 26415 41474 26424
rect 40040 26182 40092 26188
rect 39854 25936 39910 25945
rect 39854 25871 39910 25880
rect 39672 24744 39724 24750
rect 39672 24686 39724 24692
rect 39488 22704 39540 22710
rect 39488 22646 39540 22652
rect 39580 22704 39632 22710
rect 39580 22646 39632 22652
rect 39684 22438 39712 24686
rect 40052 24410 40080 26182
rect 40236 24818 40264 26200
rect 40592 25628 40644 25634
rect 40592 25570 40644 25576
rect 40224 24812 40276 24818
rect 40224 24754 40276 24760
rect 40316 24676 40368 24682
rect 40316 24618 40368 24624
rect 40040 24404 40092 24410
rect 40040 24346 40092 24352
rect 40224 24200 40276 24206
rect 40224 24142 40276 24148
rect 39948 24064 40000 24070
rect 39948 24006 40000 24012
rect 39764 23724 39816 23730
rect 39764 23666 39816 23672
rect 39776 23322 39804 23666
rect 39856 23656 39908 23662
rect 39856 23598 39908 23604
rect 39764 23316 39816 23322
rect 39764 23258 39816 23264
rect 39764 23180 39816 23186
rect 39764 23122 39816 23128
rect 39776 22982 39804 23122
rect 39764 22976 39816 22982
rect 39764 22918 39816 22924
rect 39672 22432 39724 22438
rect 39672 22374 39724 22380
rect 39764 22228 39816 22234
rect 39764 22170 39816 22176
rect 39394 22128 39450 22137
rect 39394 22063 39450 22072
rect 39408 22030 39436 22063
rect 39396 22024 39448 22030
rect 39396 21966 39448 21972
rect 39578 21992 39634 22001
rect 39578 21927 39580 21936
rect 39632 21927 39634 21936
rect 39580 21898 39632 21904
rect 39316 21542 39436 21570
rect 39304 21480 39356 21486
rect 39224 21440 39304 21468
rect 39040 21026 39068 21422
rect 39224 21146 39252 21440
rect 39304 21422 39356 21428
rect 39408 21418 39436 21542
rect 39396 21412 39448 21418
rect 39396 21354 39448 21360
rect 39212 21140 39264 21146
rect 39212 21082 39264 21088
rect 39304 21072 39356 21078
rect 39040 20998 39252 21026
rect 39408 21060 39436 21354
rect 39356 21032 39436 21060
rect 39304 21014 39356 21020
rect 39224 20942 39252 20998
rect 39212 20936 39264 20942
rect 39212 20878 39264 20884
rect 39776 20534 39804 22170
rect 38752 20528 38804 20534
rect 39764 20528 39816 20534
rect 38752 20470 38804 20476
rect 38842 20496 38898 20505
rect 38764 19990 38792 20470
rect 39764 20470 39816 20476
rect 38842 20431 38898 20440
rect 38752 19984 38804 19990
rect 38752 19926 38804 19932
rect 38384 19712 38436 19718
rect 38384 19654 38436 19660
rect 38568 19712 38620 19718
rect 38568 19654 38620 19660
rect 38660 19712 38712 19718
rect 38660 19654 38712 19660
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 37832 19304 37884 19310
rect 37832 19246 37884 19252
rect 37738 19000 37794 19009
rect 37738 18935 37794 18944
rect 37752 18630 37780 18935
rect 38200 18896 38252 18902
rect 38200 18838 38252 18844
rect 37832 18692 37884 18698
rect 37832 18634 37884 18640
rect 37740 18624 37792 18630
rect 37738 18592 37740 18601
rect 37792 18592 37794 18601
rect 37738 18527 37794 18536
rect 37740 18216 37792 18222
rect 37740 18158 37792 18164
rect 37648 17332 37700 17338
rect 37648 17274 37700 17280
rect 37752 17218 37780 18158
rect 37844 18154 37872 18634
rect 38212 18612 38240 18838
rect 38212 18584 38332 18612
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 37922 18320 37978 18329
rect 38304 18306 38332 18584
rect 37922 18255 37924 18264
rect 37976 18255 37978 18264
rect 38212 18278 38332 18306
rect 37924 18226 37976 18232
rect 37832 18148 37884 18154
rect 37832 18090 37884 18096
rect 37936 18057 37964 18226
rect 37922 18048 37978 18057
rect 37922 17983 37978 17992
rect 37832 17536 37884 17542
rect 38212 17524 38240 18278
rect 38396 18222 38424 19654
rect 38476 19440 38528 19446
rect 38476 19382 38528 19388
rect 38488 18986 38516 19382
rect 38580 19122 38608 19654
rect 38764 19446 38792 19926
rect 38856 19854 38884 20431
rect 39028 20324 39080 20330
rect 39028 20266 39080 20272
rect 39040 19922 39068 20266
rect 39764 20256 39816 20262
rect 39764 20198 39816 20204
rect 39028 19916 39080 19922
rect 39028 19858 39080 19864
rect 39580 19916 39632 19922
rect 39580 19858 39632 19864
rect 38844 19848 38896 19854
rect 38844 19790 38896 19796
rect 38752 19440 38804 19446
rect 38752 19382 38804 19388
rect 38764 19258 38792 19382
rect 38764 19230 38884 19258
rect 38752 19168 38804 19174
rect 38580 19094 38700 19122
rect 38752 19110 38804 19116
rect 38488 18958 38608 18986
rect 38474 18864 38530 18873
rect 38474 18799 38476 18808
rect 38528 18799 38530 18808
rect 38476 18770 38528 18776
rect 38476 18624 38528 18630
rect 38474 18592 38476 18601
rect 38528 18592 38530 18601
rect 38474 18527 38530 18536
rect 38476 18420 38528 18426
rect 38476 18362 38528 18368
rect 38292 18216 38344 18222
rect 38292 18158 38344 18164
rect 38384 18216 38436 18222
rect 38384 18158 38436 18164
rect 38304 18057 38332 18158
rect 38290 18048 38346 18057
rect 38290 17983 38346 17992
rect 38212 17496 38332 17524
rect 37832 17478 37884 17484
rect 37660 17190 37780 17218
rect 37660 15978 37688 17190
rect 37740 17060 37792 17066
rect 37740 17002 37792 17008
rect 37752 16590 37780 17002
rect 37740 16584 37792 16590
rect 37740 16526 37792 16532
rect 37844 16153 37872 17478
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 37830 16144 37886 16153
rect 37830 16079 37886 16088
rect 37648 15972 37700 15978
rect 37648 15914 37700 15920
rect 37648 15700 37700 15706
rect 37648 15642 37700 15648
rect 37554 14784 37610 14793
rect 37554 14719 37610 14728
rect 37464 14476 37516 14482
rect 37464 14418 37516 14424
rect 37660 12594 37688 15642
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 38304 14822 38332 17496
rect 38382 17368 38438 17377
rect 38382 17303 38384 17312
rect 38436 17303 38438 17312
rect 38384 17274 38436 17280
rect 38384 17196 38436 17202
rect 38384 17138 38436 17144
rect 38396 15366 38424 17138
rect 38488 17105 38516 18362
rect 38580 17882 38608 18958
rect 38568 17876 38620 17882
rect 38568 17818 38620 17824
rect 38568 17740 38620 17746
rect 38568 17682 38620 17688
rect 38580 17202 38608 17682
rect 38568 17196 38620 17202
rect 38568 17138 38620 17144
rect 38474 17096 38530 17105
rect 38474 17031 38530 17040
rect 38568 16992 38620 16998
rect 38568 16934 38620 16940
rect 38476 16516 38528 16522
rect 38476 16458 38528 16464
rect 38488 15994 38516 16458
rect 38580 16182 38608 16934
rect 38672 16250 38700 19094
rect 38764 17134 38792 19110
rect 38856 18358 38884 19230
rect 39486 19136 39542 19145
rect 39486 19071 39542 19080
rect 39210 18728 39266 18737
rect 39210 18663 39266 18672
rect 39224 18630 39252 18663
rect 39212 18624 39264 18630
rect 39212 18566 39264 18572
rect 38844 18352 38896 18358
rect 38844 18294 38896 18300
rect 38856 18086 38884 18294
rect 39500 18193 39528 19071
rect 39210 18184 39266 18193
rect 39210 18119 39266 18128
rect 39486 18184 39542 18193
rect 39486 18119 39542 18128
rect 38844 18080 38896 18086
rect 38844 18022 38896 18028
rect 39224 17746 39252 18119
rect 39212 17740 39264 17746
rect 39212 17682 39264 17688
rect 38844 17536 38896 17542
rect 38844 17478 38896 17484
rect 38752 17128 38804 17134
rect 38752 17070 38804 17076
rect 38856 16697 38884 17478
rect 38842 16688 38898 16697
rect 38842 16623 38898 16632
rect 38660 16244 38712 16250
rect 38660 16186 38712 16192
rect 38568 16176 38620 16182
rect 38568 16118 38620 16124
rect 38752 16176 38804 16182
rect 38752 16118 38804 16124
rect 38764 15994 38792 16118
rect 38488 15966 38792 15994
rect 39486 16008 39542 16017
rect 38488 15434 38516 15966
rect 39486 15943 39542 15952
rect 38568 15904 38620 15910
rect 38568 15846 38620 15852
rect 38476 15428 38528 15434
rect 38476 15370 38528 15376
rect 38384 15360 38436 15366
rect 38384 15302 38436 15308
rect 38488 15094 38516 15370
rect 38580 15337 38608 15846
rect 39500 15638 39528 15943
rect 39592 15910 39620 19858
rect 39776 19242 39804 20198
rect 39868 20097 39896 23598
rect 39960 21010 39988 24006
rect 40040 23520 40092 23526
rect 40040 23462 40092 23468
rect 40132 23520 40184 23526
rect 40132 23462 40184 23468
rect 40052 23322 40080 23462
rect 40040 23316 40092 23322
rect 40040 23258 40092 23264
rect 40144 23254 40172 23462
rect 40132 23248 40184 23254
rect 40132 23190 40184 23196
rect 40040 22636 40092 22642
rect 40040 22578 40092 22584
rect 40052 22234 40080 22578
rect 40236 22574 40264 24142
rect 40132 22568 40184 22574
rect 40132 22510 40184 22516
rect 40224 22568 40276 22574
rect 40224 22510 40276 22516
rect 40040 22228 40092 22234
rect 40040 22170 40092 22176
rect 40040 21888 40092 21894
rect 40040 21830 40092 21836
rect 40052 21690 40080 21830
rect 40144 21690 40172 22510
rect 40040 21684 40092 21690
rect 40040 21626 40092 21632
rect 40132 21684 40184 21690
rect 40132 21626 40184 21632
rect 40328 21146 40356 24618
rect 40408 23248 40460 23254
rect 40408 23190 40460 23196
rect 40420 22506 40448 23190
rect 40500 23044 40552 23050
rect 40500 22986 40552 22992
rect 40512 22710 40540 22986
rect 40500 22704 40552 22710
rect 40500 22646 40552 22652
rect 40408 22500 40460 22506
rect 40408 22442 40460 22448
rect 40604 21962 40632 25570
rect 41144 24404 41196 24410
rect 41144 24346 41196 24352
rect 41156 24274 41184 24346
rect 41432 24274 41460 26415
rect 42154 26200 42210 27000
rect 42798 26200 42854 27000
rect 43442 26200 43498 27000
rect 43904 26376 43956 26382
rect 43904 26318 43956 26324
rect 41602 25120 41658 25129
rect 41602 25055 41658 25064
rect 41144 24268 41196 24274
rect 41144 24210 41196 24216
rect 41420 24268 41472 24274
rect 41420 24210 41472 24216
rect 41050 24168 41106 24177
rect 41050 24103 41106 24112
rect 41064 23322 41092 24103
rect 41510 23896 41566 23905
rect 41510 23831 41566 23840
rect 41144 23656 41196 23662
rect 41144 23598 41196 23604
rect 41052 23316 41104 23322
rect 41052 23258 41104 23264
rect 40774 23216 40830 23225
rect 40774 23151 40830 23160
rect 40788 23118 40816 23151
rect 40776 23112 40828 23118
rect 40776 23054 40828 23060
rect 41064 22964 41092 23258
rect 41156 23089 41184 23598
rect 41524 23186 41552 23831
rect 41512 23180 41564 23186
rect 41512 23122 41564 23128
rect 41142 23080 41198 23089
rect 41142 23015 41198 23024
rect 41064 22936 41184 22964
rect 41052 22636 41104 22642
rect 41052 22578 41104 22584
rect 41064 22166 41092 22578
rect 40776 22160 40828 22166
rect 40776 22102 40828 22108
rect 41052 22160 41104 22166
rect 41052 22102 41104 22108
rect 40592 21956 40644 21962
rect 40592 21898 40644 21904
rect 40500 21888 40552 21894
rect 40500 21830 40552 21836
rect 40512 21146 40540 21830
rect 40788 21486 40816 22102
rect 40868 22092 40920 22098
rect 40868 22034 40920 22040
rect 40880 22001 40908 22034
rect 40866 21992 40922 22001
rect 40866 21927 40922 21936
rect 40684 21480 40736 21486
rect 40684 21422 40736 21428
rect 40776 21480 40828 21486
rect 40776 21422 40828 21428
rect 40592 21344 40644 21350
rect 40592 21286 40644 21292
rect 40316 21140 40368 21146
rect 40316 21082 40368 21088
rect 40500 21140 40552 21146
rect 40500 21082 40552 21088
rect 40604 21010 40632 21286
rect 39948 21004 40000 21010
rect 39948 20946 40000 20952
rect 40592 21004 40644 21010
rect 40592 20946 40644 20952
rect 40696 20777 40724 21422
rect 40788 20806 40816 21422
rect 40776 20800 40828 20806
rect 40682 20768 40738 20777
rect 40512 20726 40682 20754
rect 40316 20528 40368 20534
rect 40314 20496 40316 20505
rect 40368 20496 40370 20505
rect 40314 20431 40370 20440
rect 39948 20256 40000 20262
rect 39948 20198 40000 20204
rect 39854 20088 39910 20097
rect 39854 20023 39910 20032
rect 39856 19712 39908 19718
rect 39856 19654 39908 19660
rect 39868 19446 39896 19654
rect 39856 19440 39908 19446
rect 39856 19382 39908 19388
rect 39764 19236 39816 19242
rect 39764 19178 39816 19184
rect 39672 19168 39724 19174
rect 39672 19110 39724 19116
rect 39684 18290 39712 19110
rect 39764 18420 39816 18426
rect 39764 18362 39816 18368
rect 39672 18284 39724 18290
rect 39672 18226 39724 18232
rect 39776 17814 39804 18362
rect 39764 17808 39816 17814
rect 39764 17750 39816 17756
rect 39960 17746 39988 20198
rect 40132 19916 40184 19922
rect 40132 19858 40184 19864
rect 40040 19712 40092 19718
rect 40040 19654 40092 19660
rect 40052 18426 40080 19654
rect 40144 18970 40172 19858
rect 40512 19854 40540 20726
rect 40776 20742 40828 20748
rect 40682 20703 40738 20712
rect 40960 20460 41012 20466
rect 40960 20402 41012 20408
rect 40972 20233 41000 20402
rect 41052 20392 41104 20398
rect 41052 20334 41104 20340
rect 40958 20224 41014 20233
rect 40958 20159 41014 20168
rect 40776 19984 40828 19990
rect 40604 19932 40776 19938
rect 40604 19926 40828 19932
rect 40604 19910 40816 19926
rect 40316 19848 40368 19854
rect 40316 19790 40368 19796
rect 40500 19848 40552 19854
rect 40500 19790 40552 19796
rect 40132 18964 40184 18970
rect 40132 18906 40184 18912
rect 40328 18850 40356 19790
rect 40500 19508 40552 19514
rect 40500 19450 40552 19456
rect 40512 19281 40540 19450
rect 40498 19272 40554 19281
rect 40498 19207 40554 19216
rect 40604 18850 40632 19910
rect 40684 19712 40736 19718
rect 40684 19654 40736 19660
rect 40960 19712 41012 19718
rect 40960 19654 41012 19660
rect 40696 19514 40724 19654
rect 40684 19508 40736 19514
rect 40684 19450 40736 19456
rect 40972 19394 41000 19654
rect 40696 19366 41000 19394
rect 40696 19310 40724 19366
rect 40684 19304 40736 19310
rect 40684 19246 40736 19252
rect 41064 18970 41092 20334
rect 41156 20330 41184 22936
rect 41328 22704 41380 22710
rect 41328 22646 41380 22652
rect 41340 20874 41368 22646
rect 41420 22092 41472 22098
rect 41420 22034 41472 22040
rect 41432 21434 41460 22034
rect 41512 21888 41564 21894
rect 41512 21830 41564 21836
rect 41524 21622 41552 21830
rect 41512 21616 41564 21622
rect 41512 21558 41564 21564
rect 41512 21480 41564 21486
rect 41432 21428 41512 21434
rect 41432 21422 41564 21428
rect 41432 21406 41552 21422
rect 41328 20868 41380 20874
rect 41328 20810 41380 20816
rect 41144 20324 41196 20330
rect 41144 20266 41196 20272
rect 41340 19334 41368 20810
rect 41512 20392 41564 20398
rect 41512 20334 41564 20340
rect 41616 20346 41644 25055
rect 42168 24138 42196 26200
rect 43534 25800 43590 25809
rect 43534 25735 43590 25744
rect 42798 25664 42854 25673
rect 42798 25599 42854 25608
rect 42616 25560 42668 25566
rect 42616 25502 42668 25508
rect 42524 25152 42576 25158
rect 42524 25094 42576 25100
rect 42340 25016 42392 25022
rect 42340 24958 42392 24964
rect 42156 24132 42208 24138
rect 42156 24074 42208 24080
rect 41788 24064 41840 24070
rect 41788 24006 41840 24012
rect 41696 23044 41748 23050
rect 41696 22986 41748 22992
rect 41708 22778 41736 22986
rect 41696 22772 41748 22778
rect 41696 22714 41748 22720
rect 41800 22094 41828 24006
rect 41880 23520 41932 23526
rect 41880 23462 41932 23468
rect 41972 23520 42024 23526
rect 41972 23462 42024 23468
rect 41892 22710 41920 23462
rect 41880 22704 41932 22710
rect 41880 22646 41932 22652
rect 41708 22066 41828 22094
rect 41708 21894 41736 22066
rect 41696 21888 41748 21894
rect 41696 21830 41748 21836
rect 41524 19990 41552 20334
rect 41616 20318 41920 20346
rect 41984 20330 42012 23462
rect 42156 22704 42208 22710
rect 42156 22646 42208 22652
rect 42064 21344 42116 21350
rect 42064 21286 42116 21292
rect 42076 20602 42104 21286
rect 42168 20602 42196 22646
rect 42352 22098 42380 24958
rect 42432 24676 42484 24682
rect 42432 24618 42484 24624
rect 42444 24070 42472 24618
rect 42432 24064 42484 24070
rect 42432 24006 42484 24012
rect 42430 23488 42486 23497
rect 42430 23423 42486 23432
rect 42340 22092 42392 22098
rect 42340 22034 42392 22040
rect 42248 21684 42300 21690
rect 42248 21626 42300 21632
rect 42260 21486 42288 21626
rect 42248 21480 42300 21486
rect 42248 21422 42300 21428
rect 42260 20890 42288 21422
rect 42340 21344 42392 21350
rect 42340 21286 42392 21292
rect 42352 21078 42380 21286
rect 42340 21072 42392 21078
rect 42340 21014 42392 21020
rect 42444 21010 42472 23423
rect 42432 21004 42484 21010
rect 42432 20946 42484 20952
rect 42536 20890 42564 25094
rect 42628 22506 42656 25502
rect 42812 24392 42840 25599
rect 43352 25492 43404 25498
rect 43352 25434 43404 25440
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 42812 24364 42932 24392
rect 42798 24304 42854 24313
rect 42798 24239 42854 24248
rect 42812 23730 42840 24239
rect 42800 23724 42852 23730
rect 42800 23666 42852 23672
rect 42904 23662 42932 24364
rect 42892 23656 42944 23662
rect 42892 23598 42944 23604
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 43260 23316 43312 23322
rect 43260 23258 43312 23264
rect 42892 23248 42944 23254
rect 42892 23190 42944 23196
rect 42706 22944 42762 22953
rect 42706 22879 42762 22888
rect 42616 22500 42668 22506
rect 42616 22442 42668 22448
rect 42720 21010 42748 22879
rect 42904 22420 42932 23190
rect 43076 23112 43128 23118
rect 43076 23054 43128 23060
rect 43088 22710 43116 23054
rect 43076 22704 43128 22710
rect 43076 22646 43128 22652
rect 43272 22522 43300 23258
rect 43364 22642 43392 25434
rect 43444 25288 43496 25294
rect 43444 25230 43496 25236
rect 43352 22636 43404 22642
rect 43352 22578 43404 22584
rect 43272 22494 43392 22522
rect 42812 22392 42932 22420
rect 42812 22114 42840 22392
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 42892 22160 42944 22166
rect 42812 22108 42892 22114
rect 42812 22102 42944 22108
rect 42812 22086 42932 22102
rect 42904 21690 42932 22086
rect 43364 22030 43392 22494
rect 43456 22094 43484 25230
rect 43548 23322 43576 25735
rect 43718 25392 43774 25401
rect 43718 25327 43774 25336
rect 43628 24608 43680 24614
rect 43628 24550 43680 24556
rect 43536 23316 43588 23322
rect 43536 23258 43588 23264
rect 43640 23254 43668 24550
rect 43628 23248 43680 23254
rect 43628 23190 43680 23196
rect 43732 23066 43760 25327
rect 43812 24744 43864 24750
rect 43812 24686 43864 24692
rect 43824 23594 43852 24686
rect 43916 23662 43944 26318
rect 44086 26200 44142 27000
rect 44730 26330 44786 27000
rect 44730 26302 45048 26330
rect 44730 26200 44786 26302
rect 43996 24880 44048 24886
rect 43996 24822 44048 24828
rect 43904 23656 43956 23662
rect 43904 23598 43956 23604
rect 43812 23588 43864 23594
rect 43812 23530 43864 23536
rect 43902 23352 43958 23361
rect 43902 23287 43904 23296
rect 43956 23287 43958 23296
rect 43904 23258 43956 23264
rect 43902 23216 43958 23225
rect 43902 23151 43904 23160
rect 43956 23151 43958 23160
rect 43904 23122 43956 23128
rect 43628 23044 43680 23050
rect 43732 23038 43852 23066
rect 43628 22986 43680 22992
rect 43534 22672 43590 22681
rect 43534 22607 43536 22616
rect 43588 22607 43590 22616
rect 43536 22578 43588 22584
rect 43640 22234 43668 22986
rect 43720 22976 43772 22982
rect 43824 22953 43852 23038
rect 44008 22982 44036 24822
rect 44100 23254 44128 26200
rect 44640 26036 44692 26042
rect 44640 25978 44692 25984
rect 44546 25936 44602 25945
rect 44546 25871 44602 25880
rect 44270 25256 44326 25265
rect 44270 25191 44326 25200
rect 44180 24064 44232 24070
rect 44180 24006 44232 24012
rect 44192 23474 44220 24006
rect 44284 23730 44312 25191
rect 44364 25084 44416 25090
rect 44364 25026 44416 25032
rect 44272 23724 44324 23730
rect 44272 23666 44324 23672
rect 44192 23446 44312 23474
rect 44284 23361 44312 23446
rect 44270 23352 44326 23361
rect 44180 23316 44232 23322
rect 44270 23287 44326 23296
rect 44180 23258 44232 23264
rect 44088 23248 44140 23254
rect 44088 23190 44140 23196
rect 44100 23118 44128 23190
rect 44088 23112 44140 23118
rect 44088 23054 44140 23060
rect 43996 22976 44048 22982
rect 43720 22918 43772 22924
rect 43810 22944 43866 22953
rect 43628 22228 43680 22234
rect 43628 22170 43680 22176
rect 43536 22094 43588 22098
rect 43456 22092 43588 22094
rect 43456 22066 43536 22092
rect 43536 22034 43588 22040
rect 43732 22030 43760 22918
rect 43996 22918 44048 22924
rect 44086 22944 44142 22953
rect 43810 22879 43866 22888
rect 44086 22879 44142 22888
rect 43902 22672 43958 22681
rect 43902 22607 43958 22616
rect 43352 22024 43404 22030
rect 43352 21966 43404 21972
rect 43720 22024 43772 22030
rect 43720 21966 43772 21972
rect 42892 21684 42944 21690
rect 42892 21626 42944 21632
rect 43260 21684 43312 21690
rect 43260 21626 43312 21632
rect 43272 21457 43300 21626
rect 43258 21448 43314 21457
rect 43258 21383 43314 21392
rect 42798 21312 42854 21321
rect 42798 21247 42854 21256
rect 42812 21078 42840 21247
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 42800 21072 42852 21078
rect 42800 21014 42852 21020
rect 42708 21004 42760 21010
rect 42708 20946 42760 20952
rect 42892 20936 42944 20942
rect 42260 20862 42472 20890
rect 42536 20884 42892 20890
rect 42536 20878 42944 20884
rect 42536 20862 42932 20878
rect 42984 20868 43036 20874
rect 42338 20768 42394 20777
rect 42338 20703 42394 20712
rect 42064 20596 42116 20602
rect 42064 20538 42116 20544
rect 42156 20596 42208 20602
rect 42156 20538 42208 20544
rect 41788 20256 41840 20262
rect 41788 20198 41840 20204
rect 41512 19984 41564 19990
rect 41512 19926 41564 19932
rect 41156 19306 41368 19334
rect 41052 18964 41104 18970
rect 41052 18906 41104 18912
rect 40328 18822 40632 18850
rect 40040 18420 40092 18426
rect 40040 18362 40092 18368
rect 39948 17740 40000 17746
rect 39948 17682 40000 17688
rect 40316 17604 40368 17610
rect 40316 17546 40368 17552
rect 40224 17536 40276 17542
rect 40224 17478 40276 17484
rect 40236 17377 40264 17478
rect 40222 17368 40278 17377
rect 40222 17303 40278 17312
rect 39854 17096 39910 17105
rect 39854 17031 39910 17040
rect 39672 16448 39724 16454
rect 39672 16390 39724 16396
rect 39580 15904 39632 15910
rect 39684 15881 39712 16390
rect 39764 16108 39816 16114
rect 39764 16050 39816 16056
rect 39776 16017 39804 16050
rect 39762 16008 39818 16017
rect 39868 15978 39896 17031
rect 39762 15943 39818 15952
rect 39856 15972 39908 15978
rect 39856 15914 39908 15920
rect 39580 15846 39632 15852
rect 39670 15872 39726 15881
rect 39670 15807 39726 15816
rect 40130 15736 40186 15745
rect 40130 15671 40186 15680
rect 39488 15632 39540 15638
rect 39488 15574 39540 15580
rect 40040 15360 40092 15366
rect 38566 15328 38622 15337
rect 40040 15302 40092 15308
rect 38566 15263 38622 15272
rect 38476 15088 38528 15094
rect 38476 15030 38528 15036
rect 38200 14816 38252 14822
rect 38200 14758 38252 14764
rect 38292 14816 38344 14822
rect 38292 14758 38344 14764
rect 37740 14612 37792 14618
rect 37740 14554 37792 14560
rect 37752 14074 37780 14554
rect 37832 14476 37884 14482
rect 37832 14418 37884 14424
rect 37740 14068 37792 14074
rect 37740 14010 37792 14016
rect 37740 13932 37792 13938
rect 37844 13920 37872 14418
rect 38212 14260 38240 14758
rect 38488 14414 38516 15030
rect 39856 15020 39908 15026
rect 39856 14962 39908 14968
rect 39868 14793 39896 14962
rect 40052 14958 40080 15302
rect 40144 15162 40172 15671
rect 40132 15156 40184 15162
rect 40132 15098 40184 15104
rect 40236 15042 40264 17303
rect 40328 16590 40356 17546
rect 40316 16584 40368 16590
rect 40316 16526 40368 16532
rect 40316 15428 40368 15434
rect 40316 15370 40368 15376
rect 40144 15014 40264 15042
rect 40328 15026 40356 15370
rect 40316 15020 40368 15026
rect 40040 14952 40092 14958
rect 40040 14894 40092 14900
rect 39948 14884 40000 14890
rect 39948 14826 40000 14832
rect 39854 14784 39910 14793
rect 39854 14719 39910 14728
rect 39856 14544 39908 14550
rect 39486 14512 39542 14521
rect 38936 14476 38988 14482
rect 39856 14486 39908 14492
rect 39486 14447 39542 14456
rect 38936 14418 38988 14424
rect 38476 14408 38528 14414
rect 38476 14350 38528 14356
rect 38212 14232 38332 14260
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 37792 13892 37872 13920
rect 37740 13874 37792 13880
rect 37476 12566 37688 12594
rect 37476 12238 37504 12566
rect 37554 12336 37610 12345
rect 37752 12306 37780 13874
rect 38304 13870 38332 14232
rect 37924 13864 37976 13870
rect 37922 13832 37924 13841
rect 38292 13864 38344 13870
rect 37976 13832 37978 13841
rect 38292 13806 38344 13812
rect 37922 13767 37978 13776
rect 38200 13796 38252 13802
rect 38200 13738 38252 13744
rect 38212 13530 38240 13738
rect 38200 13524 38252 13530
rect 38200 13466 38252 13472
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 38488 12918 38516 14350
rect 38948 14278 38976 14418
rect 39500 14414 39528 14447
rect 39488 14408 39540 14414
rect 39488 14350 39540 14356
rect 38936 14272 38988 14278
rect 38936 14214 38988 14220
rect 39304 14272 39356 14278
rect 39304 14214 39356 14220
rect 38568 13388 38620 13394
rect 38568 13330 38620 13336
rect 38476 12912 38528 12918
rect 38212 12872 38476 12900
rect 38212 12442 38240 12872
rect 38476 12854 38528 12860
rect 38476 12640 38528 12646
rect 38476 12582 38528 12588
rect 38200 12436 38252 12442
rect 38200 12378 38252 12384
rect 37554 12271 37556 12280
rect 37608 12271 37610 12280
rect 37740 12300 37792 12306
rect 37556 12242 37608 12248
rect 37740 12242 37792 12248
rect 38488 12238 38516 12582
rect 38580 12481 38608 13330
rect 38750 13288 38806 13297
rect 38750 13223 38752 13232
rect 38804 13223 38806 13232
rect 38752 13194 38804 13200
rect 38752 12640 38804 12646
rect 38750 12608 38752 12617
rect 38804 12608 38806 12617
rect 38750 12543 38806 12552
rect 38566 12472 38622 12481
rect 38566 12407 38622 12416
rect 38948 12374 38976 14214
rect 39120 14068 39172 14074
rect 39120 14010 39172 14016
rect 39132 13920 39160 14010
rect 39316 14006 39344 14214
rect 39304 14000 39356 14006
rect 39304 13942 39356 13948
rect 39868 13938 39896 14486
rect 39960 14482 39988 14826
rect 39948 14476 40000 14482
rect 39948 14418 40000 14424
rect 39212 13932 39264 13938
rect 39132 13892 39212 13920
rect 39212 13874 39264 13880
rect 39856 13932 39908 13938
rect 39856 13874 39908 13880
rect 39854 13696 39910 13705
rect 39854 13631 39910 13640
rect 40038 13696 40094 13705
rect 40038 13631 40094 13640
rect 39028 13184 39080 13190
rect 39028 13126 39080 13132
rect 39304 13184 39356 13190
rect 39304 13126 39356 13132
rect 39580 13184 39632 13190
rect 39580 13126 39632 13132
rect 39040 12850 39068 13126
rect 39316 12889 39344 13126
rect 39302 12880 39358 12889
rect 39028 12844 39080 12850
rect 39302 12815 39358 12824
rect 39028 12786 39080 12792
rect 39592 12442 39620 13126
rect 39868 12918 39896 13631
rect 39856 12912 39908 12918
rect 39856 12854 39908 12860
rect 40052 12753 40080 13631
rect 40038 12744 40094 12753
rect 40038 12679 40094 12688
rect 39580 12436 39632 12442
rect 40144 12434 40172 15014
rect 40316 14962 40368 14968
rect 40420 14906 40448 18822
rect 41064 18222 41092 18906
rect 41052 18216 41104 18222
rect 41052 18158 41104 18164
rect 41156 18068 41184 19306
rect 41696 18760 41748 18766
rect 41696 18702 41748 18708
rect 41604 18692 41656 18698
rect 41604 18634 41656 18640
rect 41616 18306 41644 18634
rect 41524 18278 41644 18306
rect 41708 18290 41736 18702
rect 41696 18284 41748 18290
rect 41524 18086 41552 18278
rect 41696 18226 41748 18232
rect 41602 18184 41658 18193
rect 41602 18119 41604 18128
rect 41656 18119 41658 18128
rect 41604 18090 41656 18096
rect 41064 18040 41184 18068
rect 41512 18080 41564 18086
rect 41064 17785 41092 18040
rect 41512 18022 41564 18028
rect 41800 17921 41828 20198
rect 41892 18290 41920 20318
rect 41972 20324 42024 20330
rect 41972 20266 42024 20272
rect 41984 19990 42012 20266
rect 41972 19984 42024 19990
rect 41972 19926 42024 19932
rect 42352 19786 42380 20703
rect 42340 19780 42392 19786
rect 42340 19722 42392 19728
rect 42156 19508 42208 19514
rect 42156 19450 42208 19456
rect 41972 19372 42024 19378
rect 41972 19314 42024 19320
rect 41984 18873 42012 19314
rect 42168 19122 42196 19450
rect 42444 19174 42472 20862
rect 42984 20810 43036 20816
rect 42800 20800 42852 20806
rect 42800 20742 42852 20748
rect 42614 20632 42670 20641
rect 42614 20567 42670 20576
rect 42708 20596 42760 20602
rect 42628 20398 42656 20567
rect 42708 20538 42760 20544
rect 42616 20392 42668 20398
rect 42616 20334 42668 20340
rect 42628 20058 42656 20334
rect 42616 20052 42668 20058
rect 42616 19994 42668 20000
rect 42720 19514 42748 20538
rect 42708 19508 42760 19514
rect 42708 19450 42760 19456
rect 42812 19417 42840 20742
rect 42996 20398 43024 20810
rect 43258 20496 43314 20505
rect 43258 20431 43314 20440
rect 42984 20392 43036 20398
rect 42984 20334 43036 20340
rect 43272 20330 43300 20431
rect 43260 20324 43312 20330
rect 43260 20266 43312 20272
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 43364 20058 43392 21966
rect 43444 21888 43496 21894
rect 43444 21830 43496 21836
rect 43352 20052 43404 20058
rect 43352 19994 43404 20000
rect 43456 19854 43484 21830
rect 43916 21554 43944 22607
rect 44100 22574 44128 22879
rect 44088 22568 44140 22574
rect 44088 22510 44140 22516
rect 44192 22094 44220 23258
rect 44272 22772 44324 22778
rect 44272 22714 44324 22720
rect 44100 22066 44220 22094
rect 43904 21548 43956 21554
rect 43904 21490 43956 21496
rect 43720 21344 43772 21350
rect 43720 21286 43772 21292
rect 43732 19990 43760 21286
rect 43812 20936 43864 20942
rect 43812 20878 43864 20884
rect 43824 20602 43852 20878
rect 43812 20596 43864 20602
rect 43812 20538 43864 20544
rect 43916 20534 43944 21490
rect 43904 20528 43956 20534
rect 43904 20470 43956 20476
rect 44100 20466 44128 22066
rect 44284 21622 44312 22714
rect 44376 22642 44404 25026
rect 44456 24948 44508 24954
rect 44456 24890 44508 24896
rect 44364 22636 44416 22642
rect 44364 22578 44416 22584
rect 44362 21720 44418 21729
rect 44362 21655 44418 21664
rect 44272 21616 44324 21622
rect 44272 21558 44324 21564
rect 44376 21350 44404 21655
rect 44364 21344 44416 21350
rect 44364 21286 44416 21292
rect 44272 21140 44324 21146
rect 44272 21082 44324 21088
rect 44284 20806 44312 21082
rect 44468 20942 44496 24890
rect 44560 23118 44588 25871
rect 44652 23168 44680 25978
rect 44914 24712 44970 24721
rect 44914 24647 44970 24656
rect 44732 24336 44784 24342
rect 44732 24278 44784 24284
rect 44824 24336 44876 24342
rect 44824 24278 44876 24284
rect 44744 24070 44772 24278
rect 44732 24064 44784 24070
rect 44732 24006 44784 24012
rect 44744 23866 44772 24006
rect 44732 23860 44784 23866
rect 44732 23802 44784 23808
rect 44836 23322 44864 24278
rect 44824 23316 44876 23322
rect 44824 23258 44876 23264
rect 44652 23140 44772 23168
rect 44548 23112 44600 23118
rect 44548 23054 44600 23060
rect 44640 23044 44692 23050
rect 44640 22986 44692 22992
rect 44548 21956 44600 21962
rect 44548 21898 44600 21904
rect 44560 21729 44588 21898
rect 44546 21720 44602 21729
rect 44546 21655 44602 21664
rect 44548 21548 44600 21554
rect 44548 21490 44600 21496
rect 44456 20936 44508 20942
rect 44456 20878 44508 20884
rect 44272 20800 44324 20806
rect 44272 20742 44324 20748
rect 44468 20602 44496 20878
rect 44456 20596 44508 20602
rect 44456 20538 44508 20544
rect 44088 20460 44140 20466
rect 44088 20402 44140 20408
rect 44560 20369 44588 21490
rect 44546 20360 44602 20369
rect 44546 20295 44602 20304
rect 43720 19984 43772 19990
rect 43720 19926 43772 19932
rect 43444 19848 43496 19854
rect 43444 19790 43496 19796
rect 44652 19786 44680 22986
rect 44744 22574 44772 23140
rect 44824 23044 44876 23050
rect 44824 22986 44876 22992
rect 44732 22568 44784 22574
rect 44836 22545 44864 22986
rect 44732 22510 44784 22516
rect 44822 22536 44878 22545
rect 44822 22471 44878 22480
rect 44824 21616 44876 21622
rect 44824 21558 44876 21564
rect 44732 21548 44784 21554
rect 44732 21490 44784 21496
rect 44744 20602 44772 21490
rect 44836 20602 44864 21558
rect 44928 21146 44956 24647
rect 45020 24070 45048 26302
rect 45100 26308 45152 26314
rect 45100 26250 45152 26256
rect 45008 24064 45060 24070
rect 45008 24006 45060 24012
rect 45112 23798 45140 26250
rect 45374 26200 45430 27000
rect 46018 26330 46074 27000
rect 46662 26330 46718 27000
rect 46018 26302 46336 26330
rect 45926 26208 45982 26217
rect 45284 26172 45336 26178
rect 45284 26114 45336 26120
rect 45192 24200 45244 24206
rect 45192 24142 45244 24148
rect 45100 23792 45152 23798
rect 45100 23734 45152 23740
rect 45112 23662 45140 23734
rect 45100 23656 45152 23662
rect 45100 23598 45152 23604
rect 45100 23316 45152 23322
rect 45100 23258 45152 23264
rect 45008 22568 45060 22574
rect 45008 22510 45060 22516
rect 45020 21554 45048 22510
rect 45008 21548 45060 21554
rect 45008 21490 45060 21496
rect 45008 21344 45060 21350
rect 45008 21286 45060 21292
rect 44916 21140 44968 21146
rect 44916 21082 44968 21088
rect 45020 21049 45048 21286
rect 45006 21040 45062 21049
rect 45006 20975 45062 20984
rect 45112 20942 45140 23258
rect 45204 21434 45232 24142
rect 45296 23322 45324 26114
rect 45388 23746 45416 26200
rect 46018 26200 46074 26302
rect 45926 26143 45982 26152
rect 45836 26104 45888 26110
rect 45836 26046 45888 26052
rect 45466 24984 45522 24993
rect 45466 24919 45522 24928
rect 45480 24274 45508 24919
rect 45652 24812 45704 24818
rect 45652 24754 45704 24760
rect 45468 24268 45520 24274
rect 45468 24210 45520 24216
rect 45388 23730 45600 23746
rect 45388 23724 45612 23730
rect 45388 23718 45560 23724
rect 45560 23666 45612 23672
rect 45560 23588 45612 23594
rect 45560 23530 45612 23536
rect 45284 23316 45336 23322
rect 45284 23258 45336 23264
rect 45572 23186 45600 23530
rect 45560 23180 45612 23186
rect 45560 23122 45612 23128
rect 45664 22234 45692 24754
rect 45848 22642 45876 26046
rect 45836 22636 45888 22642
rect 45836 22578 45888 22584
rect 45560 22228 45612 22234
rect 45560 22170 45612 22176
rect 45652 22228 45704 22234
rect 45652 22170 45704 22176
rect 45284 22024 45336 22030
rect 45284 21966 45336 21972
rect 45296 21690 45324 21966
rect 45468 21956 45520 21962
rect 45468 21898 45520 21904
rect 45480 21729 45508 21898
rect 45572 21842 45600 22170
rect 45664 22030 45692 22170
rect 45652 22024 45704 22030
rect 45652 21966 45704 21972
rect 45744 22024 45796 22030
rect 45744 21966 45796 21972
rect 45756 21865 45784 21966
rect 45742 21856 45798 21865
rect 45572 21814 45692 21842
rect 45466 21720 45522 21729
rect 45284 21684 45336 21690
rect 45466 21655 45522 21664
rect 45560 21684 45612 21690
rect 45284 21626 45336 21632
rect 45560 21626 45612 21632
rect 45572 21593 45600 21626
rect 45558 21584 45614 21593
rect 45558 21519 45614 21528
rect 45204 21406 45324 21434
rect 45192 21344 45244 21350
rect 45192 21286 45244 21292
rect 45100 20936 45152 20942
rect 45100 20878 45152 20884
rect 44732 20596 44784 20602
rect 44732 20538 44784 20544
rect 44824 20596 44876 20602
rect 44824 20538 44876 20544
rect 45204 19961 45232 21286
rect 45190 19952 45246 19961
rect 45190 19887 45246 19896
rect 44640 19780 44692 19786
rect 44640 19722 44692 19728
rect 45296 19718 45324 21406
rect 45560 21412 45612 21418
rect 45664 21400 45692 21814
rect 45742 21791 45798 21800
rect 45834 21584 45890 21593
rect 45940 21554 45968 26143
rect 46020 25968 46072 25974
rect 46020 25910 46072 25916
rect 46032 22166 46060 25910
rect 46308 24274 46336 26302
rect 46662 26302 46888 26330
rect 46662 26200 46718 26302
rect 46572 24744 46624 24750
rect 46572 24686 46624 24692
rect 46296 24268 46348 24274
rect 46296 24210 46348 24216
rect 46386 23760 46442 23769
rect 46204 23724 46256 23730
rect 46386 23695 46442 23704
rect 46204 23666 46256 23672
rect 46112 22568 46164 22574
rect 46112 22510 46164 22516
rect 46020 22160 46072 22166
rect 46020 22102 46072 22108
rect 45834 21519 45836 21528
rect 45888 21519 45890 21528
rect 45928 21548 45980 21554
rect 45836 21490 45888 21496
rect 45928 21490 45980 21496
rect 45612 21372 45692 21400
rect 45560 21354 45612 21360
rect 45572 20398 45600 21354
rect 45744 21344 45796 21350
rect 45744 21286 45796 21292
rect 45756 20913 45784 21286
rect 45848 21146 45876 21490
rect 46032 21146 46060 22102
rect 45836 21140 45888 21146
rect 45836 21082 45888 21088
rect 46020 21140 46072 21146
rect 46020 21082 46072 21088
rect 45742 20904 45798 20913
rect 45742 20839 45798 20848
rect 45560 20392 45612 20398
rect 45560 20334 45612 20340
rect 45284 19712 45336 19718
rect 45284 19654 45336 19660
rect 42798 19408 42854 19417
rect 42798 19343 42854 19352
rect 42432 19168 42484 19174
rect 42168 19094 42288 19122
rect 42432 19110 42484 19116
rect 42154 19000 42210 19009
rect 42154 18935 42156 18944
rect 42208 18935 42210 18944
rect 42156 18906 42208 18912
rect 41970 18864 42026 18873
rect 41970 18799 42026 18808
rect 42168 18426 42196 18906
rect 42260 18902 42288 19094
rect 42248 18896 42300 18902
rect 42248 18838 42300 18844
rect 42340 18828 42392 18834
rect 42340 18770 42392 18776
rect 42156 18420 42208 18426
rect 42156 18362 42208 18368
rect 41880 18284 41932 18290
rect 41880 18226 41932 18232
rect 41786 17912 41842 17921
rect 41786 17847 41842 17856
rect 41892 17814 41920 18226
rect 42352 17882 42380 18770
rect 42444 18601 42472 19110
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 42616 18692 42668 18698
rect 42616 18634 42668 18640
rect 42430 18592 42486 18601
rect 42430 18527 42486 18536
rect 42628 17882 42656 18634
rect 42800 18624 42852 18630
rect 42800 18566 42852 18572
rect 42812 18057 42840 18566
rect 43352 18080 43404 18086
rect 42798 18048 42854 18057
rect 43352 18022 43404 18028
rect 42798 17983 42854 17992
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 42340 17876 42392 17882
rect 42340 17818 42392 17824
rect 42616 17876 42668 17882
rect 42616 17818 42668 17824
rect 41880 17808 41932 17814
rect 41050 17776 41106 17785
rect 41880 17750 41932 17756
rect 41050 17711 41106 17720
rect 40592 17672 40644 17678
rect 40592 17614 40644 17620
rect 40604 16998 40632 17614
rect 42064 17536 42116 17542
rect 42064 17478 42116 17484
rect 41604 17332 41656 17338
rect 41604 17274 41656 17280
rect 41052 17196 41104 17202
rect 41052 17138 41104 17144
rect 40592 16992 40644 16998
rect 40592 16934 40644 16940
rect 40604 16658 40632 16934
rect 41064 16794 41092 17138
rect 41052 16788 41104 16794
rect 41052 16730 41104 16736
rect 40592 16652 40644 16658
rect 40592 16594 40644 16600
rect 41328 16584 41380 16590
rect 40682 16552 40738 16561
rect 41328 16526 41380 16532
rect 40682 16487 40684 16496
rect 40736 16487 40738 16496
rect 40684 16458 40736 16464
rect 41052 16040 41104 16046
rect 41052 15982 41104 15988
rect 41064 15586 41092 15982
rect 41340 15638 41368 16526
rect 41616 16250 41644 17274
rect 41604 16244 41656 16250
rect 41604 16186 41656 16192
rect 41328 15632 41380 15638
rect 41064 15580 41328 15586
rect 41064 15574 41380 15580
rect 41064 15558 41368 15574
rect 40866 15328 40922 15337
rect 40866 15263 40922 15272
rect 39580 12378 39632 12384
rect 40052 12406 40172 12434
rect 40236 14878 40448 14906
rect 38936 12368 38988 12374
rect 38936 12310 38988 12316
rect 37464 12232 37516 12238
rect 37464 12174 37516 12180
rect 38476 12232 38528 12238
rect 38476 12174 38528 12180
rect 38936 12096 38988 12102
rect 38936 12038 38988 12044
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 37372 11824 37424 11830
rect 38948 11801 38976 12038
rect 37372 11766 37424 11772
rect 38934 11792 38990 11801
rect 38384 11756 38436 11762
rect 38934 11727 38990 11736
rect 38384 11698 38436 11704
rect 37372 11620 37424 11626
rect 37372 11562 37424 11568
rect 37384 11286 37412 11562
rect 37372 11280 37424 11286
rect 37200 11206 37320 11234
rect 37372 11222 37424 11228
rect 37292 11150 37320 11206
rect 37280 11144 37332 11150
rect 37280 11086 37332 11092
rect 37740 11076 37792 11082
rect 37740 11018 37792 11024
rect 37752 10985 37780 11018
rect 37738 10976 37794 10985
rect 37738 10911 37794 10920
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 37280 10668 37332 10674
rect 37280 10610 37332 10616
rect 37292 9722 37320 10610
rect 38290 10024 38346 10033
rect 38290 9959 38292 9968
rect 38344 9959 38346 9968
rect 38292 9930 38344 9936
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 37280 9716 37332 9722
rect 37280 9658 37332 9664
rect 38396 9518 38424 11698
rect 39120 11688 39172 11694
rect 39120 11630 39172 11636
rect 39212 11688 39264 11694
rect 39212 11630 39264 11636
rect 39132 11218 39160 11630
rect 39120 11212 39172 11218
rect 39120 11154 39172 11160
rect 39224 11150 39252 11630
rect 40052 11393 40080 12406
rect 40132 12164 40184 12170
rect 40132 12106 40184 12112
rect 40144 11694 40172 12106
rect 40132 11688 40184 11694
rect 40130 11656 40132 11665
rect 40184 11656 40186 11665
rect 40130 11591 40186 11600
rect 40038 11384 40094 11393
rect 40038 11319 40094 11328
rect 40130 11248 40186 11257
rect 40130 11183 40186 11192
rect 39212 11144 39264 11150
rect 39212 11086 39264 11092
rect 40040 11144 40092 11150
rect 40040 11086 40092 11092
rect 39304 11008 39356 11014
rect 39304 10950 39356 10956
rect 39316 10062 39344 10950
rect 39488 10668 39540 10674
rect 39488 10610 39540 10616
rect 39500 10169 39528 10610
rect 40052 10538 40080 11086
rect 40144 11082 40172 11183
rect 40132 11076 40184 11082
rect 40132 11018 40184 11024
rect 40144 10810 40172 11018
rect 40132 10804 40184 10810
rect 40132 10746 40184 10752
rect 40236 10713 40264 14878
rect 40684 14272 40736 14278
rect 40684 14214 40736 14220
rect 40696 13569 40724 14214
rect 40880 13938 40908 15263
rect 40958 13968 41014 13977
rect 40868 13932 40920 13938
rect 40958 13903 40960 13912
rect 40868 13874 40920 13880
rect 41012 13903 41014 13912
rect 40960 13874 41012 13880
rect 40682 13560 40738 13569
rect 40682 13495 40738 13504
rect 40776 12096 40828 12102
rect 40776 12038 40828 12044
rect 40788 11830 40816 12038
rect 40776 11824 40828 11830
rect 40776 11766 40828 11772
rect 40314 11384 40370 11393
rect 40314 11319 40370 11328
rect 40222 10704 40278 10713
rect 40222 10639 40278 10648
rect 40040 10532 40092 10538
rect 40040 10474 40092 10480
rect 39486 10160 39542 10169
rect 39486 10095 39488 10104
rect 39540 10095 39542 10104
rect 39488 10066 39540 10072
rect 39304 10056 39356 10062
rect 39304 9998 39356 10004
rect 40328 9994 40356 11319
rect 40774 11112 40830 11121
rect 40774 11047 40776 11056
rect 40828 11047 40830 11056
rect 40776 11018 40828 11024
rect 40788 10810 40816 11018
rect 40776 10804 40828 10810
rect 40776 10746 40828 10752
rect 40316 9988 40368 9994
rect 40316 9930 40368 9936
rect 38384 9512 38436 9518
rect 38384 9454 38436 9460
rect 40040 9104 40092 9110
rect 40040 9046 40092 9052
rect 37280 8900 37332 8906
rect 37280 8842 37332 8848
rect 37292 5370 37320 8842
rect 39580 8832 39632 8838
rect 39580 8774 39632 8780
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 39592 8566 39620 8774
rect 39580 8560 39632 8566
rect 39580 8502 39632 8508
rect 38660 7744 38712 7750
rect 38660 7686 38712 7692
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37370 7576 37426 7585
rect 37950 7579 38258 7588
rect 37370 7511 37372 7520
rect 37424 7511 37426 7520
rect 37372 7482 37424 7488
rect 38672 7342 38700 7686
rect 38660 7336 38712 7342
rect 38660 7278 38712 7284
rect 37924 7200 37976 7206
rect 37924 7142 37976 7148
rect 37936 6934 37964 7142
rect 37924 6928 37976 6934
rect 37924 6870 37976 6876
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 37648 6112 37700 6118
rect 37648 6054 37700 6060
rect 37660 5914 37688 6054
rect 37648 5908 37700 5914
rect 37648 5850 37700 5856
rect 40052 5710 40080 9046
rect 40592 7812 40644 7818
rect 40592 7754 40644 7760
rect 40604 6798 40632 7754
rect 40592 6792 40644 6798
rect 40592 6734 40644 6740
rect 40040 5704 40092 5710
rect 40040 5646 40092 5652
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 37280 5364 37332 5370
rect 37280 5306 37332 5312
rect 37292 5234 37320 5306
rect 37280 5228 37332 5234
rect 37280 5170 37332 5176
rect 40040 5092 40092 5098
rect 40040 5034 40092 5040
rect 37924 5024 37976 5030
rect 37924 4966 37976 4972
rect 37936 4826 37964 4966
rect 37924 4820 37976 4826
rect 37924 4762 37976 4768
rect 39396 4480 39448 4486
rect 39396 4422 39448 4428
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 39212 4140 39264 4146
rect 39212 4082 39264 4088
rect 39304 4140 39356 4146
rect 39304 4082 39356 4088
rect 37004 3664 37056 3670
rect 37004 3606 37056 3612
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 31668 2644 31720 2650
rect 31668 2586 31720 2592
rect 33600 2644 33652 2650
rect 33600 2586 33652 2592
rect 30840 2576 30892 2582
rect 30840 2518 30892 2524
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 33140 2440 33192 2446
rect 33140 2382 33192 2388
rect 34980 2440 35032 2446
rect 34980 2382 35032 2388
rect 30656 2304 30708 2310
rect 30656 2246 30708 2252
rect 30760 800 30788 2382
rect 33152 1578 33180 2382
rect 32876 1550 33180 1578
rect 32876 800 32904 1550
rect 34992 800 35020 2382
rect 37096 2304 37148 2310
rect 37096 2246 37148 2252
rect 37108 800 37136 2246
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 39224 800 39252 4082
rect 39316 3738 39344 4082
rect 39304 3732 39356 3738
rect 39304 3674 39356 3680
rect 39408 3058 39436 4422
rect 40052 3534 40080 5034
rect 40040 3528 40092 3534
rect 40040 3470 40092 3476
rect 40880 3466 40908 13874
rect 40868 3460 40920 3466
rect 40868 3402 40920 3408
rect 40972 3398 41000 13874
rect 41064 13734 41092 15558
rect 41616 15434 41644 16186
rect 41604 15428 41656 15434
rect 41604 15370 41656 15376
rect 41616 15162 41644 15370
rect 41604 15156 41656 15162
rect 41604 15098 41656 15104
rect 41144 14816 41196 14822
rect 41144 14758 41196 14764
rect 41156 14414 41184 14758
rect 41616 14618 41644 15098
rect 42076 15026 42104 17478
rect 42628 17338 42656 17818
rect 42616 17332 42668 17338
rect 42616 17274 42668 17280
rect 43364 17134 43392 18022
rect 43352 17128 43404 17134
rect 43352 17070 43404 17076
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 42156 16448 42208 16454
rect 42156 16390 42208 16396
rect 42168 15706 42196 16390
rect 42248 16108 42300 16114
rect 42248 16050 42300 16056
rect 42156 15700 42208 15706
rect 42156 15642 42208 15648
rect 42260 15502 42288 16050
rect 42340 15904 42392 15910
rect 42340 15846 42392 15852
rect 42352 15570 42380 15846
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 42340 15564 42392 15570
rect 42340 15506 42392 15512
rect 42248 15496 42300 15502
rect 42248 15438 42300 15444
rect 42064 15020 42116 15026
rect 42064 14962 42116 14968
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 41604 14612 41656 14618
rect 41604 14554 41656 14560
rect 41144 14408 41196 14414
rect 41144 14350 41196 14356
rect 41420 14272 41472 14278
rect 41420 14214 41472 14220
rect 41432 14074 41460 14214
rect 41420 14068 41472 14074
rect 41420 14010 41472 14016
rect 41512 14068 41564 14074
rect 41512 14010 41564 14016
rect 41524 13920 41552 14010
rect 41340 13892 41552 13920
rect 41340 13841 41368 13892
rect 41326 13832 41382 13841
rect 41144 13796 41196 13802
rect 41326 13767 41382 13776
rect 41144 13738 41196 13744
rect 41052 13728 41104 13734
rect 41052 13670 41104 13676
rect 41156 13326 41184 13738
rect 41144 13320 41196 13326
rect 41144 13262 41196 13268
rect 41340 8498 41368 13767
rect 41616 12850 41644 14554
rect 44180 14272 44232 14278
rect 44180 14214 44232 14220
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 41788 13184 41840 13190
rect 41788 13126 41840 13132
rect 41800 12986 41828 13126
rect 41788 12980 41840 12986
rect 41788 12922 41840 12928
rect 44192 12850 44220 14214
rect 45296 13705 45324 19654
rect 46124 17241 46152 22510
rect 46216 20058 46244 23666
rect 46400 20942 46428 23695
rect 46480 22976 46532 22982
rect 46480 22918 46532 22924
rect 46492 22710 46520 22918
rect 46480 22704 46532 22710
rect 46480 22646 46532 22652
rect 46584 21146 46612 24686
rect 46756 24132 46808 24138
rect 46756 24074 46808 24080
rect 46572 21140 46624 21146
rect 46572 21082 46624 21088
rect 46388 20936 46440 20942
rect 46388 20878 46440 20884
rect 46400 20534 46428 20878
rect 46768 20602 46796 24074
rect 46860 23882 46888 26302
rect 47306 26200 47362 27000
rect 47950 26330 48006 27000
rect 47872 26302 48006 26330
rect 47030 25120 47086 25129
rect 47030 25055 47086 25064
rect 46860 23854 46980 23882
rect 46952 23798 46980 23854
rect 46940 23792 46992 23798
rect 46940 23734 46992 23740
rect 46938 23080 46994 23089
rect 46938 23015 46994 23024
rect 46846 22944 46902 22953
rect 46846 22879 46902 22888
rect 46860 22642 46888 22879
rect 46952 22778 46980 23015
rect 46940 22772 46992 22778
rect 46940 22714 46992 22720
rect 46848 22636 46900 22642
rect 46848 22578 46900 22584
rect 46848 22500 46900 22506
rect 46848 22442 46900 22448
rect 46860 21554 46888 22442
rect 46848 21548 46900 21554
rect 46848 21490 46900 21496
rect 47044 20942 47072 25055
rect 47216 24336 47268 24342
rect 47216 24278 47268 24284
rect 47124 24132 47176 24138
rect 47124 24074 47176 24080
rect 47032 20936 47084 20942
rect 47032 20878 47084 20884
rect 46756 20596 46808 20602
rect 46756 20538 46808 20544
rect 46388 20528 46440 20534
rect 46388 20470 46440 20476
rect 47044 20466 47072 20878
rect 47136 20602 47164 24074
rect 47124 20596 47176 20602
rect 47124 20538 47176 20544
rect 47032 20460 47084 20466
rect 47032 20402 47084 20408
rect 46204 20052 46256 20058
rect 46204 19994 46256 20000
rect 47228 19242 47256 24278
rect 47320 23050 47348 26200
rect 47398 24712 47454 24721
rect 47398 24647 47454 24656
rect 47584 24676 47636 24682
rect 47308 23044 47360 23050
rect 47308 22986 47360 22992
rect 47320 22778 47348 22986
rect 47308 22772 47360 22778
rect 47308 22714 47360 22720
rect 47308 22228 47360 22234
rect 47308 22170 47360 22176
rect 47320 22030 47348 22170
rect 47308 22024 47360 22030
rect 47308 21966 47360 21972
rect 47412 21690 47440 24647
rect 47584 24618 47636 24624
rect 47492 23792 47544 23798
rect 47492 23734 47544 23740
rect 47400 21684 47452 21690
rect 47400 21626 47452 21632
rect 47504 20058 47532 23734
rect 47596 23526 47624 24618
rect 47766 24304 47822 24313
rect 47766 24239 47822 24248
rect 47584 23520 47636 23526
rect 47584 23462 47636 23468
rect 47674 23488 47730 23497
rect 47674 23423 47730 23432
rect 47582 23352 47638 23361
rect 47582 23287 47584 23296
rect 47636 23287 47638 23296
rect 47584 23258 47636 23264
rect 47584 21480 47636 21486
rect 47584 21422 47636 21428
rect 47596 21146 47624 21422
rect 47584 21140 47636 21146
rect 47584 21082 47636 21088
rect 47688 20942 47716 23423
rect 47780 23322 47808 24239
rect 47872 23746 47900 26302
rect 47950 26200 48006 26302
rect 48594 26200 48650 27000
rect 49238 26200 49294 27000
rect 48502 26072 48558 26081
rect 48502 26007 48558 26016
rect 48226 25528 48282 25537
rect 48226 25463 48282 25472
rect 47952 24608 48004 24614
rect 47952 24550 48004 24556
rect 47964 24410 47992 24550
rect 47952 24404 48004 24410
rect 47952 24346 48004 24352
rect 48240 24274 48268 25463
rect 48412 25424 48464 25430
rect 48412 25366 48464 25372
rect 48228 24268 48280 24274
rect 48228 24210 48280 24216
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 47872 23730 47992 23746
rect 47872 23724 48004 23730
rect 47872 23718 47952 23724
rect 47768 23316 47820 23322
rect 47768 23258 47820 23264
rect 47780 22642 47808 23258
rect 47768 22636 47820 22642
rect 47768 22578 47820 22584
rect 47872 22094 47900 23718
rect 47952 23666 48004 23672
rect 48424 23202 48452 25366
rect 48516 23322 48544 26007
rect 48504 23316 48556 23322
rect 48504 23258 48556 23264
rect 48424 23174 48544 23202
rect 48320 23112 48372 23118
rect 48318 23080 48320 23089
rect 48372 23080 48374 23089
rect 48374 23038 48452 23066
rect 48318 23015 48374 23024
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 48320 22432 48372 22438
rect 48320 22374 48372 22380
rect 47780 22066 47900 22094
rect 47676 20936 47728 20942
rect 47676 20878 47728 20884
rect 47688 20602 47716 20878
rect 47676 20596 47728 20602
rect 47676 20538 47728 20544
rect 47492 20052 47544 20058
rect 47492 19994 47544 20000
rect 47780 19310 47808 22066
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 48228 21684 48280 21690
rect 48228 21626 48280 21632
rect 48240 20942 48268 21626
rect 48332 21146 48360 22374
rect 48320 21140 48372 21146
rect 48320 21082 48372 21088
rect 48228 20936 48280 20942
rect 48228 20878 48280 20884
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 48320 20256 48372 20262
rect 48320 20198 48372 20204
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 47768 19304 47820 19310
rect 48332 19281 48360 20198
rect 48424 19310 48452 23038
rect 48516 22778 48544 23174
rect 48504 22772 48556 22778
rect 48504 22714 48556 22720
rect 48608 22098 48636 26200
rect 48780 25356 48832 25362
rect 48780 25298 48832 25304
rect 48792 24274 48820 25298
rect 48964 25220 49016 25226
rect 48964 25162 49016 25168
rect 48780 24268 48832 24274
rect 48780 24210 48832 24216
rect 48976 23322 49004 25162
rect 49146 23624 49202 23633
rect 49146 23559 49202 23568
rect 49056 23520 49108 23526
rect 49056 23462 49108 23468
rect 48964 23316 49016 23322
rect 48964 23258 49016 23264
rect 49068 22681 49096 23462
rect 49160 22778 49188 23559
rect 49148 22772 49200 22778
rect 49148 22714 49200 22720
rect 49054 22672 49110 22681
rect 49054 22607 49110 22616
rect 48596 22092 48648 22098
rect 48596 22034 48648 22040
rect 48608 21622 48636 22034
rect 49068 22030 49096 22607
rect 49148 22500 49200 22506
rect 49148 22442 49200 22448
rect 49056 22024 49108 22030
rect 49056 21966 49108 21972
rect 49160 21962 49188 22442
rect 49252 22234 49280 26200
rect 49332 22636 49384 22642
rect 49332 22578 49384 22584
rect 49344 22273 49372 22578
rect 49330 22264 49386 22273
rect 49240 22228 49292 22234
rect 49330 22199 49386 22208
rect 49240 22170 49292 22176
rect 49148 21956 49200 21962
rect 49148 21898 49200 21904
rect 48686 21856 48742 21865
rect 48686 21791 48742 21800
rect 48596 21616 48648 21622
rect 48596 21558 48648 21564
rect 48504 21548 48556 21554
rect 48504 21490 48556 21496
rect 48516 21049 48544 21490
rect 48502 21040 48558 21049
rect 48502 20975 48558 20984
rect 48412 19304 48464 19310
rect 47768 19246 47820 19252
rect 48318 19272 48374 19281
rect 47216 19236 47268 19242
rect 48412 19246 48464 19252
rect 48318 19207 48374 19216
rect 47216 19178 47268 19184
rect 48516 19174 48544 20975
rect 48596 20460 48648 20466
rect 48596 20402 48648 20408
rect 48608 20233 48636 20402
rect 48594 20224 48650 20233
rect 48594 20159 48650 20168
rect 48700 19854 48728 21791
rect 49160 21457 49188 21898
rect 49146 21448 49202 21457
rect 49146 21383 49202 21392
rect 48872 21344 48924 21350
rect 48872 21286 48924 21292
rect 48780 21004 48832 21010
rect 48780 20946 48832 20952
rect 48792 19990 48820 20946
rect 48780 19984 48832 19990
rect 48780 19926 48832 19932
rect 48688 19848 48740 19854
rect 48688 19790 48740 19796
rect 48884 19514 48912 21286
rect 49056 20936 49108 20942
rect 49056 20878 49108 20884
rect 49238 20904 49294 20913
rect 49068 20641 49096 20878
rect 49238 20839 49294 20848
rect 49252 20806 49280 20839
rect 49240 20800 49292 20806
rect 49240 20742 49292 20748
rect 49054 20632 49110 20641
rect 48976 20590 49054 20618
rect 48976 20058 49004 20590
rect 49054 20567 49110 20576
rect 49344 20534 49372 22199
rect 49424 21956 49476 21962
rect 49424 21898 49476 21904
rect 49332 20528 49384 20534
rect 49332 20470 49384 20476
rect 49056 20460 49108 20466
rect 49056 20402 49108 20408
rect 48964 20052 49016 20058
rect 48964 19994 49016 20000
rect 49068 19825 49096 20402
rect 49054 19816 49110 19825
rect 49054 19751 49110 19760
rect 49332 19780 49384 19786
rect 49332 19722 49384 19728
rect 48872 19508 48924 19514
rect 48872 19450 48924 19456
rect 49344 19417 49372 19722
rect 49330 19408 49386 19417
rect 49148 19372 49200 19378
rect 49330 19343 49386 19352
rect 49148 19314 49200 19320
rect 48504 19168 48556 19174
rect 48504 19110 48556 19116
rect 49056 19168 49108 19174
rect 49056 19110 49108 19116
rect 49068 18850 49096 19110
rect 49160 19009 49188 19314
rect 49240 19168 49292 19174
rect 49240 19110 49292 19116
rect 49146 19000 49202 19009
rect 49252 18970 49280 19110
rect 49146 18935 49202 18944
rect 49240 18964 49292 18970
rect 49240 18906 49292 18912
rect 49068 18822 49188 18850
rect 49160 18766 49188 18822
rect 48780 18760 48832 18766
rect 48780 18702 48832 18708
rect 49148 18760 49200 18766
rect 49148 18702 49200 18708
rect 48412 18624 48464 18630
rect 48792 18601 48820 18702
rect 48872 18624 48924 18630
rect 48412 18566 48464 18572
rect 48778 18592 48834 18601
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 48424 18358 48452 18566
rect 48872 18566 48924 18572
rect 48778 18527 48834 18536
rect 48792 18426 48820 18527
rect 48780 18420 48832 18426
rect 48780 18362 48832 18368
rect 48412 18352 48464 18358
rect 48412 18294 48464 18300
rect 48320 18080 48372 18086
rect 48320 18022 48372 18028
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 46110 17232 46166 17241
rect 46110 17167 46166 17176
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 48332 15609 48360 18022
rect 48412 17604 48464 17610
rect 48412 17546 48464 17552
rect 48424 17338 48452 17546
rect 48412 17332 48464 17338
rect 48412 17274 48464 17280
rect 48780 17196 48832 17202
rect 48780 17138 48832 17144
rect 48688 16992 48740 16998
rect 48792 16969 48820 17138
rect 48688 16934 48740 16940
rect 48778 16960 48834 16969
rect 48596 15904 48648 15910
rect 48596 15846 48648 15852
rect 48318 15600 48374 15609
rect 48318 15535 48374 15544
rect 47950 15260 48258 15269
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 48412 15088 48464 15094
rect 48412 15030 48464 15036
rect 48502 15056 48558 15065
rect 48318 14920 48374 14929
rect 48318 14855 48320 14864
rect 48372 14855 48374 14864
rect 48320 14826 48372 14832
rect 45836 14816 45888 14822
rect 45836 14758 45888 14764
rect 45560 14544 45612 14550
rect 45560 14486 45612 14492
rect 45282 13696 45338 13705
rect 45282 13631 45338 13640
rect 45572 13433 45600 14486
rect 45848 13938 45876 14758
rect 48320 14272 48372 14278
rect 48320 14214 48372 14220
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 47860 14068 47912 14074
rect 47860 14010 47912 14016
rect 45836 13932 45888 13938
rect 45836 13874 45888 13880
rect 46572 13864 46624 13870
rect 46572 13806 46624 13812
rect 45558 13424 45614 13433
rect 45558 13359 45614 13368
rect 46584 13326 46612 13806
rect 46572 13320 46624 13326
rect 46572 13262 46624 13268
rect 47872 12850 47900 14010
rect 48332 13954 48360 14214
rect 48424 14074 48452 15030
rect 48502 14991 48558 15000
rect 48516 14074 48544 14991
rect 48608 14550 48636 15846
rect 48596 14544 48648 14550
rect 48596 14486 48648 14492
rect 48412 14068 48464 14074
rect 48412 14010 48464 14016
rect 48504 14068 48556 14074
rect 48504 14010 48556 14016
rect 48240 13938 48360 13954
rect 48228 13932 48360 13938
rect 48280 13926 48360 13932
rect 48228 13874 48280 13880
rect 48240 13705 48268 13874
rect 48226 13696 48282 13705
rect 48226 13631 48282 13640
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 41604 12844 41656 12850
rect 41604 12786 41656 12792
rect 44180 12844 44232 12850
rect 44180 12786 44232 12792
rect 47860 12844 47912 12850
rect 47860 12786 47912 12792
rect 44180 12708 44232 12714
rect 44180 12650 44232 12656
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 41604 12232 41656 12238
rect 41604 12174 41656 12180
rect 41616 11626 41644 12174
rect 41604 11620 41656 11626
rect 41604 11562 41656 11568
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 44192 11286 44220 12650
rect 47952 12640 48004 12646
rect 47952 12582 48004 12588
rect 47964 12238 47992 12582
rect 47952 12232 48004 12238
rect 48700 12209 48728 16934
rect 48778 16895 48834 16904
rect 48792 16794 48820 16895
rect 48780 16788 48832 16794
rect 48780 16730 48832 16736
rect 48884 12434 48912 18566
rect 49056 18284 49108 18290
rect 49056 18226 49108 18232
rect 49068 17785 49096 18226
rect 49160 18193 49188 18702
rect 49146 18184 49202 18193
rect 49146 18119 49202 18128
rect 49054 17776 49110 17785
rect 49054 17711 49110 17720
rect 49056 17672 49108 17678
rect 49056 17614 49108 17620
rect 49238 17640 49294 17649
rect 49068 17377 49096 17614
rect 49238 17575 49294 17584
rect 49252 17542 49280 17575
rect 49148 17536 49200 17542
rect 49148 17478 49200 17484
rect 49240 17536 49292 17542
rect 49240 17478 49292 17484
rect 49054 17368 49110 17377
rect 49054 17303 49110 17312
rect 49160 17184 49188 17478
rect 49240 17196 49292 17202
rect 49160 17156 49240 17184
rect 49240 17138 49292 17144
rect 49148 16584 49200 16590
rect 49252 16561 49280 17138
rect 49148 16526 49200 16532
rect 49238 16552 49294 16561
rect 48964 16176 49016 16182
rect 49160 16153 49188 16526
rect 49238 16487 49294 16496
rect 49240 16448 49292 16454
rect 49240 16390 49292 16396
rect 48964 16118 49016 16124
rect 49146 16144 49202 16153
rect 48976 15706 49004 16118
rect 49056 16108 49108 16114
rect 49146 16079 49202 16088
rect 49056 16050 49108 16056
rect 49068 15745 49096 16050
rect 49054 15736 49110 15745
rect 48964 15700 49016 15706
rect 49054 15671 49110 15680
rect 48964 15642 49016 15648
rect 49252 15473 49280 16390
rect 49332 15496 49384 15502
rect 49238 15464 49294 15473
rect 49332 15438 49384 15444
rect 49238 15399 49294 15408
rect 49344 15337 49372 15438
rect 49330 15328 49386 15337
rect 49330 15263 49386 15272
rect 49436 15178 49464 21898
rect 48792 12406 48912 12434
rect 48976 15150 49464 15178
rect 47952 12174 48004 12180
rect 48686 12200 48742 12209
rect 47216 12164 47268 12170
rect 48686 12135 48742 12144
rect 47216 12106 47268 12112
rect 45928 12096 45980 12102
rect 45928 12038 45980 12044
rect 45940 11762 45968 12038
rect 45928 11756 45980 11762
rect 45928 11698 45980 11704
rect 46664 11620 46716 11626
rect 46664 11562 46716 11568
rect 44180 11280 44232 11286
rect 44180 11222 44232 11228
rect 44180 11076 44232 11082
rect 44180 11018 44232 11024
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 44192 10062 44220 11018
rect 45836 10124 45888 10130
rect 45836 10066 45888 10072
rect 44180 10056 44232 10062
rect 44180 9998 44232 10004
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 42708 8900 42760 8906
rect 42708 8842 42760 8848
rect 41328 8492 41380 8498
rect 41328 8434 41380 8440
rect 41420 8356 41472 8362
rect 41420 8298 41472 8304
rect 41432 6390 41460 8298
rect 41420 6384 41472 6390
rect 41420 6326 41472 6332
rect 42720 6322 42748 8842
rect 44824 8628 44876 8634
rect 44824 8570 44876 8576
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 44836 7478 44864 8570
rect 45848 8498 45876 10066
rect 46676 10062 46704 11562
rect 47124 11348 47176 11354
rect 47124 11290 47176 11296
rect 46940 11076 46992 11082
rect 46940 11018 46992 11024
rect 46952 10674 46980 11018
rect 46940 10668 46992 10674
rect 46940 10610 46992 10616
rect 47032 10600 47084 10606
rect 47032 10542 47084 10548
rect 46940 10192 46992 10198
rect 46940 10134 46992 10140
rect 46664 10056 46716 10062
rect 46664 9998 46716 10004
rect 46756 9988 46808 9994
rect 46756 9930 46808 9936
rect 46768 8498 46796 9930
rect 45836 8492 45888 8498
rect 45836 8434 45888 8440
rect 46756 8492 46808 8498
rect 46756 8434 46808 8440
rect 46848 8424 46900 8430
rect 46848 8366 46900 8372
rect 46860 7993 46888 8366
rect 46846 7984 46902 7993
rect 46846 7919 46902 7928
rect 44824 7472 44876 7478
rect 44824 7414 44876 7420
rect 46952 7410 46980 10134
rect 47044 7886 47072 10542
rect 47136 8974 47164 11290
rect 47228 9586 47256 12106
rect 47950 11996 48258 12005
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 48792 10577 48820 12406
rect 48976 11801 49004 15150
rect 49056 15020 49108 15026
rect 49056 14962 49108 14968
rect 49068 14929 49096 14962
rect 49054 14920 49110 14929
rect 49054 14855 49110 14864
rect 49054 14512 49110 14521
rect 49054 14447 49110 14456
rect 49068 14414 49096 14447
rect 49056 14408 49108 14414
rect 49056 14350 49108 14356
rect 49238 14376 49294 14385
rect 49238 14311 49294 14320
rect 49252 14278 49280 14311
rect 49240 14272 49292 14278
rect 49240 14214 49292 14220
rect 49146 14104 49202 14113
rect 49146 14039 49202 14048
rect 49160 14006 49188 14039
rect 49148 14000 49200 14006
rect 49148 13942 49200 13948
rect 49148 13320 49200 13326
rect 49146 13288 49148 13297
rect 49200 13288 49202 13297
rect 49146 13223 49202 13232
rect 49146 12880 49202 12889
rect 49146 12815 49148 12824
rect 49200 12815 49202 12824
rect 49148 12786 49200 12792
rect 49146 12472 49202 12481
rect 49146 12407 49202 12416
rect 49160 12306 49188 12407
rect 49148 12300 49200 12306
rect 49148 12242 49200 12248
rect 49146 12064 49202 12073
rect 49146 11999 49202 12008
rect 49160 11830 49188 11999
rect 49148 11824 49200 11830
rect 48962 11792 49018 11801
rect 49148 11766 49200 11772
rect 48962 11727 49018 11736
rect 49146 11656 49202 11665
rect 49146 11591 49202 11600
rect 49160 11218 49188 11591
rect 49238 11248 49294 11257
rect 49148 11212 49200 11218
rect 49238 11183 49294 11192
rect 49148 11154 49200 11160
rect 49146 10840 49202 10849
rect 49146 10775 49202 10784
rect 48778 10568 48834 10577
rect 48778 10503 48834 10512
rect 49160 10130 49188 10775
rect 49252 10742 49280 11183
rect 49240 10736 49292 10742
rect 49240 10678 49292 10684
rect 49330 10432 49386 10441
rect 49330 10367 49386 10376
rect 49148 10124 49200 10130
rect 49148 10066 49200 10072
rect 49238 10024 49294 10033
rect 47308 9988 47360 9994
rect 49238 9959 49294 9968
rect 47308 9930 47360 9936
rect 47320 9625 47348 9930
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 47306 9616 47362 9625
rect 47216 9580 47268 9586
rect 47306 9551 47362 9560
rect 47216 9522 47268 9528
rect 49146 9208 49202 9217
rect 49146 9143 49202 9152
rect 47124 8968 47176 8974
rect 47124 8910 47176 8916
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 49160 8566 49188 9143
rect 49252 9042 49280 9959
rect 49344 9654 49372 10367
rect 49332 9648 49384 9654
rect 49332 9590 49384 9596
rect 49240 9036 49292 9042
rect 49240 8978 49292 8984
rect 49238 8800 49294 8809
rect 49238 8735 49294 8744
rect 47676 8560 47728 8566
rect 47676 8502 47728 8508
rect 49148 8560 49200 8566
rect 49148 8502 49200 8508
rect 47584 8356 47636 8362
rect 47584 8298 47636 8304
rect 47032 7880 47084 7886
rect 47032 7822 47084 7828
rect 46940 7404 46992 7410
rect 46940 7346 46992 7352
rect 47032 7336 47084 7342
rect 47032 7278 47084 7284
rect 45744 7200 45796 7206
rect 45744 7142 45796 7148
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 42708 6316 42760 6322
rect 42708 6258 42760 6264
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 45756 5234 45784 7142
rect 46940 6180 46992 6186
rect 46940 6122 46992 6128
rect 45836 5636 45888 5642
rect 45836 5578 45888 5584
rect 45744 5228 45796 5234
rect 45744 5170 45796 5176
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 44456 4480 44508 4486
rect 44456 4422 44508 4428
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 43444 3460 43496 3466
rect 43444 3402 43496 3408
rect 40960 3392 41012 3398
rect 40960 3334 41012 3340
rect 39396 3052 39448 3058
rect 39396 2994 39448 3000
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 41328 2508 41380 2514
rect 41328 2450 41380 2456
rect 41340 800 41368 2450
rect 43456 800 43484 3402
rect 44468 2446 44496 4422
rect 45560 3664 45612 3670
rect 45560 3606 45612 3612
rect 44456 2440 44508 2446
rect 44456 2382 44508 2388
rect 45572 800 45600 3606
rect 45848 3058 45876 5578
rect 46664 4072 46716 4078
rect 46664 4014 46716 4020
rect 45836 3052 45888 3058
rect 45836 2994 45888 3000
rect 46676 1465 46704 4014
rect 46952 3534 46980 6122
rect 47044 4622 47072 7278
rect 47216 7268 47268 7274
rect 47216 7210 47268 7216
rect 47124 6928 47176 6934
rect 47124 6870 47176 6876
rect 47032 4616 47084 4622
rect 47032 4558 47084 4564
rect 47136 4146 47164 6870
rect 47228 5234 47256 7210
rect 47308 5908 47360 5914
rect 47308 5850 47360 5856
rect 47216 5228 47268 5234
rect 47216 5170 47268 5176
rect 47216 4820 47268 4826
rect 47216 4762 47268 4768
rect 47124 4140 47176 4146
rect 47124 4082 47176 4088
rect 46940 3528 46992 3534
rect 46940 3470 46992 3476
rect 46756 2984 46808 2990
rect 46756 2926 46808 2932
rect 46848 2984 46900 2990
rect 46848 2926 46900 2932
rect 46768 1873 46796 2926
rect 46860 2689 46888 2926
rect 46846 2680 46902 2689
rect 46846 2615 46902 2624
rect 47228 2446 47256 4762
rect 47320 3058 47348 5850
rect 47596 5710 47624 8298
rect 47688 6798 47716 8502
rect 49252 7954 49280 8735
rect 49330 8392 49386 8401
rect 49330 8327 49386 8336
rect 49240 7948 49292 7954
rect 49240 7890 49292 7896
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 49146 7576 49202 7585
rect 49146 7511 49202 7520
rect 49160 6866 49188 7511
rect 49344 7478 49372 8327
rect 49332 7472 49384 7478
rect 49332 7414 49384 7420
rect 49330 7168 49386 7177
rect 49330 7103 49386 7112
rect 49148 6860 49200 6866
rect 49148 6802 49200 6808
rect 47676 6792 47728 6798
rect 47676 6734 47728 6740
rect 49238 6760 49294 6769
rect 48872 6724 48924 6730
rect 49238 6695 49294 6704
rect 48872 6666 48924 6672
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 48884 6361 48912 6666
rect 48870 6352 48926 6361
rect 48870 6287 48926 6296
rect 49146 5944 49202 5953
rect 49146 5879 49202 5888
rect 47584 5704 47636 5710
rect 47584 5646 47636 5652
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 49160 5302 49188 5879
rect 49252 5778 49280 6695
rect 49344 6390 49372 7103
rect 49332 6384 49384 6390
rect 49332 6326 49384 6332
rect 49240 5772 49292 5778
rect 49240 5714 49292 5720
rect 49422 5536 49478 5545
rect 49422 5471 49478 5480
rect 49148 5296 49200 5302
rect 49148 5238 49200 5244
rect 48320 5160 48372 5166
rect 48320 5102 48372 5108
rect 49330 5128 49386 5137
rect 48332 4729 48360 5102
rect 49330 5063 49386 5072
rect 48318 4720 48374 4729
rect 48318 4655 48374 4664
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 49146 4312 49202 4321
rect 49146 4247 49202 4256
rect 49160 3602 49188 4247
rect 49344 4146 49372 5063
rect 49436 4690 49464 5471
rect 49424 4684 49476 4690
rect 49424 4626 49476 4632
rect 49332 4140 49384 4146
rect 49332 4082 49384 4088
rect 49238 3904 49294 3913
rect 49238 3839 49294 3848
rect 47676 3596 47728 3602
rect 47676 3538 47728 3544
rect 49148 3596 49200 3602
rect 49148 3538 49200 3544
rect 47308 3052 47360 3058
rect 47308 2994 47360 3000
rect 47216 2440 47268 2446
rect 47216 2382 47268 2388
rect 46754 1864 46810 1873
rect 46754 1799 46810 1808
rect 46662 1456 46718 1465
rect 46662 1391 46718 1400
rect 47688 800 47716 3538
rect 49146 3496 49202 3505
rect 48688 3460 48740 3466
rect 49146 3431 49202 3440
rect 48688 3402 48740 3408
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 48700 3097 48728 3402
rect 48686 3088 48742 3097
rect 48686 3023 48742 3032
rect 49160 2514 49188 3431
rect 49252 3126 49280 3839
rect 49792 3392 49844 3398
rect 49792 3334 49844 3340
rect 49240 3120 49292 3126
rect 49240 3062 49292 3068
rect 49148 2508 49200 2514
rect 49148 2450 49200 2456
rect 48504 2372 48556 2378
rect 48504 2314 48556 2320
rect 48516 2281 48544 2314
rect 48502 2272 48558 2281
rect 47950 2204 48258 2213
rect 48502 2207 48558 2216
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 49804 800 49832 3334
rect 18156 734 18368 762
rect 20166 0 20222 800
rect 22282 0 22338 800
rect 24398 0 24454 800
rect 26514 0 26570 800
rect 28630 0 28686 800
rect 30746 0 30802 800
rect 32862 0 32918 800
rect 34978 0 35034 800
rect 37094 0 37150 800
rect 39210 0 39266 800
rect 41326 0 41382 800
rect 43442 0 43498 800
rect 45558 0 45614 800
rect 47674 0 47730 800
rect 49790 0 49846 800
<< via2 >>
rect 2778 24404 2834 24440
rect 2778 24384 2780 24404
rect 2780 24384 2832 24404
rect 2832 24384 2834 24404
rect 1306 20712 1362 20768
rect 1398 19896 1454 19952
rect 1766 19896 1822 19952
rect 1858 19760 1914 19816
rect 3054 25608 3110 25664
rect 3422 24812 3478 24848
rect 3422 24792 3424 24812
rect 3424 24792 3476 24812
rect 3476 24792 3478 24812
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 3606 25200 3662 25256
rect 3514 23976 3570 24032
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 3146 22772 3202 22808
rect 3146 22752 3148 22772
rect 3148 22752 3200 22772
rect 3200 22752 3202 22772
rect 2686 21528 2742 21584
rect 2778 21120 2834 21176
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2686 19488 2742 19544
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2778 18808 2834 18864
rect 2962 19216 3018 19272
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2870 18264 2926 18320
rect 2686 17856 2742 17912
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 3422 23568 3478 23624
rect 3422 23160 3478 23216
rect 3882 24792 3938 24848
rect 3974 22208 4030 22264
rect 3790 21936 3846 21992
rect 3882 20340 3884 20360
rect 3884 20340 3936 20360
rect 3936 20340 3938 20360
rect 3882 20304 3938 20340
rect 4158 22516 4160 22536
rect 4160 22516 4212 22536
rect 4212 22516 4214 22536
rect 4158 22480 4214 22516
rect 4158 22072 4214 22128
rect 2778 17448 2834 17504
rect 1214 17040 1270 17096
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 1306 16632 1362 16688
rect 1306 16224 1362 16280
rect 1306 15816 1362 15872
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 4710 18284 4766 18320
rect 4710 18264 4712 18284
rect 4712 18264 4764 18284
rect 4764 18264 4766 18284
rect 4802 16532 4804 16552
rect 4804 16532 4856 16552
rect 4856 16532 4858 16552
rect 4802 16496 4858 16532
rect 1306 15408 1362 15464
rect 1306 15000 1362 15056
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 1306 14592 1362 14648
rect 938 14184 994 14240
rect 2778 13776 2834 13832
rect 1766 13368 1822 13424
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 3514 13232 3570 13288
rect 1214 12960 1270 13016
rect 1306 12552 1362 12608
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 1214 12144 1270 12200
rect 1306 11736 1362 11792
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 1306 11328 1362 11384
rect 1766 11056 1822 11112
rect 1582 10920 1638 10976
rect 1306 10512 1362 10568
rect 1214 10104 1270 10160
rect 2502 10512 2558 10568
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 1306 9716 1362 9752
rect 1306 9696 1308 9716
rect 1308 9696 1360 9716
rect 1360 9696 1362 9716
rect 1858 9460 1860 9480
rect 1860 9460 1912 9480
rect 1912 9460 1914 9480
rect 1858 9424 1914 9460
rect 1306 9288 1362 9344
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 1306 8900 1362 8936
rect 1306 8880 1308 8900
rect 1308 8880 1360 8900
rect 1360 8880 1362 8900
rect 1214 8472 1270 8528
rect 1398 8084 1454 8120
rect 1398 8064 1400 8084
rect 1400 8064 1452 8084
rect 1452 8064 1454 8084
rect 1306 7656 1362 7712
rect 1306 7248 1362 7304
rect 1214 6840 1270 6896
rect 2502 8880 2558 8936
rect 5446 21412 5502 21448
rect 5446 21392 5448 21412
rect 5448 21392 5500 21412
rect 5500 21392 5502 21412
rect 6090 18808 6146 18864
rect 6826 19352 6882 19408
rect 6642 19116 6644 19136
rect 6644 19116 6696 19136
rect 6696 19116 6698 19136
rect 6642 19080 6698 19116
rect 6550 18944 6606 19000
rect 7378 24248 7434 24304
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7930 21972 7932 21992
rect 7932 21972 7984 21992
rect 7984 21972 7986 21992
rect 7930 21936 7986 21972
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7286 18264 7342 18320
rect 7838 21428 7840 21448
rect 7840 21428 7892 21448
rect 7892 21428 7894 21448
rect 7838 21392 7894 21428
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7838 20440 7894 20496
rect 9402 23180 9458 23216
rect 9402 23160 9404 23180
rect 9404 23160 9456 23180
rect 9456 23160 9458 23180
rect 9218 23060 9220 23080
rect 9220 23060 9272 23080
rect 9272 23060 9274 23080
rect 9218 23024 9274 23060
rect 9034 21528 9090 21584
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 8574 17720 8630 17776
rect 10322 21800 10378 21856
rect 9218 18672 9274 18728
rect 9126 18128 9182 18184
rect 9678 18828 9734 18864
rect 9678 18808 9680 18828
rect 9680 18808 9732 18828
rect 9732 18808 9734 18828
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 9402 17040 9458 17096
rect 9310 16360 9366 16416
rect 10046 19216 10102 19272
rect 10138 19080 10194 19136
rect 10138 17584 10194 17640
rect 10690 21664 10746 21720
rect 10230 17448 10286 17504
rect 9862 16224 9918 16280
rect 9402 15428 9458 15464
rect 9402 15408 9404 15428
rect 9404 15408 9456 15428
rect 9456 15408 9458 15428
rect 9862 14068 9918 14104
rect 9862 14048 9864 14068
rect 9864 14048 9916 14068
rect 9916 14048 9918 14068
rect 10138 16652 10194 16688
rect 10138 16632 10140 16652
rect 10140 16632 10192 16652
rect 10192 16632 10194 16652
rect 10598 18944 10654 19000
rect 10322 13912 10378 13968
rect 10230 13776 10286 13832
rect 9954 13640 10010 13696
rect 9954 13252 10010 13288
rect 9954 13232 9956 13252
rect 9956 13232 10008 13252
rect 10008 13232 10010 13252
rect 10322 13096 10378 13152
rect 9218 12688 9274 12744
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 1306 6432 1362 6488
rect 1306 6024 1362 6080
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 1306 5652 1308 5672
rect 1308 5652 1360 5672
rect 1360 5652 1362 5672
rect 1306 5616 1362 5652
rect 2778 5208 2834 5264
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 1306 4820 1362 4856
rect 1306 4800 1308 4820
rect 1308 4800 1360 4820
rect 1360 4800 1362 4820
rect 1306 4392 1362 4448
rect 1398 3984 1454 4040
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 1306 3576 1362 3632
rect 1306 3188 1362 3224
rect 1306 3168 1308 3188
rect 1308 3168 1360 3188
rect 1360 3168 1362 3188
rect 1306 2760 1362 2816
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 1306 2388 1308 2408
rect 1308 2388 1360 2408
rect 1360 2388 1362 2408
rect 1306 2352 1362 2388
rect 1214 1944 1270 2000
rect 1306 1536 1362 1592
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 10598 17312 10654 17368
rect 10598 16224 10654 16280
rect 10598 15816 10654 15872
rect 11518 22752 11574 22808
rect 11702 22616 11758 22672
rect 11518 22208 11574 22264
rect 11150 21428 11152 21448
rect 11152 21428 11204 21448
rect 11204 21428 11206 21448
rect 11150 21392 11206 21428
rect 11794 22516 11796 22536
rect 11796 22516 11848 22536
rect 11848 22516 11850 22536
rect 11794 22480 11850 22516
rect 11978 24656 12034 24712
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12070 23724 12126 23760
rect 12070 23704 12072 23724
rect 12072 23704 12124 23724
rect 12124 23704 12126 23724
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 11702 20476 11704 20496
rect 11704 20476 11756 20496
rect 11756 20476 11758 20496
rect 11702 20440 11758 20476
rect 11058 16088 11114 16144
rect 11794 19372 11850 19408
rect 11794 19352 11796 19372
rect 11796 19352 11848 19372
rect 11848 19352 11850 19372
rect 10966 14864 11022 14920
rect 10690 14184 10746 14240
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 8850 5072 8906 5128
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12070 20304 12126 20360
rect 12714 20712 12770 20768
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12162 17196 12218 17232
rect 12162 17176 12164 17196
rect 12164 17176 12216 17196
rect 12216 17176 12218 17196
rect 12070 15852 12072 15872
rect 12072 15852 12124 15872
rect 12124 15852 12126 15872
rect 12070 15816 12126 15852
rect 11978 15136 12034 15192
rect 12070 15000 12126 15056
rect 13634 19080 13690 19136
rect 14186 21256 14242 21312
rect 13726 18944 13782 19000
rect 13542 18264 13598 18320
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 13358 17856 13414 17912
rect 14738 21684 14794 21720
rect 14738 21664 14740 21684
rect 14740 21664 14792 21684
rect 14792 21664 14794 21684
rect 14646 19760 14702 19816
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 11794 11600 11850 11656
rect 11334 9968 11390 10024
rect 12070 11500 12072 11520
rect 12072 11500 12124 11520
rect 12124 11500 12126 11520
rect 12070 11464 12126 11500
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 13450 14320 13506 14376
rect 12622 13812 12624 13832
rect 12624 13812 12676 13832
rect 12676 13812 12678 13832
rect 12622 13776 12678 13812
rect 12438 11464 12494 11520
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12898 11736 12954 11792
rect 13450 11736 13506 11792
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 13910 12144 13966 12200
rect 13910 12008 13966 12064
rect 13726 10648 13782 10704
rect 14370 18128 14426 18184
rect 15106 20848 15162 20904
rect 17774 24148 17776 24168
rect 17776 24148 17828 24168
rect 17828 24148 17830 24168
rect 16486 22752 16542 22808
rect 16026 22072 16082 22128
rect 15750 20032 15806 20088
rect 15474 17856 15530 17912
rect 14922 17584 14978 17640
rect 14646 17040 14702 17096
rect 14186 15544 14242 15600
rect 14278 14456 14334 14512
rect 14462 13368 14518 13424
rect 14370 13252 14426 13288
rect 14370 13232 14372 13252
rect 14372 13232 14424 13252
rect 14424 13232 14426 13252
rect 15198 16496 15254 16552
rect 14646 14864 14702 14920
rect 14922 14220 14924 14240
rect 14924 14220 14976 14240
rect 14976 14220 14978 14240
rect 14922 14184 14978 14220
rect 15290 14320 15346 14376
rect 15106 13504 15162 13560
rect 15014 13368 15070 13424
rect 14830 13132 14832 13152
rect 14832 13132 14884 13152
rect 14884 13132 14886 13152
rect 14830 13096 14886 13132
rect 14830 11500 14832 11520
rect 14832 11500 14884 11520
rect 14884 11500 14886 11520
rect 14830 11464 14886 11500
rect 14646 11056 14702 11112
rect 15106 11076 15162 11112
rect 15106 11056 15108 11076
rect 15108 11056 15160 11076
rect 15160 11056 15162 11076
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 15382 13096 15438 13152
rect 15014 10240 15070 10296
rect 16118 21548 16174 21584
rect 16118 21528 16120 21548
rect 16120 21528 16172 21548
rect 16172 21528 16174 21548
rect 16394 20748 16396 20768
rect 16396 20748 16448 20768
rect 16448 20748 16450 20768
rect 16394 20712 16450 20748
rect 16118 20460 16174 20496
rect 16118 20440 16120 20460
rect 16120 20440 16172 20460
rect 16172 20440 16174 20460
rect 16210 19896 16266 19952
rect 16210 19624 16266 19680
rect 15934 17484 15936 17504
rect 15936 17484 15988 17504
rect 15988 17484 15990 17504
rect 15934 17448 15990 17484
rect 16302 18964 16358 19000
rect 16302 18944 16304 18964
rect 16304 18944 16356 18964
rect 16356 18944 16358 18964
rect 16578 22072 16634 22128
rect 17774 24112 17830 24148
rect 17130 23316 17186 23352
rect 17130 23296 17132 23316
rect 17132 23296 17184 23316
rect 17184 23296 17186 23316
rect 16946 21800 17002 21856
rect 16854 20984 16910 21040
rect 17130 21120 17186 21176
rect 17130 20576 17186 20632
rect 16578 18944 16634 19000
rect 16762 18808 16818 18864
rect 17038 19080 17094 19136
rect 16394 17040 16450 17096
rect 15934 15952 15990 16008
rect 15934 15136 15990 15192
rect 16302 15680 16358 15736
rect 16210 14320 16266 14376
rect 16118 13912 16174 13968
rect 15658 13096 15714 13152
rect 15474 11756 15530 11792
rect 15474 11736 15476 11756
rect 15476 11736 15528 11756
rect 15528 11736 15530 11756
rect 15106 9288 15162 9344
rect 16026 12844 16082 12880
rect 16026 12824 16028 12844
rect 16028 12824 16080 12844
rect 16080 12824 16082 12844
rect 16394 13912 16450 13968
rect 16946 18128 17002 18184
rect 17130 16632 17186 16688
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17590 20984 17646 21040
rect 19062 23432 19118 23488
rect 21270 25472 21326 25528
rect 21178 24792 21234 24848
rect 20166 23296 20222 23352
rect 17958 20868 18014 20904
rect 17958 20848 17960 20868
rect 17960 20848 18012 20868
rect 18012 20848 18014 20868
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 18602 21936 18658 21992
rect 18878 21936 18934 21992
rect 18878 20984 18934 21040
rect 19338 20984 19394 21040
rect 17406 17312 17462 17368
rect 16762 14864 16818 14920
rect 16578 14048 16634 14104
rect 16118 12552 16174 12608
rect 16026 12144 16082 12200
rect 15658 10512 15714 10568
rect 15842 10240 15898 10296
rect 16486 10104 16542 10160
rect 16854 14320 16910 14376
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18326 19216 18382 19272
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 19890 22616 19946 22672
rect 20166 22616 20222 22672
rect 19982 21120 20038 21176
rect 19614 20712 19670 20768
rect 18510 18400 18566 18456
rect 17774 17176 17830 17232
rect 17682 16108 17738 16144
rect 17682 16088 17684 16108
rect 17684 16088 17736 16108
rect 17736 16088 17738 16108
rect 17222 14184 17278 14240
rect 17130 13096 17186 13152
rect 17682 14456 17738 14512
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17774 14184 17830 14240
rect 17590 13912 17646 13968
rect 17406 13776 17462 13832
rect 17314 13504 17370 13560
rect 17222 12144 17278 12200
rect 17130 12044 17132 12064
rect 17132 12044 17184 12064
rect 17184 12044 17186 12064
rect 17130 12008 17186 12044
rect 17222 11872 17278 11928
rect 16946 11600 17002 11656
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 16578 8200 16634 8256
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18694 19352 18750 19408
rect 18510 17992 18566 18048
rect 19706 20032 19762 20088
rect 19154 17992 19210 18048
rect 18878 15680 18934 15736
rect 18602 14476 18658 14512
rect 18602 14456 18604 14476
rect 18604 14456 18656 14476
rect 18656 14456 18658 14476
rect 18878 14728 18934 14784
rect 18878 14048 18934 14104
rect 18786 13776 18842 13832
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18602 11464 18658 11520
rect 18510 11092 18512 11112
rect 18512 11092 18564 11112
rect 18564 11092 18566 11112
rect 18510 11056 18566 11092
rect 18602 10004 18604 10024
rect 18604 10004 18656 10024
rect 18656 10004 18658 10024
rect 18602 9968 18658 10004
rect 19062 14320 19118 14376
rect 19614 18708 19616 18728
rect 19616 18708 19668 18728
rect 19668 18708 19670 18728
rect 19614 18672 19670 18708
rect 19430 16496 19486 16552
rect 19338 15680 19394 15736
rect 19154 13640 19210 13696
rect 19522 15136 19578 15192
rect 19890 18672 19946 18728
rect 20350 20712 20406 20768
rect 20166 17584 20222 17640
rect 19798 17176 19854 17232
rect 20994 21256 21050 21312
rect 22098 22924 22100 22944
rect 22100 22924 22152 22944
rect 22152 22924 22154 22944
rect 22098 22888 22154 22924
rect 21730 21800 21786 21856
rect 21270 21664 21326 21720
rect 22098 21392 22154 21448
rect 21454 20984 21510 21040
rect 22098 21120 22154 21176
rect 20902 17604 20958 17640
rect 20902 17584 20904 17604
rect 20904 17584 20956 17604
rect 20956 17584 20958 17604
rect 21454 20304 21510 20360
rect 21178 17176 21234 17232
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 20258 12588 20260 12608
rect 20260 12588 20312 12608
rect 20312 12588 20314 12608
rect 20258 12552 20314 12588
rect 19890 11872 19946 11928
rect 20626 12708 20682 12744
rect 20626 12688 20628 12708
rect 20628 12688 20680 12708
rect 20680 12688 20682 12708
rect 20994 11600 21050 11656
rect 19890 10784 19946 10840
rect 19890 10240 19946 10296
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 20718 10648 20774 10704
rect 20534 8880 20590 8936
rect 22006 20596 22062 20632
rect 22006 20576 22008 20596
rect 22008 20576 22060 20596
rect 22060 20576 22062 20596
rect 22006 18944 22062 19000
rect 21270 13096 21326 13152
rect 21638 14864 21694 14920
rect 22742 23704 22798 23760
rect 22466 23432 22522 23488
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22834 23024 22890 23080
rect 23110 22888 23166 22944
rect 23570 23160 23626 23216
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22374 21256 22430 21312
rect 22374 15580 22376 15600
rect 22376 15580 22428 15600
rect 22428 15580 22430 15600
rect 22374 15544 22430 15580
rect 22834 22072 22890 22128
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22834 20884 22836 20904
rect 22836 20884 22888 20904
rect 22888 20884 22890 20904
rect 22834 20848 22890 20884
rect 23846 23060 23848 23080
rect 23848 23060 23900 23080
rect 23900 23060 23902 23080
rect 23846 23024 23902 23060
rect 24858 24248 24914 24304
rect 24122 23432 24178 23488
rect 23938 22480 23994 22536
rect 23754 21120 23810 21176
rect 23662 20748 23664 20768
rect 23664 20748 23716 20768
rect 23716 20748 23718 20768
rect 23662 20712 23718 20748
rect 22742 19216 22798 19272
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 23846 20576 23902 20632
rect 24582 22072 24638 22128
rect 23478 19116 23480 19136
rect 23480 19116 23532 19136
rect 23532 19116 23534 19136
rect 23478 19080 23534 19116
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22466 14184 22522 14240
rect 21638 13132 21640 13152
rect 21640 13132 21692 13152
rect 21692 13132 21694 13152
rect 21638 13096 21694 13132
rect 21546 12552 21602 12608
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 21546 8372 21548 8392
rect 21548 8372 21600 8392
rect 21600 8372 21602 8392
rect 21546 8336 21602 8372
rect 22190 10648 22246 10704
rect 23938 16904 23994 16960
rect 23846 16632 23902 16688
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22834 15408 22890 15464
rect 23294 15136 23350 15192
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 23110 13404 23112 13424
rect 23112 13404 23164 13424
rect 23164 13404 23166 13424
rect 23110 13368 23166 13404
rect 22374 11892 22430 11928
rect 22374 11872 22376 11892
rect 22376 11872 22428 11892
rect 22428 11872 22430 11892
rect 22466 9016 22522 9072
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 24214 17332 24270 17368
rect 24214 17312 24216 17332
rect 24216 17312 24268 17332
rect 24268 17312 24270 17332
rect 25134 22072 25190 22128
rect 24582 20984 24638 21040
rect 24674 20032 24730 20088
rect 24490 19660 24492 19680
rect 24492 19660 24544 19680
rect 24544 19660 24546 19680
rect 24490 19624 24546 19660
rect 24306 17040 24362 17096
rect 23754 12144 23810 12200
rect 23294 11056 23350 11112
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 23754 11076 23810 11112
rect 23754 11056 23756 11076
rect 23756 11056 23808 11076
rect 23808 11056 23810 11076
rect 23386 9424 23442 9480
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 23478 8916 23480 8936
rect 23480 8916 23532 8936
rect 23532 8916 23534 8936
rect 23478 8880 23534 8916
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 24950 19760 25006 19816
rect 25134 18420 25190 18456
rect 25134 18400 25136 18420
rect 25136 18400 25188 18420
rect 25188 18400 25190 18420
rect 25042 18284 25098 18320
rect 25042 18264 25044 18284
rect 25044 18264 25096 18284
rect 25096 18264 25098 18284
rect 25778 23432 25834 23488
rect 25594 20984 25650 21040
rect 25410 20032 25466 20088
rect 25686 19252 25688 19272
rect 25688 19252 25740 19272
rect 25740 19252 25742 19272
rect 25686 19216 25742 19252
rect 26054 21528 26110 21584
rect 26698 22616 26754 22672
rect 26330 21004 26386 21040
rect 26330 20984 26332 21004
rect 26332 20984 26384 21004
rect 26384 20984 26386 21004
rect 26238 19660 26240 19680
rect 26240 19660 26292 19680
rect 26292 19660 26294 19680
rect 26238 19624 26294 19660
rect 25962 18944 26018 19000
rect 24674 15952 24730 16008
rect 24490 15544 24546 15600
rect 24582 13232 24638 13288
rect 24490 12824 24546 12880
rect 25134 16088 25190 16144
rect 25134 15680 25190 15736
rect 25318 17040 25374 17096
rect 25226 14728 25282 14784
rect 25410 15408 25466 15464
rect 26238 19216 26294 19272
rect 26698 19080 26754 19136
rect 27158 21684 27214 21720
rect 27158 21664 27160 21684
rect 27160 21664 27212 21684
rect 27212 21664 27214 21684
rect 27342 21836 27344 21856
rect 27344 21836 27396 21856
rect 27396 21836 27398 21856
rect 27342 21800 27398 21836
rect 27342 20304 27398 20360
rect 27066 19352 27122 19408
rect 27250 19352 27306 19408
rect 26882 18808 26938 18864
rect 26146 17720 26202 17776
rect 25410 14048 25466 14104
rect 25410 10512 25466 10568
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 25962 15272 26018 15328
rect 27066 17040 27122 17096
rect 27158 16632 27214 16688
rect 27066 16088 27122 16144
rect 26238 15544 26294 15600
rect 26146 12824 26202 12880
rect 26238 12280 26294 12336
rect 26974 15544 27030 15600
rect 26974 15308 26976 15328
rect 26976 15308 27028 15328
rect 27028 15308 27030 15328
rect 26974 15272 27030 15308
rect 27066 15000 27122 15056
rect 27342 18128 27398 18184
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 30102 26152 30158 26208
rect 29550 25744 29606 25800
rect 28446 23160 28502 23216
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 28354 21528 28410 21584
rect 28262 21120 28318 21176
rect 28354 20712 28410 20768
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 27802 20576 27858 20632
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 27710 18944 27766 19000
rect 28078 18944 28134 19000
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 27618 16904 27674 16960
rect 27434 15952 27490 16008
rect 27250 15020 27306 15056
rect 27250 15000 27252 15020
rect 27252 15000 27304 15020
rect 27304 15000 27306 15020
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 27802 17332 27858 17368
rect 27802 17312 27804 17332
rect 27804 17312 27856 17332
rect 27856 17312 27858 17332
rect 27802 17196 27858 17232
rect 27802 17176 27804 17196
rect 27804 17176 27856 17196
rect 27856 17176 27858 17196
rect 28078 17176 28134 17232
rect 27986 17040 28042 17096
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 28630 21836 28632 21856
rect 28632 21836 28684 21856
rect 28684 21836 28686 21856
rect 28630 21800 28686 21836
rect 28814 21664 28870 21720
rect 28814 21428 28816 21448
rect 28816 21428 28868 21448
rect 28868 21428 28870 21448
rect 28814 21392 28870 21428
rect 29090 22924 29092 22944
rect 29092 22924 29144 22944
rect 29144 22924 29146 22944
rect 29090 22888 29146 22924
rect 29918 24112 29974 24168
rect 30378 25336 30434 25392
rect 28814 20440 28870 20496
rect 28998 20440 29054 20496
rect 28814 19488 28870 19544
rect 28538 17448 28594 17504
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 28814 17620 28816 17640
rect 28816 17620 28868 17640
rect 28868 17620 28870 17640
rect 28814 17584 28870 17620
rect 29090 17584 29146 17640
rect 29090 17332 29146 17368
rect 29090 17312 29092 17332
rect 29092 17312 29144 17332
rect 29144 17312 29146 17332
rect 29090 17076 29092 17096
rect 29092 17076 29144 17096
rect 29144 17076 29146 17096
rect 29090 17040 29146 17076
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 27618 13096 27674 13152
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 27066 10104 27122 10160
rect 26054 9596 26056 9616
rect 26056 9596 26108 9616
rect 26108 9596 26110 9616
rect 26054 9560 26110 9596
rect 26146 9016 26202 9072
rect 26238 5072 26294 5128
rect 27434 11636 27436 11656
rect 27436 11636 27488 11656
rect 27488 11636 27490 11656
rect 27434 11600 27490 11636
rect 27342 10784 27398 10840
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 28722 13640 28778 13696
rect 28814 11736 28870 11792
rect 28630 11056 28686 11112
rect 29826 21800 29882 21856
rect 29734 20848 29790 20904
rect 29458 17040 29514 17096
rect 29274 14220 29276 14240
rect 29276 14220 29328 14240
rect 29328 14220 29330 14240
rect 29274 14184 29330 14220
rect 29182 11872 29238 11928
rect 28998 11600 29054 11656
rect 29458 12280 29514 12336
rect 28998 11192 29054 11248
rect 29734 16224 29790 16280
rect 30194 21800 30250 21856
rect 30378 21528 30434 21584
rect 30194 19896 30250 19952
rect 30286 19760 30342 19816
rect 30194 19624 30250 19680
rect 29918 18400 29974 18456
rect 29918 17176 29974 17232
rect 30378 18808 30434 18864
rect 30562 20712 30618 20768
rect 31482 26288 31538 26344
rect 31942 25880 31998 25936
rect 30746 22752 30802 22808
rect 30562 20168 30618 20224
rect 30102 15816 30158 15872
rect 30194 13912 30250 13968
rect 30010 12824 30066 12880
rect 29918 11872 29974 11928
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 30746 19896 30802 19952
rect 30746 19488 30802 19544
rect 31114 21392 31170 21448
rect 31390 22072 31446 22128
rect 31206 20168 31262 20224
rect 31390 20576 31446 20632
rect 30838 17720 30894 17776
rect 30562 10512 30618 10568
rect 31390 20032 31446 20088
rect 31298 19896 31354 19952
rect 31850 22888 31906 22944
rect 31666 21392 31722 21448
rect 31482 19080 31538 19136
rect 31022 17312 31078 17368
rect 31114 15816 31170 15872
rect 31022 15272 31078 15328
rect 30746 14728 30802 14784
rect 31114 13776 31170 13832
rect 31022 12280 31078 12336
rect 30930 12008 30986 12064
rect 30562 9988 30618 10024
rect 30562 9968 30564 9988
rect 30564 9968 30616 9988
rect 30616 9968 30618 9988
rect 31390 16224 31446 16280
rect 31850 19624 31906 19680
rect 31666 18536 31722 18592
rect 32586 26152 32642 26208
rect 32126 25064 32182 25120
rect 32218 24656 32274 24712
rect 32126 23840 32182 23896
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32586 22888 32642 22944
rect 32218 21800 32274 21856
rect 32126 20848 32182 20904
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 31482 13252 31538 13288
rect 31482 13232 31484 13252
rect 31484 13232 31536 13252
rect 31536 13232 31538 13252
rect 31758 17856 31814 17912
rect 31758 16516 31814 16552
rect 31758 16496 31760 16516
rect 31760 16496 31812 16516
rect 31812 16496 31814 16516
rect 31758 15272 31814 15328
rect 31666 14184 31722 14240
rect 31574 12724 31576 12744
rect 31576 12724 31628 12744
rect 31628 12724 31630 12744
rect 31574 12688 31630 12724
rect 32770 20984 32826 21040
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 33414 24248 33470 24304
rect 33598 23704 33654 23760
rect 34242 23840 34298 23896
rect 33414 21664 33470 21720
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 33046 20868 33102 20904
rect 33046 20848 33048 20868
rect 33048 20848 33100 20868
rect 33100 20848 33102 20868
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 32678 19760 32734 19816
rect 32678 19352 32734 19408
rect 33874 21664 33930 21720
rect 33690 21428 33692 21448
rect 33692 21428 33744 21448
rect 33744 21428 33746 21448
rect 33690 21392 33746 21428
rect 33598 21256 33654 21312
rect 33874 20848 33930 20904
rect 34058 22616 34114 22672
rect 33230 19252 33232 19272
rect 33232 19252 33284 19272
rect 33284 19252 33286 19272
rect 33230 19216 33286 19252
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 33138 18284 33194 18320
rect 33138 18264 33140 18284
rect 33140 18264 33192 18284
rect 33192 18264 33194 18284
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 33414 18420 33470 18456
rect 33414 18400 33416 18420
rect 33416 18400 33468 18420
rect 33468 18400 33470 18420
rect 33598 18400 33654 18456
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 32494 15680 32550 15736
rect 32862 16088 32918 16144
rect 33874 20032 33930 20088
rect 33874 19216 33930 19272
rect 33782 18808 33838 18864
rect 33966 18808 34022 18864
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 31850 12824 31906 12880
rect 31758 12144 31814 12200
rect 32218 14184 32274 14240
rect 32586 13368 32642 13424
rect 32034 11600 32090 11656
rect 31574 11056 31630 11112
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 33230 15136 33286 15192
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 33230 14456 33286 14512
rect 32954 14184 33010 14240
rect 33506 14456 33562 14512
rect 34518 21528 34574 21584
rect 34334 20304 34390 20360
rect 33966 17992 34022 18048
rect 33690 14728 33746 14784
rect 34058 15136 34114 15192
rect 34150 14728 34206 14784
rect 33322 14184 33378 14240
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 32770 11872 32826 11928
rect 32678 9424 32734 9480
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 34058 14184 34114 14240
rect 34150 12552 34206 12608
rect 33966 11056 34022 11112
rect 33690 10104 33746 10160
rect 33414 8916 33416 8936
rect 33416 8916 33468 8936
rect 33468 8916 33470 8936
rect 33414 8880 33470 8916
rect 33966 8916 33968 8936
rect 33968 8916 34020 8936
rect 34020 8916 34022 8936
rect 33966 8880 34022 8916
rect 34794 21120 34850 21176
rect 34794 18808 34850 18864
rect 34426 13368 34482 13424
rect 34978 20848 35034 20904
rect 35346 24112 35402 24168
rect 35714 25200 35770 25256
rect 35622 23860 35678 23896
rect 35622 23840 35624 23860
rect 35624 23840 35676 23860
rect 35676 23840 35678 23860
rect 35438 23296 35494 23352
rect 35346 22480 35402 22536
rect 37186 24928 37242 24984
rect 36082 23432 36138 23488
rect 35254 21936 35310 21992
rect 35070 20440 35126 20496
rect 34794 16124 34796 16144
rect 34796 16124 34848 16144
rect 34848 16124 34850 16144
rect 34794 16088 34850 16124
rect 35898 22072 35954 22128
rect 35346 19660 35348 19680
rect 35348 19660 35400 19680
rect 35400 19660 35402 19680
rect 35346 19624 35402 19660
rect 35254 19080 35310 19136
rect 35254 18944 35310 19000
rect 35070 16224 35126 16280
rect 35622 20984 35678 21040
rect 36450 22888 36506 22944
rect 36266 20476 36268 20496
rect 36268 20476 36320 20496
rect 36320 20476 36322 20496
rect 36266 20440 36322 20476
rect 35070 16088 35126 16144
rect 34978 15136 35034 15192
rect 35162 15816 35218 15872
rect 35346 15680 35402 15736
rect 35622 20032 35678 20088
rect 35898 19896 35954 19952
rect 35806 18808 35862 18864
rect 35806 16360 35862 16416
rect 34426 12008 34482 12064
rect 34702 12688 34758 12744
rect 34794 11872 34850 11928
rect 34702 11192 34758 11248
rect 34334 10920 34390 10976
rect 34426 10124 34482 10160
rect 34426 10104 34428 10124
rect 34428 10104 34480 10124
rect 34480 10104 34482 10124
rect 35254 11076 35310 11112
rect 35254 11056 35256 11076
rect 35256 11056 35308 11076
rect 35308 11056 35310 11076
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 34242 5616 34298 5672
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 35530 9424 35586 9480
rect 36634 20168 36690 20224
rect 36910 19216 36966 19272
rect 36910 18400 36966 18456
rect 36910 18264 36966 18320
rect 36726 17448 36782 17504
rect 36634 16632 36690 16688
rect 37830 24384 37886 24440
rect 37922 24112 37978 24168
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 37738 23568 37794 23624
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 38474 22752 38530 22808
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 37278 20304 37334 20360
rect 37094 18128 37150 18184
rect 37554 18944 37610 19000
rect 36910 16360 36966 16416
rect 36818 15952 36874 16008
rect 36450 12436 36506 12472
rect 36450 12416 36452 12436
rect 36452 12416 36504 12436
rect 36504 12416 36506 12436
rect 37278 13912 37334 13968
rect 36266 9560 36322 9616
rect 38474 21528 38530 21584
rect 38474 21120 38530 21176
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 39026 23840 39082 23896
rect 38934 23704 38990 23760
rect 39118 22072 39174 22128
rect 39854 26560 39910 26616
rect 39486 25880 39542 25936
rect 39394 24404 39450 24440
rect 39394 24384 39396 24404
rect 39396 24384 39448 24404
rect 39448 24384 39450 24404
rect 39394 23196 39396 23216
rect 39396 23196 39448 23216
rect 39448 23196 39450 23216
rect 39394 23160 39450 23196
rect 41418 26424 41474 26480
rect 39854 25880 39910 25936
rect 39394 22072 39450 22128
rect 39578 21956 39634 21992
rect 39578 21936 39580 21956
rect 39580 21936 39632 21956
rect 39632 21936 39634 21956
rect 38842 20440 38898 20496
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 37738 18944 37794 19000
rect 37738 18572 37740 18592
rect 37740 18572 37792 18592
rect 37792 18572 37794 18592
rect 37738 18536 37794 18572
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 37922 18284 37978 18320
rect 37922 18264 37924 18284
rect 37924 18264 37976 18284
rect 37976 18264 37978 18284
rect 37922 17992 37978 18048
rect 38474 18828 38530 18864
rect 38474 18808 38476 18828
rect 38476 18808 38528 18828
rect 38528 18808 38530 18828
rect 38474 18572 38476 18592
rect 38476 18572 38528 18592
rect 38528 18572 38530 18592
rect 38474 18536 38530 18572
rect 38290 17992 38346 18048
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 37830 16088 37886 16144
rect 37554 14728 37610 14784
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 38382 17332 38438 17368
rect 38382 17312 38384 17332
rect 38384 17312 38436 17332
rect 38436 17312 38438 17332
rect 38474 17040 38530 17096
rect 39486 19080 39542 19136
rect 39210 18672 39266 18728
rect 39210 18128 39266 18184
rect 39486 18128 39542 18184
rect 38842 16632 38898 16688
rect 39486 15952 39542 16008
rect 41602 25064 41658 25120
rect 41050 24112 41106 24168
rect 41510 23840 41566 23896
rect 40774 23160 40830 23216
rect 41142 23024 41198 23080
rect 40866 21936 40922 21992
rect 40314 20476 40316 20496
rect 40316 20476 40368 20496
rect 40368 20476 40370 20496
rect 40314 20440 40370 20476
rect 39854 20032 39910 20088
rect 40682 20712 40738 20768
rect 40958 20168 41014 20224
rect 40498 19216 40554 19272
rect 43534 25744 43590 25800
rect 42798 25608 42854 25664
rect 42430 23432 42486 23488
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 42798 24248 42854 24304
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 42706 22888 42762 22944
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 43718 25336 43774 25392
rect 43902 23316 43958 23352
rect 43902 23296 43904 23316
rect 43904 23296 43956 23316
rect 43956 23296 43958 23316
rect 43902 23180 43958 23216
rect 43902 23160 43904 23180
rect 43904 23160 43956 23180
rect 43956 23160 43958 23180
rect 43534 22636 43590 22672
rect 43534 22616 43536 22636
rect 43536 22616 43588 22636
rect 43588 22616 43590 22636
rect 44546 25880 44602 25936
rect 44270 25200 44326 25256
rect 44270 23296 44326 23352
rect 43810 22888 43866 22944
rect 44086 22888 44142 22944
rect 43902 22616 43958 22672
rect 43258 21392 43314 21448
rect 42798 21256 42854 21312
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 42338 20712 42394 20768
rect 40222 17312 40278 17368
rect 39854 17040 39910 17096
rect 39762 15952 39818 16008
rect 39670 15816 39726 15872
rect 40130 15680 40186 15736
rect 38566 15272 38622 15328
rect 39854 14728 39910 14784
rect 39486 14456 39542 14512
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 37554 12300 37610 12336
rect 37922 13812 37924 13832
rect 37924 13812 37976 13832
rect 37976 13812 37978 13832
rect 37922 13776 37978 13812
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 37554 12280 37556 12300
rect 37556 12280 37608 12300
rect 37608 12280 37610 12300
rect 38750 13252 38806 13288
rect 38750 13232 38752 13252
rect 38752 13232 38804 13252
rect 38804 13232 38806 13252
rect 38750 12588 38752 12608
rect 38752 12588 38804 12608
rect 38804 12588 38806 12608
rect 38750 12552 38806 12588
rect 38566 12416 38622 12472
rect 39854 13640 39910 13696
rect 40038 13640 40094 13696
rect 39302 12824 39358 12880
rect 40038 12688 40094 12744
rect 41602 18148 41658 18184
rect 41602 18128 41604 18148
rect 41604 18128 41656 18148
rect 41656 18128 41658 18148
rect 42614 20576 42670 20632
rect 43258 20440 43314 20496
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 44362 21664 44418 21720
rect 44914 24656 44970 24712
rect 44546 21664 44602 21720
rect 44546 20304 44602 20360
rect 44822 22480 44878 22536
rect 45006 20984 45062 21040
rect 45926 26152 45982 26208
rect 45466 24928 45522 24984
rect 45466 21664 45522 21720
rect 45558 21528 45614 21584
rect 45190 19896 45246 19952
rect 45742 21800 45798 21856
rect 45834 21548 45890 21584
rect 46386 23704 46442 23760
rect 45834 21528 45836 21548
rect 45836 21528 45888 21548
rect 45888 21528 45890 21548
rect 45742 20848 45798 20904
rect 42798 19352 42854 19408
rect 42154 18964 42210 19000
rect 42154 18944 42156 18964
rect 42156 18944 42208 18964
rect 42208 18944 42210 18964
rect 41970 18808 42026 18864
rect 41786 17856 41842 17912
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 42430 18536 42486 18592
rect 42798 17992 42854 18048
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 41050 17720 41106 17776
rect 40682 16516 40738 16552
rect 40682 16496 40684 16516
rect 40684 16496 40736 16516
rect 40736 16496 40738 16516
rect 40866 15272 40922 15328
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 38934 11736 38990 11792
rect 37738 10920 37794 10976
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 38290 9988 38346 10024
rect 38290 9968 38292 9988
rect 38292 9968 38344 9988
rect 38344 9968 38346 9988
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 40130 11636 40132 11656
rect 40132 11636 40184 11656
rect 40184 11636 40186 11656
rect 40130 11600 40186 11636
rect 40038 11328 40094 11384
rect 40130 11192 40186 11248
rect 40958 13932 41014 13968
rect 40958 13912 40960 13932
rect 40960 13912 41012 13932
rect 41012 13912 41014 13932
rect 40682 13504 40738 13560
rect 40314 11328 40370 11384
rect 40222 10648 40278 10704
rect 39486 10124 39542 10160
rect 39486 10104 39488 10124
rect 39488 10104 39540 10124
rect 39540 10104 39542 10124
rect 40774 11076 40830 11112
rect 40774 11056 40776 11076
rect 40776 11056 40828 11076
rect 40828 11056 40830 11076
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 37370 7540 37426 7576
rect 37370 7520 37372 7540
rect 37372 7520 37424 7540
rect 37424 7520 37426 7540
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 41326 13776 41382 13832
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 47030 25064 47086 25120
rect 46938 23024 46994 23080
rect 46846 22888 46902 22944
rect 47398 24656 47454 24712
rect 47766 24248 47822 24304
rect 47674 23432 47730 23488
rect 47582 23316 47638 23352
rect 47582 23296 47584 23316
rect 47584 23296 47636 23316
rect 47636 23296 47638 23316
rect 48502 26016 48558 26072
rect 48226 25472 48282 25528
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 48318 23060 48320 23080
rect 48320 23060 48372 23080
rect 48372 23060 48374 23080
rect 48318 23024 48374 23060
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 49146 23568 49202 23624
rect 49054 22616 49110 22672
rect 49330 22208 49386 22264
rect 48686 21800 48742 21856
rect 48502 20984 48558 21040
rect 48318 19216 48374 19272
rect 48594 20168 48650 20224
rect 49146 21392 49202 21448
rect 49238 20848 49294 20904
rect 49054 20576 49110 20632
rect 49054 19760 49110 19816
rect 49330 19352 49386 19408
rect 49146 18944 49202 19000
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 48778 18536 48834 18592
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 46110 17176 46166 17232
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 48318 15544 48374 15600
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 48318 14884 48374 14920
rect 48318 14864 48320 14884
rect 48320 14864 48372 14884
rect 48372 14864 48374 14884
rect 45282 13640 45338 13696
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 45558 13368 45614 13424
rect 48502 15000 48558 15056
rect 48226 13640 48282 13696
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 48778 16904 48834 16960
rect 49146 18128 49202 18184
rect 49054 17720 49110 17776
rect 49238 17584 49294 17640
rect 49054 17312 49110 17368
rect 49238 16496 49294 16552
rect 49146 16088 49202 16144
rect 49054 15680 49110 15736
rect 49238 15408 49294 15464
rect 49330 15272 49386 15328
rect 48686 12144 48742 12200
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 46846 7928 46902 7984
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 49054 14864 49110 14920
rect 49054 14456 49110 14512
rect 49238 14320 49294 14376
rect 49146 14048 49202 14104
rect 49146 13268 49148 13288
rect 49148 13268 49200 13288
rect 49200 13268 49202 13288
rect 49146 13232 49202 13268
rect 49146 12844 49202 12880
rect 49146 12824 49148 12844
rect 49148 12824 49200 12844
rect 49200 12824 49202 12844
rect 49146 12416 49202 12472
rect 49146 12008 49202 12064
rect 48962 11736 49018 11792
rect 49146 11600 49202 11656
rect 49238 11192 49294 11248
rect 49146 10784 49202 10840
rect 48778 10512 48834 10568
rect 49330 10376 49386 10432
rect 49238 9968 49294 10024
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 47306 9560 47362 9616
rect 49146 9152 49202 9208
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 49238 8744 49294 8800
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 46846 2624 46902 2680
rect 49330 8336 49386 8392
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 49146 7520 49202 7576
rect 49330 7112 49386 7168
rect 49238 6704 49294 6760
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 48870 6296 48926 6352
rect 49146 5888 49202 5944
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 49422 5480 49478 5536
rect 49330 5072 49386 5128
rect 48318 4664 48374 4720
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 49146 4256 49202 4312
rect 49238 3848 49294 3904
rect 46754 1808 46810 1864
rect 46662 1400 46718 1456
rect 49146 3440 49202 3496
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 48686 3032 48742 3088
rect 48502 2216 48558 2272
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
<< metal3 >>
rect 33542 26556 33548 26620
rect 33612 26618 33618 26620
rect 39849 26618 39915 26621
rect 33612 26616 39915 26618
rect 33612 26560 39854 26616
rect 39910 26560 39915 26616
rect 33612 26558 39915 26560
rect 33612 26556 33618 26558
rect 39849 26555 39915 26558
rect 41413 26482 41479 26485
rect 30238 26480 41479 26482
rect 30238 26424 41418 26480
rect 41474 26424 41479 26480
rect 30238 26422 41479 26424
rect 30097 26210 30163 26213
rect 30238 26210 30298 26422
rect 41413 26419 41479 26422
rect 31477 26346 31543 26349
rect 45686 26346 45692 26348
rect 31477 26344 45692 26346
rect 31477 26288 31482 26344
rect 31538 26288 45692 26344
rect 31477 26286 45692 26288
rect 31477 26283 31543 26286
rect 45686 26284 45692 26286
rect 45756 26284 45762 26348
rect 30097 26208 30298 26210
rect 30097 26152 30102 26208
rect 30158 26152 30298 26208
rect 30097 26150 30298 26152
rect 32581 26210 32647 26213
rect 45921 26210 45987 26213
rect 32581 26208 45987 26210
rect 32581 26152 32586 26208
rect 32642 26152 45926 26208
rect 45982 26152 45987 26208
rect 32581 26150 45987 26152
rect 30097 26147 30163 26150
rect 32581 26147 32647 26150
rect 45921 26147 45987 26150
rect 34278 26012 34284 26076
rect 34348 26074 34354 26076
rect 48497 26074 48563 26077
rect 34348 26072 48563 26074
rect 34348 26016 48502 26072
rect 48558 26016 48563 26072
rect 34348 26014 48563 26016
rect 34348 26012 34354 26014
rect 48497 26011 48563 26014
rect 31937 25938 32003 25941
rect 39481 25938 39547 25941
rect 31937 25936 39547 25938
rect 31937 25880 31942 25936
rect 31998 25880 39486 25936
rect 39542 25880 39547 25936
rect 31937 25878 39547 25880
rect 31937 25875 32003 25878
rect 39481 25875 39547 25878
rect 39849 25938 39915 25941
rect 44541 25938 44607 25941
rect 39849 25936 44607 25938
rect 39849 25880 39854 25936
rect 39910 25880 44546 25936
rect 44602 25880 44607 25936
rect 39849 25878 44607 25880
rect 39849 25875 39915 25878
rect 44541 25875 44607 25878
rect 29545 25802 29611 25805
rect 43529 25802 43595 25805
rect 29545 25800 43595 25802
rect 29545 25744 29550 25800
rect 29606 25744 43534 25800
rect 43590 25744 43595 25800
rect 29545 25742 43595 25744
rect 29545 25739 29611 25742
rect 43529 25739 43595 25742
rect 0 25666 800 25696
rect 3049 25666 3115 25669
rect 0 25664 3115 25666
rect 0 25608 3054 25664
rect 3110 25608 3115 25664
rect 0 25606 3115 25608
rect 0 25576 800 25606
rect 3049 25603 3115 25606
rect 19926 25604 19932 25668
rect 19996 25666 20002 25668
rect 42793 25666 42859 25669
rect 19996 25664 42859 25666
rect 19996 25608 42798 25664
rect 42854 25608 42859 25664
rect 19996 25606 42859 25608
rect 19996 25604 20002 25606
rect 42793 25603 42859 25606
rect 21265 25530 21331 25533
rect 44214 25530 44220 25532
rect 21265 25528 44220 25530
rect 21265 25472 21270 25528
rect 21326 25472 44220 25528
rect 21265 25470 44220 25472
rect 21265 25467 21331 25470
rect 44214 25468 44220 25470
rect 44284 25468 44290 25532
rect 48221 25530 48287 25533
rect 50200 25530 51000 25560
rect 48221 25528 51000 25530
rect 48221 25472 48226 25528
rect 48282 25472 51000 25528
rect 48221 25470 51000 25472
rect 48221 25467 48287 25470
rect 50200 25440 51000 25470
rect 30373 25394 30439 25397
rect 43713 25394 43779 25397
rect 30373 25392 43779 25394
rect 30373 25336 30378 25392
rect 30434 25336 43718 25392
rect 43774 25336 43779 25392
rect 30373 25334 43779 25336
rect 30373 25331 30439 25334
rect 43713 25331 43779 25334
rect 0 25258 800 25288
rect 3601 25258 3667 25261
rect 0 25256 3667 25258
rect 0 25200 3606 25256
rect 3662 25200 3667 25256
rect 0 25198 3667 25200
rect 0 25168 800 25198
rect 3601 25195 3667 25198
rect 35709 25258 35775 25261
rect 44265 25258 44331 25261
rect 35709 25256 44331 25258
rect 35709 25200 35714 25256
rect 35770 25200 44270 25256
rect 44326 25200 44331 25256
rect 35709 25198 44331 25200
rect 35709 25195 35775 25198
rect 44265 25195 44331 25198
rect 32121 25122 32187 25125
rect 41597 25122 41663 25125
rect 32121 25120 41663 25122
rect 32121 25064 32126 25120
rect 32182 25064 41602 25120
rect 41658 25064 41663 25120
rect 32121 25062 41663 25064
rect 32121 25059 32187 25062
rect 41597 25059 41663 25062
rect 47025 25122 47091 25125
rect 50200 25122 51000 25152
rect 47025 25120 51000 25122
rect 47025 25064 47030 25120
rect 47086 25064 51000 25120
rect 47025 25062 51000 25064
rect 47025 25059 47091 25062
rect 50200 25032 51000 25062
rect 37181 24986 37247 24989
rect 45461 24986 45527 24989
rect 37181 24984 45527 24986
rect 37181 24928 37186 24984
rect 37242 24928 45466 24984
rect 45522 24928 45527 24984
rect 37181 24926 45527 24928
rect 37181 24923 37247 24926
rect 45461 24923 45527 24926
rect 0 24850 800 24880
rect 3417 24850 3483 24853
rect 0 24848 3483 24850
rect 0 24792 3422 24848
rect 3478 24792 3483 24848
rect 0 24790 3483 24792
rect 0 24760 800 24790
rect 3417 24787 3483 24790
rect 3877 24850 3943 24853
rect 21173 24850 21239 24853
rect 3877 24848 21239 24850
rect 3877 24792 3882 24848
rect 3938 24792 21178 24848
rect 21234 24792 21239 24848
rect 3877 24790 21239 24792
rect 3877 24787 3943 24790
rect 21173 24787 21239 24790
rect 11973 24714 12039 24717
rect 30046 24714 30052 24716
rect 11973 24712 30052 24714
rect 11973 24656 11978 24712
rect 12034 24656 30052 24712
rect 11973 24654 30052 24656
rect 11973 24651 12039 24654
rect 30046 24652 30052 24654
rect 30116 24652 30122 24716
rect 32213 24714 32279 24717
rect 44909 24714 44975 24717
rect 32213 24712 44975 24714
rect 32213 24656 32218 24712
rect 32274 24656 44914 24712
rect 44970 24656 44975 24712
rect 32213 24654 44975 24656
rect 32213 24651 32279 24654
rect 44909 24651 44975 24654
rect 47393 24714 47459 24717
rect 50200 24714 51000 24744
rect 47393 24712 51000 24714
rect 47393 24656 47398 24712
rect 47454 24656 51000 24712
rect 47393 24654 51000 24656
rect 47393 24651 47459 24654
rect 50200 24624 51000 24654
rect 2946 24512 3262 24513
rect 0 24442 800 24472
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 2773 24442 2839 24445
rect 0 24440 2839 24442
rect 0 24384 2778 24440
rect 2834 24384 2839 24440
rect 0 24382 2839 24384
rect 0 24352 800 24382
rect 2773 24379 2839 24382
rect 37825 24442 37891 24445
rect 39389 24442 39455 24445
rect 37825 24440 39455 24442
rect 37825 24384 37830 24440
rect 37886 24384 39394 24440
rect 39450 24384 39455 24440
rect 37825 24382 39455 24384
rect 37825 24379 37891 24382
rect 39389 24379 39455 24382
rect 7373 24306 7439 24309
rect 24853 24306 24919 24309
rect 7373 24304 24919 24306
rect 7373 24248 7378 24304
rect 7434 24248 24858 24304
rect 24914 24248 24919 24304
rect 7373 24246 24919 24248
rect 7373 24243 7439 24246
rect 24853 24243 24919 24246
rect 33409 24306 33475 24309
rect 42793 24306 42859 24309
rect 33409 24304 42859 24306
rect 33409 24248 33414 24304
rect 33470 24248 42798 24304
rect 42854 24248 42859 24304
rect 33409 24246 42859 24248
rect 33409 24243 33475 24246
rect 42793 24243 42859 24246
rect 47761 24306 47827 24309
rect 50200 24306 51000 24336
rect 47761 24304 51000 24306
rect 47761 24248 47766 24304
rect 47822 24248 51000 24304
rect 47761 24246 51000 24248
rect 47761 24243 47827 24246
rect 50200 24216 51000 24246
rect 17769 24170 17835 24173
rect 29913 24170 29979 24173
rect 17769 24168 29979 24170
rect 17769 24112 17774 24168
rect 17830 24112 29918 24168
rect 29974 24112 29979 24168
rect 17769 24110 29979 24112
rect 17769 24107 17835 24110
rect 29913 24107 29979 24110
rect 35341 24170 35407 24173
rect 37917 24170 37983 24173
rect 41045 24170 41111 24173
rect 35341 24168 41111 24170
rect 35341 24112 35346 24168
rect 35402 24112 37922 24168
rect 37978 24112 41050 24168
rect 41106 24112 41111 24168
rect 35341 24110 41111 24112
rect 35341 24107 35407 24110
rect 37917 24107 37983 24110
rect 41045 24107 41111 24110
rect 0 24034 800 24064
rect 3509 24034 3575 24037
rect 0 24032 3575 24034
rect 0 23976 3514 24032
rect 3570 23976 3575 24032
rect 0 23974 3575 23976
rect 0 23944 800 23974
rect 3509 23971 3575 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 32121 23898 32187 23901
rect 34237 23898 34303 23901
rect 35617 23898 35683 23901
rect 32121 23896 35683 23898
rect 32121 23840 32126 23896
rect 32182 23840 34242 23896
rect 34298 23840 35622 23896
rect 35678 23840 35683 23896
rect 32121 23838 35683 23840
rect 32121 23835 32187 23838
rect 34237 23835 34303 23838
rect 35617 23835 35683 23838
rect 39021 23898 39087 23901
rect 41505 23898 41571 23901
rect 50200 23898 51000 23928
rect 39021 23896 41571 23898
rect 39021 23840 39026 23896
rect 39082 23840 41510 23896
rect 41566 23840 41571 23896
rect 39021 23838 41571 23840
rect 39021 23835 39087 23838
rect 41505 23835 41571 23838
rect 48454 23838 51000 23898
rect 12065 23762 12131 23765
rect 22737 23762 22803 23765
rect 12065 23760 22803 23762
rect 12065 23704 12070 23760
rect 12126 23704 22742 23760
rect 22798 23704 22803 23760
rect 12065 23702 22803 23704
rect 12065 23699 12131 23702
rect 22737 23699 22803 23702
rect 33593 23762 33659 23765
rect 38929 23762 38995 23765
rect 33593 23760 38995 23762
rect 33593 23704 33598 23760
rect 33654 23704 38934 23760
rect 38990 23704 38995 23760
rect 33593 23702 38995 23704
rect 33593 23699 33659 23702
rect 38929 23699 38995 23702
rect 46381 23762 46447 23765
rect 48454 23762 48514 23838
rect 50200 23808 51000 23838
rect 46381 23760 48514 23762
rect 46381 23704 46386 23760
rect 46442 23704 48514 23760
rect 46381 23702 48514 23704
rect 46381 23699 46447 23702
rect 0 23626 800 23656
rect 3417 23626 3483 23629
rect 0 23624 3483 23626
rect 0 23568 3422 23624
rect 3478 23568 3483 23624
rect 0 23566 3483 23568
rect 0 23536 800 23566
rect 3417 23563 3483 23566
rect 37733 23626 37799 23629
rect 49141 23626 49207 23629
rect 37733 23624 49207 23626
rect 37733 23568 37738 23624
rect 37794 23568 49146 23624
rect 49202 23568 49207 23624
rect 37733 23566 49207 23568
rect 37733 23563 37799 23566
rect 49141 23563 49207 23566
rect 19057 23490 19123 23493
rect 22461 23490 22527 23493
rect 19057 23488 22527 23490
rect 19057 23432 19062 23488
rect 19118 23432 22466 23488
rect 22522 23432 22527 23488
rect 19057 23430 22527 23432
rect 19057 23427 19123 23430
rect 22461 23427 22527 23430
rect 24117 23490 24183 23493
rect 25773 23490 25839 23493
rect 24117 23488 25839 23490
rect 24117 23432 24122 23488
rect 24178 23432 25778 23488
rect 25834 23432 25839 23488
rect 24117 23430 25839 23432
rect 24117 23427 24183 23430
rect 25773 23427 25839 23430
rect 36077 23490 36143 23493
rect 42425 23490 42491 23493
rect 36077 23488 42491 23490
rect 36077 23432 36082 23488
rect 36138 23432 42430 23488
rect 42486 23432 42491 23488
rect 36077 23430 42491 23432
rect 36077 23427 36143 23430
rect 42425 23427 42491 23430
rect 47669 23490 47735 23493
rect 50200 23490 51000 23520
rect 47669 23488 51000 23490
rect 47669 23432 47674 23488
rect 47730 23432 51000 23488
rect 47669 23430 51000 23432
rect 47669 23427 47735 23430
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 50200 23400 51000 23430
rect 42946 23359 43262 23360
rect 17125 23354 17191 23357
rect 20161 23354 20227 23357
rect 17125 23352 20227 23354
rect 17125 23296 17130 23352
rect 17186 23296 20166 23352
rect 20222 23296 20227 23352
rect 17125 23294 20227 23296
rect 17125 23291 17191 23294
rect 20161 23291 20227 23294
rect 35433 23354 35499 23357
rect 43897 23354 43963 23357
rect 44265 23354 44331 23357
rect 47577 23354 47643 23357
rect 35433 23352 41430 23354
rect 35433 23296 35438 23352
rect 35494 23296 41430 23352
rect 35433 23294 41430 23296
rect 35433 23291 35499 23294
rect 0 23218 800 23248
rect 3417 23218 3483 23221
rect 0 23216 3483 23218
rect 0 23160 3422 23216
rect 3478 23160 3483 23216
rect 0 23158 3483 23160
rect 0 23128 800 23158
rect 3417 23155 3483 23158
rect 9397 23218 9463 23221
rect 23565 23218 23631 23221
rect 9397 23216 23631 23218
rect 9397 23160 9402 23216
rect 9458 23160 23570 23216
rect 23626 23160 23631 23216
rect 9397 23158 23631 23160
rect 9397 23155 9463 23158
rect 23565 23155 23631 23158
rect 28441 23218 28507 23221
rect 39389 23218 39455 23221
rect 40769 23218 40835 23221
rect 28441 23216 38578 23218
rect 28441 23160 28446 23216
rect 28502 23160 38578 23216
rect 28441 23158 38578 23160
rect 28441 23155 28507 23158
rect 9213 23082 9279 23085
rect 22829 23082 22895 23085
rect 9213 23080 22895 23082
rect 9213 23024 9218 23080
rect 9274 23024 22834 23080
rect 22890 23024 22895 23080
rect 9213 23022 22895 23024
rect 9213 23019 9279 23022
rect 22829 23019 22895 23022
rect 23841 23082 23907 23085
rect 38518 23082 38578 23158
rect 39389 23216 40835 23218
rect 39389 23160 39394 23216
rect 39450 23160 40774 23216
rect 40830 23160 40835 23216
rect 39389 23158 40835 23160
rect 41370 23218 41430 23294
rect 43897 23352 47643 23354
rect 43897 23296 43902 23352
rect 43958 23296 44270 23352
rect 44326 23296 47582 23352
rect 47638 23296 47643 23352
rect 43897 23294 47643 23296
rect 43897 23291 43963 23294
rect 44265 23291 44331 23294
rect 47577 23291 47643 23294
rect 43897 23218 43963 23221
rect 41370 23216 43963 23218
rect 41370 23160 43902 23216
rect 43958 23160 43963 23216
rect 41370 23158 43963 23160
rect 39389 23155 39455 23158
rect 40769 23155 40835 23158
rect 43897 23155 43963 23158
rect 41137 23082 41203 23085
rect 46933 23082 46999 23085
rect 23841 23080 38394 23082
rect 23841 23024 23846 23080
rect 23902 23024 38394 23080
rect 23841 23022 38394 23024
rect 38518 23080 46999 23082
rect 38518 23024 41142 23080
rect 41198 23024 46938 23080
rect 46994 23024 46999 23080
rect 38518 23022 46999 23024
rect 23841 23019 23907 23022
rect 22093 22946 22159 22949
rect 23105 22946 23171 22949
rect 22093 22944 23171 22946
rect 22093 22888 22098 22944
rect 22154 22888 23110 22944
rect 23166 22888 23171 22944
rect 22093 22886 23171 22888
rect 22093 22883 22159 22886
rect 23105 22883 23171 22886
rect 29085 22946 29151 22949
rect 31845 22946 31911 22949
rect 29085 22944 31911 22946
rect 29085 22888 29090 22944
rect 29146 22888 31850 22944
rect 31906 22888 31911 22944
rect 29085 22886 31911 22888
rect 29085 22883 29151 22886
rect 31845 22883 31911 22886
rect 32581 22946 32647 22949
rect 36445 22946 36511 22949
rect 32581 22944 36511 22946
rect 32581 22888 32586 22944
rect 32642 22888 36450 22944
rect 36506 22888 36511 22944
rect 32581 22886 36511 22888
rect 38334 22946 38394 23022
rect 41137 23019 41203 23022
rect 46933 23019 46999 23022
rect 48313 23082 48379 23085
rect 50200 23082 51000 23112
rect 48313 23080 51000 23082
rect 48313 23024 48318 23080
rect 48374 23024 51000 23080
rect 48313 23022 51000 23024
rect 48313 23019 48379 23022
rect 50200 22992 51000 23022
rect 42701 22946 42767 22949
rect 38334 22944 42767 22946
rect 38334 22888 42706 22944
rect 42762 22888 42767 22944
rect 38334 22886 42767 22888
rect 32581 22883 32647 22886
rect 36445 22883 36511 22886
rect 42701 22883 42767 22886
rect 43805 22946 43871 22949
rect 44081 22946 44147 22949
rect 46841 22946 46907 22949
rect 43805 22944 46907 22946
rect 43805 22888 43810 22944
rect 43866 22888 44086 22944
rect 44142 22888 46846 22944
rect 46902 22888 46907 22944
rect 43805 22886 46907 22888
rect 43805 22883 43871 22886
rect 44081 22883 44147 22886
rect 46841 22883 46907 22886
rect 7946 22880 8262 22881
rect 0 22810 800 22840
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 47946 22815 48262 22816
rect 3141 22810 3207 22813
rect 0 22808 3207 22810
rect 0 22752 3146 22808
rect 3202 22752 3207 22808
rect 0 22750 3207 22752
rect 0 22720 800 22750
rect 3141 22747 3207 22750
rect 11513 22810 11579 22813
rect 16481 22810 16547 22813
rect 11513 22808 16547 22810
rect 11513 22752 11518 22808
rect 11574 22752 16486 22808
rect 16542 22752 16547 22808
rect 11513 22750 16547 22752
rect 11513 22747 11579 22750
rect 16481 22747 16547 22750
rect 30741 22810 30807 22813
rect 36486 22810 36492 22812
rect 30741 22808 36492 22810
rect 30741 22752 30746 22808
rect 30802 22752 36492 22808
rect 30741 22750 36492 22752
rect 30741 22747 30807 22750
rect 36486 22748 36492 22750
rect 36556 22748 36562 22812
rect 38469 22810 38535 22813
rect 38469 22808 43730 22810
rect 38469 22752 38474 22808
rect 38530 22752 43730 22808
rect 38469 22750 43730 22752
rect 38469 22747 38535 22750
rect 11697 22674 11763 22677
rect 19885 22676 19951 22677
rect 19885 22674 19932 22676
rect 11697 22672 19932 22674
rect 19996 22674 20002 22676
rect 20161 22674 20227 22677
rect 26693 22674 26759 22677
rect 11697 22616 11702 22672
rect 11758 22616 19890 22672
rect 11697 22614 19932 22616
rect 11697 22611 11763 22614
rect 19885 22612 19932 22614
rect 19996 22614 20078 22674
rect 20161 22672 26759 22674
rect 20161 22616 20166 22672
rect 20222 22616 26698 22672
rect 26754 22616 26759 22672
rect 20161 22614 26759 22616
rect 19996 22612 20002 22614
rect 19885 22611 19951 22612
rect 20161 22611 20227 22614
rect 26693 22611 26759 22614
rect 34053 22674 34119 22677
rect 43529 22674 43595 22677
rect 34053 22672 43595 22674
rect 34053 22616 34058 22672
rect 34114 22616 43534 22672
rect 43590 22616 43595 22672
rect 34053 22614 43595 22616
rect 43670 22674 43730 22750
rect 43897 22674 43963 22677
rect 43670 22672 43963 22674
rect 43670 22616 43902 22672
rect 43958 22616 43963 22672
rect 43670 22614 43963 22616
rect 34053 22611 34119 22614
rect 43529 22611 43595 22614
rect 43897 22611 43963 22614
rect 49049 22674 49115 22677
rect 50200 22674 51000 22704
rect 49049 22672 51000 22674
rect 49049 22616 49054 22672
rect 49110 22616 51000 22672
rect 49049 22614 51000 22616
rect 49049 22611 49115 22614
rect 50200 22584 51000 22614
rect 4153 22538 4219 22541
rect 11789 22538 11855 22541
rect 23933 22538 23999 22541
rect 4153 22536 11714 22538
rect 4153 22480 4158 22536
rect 4214 22480 11714 22536
rect 4153 22478 11714 22480
rect 4153 22475 4219 22478
rect 0 22402 800 22432
rect 0 22342 2514 22402
rect 0 22312 800 22342
rect 2454 22130 2514 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 3969 22266 4035 22269
rect 11513 22266 11579 22269
rect 3969 22264 11579 22266
rect 3969 22208 3974 22264
rect 4030 22208 11518 22264
rect 11574 22208 11579 22264
rect 3969 22206 11579 22208
rect 3969 22203 4035 22206
rect 11513 22203 11579 22206
rect 4153 22130 4219 22133
rect 2454 22128 4219 22130
rect 2454 22072 4158 22128
rect 4214 22072 4219 22128
rect 2454 22070 4219 22072
rect 11654 22130 11714 22478
rect 11789 22536 23999 22538
rect 11789 22480 11794 22536
rect 11850 22480 23938 22536
rect 23994 22480 23999 22536
rect 11789 22478 23999 22480
rect 11789 22475 11855 22478
rect 23933 22475 23999 22478
rect 35341 22538 35407 22541
rect 44817 22538 44883 22541
rect 35341 22536 44883 22538
rect 35341 22480 35346 22536
rect 35402 22480 44822 22536
rect 44878 22480 44883 22536
rect 35341 22478 44883 22480
rect 35341 22475 35407 22478
rect 44817 22475 44883 22478
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 49325 22266 49391 22269
rect 50200 22266 51000 22296
rect 49325 22264 51000 22266
rect 49325 22208 49330 22264
rect 49386 22208 51000 22264
rect 49325 22206 51000 22208
rect 49325 22203 49391 22206
rect 50200 22176 51000 22206
rect 16021 22130 16087 22133
rect 11654 22128 16087 22130
rect 11654 22072 16026 22128
rect 16082 22072 16087 22128
rect 11654 22070 16087 22072
rect 4153 22067 4219 22070
rect 16021 22067 16087 22070
rect 16573 22130 16639 22133
rect 22829 22130 22895 22133
rect 16573 22128 22895 22130
rect 16573 22072 16578 22128
rect 16634 22072 22834 22128
rect 22890 22072 22895 22128
rect 16573 22070 22895 22072
rect 16573 22067 16639 22070
rect 22829 22067 22895 22070
rect 24577 22130 24643 22133
rect 25129 22130 25195 22133
rect 24577 22128 25195 22130
rect 24577 22072 24582 22128
rect 24638 22072 25134 22128
rect 25190 22072 25195 22128
rect 24577 22070 25195 22072
rect 24577 22067 24643 22070
rect 25129 22067 25195 22070
rect 31385 22130 31451 22133
rect 35893 22130 35959 22133
rect 39113 22130 39179 22133
rect 39389 22130 39455 22133
rect 31385 22128 39455 22130
rect 31385 22072 31390 22128
rect 31446 22072 35898 22128
rect 35954 22072 39118 22128
rect 39174 22072 39394 22128
rect 39450 22072 39455 22128
rect 31385 22070 39455 22072
rect 31385 22067 31451 22070
rect 35893 22067 35959 22070
rect 39113 22067 39179 22070
rect 39389 22067 39455 22070
rect 0 21994 800 22024
rect 3785 21994 3851 21997
rect 0 21992 3851 21994
rect 0 21936 3790 21992
rect 3846 21936 3851 21992
rect 0 21934 3851 21936
rect 0 21904 800 21934
rect 3785 21931 3851 21934
rect 7925 21994 7991 21997
rect 18597 21994 18663 21997
rect 7925 21992 18663 21994
rect 7925 21936 7930 21992
rect 7986 21936 18602 21992
rect 18658 21936 18663 21992
rect 7925 21934 18663 21936
rect 7925 21931 7991 21934
rect 18597 21931 18663 21934
rect 18873 21994 18939 21997
rect 35249 21994 35315 21997
rect 39573 21994 39639 21997
rect 40861 21994 40927 21997
rect 18873 21992 40927 21994
rect 18873 21936 18878 21992
rect 18934 21936 35254 21992
rect 35310 21936 39578 21992
rect 39634 21936 40866 21992
rect 40922 21936 40927 21992
rect 18873 21934 40927 21936
rect 18873 21931 18939 21934
rect 35249 21931 35315 21934
rect 39573 21931 39639 21934
rect 40861 21931 40927 21934
rect 10317 21858 10383 21861
rect 16941 21858 17007 21861
rect 10317 21856 17007 21858
rect 10317 21800 10322 21856
rect 10378 21800 16946 21856
rect 17002 21800 17007 21856
rect 10317 21798 17007 21800
rect 10317 21795 10383 21798
rect 16941 21795 17007 21798
rect 21725 21858 21791 21861
rect 27337 21858 27403 21861
rect 21725 21856 27403 21858
rect 21725 21800 21730 21856
rect 21786 21800 27342 21856
rect 27398 21800 27403 21856
rect 21725 21798 27403 21800
rect 21725 21795 21791 21798
rect 27337 21795 27403 21798
rect 28625 21858 28691 21861
rect 29821 21858 29887 21861
rect 28625 21856 29887 21858
rect 28625 21800 28630 21856
rect 28686 21800 29826 21856
rect 29882 21800 29887 21856
rect 28625 21798 29887 21800
rect 28625 21795 28691 21798
rect 29821 21795 29887 21798
rect 30189 21858 30255 21861
rect 32213 21858 32279 21861
rect 45737 21858 45803 21861
rect 30189 21856 32279 21858
rect 30189 21800 30194 21856
rect 30250 21800 32218 21856
rect 32274 21800 32279 21856
rect 30189 21798 32279 21800
rect 30189 21795 30255 21798
rect 32213 21795 32279 21798
rect 38334 21856 45803 21858
rect 38334 21800 45742 21856
rect 45798 21800 45803 21856
rect 38334 21798 45803 21800
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 10685 21722 10751 21725
rect 14733 21722 14799 21725
rect 10685 21720 14799 21722
rect 10685 21664 10690 21720
rect 10746 21664 14738 21720
rect 14794 21664 14799 21720
rect 10685 21662 14799 21664
rect 10685 21659 10751 21662
rect 14733 21659 14799 21662
rect 21265 21722 21331 21725
rect 27153 21722 27219 21725
rect 21265 21720 27219 21722
rect 21265 21664 21270 21720
rect 21326 21664 27158 21720
rect 27214 21664 27219 21720
rect 21265 21662 27219 21664
rect 21265 21659 21331 21662
rect 27153 21659 27219 21662
rect 28809 21722 28875 21725
rect 33409 21722 33475 21725
rect 28809 21720 33475 21722
rect 28809 21664 28814 21720
rect 28870 21664 33414 21720
rect 33470 21664 33475 21720
rect 28809 21662 33475 21664
rect 28809 21659 28875 21662
rect 33409 21659 33475 21662
rect 33869 21722 33935 21725
rect 34278 21722 34284 21724
rect 33869 21720 34284 21722
rect 33869 21664 33874 21720
rect 33930 21664 34284 21720
rect 33869 21662 34284 21664
rect 33869 21659 33935 21662
rect 34278 21660 34284 21662
rect 34348 21660 34354 21724
rect 0 21586 800 21616
rect 2681 21586 2747 21589
rect 0 21584 2747 21586
rect 0 21528 2686 21584
rect 2742 21528 2747 21584
rect 0 21526 2747 21528
rect 0 21496 800 21526
rect 2681 21523 2747 21526
rect 9029 21586 9095 21589
rect 16113 21586 16179 21589
rect 26049 21586 26115 21589
rect 9029 21584 26115 21586
rect 9029 21528 9034 21584
rect 9090 21528 16118 21584
rect 16174 21528 26054 21584
rect 26110 21528 26115 21584
rect 9029 21526 26115 21528
rect 9029 21523 9095 21526
rect 16113 21523 16179 21526
rect 26049 21523 26115 21526
rect 28349 21586 28415 21589
rect 30373 21586 30439 21589
rect 34513 21586 34579 21589
rect 38334 21586 38394 21798
rect 45737 21795 45803 21798
rect 48681 21858 48747 21861
rect 50200 21858 51000 21888
rect 48681 21856 51000 21858
rect 48681 21800 48686 21856
rect 48742 21800 51000 21856
rect 48681 21798 51000 21800
rect 48681 21795 48747 21798
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 50200 21768 51000 21798
rect 47946 21727 48262 21728
rect 44214 21660 44220 21724
rect 44284 21722 44290 21724
rect 44357 21722 44423 21725
rect 44284 21720 44423 21722
rect 44284 21664 44362 21720
rect 44418 21664 44423 21720
rect 44284 21662 44423 21664
rect 44284 21660 44290 21662
rect 44357 21659 44423 21662
rect 44541 21722 44607 21725
rect 45461 21722 45527 21725
rect 44541 21720 45527 21722
rect 44541 21664 44546 21720
rect 44602 21664 45466 21720
rect 45522 21664 45527 21720
rect 44541 21662 45527 21664
rect 44541 21659 44607 21662
rect 45461 21659 45527 21662
rect 28349 21584 38394 21586
rect 28349 21528 28354 21584
rect 28410 21528 30378 21584
rect 30434 21528 34518 21584
rect 34574 21528 38394 21584
rect 28349 21526 38394 21528
rect 38469 21586 38535 21589
rect 45553 21586 45619 21589
rect 38469 21584 45619 21586
rect 38469 21528 38474 21584
rect 38530 21528 45558 21584
rect 45614 21528 45619 21584
rect 38469 21526 45619 21528
rect 28349 21523 28415 21526
rect 30373 21523 30439 21526
rect 34513 21523 34579 21526
rect 38469 21523 38535 21526
rect 45553 21523 45619 21526
rect 45686 21524 45692 21588
rect 45756 21586 45762 21588
rect 45829 21586 45895 21589
rect 45756 21584 45895 21586
rect 45756 21528 45834 21584
rect 45890 21528 45895 21584
rect 45756 21526 45895 21528
rect 45756 21524 45762 21526
rect 45829 21523 45895 21526
rect 5441 21450 5507 21453
rect 7833 21450 7899 21453
rect 5441 21448 7899 21450
rect 5441 21392 5446 21448
rect 5502 21392 7838 21448
rect 7894 21392 7899 21448
rect 5441 21390 7899 21392
rect 5441 21387 5507 21390
rect 7833 21387 7899 21390
rect 11145 21450 11211 21453
rect 22093 21450 22159 21453
rect 28809 21450 28875 21453
rect 31109 21450 31175 21453
rect 31661 21450 31727 21453
rect 11145 21448 21236 21450
rect 11145 21392 11150 21448
rect 11206 21392 21236 21448
rect 11145 21390 21236 21392
rect 11145 21387 11211 21390
rect 14181 21314 14247 21317
rect 20989 21314 21055 21317
rect 14181 21312 21055 21314
rect 14181 21256 14186 21312
rect 14242 21256 20994 21312
rect 21050 21256 21055 21312
rect 14181 21254 21055 21256
rect 21176 21314 21236 21390
rect 22093 21448 23812 21450
rect 22093 21392 22098 21448
rect 22154 21392 23812 21448
rect 22093 21390 23812 21392
rect 22093 21387 22159 21390
rect 22369 21314 22435 21317
rect 21176 21312 22435 21314
rect 21176 21256 22374 21312
rect 22430 21256 22435 21312
rect 21176 21254 22435 21256
rect 14181 21251 14247 21254
rect 20989 21251 21055 21254
rect 22369 21251 22435 21254
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 23752 21181 23812 21390
rect 28809 21448 31727 21450
rect 28809 21392 28814 21448
rect 28870 21392 31114 21448
rect 31170 21392 31666 21448
rect 31722 21392 31727 21448
rect 28809 21390 31727 21392
rect 28809 21387 28875 21390
rect 31109 21387 31175 21390
rect 31661 21387 31727 21390
rect 33685 21450 33751 21453
rect 43253 21450 43319 21453
rect 33685 21448 43319 21450
rect 33685 21392 33690 21448
rect 33746 21392 43258 21448
rect 43314 21392 43319 21448
rect 33685 21390 43319 21392
rect 33685 21387 33751 21390
rect 43253 21387 43319 21390
rect 49141 21450 49207 21453
rect 50200 21450 51000 21480
rect 49141 21448 51000 21450
rect 49141 21392 49146 21448
rect 49202 21392 51000 21448
rect 49141 21390 51000 21392
rect 49141 21387 49207 21390
rect 50200 21360 51000 21390
rect 33593 21314 33659 21317
rect 42793 21314 42859 21317
rect 33593 21312 42859 21314
rect 33593 21256 33598 21312
rect 33654 21256 42798 21312
rect 42854 21256 42859 21312
rect 33593 21254 42859 21256
rect 33593 21251 33659 21254
rect 42793 21251 42859 21254
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 0 21088 800 21118
rect 2773 21115 2839 21118
rect 17125 21178 17191 21181
rect 19977 21178 20043 21181
rect 22093 21178 22159 21181
rect 17125 21176 20043 21178
rect 17125 21120 17130 21176
rect 17186 21120 19982 21176
rect 20038 21120 20043 21176
rect 17125 21118 20043 21120
rect 17125 21115 17191 21118
rect 19977 21115 20043 21118
rect 20118 21176 22159 21178
rect 20118 21120 22098 21176
rect 22154 21120 22159 21176
rect 20118 21118 22159 21120
rect 7782 20980 7788 21044
rect 7852 21042 7858 21044
rect 16849 21042 16915 21045
rect 7852 21040 16915 21042
rect 7852 20984 16854 21040
rect 16910 20984 16915 21040
rect 7852 20982 16915 20984
rect 7852 20980 7858 20982
rect 16849 20979 16915 20982
rect 17585 21042 17651 21045
rect 18873 21042 18939 21045
rect 17585 21040 18939 21042
rect 17585 20984 17590 21040
rect 17646 20984 18878 21040
rect 18934 20984 18939 21040
rect 17585 20982 18939 20984
rect 17585 20979 17651 20982
rect 18873 20979 18939 20982
rect 19333 21042 19399 21045
rect 20118 21042 20178 21118
rect 22093 21115 22159 21118
rect 23749 21178 23815 21181
rect 28257 21178 28323 21181
rect 23749 21176 28323 21178
rect 23749 21120 23754 21176
rect 23810 21120 28262 21176
rect 28318 21120 28323 21176
rect 23749 21118 28323 21120
rect 23749 21115 23815 21118
rect 28257 21115 28323 21118
rect 34789 21178 34855 21181
rect 38469 21178 38535 21181
rect 34789 21176 38535 21178
rect 34789 21120 34794 21176
rect 34850 21120 38474 21176
rect 38530 21120 38535 21176
rect 34789 21118 38535 21120
rect 34789 21115 34855 21118
rect 38469 21115 38535 21118
rect 19333 21040 20178 21042
rect 19333 20984 19338 21040
rect 19394 20984 20178 21040
rect 19333 20982 20178 20984
rect 21449 21042 21515 21045
rect 24577 21042 24643 21045
rect 21449 21040 24643 21042
rect 21449 20984 21454 21040
rect 21510 20984 24582 21040
rect 24638 20984 24643 21040
rect 21449 20982 24643 20984
rect 19333 20979 19399 20982
rect 21449 20979 21515 20982
rect 24577 20979 24643 20982
rect 25589 21042 25655 21045
rect 26325 21042 26391 21045
rect 25589 21040 26391 21042
rect 25589 20984 25594 21040
rect 25650 20984 26330 21040
rect 26386 20984 26391 21040
rect 25589 20982 26391 20984
rect 25589 20979 25655 20982
rect 26325 20979 26391 20982
rect 32765 21042 32831 21045
rect 35617 21042 35683 21045
rect 45001 21042 45067 21045
rect 32765 21040 45067 21042
rect 32765 20984 32770 21040
rect 32826 20984 35622 21040
rect 35678 20984 45006 21040
rect 45062 20984 45067 21040
rect 32765 20982 45067 20984
rect 32765 20979 32831 20982
rect 35617 20979 35683 20982
rect 45001 20979 45067 20982
rect 48497 21042 48563 21045
rect 50200 21042 51000 21072
rect 48497 21040 51000 21042
rect 48497 20984 48502 21040
rect 48558 20984 51000 21040
rect 48497 20982 51000 20984
rect 48497 20979 48563 20982
rect 50200 20952 51000 20982
rect 15101 20906 15167 20909
rect 17953 20906 18019 20909
rect 15101 20904 18019 20906
rect 15101 20848 15106 20904
rect 15162 20848 17958 20904
rect 18014 20848 18019 20904
rect 15101 20846 18019 20848
rect 15101 20843 15167 20846
rect 17953 20843 18019 20846
rect 22829 20906 22895 20909
rect 29729 20906 29795 20909
rect 22829 20904 29795 20906
rect 22829 20848 22834 20904
rect 22890 20848 29734 20904
rect 29790 20848 29795 20904
rect 22829 20846 29795 20848
rect 22829 20843 22895 20846
rect 29729 20843 29795 20846
rect 32121 20906 32187 20909
rect 33041 20906 33107 20909
rect 33869 20906 33935 20909
rect 32121 20904 33107 20906
rect 32121 20848 32126 20904
rect 32182 20848 33046 20904
rect 33102 20848 33107 20904
rect 32121 20846 33107 20848
rect 32121 20843 32187 20846
rect 33041 20843 33107 20846
rect 33734 20904 33935 20906
rect 33734 20848 33874 20904
rect 33930 20848 33935 20904
rect 33734 20846 33935 20848
rect 0 20770 800 20800
rect 1301 20770 1367 20773
rect 0 20768 1367 20770
rect 0 20712 1306 20768
rect 1362 20712 1367 20768
rect 0 20710 1367 20712
rect 0 20680 800 20710
rect 1301 20707 1367 20710
rect 12709 20770 12775 20773
rect 16389 20770 16455 20773
rect 12709 20768 16455 20770
rect 12709 20712 12714 20768
rect 12770 20712 16394 20768
rect 16450 20712 16455 20768
rect 12709 20710 16455 20712
rect 12709 20707 12775 20710
rect 16389 20707 16455 20710
rect 19609 20770 19675 20773
rect 20345 20770 20411 20773
rect 23657 20770 23723 20773
rect 19609 20768 23723 20770
rect 19609 20712 19614 20768
rect 19670 20712 20350 20768
rect 20406 20712 23662 20768
rect 23718 20712 23723 20768
rect 19609 20710 23723 20712
rect 19609 20707 19675 20710
rect 20345 20707 20411 20710
rect 23657 20707 23723 20710
rect 28349 20770 28415 20773
rect 30557 20770 30623 20773
rect 28349 20768 30623 20770
rect 28349 20712 28354 20768
rect 28410 20712 30562 20768
rect 30618 20712 30623 20768
rect 28349 20710 30623 20712
rect 28349 20707 28415 20710
rect 30557 20707 30623 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 17125 20634 17191 20637
rect 10182 20632 17191 20634
rect 10182 20576 17130 20632
rect 17186 20576 17191 20632
rect 10182 20574 17191 20576
rect 7833 20498 7899 20501
rect 10182 20498 10242 20574
rect 17125 20571 17191 20574
rect 22001 20634 22067 20637
rect 23841 20634 23907 20637
rect 27797 20634 27863 20637
rect 22001 20632 27863 20634
rect 22001 20576 22006 20632
rect 22062 20576 23846 20632
rect 23902 20576 27802 20632
rect 27858 20576 27863 20632
rect 22001 20574 27863 20576
rect 22001 20571 22067 20574
rect 23841 20571 23907 20574
rect 27797 20571 27863 20574
rect 31385 20634 31451 20637
rect 33734 20634 33794 20846
rect 33869 20843 33935 20846
rect 34973 20906 35039 20909
rect 45737 20906 45803 20909
rect 49233 20906 49299 20909
rect 34973 20904 45803 20906
rect 34973 20848 34978 20904
rect 35034 20848 45742 20904
rect 45798 20848 45803 20904
rect 34973 20846 45803 20848
rect 34973 20843 35039 20846
rect 45737 20843 45803 20846
rect 46982 20904 49299 20906
rect 46982 20848 49238 20904
rect 49294 20848 49299 20904
rect 46982 20846 49299 20848
rect 40677 20770 40743 20773
rect 42333 20770 42399 20773
rect 40677 20768 42399 20770
rect 40677 20712 40682 20768
rect 40738 20712 42338 20768
rect 42394 20712 42399 20768
rect 40677 20710 42399 20712
rect 40677 20707 40743 20710
rect 42333 20707 42399 20710
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 31385 20632 33794 20634
rect 31385 20576 31390 20632
rect 31446 20576 33794 20632
rect 31385 20574 33794 20576
rect 42609 20634 42675 20637
rect 46982 20634 47042 20846
rect 49233 20843 49299 20846
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 42609 20632 47042 20634
rect 42609 20576 42614 20632
rect 42670 20576 47042 20632
rect 42609 20574 47042 20576
rect 49049 20634 49115 20637
rect 50200 20634 51000 20664
rect 49049 20632 51000 20634
rect 49049 20576 49054 20632
rect 49110 20576 51000 20632
rect 49049 20574 51000 20576
rect 31385 20571 31451 20574
rect 42609 20571 42675 20574
rect 49049 20571 49115 20574
rect 50200 20544 51000 20574
rect 7833 20496 10242 20498
rect 7833 20440 7838 20496
rect 7894 20440 10242 20496
rect 7833 20438 10242 20440
rect 11697 20498 11763 20501
rect 16113 20498 16179 20501
rect 28809 20498 28875 20501
rect 11697 20496 28875 20498
rect 11697 20440 11702 20496
rect 11758 20440 16118 20496
rect 16174 20440 28814 20496
rect 28870 20440 28875 20496
rect 11697 20438 28875 20440
rect 7833 20435 7899 20438
rect 11697 20435 11763 20438
rect 16113 20435 16179 20438
rect 28809 20435 28875 20438
rect 28993 20498 29059 20501
rect 35065 20498 35131 20501
rect 28993 20496 35131 20498
rect 28993 20440 28998 20496
rect 29054 20440 35070 20496
rect 35126 20440 35131 20496
rect 28993 20438 35131 20440
rect 28993 20435 29059 20438
rect 35065 20435 35131 20438
rect 36261 20498 36327 20501
rect 38837 20498 38903 20501
rect 36261 20496 38903 20498
rect 36261 20440 36266 20496
rect 36322 20440 38842 20496
rect 38898 20440 38903 20496
rect 36261 20438 38903 20440
rect 36261 20435 36327 20438
rect 38837 20435 38903 20438
rect 40309 20498 40375 20501
rect 43253 20498 43319 20501
rect 40309 20496 43319 20498
rect 40309 20440 40314 20496
rect 40370 20440 43258 20496
rect 43314 20440 43319 20496
rect 40309 20438 43319 20440
rect 40309 20435 40375 20438
rect 43253 20435 43319 20438
rect 0 20362 800 20392
rect 3877 20362 3943 20365
rect 0 20360 3943 20362
rect 0 20304 3882 20360
rect 3938 20304 3943 20360
rect 0 20302 3943 20304
rect 0 20272 800 20302
rect 3877 20299 3943 20302
rect 12065 20362 12131 20365
rect 21449 20362 21515 20365
rect 12065 20360 21515 20362
rect 12065 20304 12070 20360
rect 12126 20304 21454 20360
rect 21510 20304 21515 20360
rect 12065 20302 21515 20304
rect 12065 20299 12131 20302
rect 21449 20299 21515 20302
rect 27337 20362 27403 20365
rect 34329 20362 34395 20365
rect 27337 20360 34395 20362
rect 27337 20304 27342 20360
rect 27398 20304 34334 20360
rect 34390 20304 34395 20360
rect 27337 20302 34395 20304
rect 27337 20299 27403 20302
rect 34329 20299 34395 20302
rect 37273 20362 37339 20365
rect 44541 20362 44607 20365
rect 37273 20360 44607 20362
rect 37273 20304 37278 20360
rect 37334 20304 44546 20360
rect 44602 20304 44607 20360
rect 37273 20302 44607 20304
rect 37273 20299 37339 20302
rect 44541 20299 44607 20302
rect 30557 20226 30623 20229
rect 31201 20226 31267 20229
rect 30557 20224 31267 20226
rect 30557 20168 30562 20224
rect 30618 20168 31206 20224
rect 31262 20168 31267 20224
rect 30557 20166 31267 20168
rect 30557 20163 30623 20166
rect 31201 20163 31267 20166
rect 36629 20226 36695 20229
rect 40953 20226 41019 20229
rect 36629 20224 41019 20226
rect 36629 20168 36634 20224
rect 36690 20168 40958 20224
rect 41014 20168 41019 20224
rect 36629 20166 41019 20168
rect 36629 20163 36695 20166
rect 40953 20163 41019 20166
rect 48589 20226 48655 20229
rect 50200 20226 51000 20256
rect 48589 20224 51000 20226
rect 48589 20168 48594 20224
rect 48650 20168 51000 20224
rect 48589 20166 51000 20168
rect 48589 20163 48655 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 50200 20136 51000 20166
rect 42946 20095 43262 20096
rect 15745 20090 15811 20093
rect 19701 20090 19767 20093
rect 24669 20090 24735 20093
rect 25405 20090 25471 20093
rect 31385 20090 31451 20093
rect 15745 20088 22110 20090
rect 15745 20032 15750 20088
rect 15806 20032 19706 20088
rect 19762 20032 22110 20088
rect 15745 20030 22110 20032
rect 15745 20027 15811 20030
rect 19701 20027 19767 20030
rect 0 19954 800 19984
rect 1393 19954 1459 19957
rect 0 19952 1459 19954
rect 0 19896 1398 19952
rect 1454 19896 1459 19952
rect 0 19894 1459 19896
rect 0 19864 800 19894
rect 1393 19891 1459 19894
rect 1761 19954 1827 19957
rect 16205 19954 16271 19957
rect 1761 19952 16271 19954
rect 1761 19896 1766 19952
rect 1822 19896 16210 19952
rect 16266 19896 16271 19952
rect 1761 19894 16271 19896
rect 22050 19954 22110 20030
rect 23430 20088 31451 20090
rect 23430 20032 24674 20088
rect 24730 20032 25410 20088
rect 25466 20032 31390 20088
rect 31446 20032 31451 20088
rect 23430 20030 31451 20032
rect 23430 19954 23490 20030
rect 24669 20027 24735 20030
rect 25405 20027 25471 20030
rect 31385 20027 31451 20030
rect 33869 20090 33935 20093
rect 35617 20090 35683 20093
rect 39849 20090 39915 20093
rect 33869 20088 35683 20090
rect 33869 20032 33874 20088
rect 33930 20032 35622 20088
rect 35678 20032 35683 20088
rect 33869 20030 35683 20032
rect 33869 20027 33935 20030
rect 35617 20027 35683 20030
rect 35758 20088 39915 20090
rect 35758 20032 39854 20088
rect 39910 20032 39915 20088
rect 35758 20030 39915 20032
rect 22050 19894 23490 19954
rect 1761 19891 1827 19894
rect 16205 19891 16271 19894
rect 30046 19892 30052 19956
rect 30116 19954 30122 19956
rect 30189 19954 30255 19957
rect 30116 19952 30255 19954
rect 30116 19896 30194 19952
rect 30250 19896 30255 19952
rect 30116 19894 30255 19896
rect 30116 19892 30122 19894
rect 30189 19891 30255 19894
rect 30741 19954 30807 19957
rect 31150 19954 31156 19956
rect 30741 19952 31156 19954
rect 30741 19896 30746 19952
rect 30802 19896 31156 19952
rect 30741 19894 31156 19896
rect 30741 19891 30807 19894
rect 31150 19892 31156 19894
rect 31220 19954 31226 19956
rect 31293 19954 31359 19957
rect 35758 19954 35818 20030
rect 39849 20027 39915 20030
rect 31220 19952 31359 19954
rect 31220 19896 31298 19952
rect 31354 19896 31359 19952
rect 31220 19894 31359 19896
rect 31220 19892 31226 19894
rect 31293 19891 31359 19894
rect 31710 19894 35818 19954
rect 35893 19954 35959 19957
rect 45185 19954 45251 19957
rect 35893 19952 45251 19954
rect 35893 19896 35898 19952
rect 35954 19896 45190 19952
rect 45246 19896 45251 19952
rect 35893 19894 45251 19896
rect 1853 19818 1919 19821
rect 14641 19818 14707 19821
rect 24945 19818 25011 19821
rect 28942 19818 28948 19820
rect 1853 19816 12450 19818
rect 1853 19760 1858 19816
rect 1914 19760 12450 19816
rect 1853 19758 12450 19760
rect 1853 19755 1919 19758
rect 12390 19682 12450 19758
rect 14641 19816 25011 19818
rect 14641 19760 14646 19816
rect 14702 19760 24950 19816
rect 25006 19760 25011 19816
rect 14641 19758 25011 19760
rect 14641 19755 14707 19758
rect 24945 19755 25011 19758
rect 27662 19758 28948 19818
rect 16205 19682 16271 19685
rect 12390 19680 16271 19682
rect 12390 19624 16210 19680
rect 16266 19624 16271 19680
rect 12390 19622 16271 19624
rect 16205 19619 16271 19622
rect 24485 19682 24551 19685
rect 26233 19682 26299 19685
rect 27662 19682 27722 19758
rect 28942 19756 28948 19758
rect 29012 19756 29018 19820
rect 30281 19818 30347 19821
rect 31710 19818 31770 19894
rect 35893 19891 35959 19894
rect 45185 19891 45251 19894
rect 30281 19816 31770 19818
rect 30281 19760 30286 19816
rect 30342 19760 31770 19816
rect 30281 19758 31770 19760
rect 32673 19818 32739 19821
rect 34462 19818 34468 19820
rect 32673 19816 34468 19818
rect 32673 19760 32678 19816
rect 32734 19760 34468 19816
rect 32673 19758 34468 19760
rect 30281 19755 30347 19758
rect 32673 19755 32739 19758
rect 34462 19756 34468 19758
rect 34532 19756 34538 19820
rect 49049 19818 49115 19821
rect 50200 19818 51000 19848
rect 49049 19816 51000 19818
rect 49049 19760 49054 19816
rect 49110 19760 51000 19816
rect 49049 19758 51000 19760
rect 49049 19755 49115 19758
rect 50200 19728 51000 19758
rect 24485 19680 27722 19682
rect 24485 19624 24490 19680
rect 24546 19624 26238 19680
rect 26294 19624 27722 19680
rect 24485 19622 27722 19624
rect 30189 19682 30255 19685
rect 31845 19682 31911 19685
rect 35341 19684 35407 19685
rect 32806 19682 32812 19684
rect 30189 19680 32812 19682
rect 30189 19624 30194 19680
rect 30250 19624 31850 19680
rect 31906 19624 32812 19680
rect 30189 19622 32812 19624
rect 24485 19619 24551 19622
rect 26233 19619 26299 19622
rect 30189 19619 30255 19622
rect 31845 19619 31911 19622
rect 32806 19620 32812 19622
rect 32876 19620 32882 19684
rect 35341 19682 35388 19684
rect 35296 19680 35388 19682
rect 35296 19624 35346 19680
rect 35296 19622 35388 19624
rect 35341 19620 35388 19622
rect 35452 19620 35458 19684
rect 35341 19619 35407 19620
rect 7946 19616 8262 19617
rect 0 19546 800 19576
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 2681 19546 2747 19549
rect 0 19544 2747 19546
rect 0 19488 2686 19544
rect 2742 19488 2747 19544
rect 0 19486 2747 19488
rect 0 19456 800 19486
rect 2681 19483 2747 19486
rect 28809 19546 28875 19549
rect 30741 19546 30807 19549
rect 28809 19544 36554 19546
rect 28809 19488 28814 19544
rect 28870 19488 30746 19544
rect 30802 19488 36554 19544
rect 28809 19486 36554 19488
rect 28809 19483 28875 19486
rect 30741 19483 30807 19486
rect 6821 19410 6887 19413
rect 11789 19410 11855 19413
rect 18689 19410 18755 19413
rect 27061 19410 27127 19413
rect 6821 19408 27127 19410
rect 6821 19352 6826 19408
rect 6882 19352 11794 19408
rect 11850 19352 18694 19408
rect 18750 19352 27066 19408
rect 27122 19352 27127 19408
rect 6821 19350 27127 19352
rect 6821 19347 6887 19350
rect 11789 19347 11855 19350
rect 18689 19347 18755 19350
rect 27061 19347 27127 19350
rect 27245 19410 27311 19413
rect 32673 19410 32739 19413
rect 27245 19408 32739 19410
rect 27245 19352 27250 19408
rect 27306 19352 32678 19408
rect 32734 19352 32739 19408
rect 27245 19350 32739 19352
rect 36494 19410 36554 19486
rect 42793 19410 42859 19413
rect 36494 19408 42859 19410
rect 36494 19352 42798 19408
rect 42854 19352 42859 19408
rect 36494 19350 42859 19352
rect 27245 19347 27311 19350
rect 32673 19347 32739 19350
rect 42793 19347 42859 19350
rect 49325 19410 49391 19413
rect 50200 19410 51000 19440
rect 49325 19408 51000 19410
rect 49325 19352 49330 19408
rect 49386 19352 51000 19408
rect 49325 19350 51000 19352
rect 49325 19347 49391 19350
rect 50200 19320 51000 19350
rect 2957 19274 3023 19277
rect 1304 19272 3023 19274
rect 1304 19216 2962 19272
rect 3018 19216 3023 19272
rect 1304 19214 3023 19216
rect 0 19138 800 19168
rect 1304 19138 1364 19214
rect 2957 19211 3023 19214
rect 10041 19274 10107 19277
rect 18321 19274 18387 19277
rect 10041 19272 18387 19274
rect 10041 19216 10046 19272
rect 10102 19216 18326 19272
rect 18382 19216 18387 19272
rect 10041 19214 18387 19216
rect 10041 19211 10107 19214
rect 18321 19211 18387 19214
rect 22737 19274 22803 19277
rect 25681 19274 25747 19277
rect 22737 19272 25747 19274
rect 22737 19216 22742 19272
rect 22798 19216 25686 19272
rect 25742 19216 25747 19272
rect 22737 19214 25747 19216
rect 22737 19211 22803 19214
rect 25681 19211 25747 19214
rect 26233 19274 26299 19277
rect 33225 19274 33291 19277
rect 26233 19272 33291 19274
rect 26233 19216 26238 19272
rect 26294 19216 33230 19272
rect 33286 19216 33291 19272
rect 26233 19214 33291 19216
rect 26233 19211 26299 19214
rect 33225 19211 33291 19214
rect 33358 19212 33364 19276
rect 33428 19274 33434 19276
rect 33869 19274 33935 19277
rect 36905 19274 36971 19277
rect 33428 19272 36971 19274
rect 33428 19216 33874 19272
rect 33930 19216 36910 19272
rect 36966 19216 36971 19272
rect 33428 19214 36971 19216
rect 33428 19212 33434 19214
rect 33869 19211 33935 19214
rect 36905 19211 36971 19214
rect 40493 19274 40559 19277
rect 48313 19274 48379 19277
rect 40493 19272 48379 19274
rect 40493 19216 40498 19272
rect 40554 19216 48318 19272
rect 48374 19216 48379 19272
rect 40493 19214 48379 19216
rect 40493 19211 40559 19214
rect 48313 19211 48379 19214
rect 0 19078 1364 19138
rect 6637 19138 6703 19141
rect 10133 19138 10199 19141
rect 6637 19136 10199 19138
rect 6637 19080 6642 19136
rect 6698 19080 10138 19136
rect 10194 19080 10199 19136
rect 6637 19078 10199 19080
rect 0 19048 800 19078
rect 6637 19075 6703 19078
rect 10133 19075 10199 19078
rect 13629 19138 13695 19141
rect 17033 19138 17099 19141
rect 13629 19136 17099 19138
rect 13629 19080 13634 19136
rect 13690 19080 17038 19136
rect 17094 19080 17099 19136
rect 13629 19078 17099 19080
rect 13629 19075 13695 19078
rect 17033 19075 17099 19078
rect 23473 19138 23539 19141
rect 26693 19138 26759 19141
rect 31477 19138 31543 19141
rect 23473 19136 31543 19138
rect 23473 19080 23478 19136
rect 23534 19080 26698 19136
rect 26754 19080 31482 19136
rect 31538 19080 31543 19136
rect 23473 19078 31543 19080
rect 23473 19075 23539 19078
rect 26693 19075 26759 19078
rect 31477 19075 31543 19078
rect 35249 19138 35315 19141
rect 39481 19138 39547 19141
rect 35249 19136 39547 19138
rect 35249 19080 35254 19136
rect 35310 19080 39486 19136
rect 39542 19080 39547 19136
rect 35249 19078 39547 19080
rect 35249 19075 35315 19078
rect 39481 19075 39547 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 6545 19002 6611 19005
rect 10593 19002 10659 19005
rect 6545 19000 10659 19002
rect 6545 18944 6550 19000
rect 6606 18944 10598 19000
rect 10654 18944 10659 19000
rect 6545 18942 10659 18944
rect 6545 18939 6611 18942
rect 10593 18939 10659 18942
rect 13721 19002 13787 19005
rect 16297 19002 16363 19005
rect 13721 19000 16363 19002
rect 13721 18944 13726 19000
rect 13782 18944 16302 19000
rect 16358 18944 16363 19000
rect 13721 18942 16363 18944
rect 13721 18939 13787 18942
rect 16297 18939 16363 18942
rect 16573 19002 16639 19005
rect 22001 19002 22067 19005
rect 16573 19000 22067 19002
rect 16573 18944 16578 19000
rect 16634 18944 22006 19000
rect 22062 18944 22067 19000
rect 16573 18942 22067 18944
rect 16573 18939 16639 18942
rect 22001 18939 22067 18942
rect 25957 19002 26023 19005
rect 27705 19002 27771 19005
rect 28073 19002 28139 19005
rect 25957 19000 28139 19002
rect 25957 18944 25962 19000
rect 26018 18944 27710 19000
rect 27766 18944 28078 19000
rect 28134 18944 28139 19000
rect 25957 18942 28139 18944
rect 25957 18939 26023 18942
rect 27705 18939 27771 18942
rect 28073 18939 28139 18942
rect 35249 19002 35315 19005
rect 37549 19002 37615 19005
rect 35249 19000 37615 19002
rect 35249 18944 35254 19000
rect 35310 18944 37554 19000
rect 37610 18944 37615 19000
rect 35249 18942 37615 18944
rect 35249 18939 35315 18942
rect 37549 18939 37615 18942
rect 37733 19002 37799 19005
rect 42149 19002 42215 19005
rect 37733 19000 42215 19002
rect 37733 18944 37738 19000
rect 37794 18944 42154 19000
rect 42210 18944 42215 19000
rect 37733 18942 42215 18944
rect 37733 18939 37799 18942
rect 42149 18939 42215 18942
rect 49141 19002 49207 19005
rect 50200 19002 51000 19032
rect 49141 19000 51000 19002
rect 49141 18944 49146 19000
rect 49202 18944 51000 19000
rect 49141 18942 51000 18944
rect 49141 18939 49207 18942
rect 50200 18912 51000 18942
rect 2773 18866 2839 18869
rect 1304 18864 2839 18866
rect 1304 18808 2778 18864
rect 2834 18808 2839 18864
rect 1304 18806 2839 18808
rect 0 18730 800 18760
rect 1304 18730 1364 18806
rect 2773 18803 2839 18806
rect 6085 18866 6151 18869
rect 7782 18866 7788 18868
rect 6085 18864 7788 18866
rect 6085 18808 6090 18864
rect 6146 18808 7788 18864
rect 6085 18806 7788 18808
rect 6085 18803 6151 18806
rect 7782 18804 7788 18806
rect 7852 18804 7858 18868
rect 9673 18866 9739 18869
rect 16757 18866 16823 18869
rect 9673 18864 16823 18866
rect 9673 18808 9678 18864
rect 9734 18808 16762 18864
rect 16818 18808 16823 18864
rect 9673 18806 16823 18808
rect 9673 18803 9739 18806
rect 16757 18803 16823 18806
rect 26877 18866 26943 18869
rect 30373 18866 30439 18869
rect 33777 18866 33843 18869
rect 26877 18864 33843 18866
rect 26877 18808 26882 18864
rect 26938 18808 30378 18864
rect 30434 18808 33782 18864
rect 33838 18808 33843 18864
rect 26877 18806 33843 18808
rect 26877 18803 26943 18806
rect 30373 18803 30439 18806
rect 33777 18803 33843 18806
rect 33961 18866 34027 18869
rect 34789 18866 34855 18869
rect 35801 18866 35867 18869
rect 33961 18864 35867 18866
rect 33961 18808 33966 18864
rect 34022 18808 34794 18864
rect 34850 18808 35806 18864
rect 35862 18808 35867 18864
rect 33961 18806 35867 18808
rect 33961 18803 34027 18806
rect 34789 18803 34855 18806
rect 35801 18803 35867 18806
rect 38469 18866 38535 18869
rect 41965 18866 42031 18869
rect 38469 18864 42031 18866
rect 38469 18808 38474 18864
rect 38530 18808 41970 18864
rect 42026 18808 42031 18864
rect 38469 18806 42031 18808
rect 38469 18803 38535 18806
rect 41965 18803 42031 18806
rect 0 18670 1364 18730
rect 9213 18730 9279 18733
rect 19609 18730 19675 18733
rect 9213 18728 19675 18730
rect 9213 18672 9218 18728
rect 9274 18672 19614 18728
rect 19670 18672 19675 18728
rect 9213 18670 19675 18672
rect 0 18640 800 18670
rect 9213 18667 9279 18670
rect 19609 18667 19675 18670
rect 19885 18730 19951 18733
rect 39205 18730 39271 18733
rect 19885 18728 39271 18730
rect 19885 18672 19890 18728
rect 19946 18672 39210 18728
rect 39266 18672 39271 18728
rect 19885 18670 39271 18672
rect 19885 18667 19951 18670
rect 39205 18667 39271 18670
rect 31661 18594 31727 18597
rect 37733 18594 37799 18597
rect 31661 18592 37799 18594
rect 31661 18536 31666 18592
rect 31722 18536 37738 18592
rect 37794 18536 37799 18592
rect 31661 18534 37799 18536
rect 31661 18531 31727 18534
rect 37733 18531 37799 18534
rect 38469 18594 38535 18597
rect 42425 18594 42491 18597
rect 38469 18592 42491 18594
rect 38469 18536 38474 18592
rect 38530 18536 42430 18592
rect 42486 18536 42491 18592
rect 38469 18534 42491 18536
rect 38469 18531 38535 18534
rect 42425 18531 42491 18534
rect 48773 18594 48839 18597
rect 50200 18594 51000 18624
rect 48773 18592 51000 18594
rect 48773 18536 48778 18592
rect 48834 18536 51000 18592
rect 48773 18534 51000 18536
rect 48773 18531 48839 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 50200 18504 51000 18534
rect 47946 18463 48262 18464
rect 18505 18458 18571 18461
rect 25129 18458 25195 18461
rect 18505 18456 25195 18458
rect 18505 18400 18510 18456
rect 18566 18400 25134 18456
rect 25190 18400 25195 18456
rect 18505 18398 25195 18400
rect 18505 18395 18571 18398
rect 25129 18395 25195 18398
rect 29913 18458 29979 18461
rect 33409 18458 33475 18461
rect 29913 18456 33475 18458
rect 29913 18400 29918 18456
rect 29974 18400 33414 18456
rect 33470 18400 33475 18456
rect 29913 18398 33475 18400
rect 29913 18395 29979 18398
rect 33409 18395 33475 18398
rect 33593 18458 33659 18461
rect 33726 18458 33732 18460
rect 33593 18456 33732 18458
rect 33593 18400 33598 18456
rect 33654 18400 33732 18456
rect 33593 18398 33732 18400
rect 33593 18395 33659 18398
rect 33726 18396 33732 18398
rect 33796 18458 33802 18460
rect 36905 18458 36971 18461
rect 33796 18456 36971 18458
rect 33796 18400 36910 18456
rect 36966 18400 36971 18456
rect 33796 18398 36971 18400
rect 33796 18396 33802 18398
rect 36905 18395 36971 18398
rect 0 18322 800 18352
rect 2865 18322 2931 18325
rect 0 18320 2931 18322
rect 0 18264 2870 18320
rect 2926 18264 2931 18320
rect 0 18262 2931 18264
rect 0 18232 800 18262
rect 2865 18259 2931 18262
rect 4705 18322 4771 18325
rect 7281 18322 7347 18325
rect 4705 18320 7347 18322
rect 4705 18264 4710 18320
rect 4766 18264 7286 18320
rect 7342 18264 7347 18320
rect 4705 18262 7347 18264
rect 4705 18259 4771 18262
rect 7281 18259 7347 18262
rect 13537 18322 13603 18325
rect 25037 18322 25103 18325
rect 13537 18320 25103 18322
rect 13537 18264 13542 18320
rect 13598 18264 25042 18320
rect 25098 18264 25103 18320
rect 13537 18262 25103 18264
rect 13537 18259 13603 18262
rect 25037 18259 25103 18262
rect 33133 18322 33199 18325
rect 36905 18322 36971 18325
rect 33133 18320 36971 18322
rect 33133 18264 33138 18320
rect 33194 18264 36910 18320
rect 36966 18264 36971 18320
rect 33133 18262 36971 18264
rect 33133 18259 33199 18262
rect 36905 18259 36971 18262
rect 37917 18322 37983 18325
rect 38326 18322 38332 18324
rect 37917 18320 38332 18322
rect 37917 18264 37922 18320
rect 37978 18264 38332 18320
rect 37917 18262 38332 18264
rect 37917 18259 37983 18262
rect 38326 18260 38332 18262
rect 38396 18260 38402 18324
rect 9121 18186 9187 18189
rect 14365 18186 14431 18189
rect 16941 18186 17007 18189
rect 27337 18186 27403 18189
rect 33542 18186 33548 18188
rect 9121 18184 14290 18186
rect 9121 18128 9126 18184
rect 9182 18128 14290 18184
rect 9121 18126 14290 18128
rect 9121 18123 9187 18126
rect 14230 18050 14290 18126
rect 14365 18184 27403 18186
rect 14365 18128 14370 18184
rect 14426 18128 16946 18184
rect 17002 18128 27342 18184
rect 27398 18128 27403 18184
rect 14365 18126 27403 18128
rect 14365 18123 14431 18126
rect 16941 18123 17007 18126
rect 27337 18123 27403 18126
rect 31756 18126 33548 18186
rect 18505 18050 18571 18053
rect 19149 18050 19215 18053
rect 14230 18048 19215 18050
rect 14230 17992 18510 18048
rect 18566 17992 19154 18048
rect 19210 17992 19215 18048
rect 14230 17990 19215 17992
rect 18505 17987 18571 17990
rect 19149 17987 19215 17990
rect 2946 17984 3262 17985
rect 0 17914 800 17944
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 31756 17917 31816 18126
rect 33542 18124 33548 18126
rect 33612 18124 33618 18188
rect 37089 18186 37155 18189
rect 39205 18186 39271 18189
rect 37089 18184 39271 18186
rect 37089 18128 37094 18184
rect 37150 18128 39210 18184
rect 39266 18128 39271 18184
rect 37089 18126 39271 18128
rect 37089 18123 37155 18126
rect 39205 18123 39271 18126
rect 39481 18186 39547 18189
rect 41597 18186 41663 18189
rect 39481 18184 41663 18186
rect 39481 18128 39486 18184
rect 39542 18128 41602 18184
rect 41658 18128 41663 18184
rect 39481 18126 41663 18128
rect 39481 18123 39547 18126
rect 41597 18123 41663 18126
rect 49141 18186 49207 18189
rect 50200 18186 51000 18216
rect 49141 18184 51000 18186
rect 49141 18128 49146 18184
rect 49202 18128 51000 18184
rect 49141 18126 51000 18128
rect 49141 18123 49207 18126
rect 50200 18096 51000 18126
rect 33961 18050 34027 18053
rect 37917 18050 37983 18053
rect 33961 18048 37983 18050
rect 33961 17992 33966 18048
rect 34022 17992 37922 18048
rect 37978 17992 37983 18048
rect 33961 17990 37983 17992
rect 33961 17987 34027 17990
rect 37917 17987 37983 17990
rect 38285 18050 38351 18053
rect 42793 18050 42859 18053
rect 38285 18048 42859 18050
rect 38285 17992 38290 18048
rect 38346 17992 42798 18048
rect 42854 17992 42859 18048
rect 38285 17990 42859 17992
rect 38285 17987 38351 17990
rect 42793 17987 42859 17990
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 2681 17914 2747 17917
rect 0 17912 2747 17914
rect 0 17856 2686 17912
rect 2742 17856 2747 17912
rect 0 17854 2747 17856
rect 0 17824 800 17854
rect 2681 17851 2747 17854
rect 13353 17914 13419 17917
rect 15469 17914 15535 17917
rect 13353 17912 15535 17914
rect 13353 17856 13358 17912
rect 13414 17856 15474 17912
rect 15530 17856 15535 17912
rect 13353 17854 15535 17856
rect 13353 17851 13419 17854
rect 15469 17851 15535 17854
rect 31753 17912 31819 17917
rect 31753 17856 31758 17912
rect 31814 17856 31819 17912
rect 31753 17851 31819 17856
rect 34462 17852 34468 17916
rect 34532 17914 34538 17916
rect 41781 17914 41847 17917
rect 34532 17912 41847 17914
rect 34532 17856 41786 17912
rect 41842 17856 41847 17912
rect 34532 17854 41847 17856
rect 34532 17852 34538 17854
rect 41781 17851 41847 17854
rect 8569 17778 8635 17781
rect 26141 17778 26207 17781
rect 8569 17776 26207 17778
rect 8569 17720 8574 17776
rect 8630 17720 26146 17776
rect 26202 17720 26207 17776
rect 8569 17718 26207 17720
rect 8569 17715 8635 17718
rect 26141 17715 26207 17718
rect 30833 17778 30899 17781
rect 41045 17778 41111 17781
rect 30833 17776 41111 17778
rect 30833 17720 30838 17776
rect 30894 17720 41050 17776
rect 41106 17720 41111 17776
rect 30833 17718 41111 17720
rect 30833 17715 30899 17718
rect 41045 17715 41111 17718
rect 49049 17778 49115 17781
rect 50200 17778 51000 17808
rect 49049 17776 51000 17778
rect 49049 17720 49054 17776
rect 49110 17720 51000 17776
rect 49049 17718 51000 17720
rect 49049 17715 49115 17718
rect 50200 17688 51000 17718
rect 10133 17642 10199 17645
rect 14917 17642 14983 17645
rect 10133 17640 14983 17642
rect 10133 17584 10138 17640
rect 10194 17584 14922 17640
rect 14978 17584 14983 17640
rect 10133 17582 14983 17584
rect 10133 17579 10199 17582
rect 14917 17579 14983 17582
rect 20161 17642 20227 17645
rect 20897 17642 20963 17645
rect 28809 17642 28875 17645
rect 20161 17640 20963 17642
rect 20161 17584 20166 17640
rect 20222 17584 20902 17640
rect 20958 17584 20963 17640
rect 20161 17582 20963 17584
rect 20161 17579 20227 17582
rect 20897 17579 20963 17582
rect 27800 17640 28875 17642
rect 27800 17584 28814 17640
rect 28870 17584 28875 17640
rect 27800 17582 28875 17584
rect 0 17506 800 17536
rect 2773 17506 2839 17509
rect 0 17504 2839 17506
rect 0 17448 2778 17504
rect 2834 17448 2839 17504
rect 0 17446 2839 17448
rect 0 17416 800 17446
rect 2773 17443 2839 17446
rect 10225 17506 10291 17509
rect 15929 17506 15995 17509
rect 10225 17504 15995 17506
rect 10225 17448 10230 17504
rect 10286 17448 15934 17504
rect 15990 17448 15995 17504
rect 10225 17446 15995 17448
rect 10225 17443 10291 17446
rect 15929 17443 15995 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27800 17373 27860 17582
rect 28809 17579 28875 17582
rect 29085 17642 29151 17645
rect 49233 17642 49299 17645
rect 29085 17640 49299 17642
rect 29085 17584 29090 17640
rect 29146 17584 49238 17640
rect 49294 17584 49299 17640
rect 29085 17582 49299 17584
rect 29085 17579 29151 17582
rect 49233 17579 49299 17582
rect 28533 17506 28599 17509
rect 36721 17506 36787 17509
rect 28533 17504 36787 17506
rect 28533 17448 28538 17504
rect 28594 17448 36726 17504
rect 36782 17448 36787 17504
rect 28533 17446 36787 17448
rect 28533 17443 28599 17446
rect 36721 17443 36787 17446
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 10593 17370 10659 17373
rect 17401 17370 17467 17373
rect 10593 17368 17467 17370
rect 10593 17312 10598 17368
rect 10654 17312 17406 17368
rect 17462 17312 17467 17368
rect 10593 17310 17467 17312
rect 10593 17307 10659 17310
rect 17401 17307 17467 17310
rect 24209 17370 24275 17373
rect 27797 17370 27863 17373
rect 24209 17368 27863 17370
rect 24209 17312 24214 17368
rect 24270 17312 27802 17368
rect 27858 17312 27863 17368
rect 24209 17310 27863 17312
rect 24209 17307 24275 17310
rect 27797 17307 27863 17310
rect 28942 17308 28948 17372
rect 29012 17370 29018 17372
rect 29085 17370 29151 17373
rect 29012 17368 29151 17370
rect 29012 17312 29090 17368
rect 29146 17312 29151 17368
rect 29012 17310 29151 17312
rect 29012 17308 29018 17310
rect 29085 17307 29151 17310
rect 31017 17370 31083 17373
rect 31150 17370 31156 17372
rect 31017 17368 31156 17370
rect 31017 17312 31022 17368
rect 31078 17312 31156 17368
rect 31017 17310 31156 17312
rect 31017 17307 31083 17310
rect 31150 17308 31156 17310
rect 31220 17308 31226 17372
rect 38377 17370 38443 17373
rect 40217 17370 40283 17373
rect 38377 17368 40283 17370
rect 38377 17312 38382 17368
rect 38438 17312 40222 17368
rect 40278 17312 40283 17368
rect 38377 17310 40283 17312
rect 38377 17307 38443 17310
rect 40217 17307 40283 17310
rect 49049 17370 49115 17373
rect 50200 17370 51000 17400
rect 49049 17368 51000 17370
rect 49049 17312 49054 17368
rect 49110 17312 51000 17368
rect 49049 17310 51000 17312
rect 49049 17307 49115 17310
rect 50200 17280 51000 17310
rect 12157 17234 12223 17237
rect 17769 17234 17835 17237
rect 19793 17234 19859 17237
rect 12157 17232 19859 17234
rect 12157 17176 12162 17232
rect 12218 17176 17774 17232
rect 17830 17176 19798 17232
rect 19854 17176 19859 17232
rect 12157 17174 19859 17176
rect 12157 17171 12223 17174
rect 17769 17171 17835 17174
rect 19793 17171 19859 17174
rect 21173 17234 21239 17237
rect 27797 17234 27863 17237
rect 28073 17234 28139 17237
rect 21173 17232 28139 17234
rect 21173 17176 21178 17232
rect 21234 17176 27802 17232
rect 27858 17176 28078 17232
rect 28134 17176 28139 17232
rect 21173 17174 28139 17176
rect 21173 17171 21239 17174
rect 27797 17171 27863 17174
rect 28073 17171 28139 17174
rect 29913 17234 29979 17237
rect 46105 17234 46171 17237
rect 29913 17232 46171 17234
rect 29913 17176 29918 17232
rect 29974 17176 46110 17232
rect 46166 17176 46171 17232
rect 29913 17174 46171 17176
rect 29913 17171 29979 17174
rect 46105 17171 46171 17174
rect 0 17098 800 17128
rect 1209 17098 1275 17101
rect 0 17096 1275 17098
rect 0 17040 1214 17096
rect 1270 17040 1275 17096
rect 0 17038 1275 17040
rect 0 17008 800 17038
rect 1209 17035 1275 17038
rect 9397 17098 9463 17101
rect 14641 17098 14707 17101
rect 9397 17096 14707 17098
rect 9397 17040 9402 17096
rect 9458 17040 14646 17096
rect 14702 17040 14707 17096
rect 9397 17038 14707 17040
rect 9397 17035 9463 17038
rect 14641 17035 14707 17038
rect 16389 17098 16455 17101
rect 24301 17098 24367 17101
rect 25313 17098 25379 17101
rect 16389 17096 25379 17098
rect 16389 17040 16394 17096
rect 16450 17040 24306 17096
rect 24362 17040 25318 17096
rect 25374 17040 25379 17096
rect 16389 17038 25379 17040
rect 16389 17035 16455 17038
rect 24301 17035 24367 17038
rect 25313 17035 25379 17038
rect 27061 17098 27127 17101
rect 27981 17098 28047 17101
rect 27061 17096 28047 17098
rect 27061 17040 27066 17096
rect 27122 17040 27986 17096
rect 28042 17040 28047 17096
rect 27061 17038 28047 17040
rect 27061 17035 27127 17038
rect 27981 17035 28047 17038
rect 29085 17098 29151 17101
rect 29453 17098 29519 17101
rect 29085 17096 29519 17098
rect 29085 17040 29090 17096
rect 29146 17040 29458 17096
rect 29514 17040 29519 17096
rect 29085 17038 29519 17040
rect 29085 17035 29151 17038
rect 29453 17035 29519 17038
rect 38469 17098 38535 17101
rect 39849 17098 39915 17101
rect 38469 17096 39915 17098
rect 38469 17040 38474 17096
rect 38530 17040 39854 17096
rect 39910 17040 39915 17096
rect 38469 17038 39915 17040
rect 38469 17035 38535 17038
rect 39849 17035 39915 17038
rect 23933 16962 23999 16965
rect 27613 16962 27679 16965
rect 23933 16960 27679 16962
rect 23933 16904 23938 16960
rect 23994 16904 27618 16960
rect 27674 16904 27679 16960
rect 23933 16902 27679 16904
rect 23933 16899 23999 16902
rect 27613 16899 27679 16902
rect 48773 16962 48839 16965
rect 50200 16962 51000 16992
rect 48773 16960 51000 16962
rect 48773 16904 48778 16960
rect 48834 16904 51000 16960
rect 48773 16902 51000 16904
rect 48773 16899 48839 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 50200 16872 51000 16902
rect 42946 16831 43262 16832
rect 0 16690 800 16720
rect 1301 16690 1367 16693
rect 0 16688 1367 16690
rect 0 16632 1306 16688
rect 1362 16632 1367 16688
rect 0 16630 1367 16632
rect 0 16600 800 16630
rect 1301 16627 1367 16630
rect 10133 16690 10199 16693
rect 17125 16690 17191 16693
rect 10133 16688 17191 16690
rect 10133 16632 10138 16688
rect 10194 16632 17130 16688
rect 17186 16632 17191 16688
rect 10133 16630 17191 16632
rect 10133 16627 10199 16630
rect 17125 16627 17191 16630
rect 23841 16690 23907 16693
rect 27153 16690 27219 16693
rect 23841 16688 27219 16690
rect 23841 16632 23846 16688
rect 23902 16632 27158 16688
rect 27214 16632 27219 16688
rect 23841 16630 27219 16632
rect 23841 16627 23907 16630
rect 27153 16627 27219 16630
rect 36629 16690 36695 16693
rect 38837 16690 38903 16693
rect 36629 16688 38903 16690
rect 36629 16632 36634 16688
rect 36690 16632 38842 16688
rect 38898 16632 38903 16688
rect 36629 16630 38903 16632
rect 36629 16627 36695 16630
rect 38837 16627 38903 16630
rect 4797 16554 4863 16557
rect 15193 16554 15259 16557
rect 19425 16554 19491 16557
rect 4797 16552 15259 16554
rect 4797 16496 4802 16552
rect 4858 16496 15198 16552
rect 15254 16496 15259 16552
rect 4797 16494 15259 16496
rect 4797 16491 4863 16494
rect 15193 16491 15259 16494
rect 15886 16552 19491 16554
rect 15886 16496 19430 16552
rect 19486 16496 19491 16552
rect 15886 16494 19491 16496
rect 9305 16418 9371 16421
rect 15886 16418 15946 16494
rect 19425 16491 19491 16494
rect 31753 16554 31819 16557
rect 40677 16554 40743 16557
rect 31753 16552 40743 16554
rect 31753 16496 31758 16552
rect 31814 16496 40682 16552
rect 40738 16496 40743 16552
rect 31753 16494 40743 16496
rect 31753 16491 31819 16494
rect 40677 16491 40743 16494
rect 49233 16554 49299 16557
rect 50200 16554 51000 16584
rect 49233 16552 51000 16554
rect 49233 16496 49238 16552
rect 49294 16496 51000 16552
rect 49233 16494 51000 16496
rect 49233 16491 49299 16494
rect 50200 16464 51000 16494
rect 9305 16416 15946 16418
rect 9305 16360 9310 16416
rect 9366 16360 15946 16416
rect 9305 16358 15946 16360
rect 35801 16418 35867 16421
rect 36905 16418 36971 16421
rect 35801 16416 36971 16418
rect 35801 16360 35806 16416
rect 35862 16360 36910 16416
rect 36966 16360 36971 16416
rect 35801 16358 36971 16360
rect 9305 16355 9371 16358
rect 35801 16355 35867 16358
rect 36905 16355 36971 16358
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 1301 16282 1367 16285
rect 0 16280 1367 16282
rect 0 16224 1306 16280
rect 1362 16224 1367 16280
rect 0 16222 1367 16224
rect 0 16192 800 16222
rect 1301 16219 1367 16222
rect 9857 16282 9923 16285
rect 10593 16282 10659 16285
rect 15326 16282 15332 16284
rect 9857 16280 15332 16282
rect 9857 16224 9862 16280
rect 9918 16224 10598 16280
rect 10654 16224 15332 16280
rect 9857 16222 15332 16224
rect 9857 16219 9923 16222
rect 10593 16219 10659 16222
rect 15326 16220 15332 16222
rect 15396 16282 15402 16284
rect 16430 16282 16436 16284
rect 15396 16222 16436 16282
rect 15396 16220 15402 16222
rect 16430 16220 16436 16222
rect 16500 16220 16506 16284
rect 29729 16282 29795 16285
rect 31385 16282 31451 16285
rect 35065 16282 35131 16285
rect 29729 16280 31451 16282
rect 29729 16224 29734 16280
rect 29790 16224 31390 16280
rect 31446 16224 31451 16280
rect 29729 16222 31451 16224
rect 29729 16219 29795 16222
rect 31385 16219 31451 16222
rect 31710 16280 35131 16282
rect 31710 16224 35070 16280
rect 35126 16224 35131 16280
rect 31710 16222 35131 16224
rect 11053 16146 11119 16149
rect 17677 16146 17743 16149
rect 25129 16146 25195 16149
rect 11053 16144 17743 16146
rect 11053 16088 11058 16144
rect 11114 16088 17682 16144
rect 17738 16088 17743 16144
rect 11053 16086 17743 16088
rect 11053 16083 11119 16086
rect 17677 16083 17743 16086
rect 17910 16144 25195 16146
rect 17910 16088 25134 16144
rect 25190 16088 25195 16144
rect 17910 16086 25195 16088
rect 15929 16010 15995 16013
rect 17910 16010 17970 16086
rect 25129 16083 25195 16086
rect 27061 16146 27127 16149
rect 31710 16146 31770 16222
rect 35065 16219 35131 16222
rect 32857 16148 32923 16149
rect 27061 16144 31770 16146
rect 27061 16088 27066 16144
rect 27122 16088 31770 16144
rect 27061 16086 31770 16088
rect 27061 16083 27127 16086
rect 32806 16084 32812 16148
rect 32876 16146 32923 16148
rect 34789 16146 34855 16149
rect 32876 16144 34855 16146
rect 32918 16088 34794 16144
rect 34850 16088 34855 16144
rect 32876 16086 34855 16088
rect 32876 16084 32923 16086
rect 32857 16083 32923 16084
rect 34789 16083 34855 16086
rect 35065 16146 35131 16149
rect 37825 16146 37891 16149
rect 35065 16144 37891 16146
rect 35065 16088 35070 16144
rect 35126 16088 37830 16144
rect 37886 16088 37891 16144
rect 35065 16086 37891 16088
rect 35065 16083 35131 16086
rect 37825 16083 37891 16086
rect 49141 16146 49207 16149
rect 50200 16146 51000 16176
rect 49141 16144 51000 16146
rect 49141 16088 49146 16144
rect 49202 16088 51000 16144
rect 49141 16086 51000 16088
rect 49141 16083 49207 16086
rect 50200 16056 51000 16086
rect 24669 16010 24735 16013
rect 27429 16010 27495 16013
rect 15929 16008 17970 16010
rect 15929 15952 15934 16008
rect 15990 15952 17970 16008
rect 15929 15950 17970 15952
rect 22050 16008 27495 16010
rect 22050 15952 24674 16008
rect 24730 15952 27434 16008
rect 27490 15952 27495 16008
rect 22050 15950 27495 15952
rect 15929 15947 15995 15950
rect 0 15874 800 15904
rect 1301 15874 1367 15877
rect 0 15872 1367 15874
rect 0 15816 1306 15872
rect 1362 15816 1367 15872
rect 0 15814 1367 15816
rect 0 15784 800 15814
rect 1301 15811 1367 15814
rect 10593 15874 10659 15877
rect 12065 15874 12131 15877
rect 10593 15872 12131 15874
rect 10593 15816 10598 15872
rect 10654 15816 12070 15872
rect 12126 15816 12131 15872
rect 10593 15814 12131 15816
rect 10593 15811 10659 15814
rect 12065 15811 12131 15814
rect 16430 15812 16436 15876
rect 16500 15874 16506 15876
rect 22050 15874 22110 15950
rect 24669 15947 24735 15950
rect 27429 15947 27495 15950
rect 36813 16010 36879 16013
rect 39481 16010 39547 16013
rect 39757 16010 39823 16013
rect 36813 16008 39823 16010
rect 36813 15952 36818 16008
rect 36874 15952 39486 16008
rect 39542 15952 39762 16008
rect 39818 15952 39823 16008
rect 36813 15950 39823 15952
rect 36813 15947 36879 15950
rect 39481 15947 39547 15950
rect 39757 15947 39823 15950
rect 16500 15814 22110 15874
rect 30097 15874 30163 15877
rect 31109 15874 31175 15877
rect 30097 15872 31175 15874
rect 30097 15816 30102 15872
rect 30158 15816 31114 15872
rect 31170 15816 31175 15872
rect 30097 15814 31175 15816
rect 16500 15812 16506 15814
rect 30097 15811 30163 15814
rect 31109 15811 31175 15814
rect 35157 15874 35223 15877
rect 39665 15874 39731 15877
rect 35157 15872 39731 15874
rect 35157 15816 35162 15872
rect 35218 15816 39670 15872
rect 39726 15816 39731 15872
rect 35157 15814 39731 15816
rect 35157 15811 35223 15814
rect 39665 15811 39731 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 16297 15738 16363 15741
rect 18873 15738 18939 15741
rect 16297 15736 18939 15738
rect 16297 15680 16302 15736
rect 16358 15680 18878 15736
rect 18934 15680 18939 15736
rect 16297 15678 18939 15680
rect 16297 15675 16363 15678
rect 18873 15675 18939 15678
rect 19333 15738 19399 15741
rect 25129 15738 25195 15741
rect 32489 15738 32555 15741
rect 19333 15736 22754 15738
rect 19333 15680 19338 15736
rect 19394 15680 22754 15736
rect 19333 15678 22754 15680
rect 19333 15675 19399 15678
rect 14181 15602 14247 15605
rect 22369 15602 22435 15605
rect 14181 15600 22435 15602
rect 14181 15544 14186 15600
rect 14242 15544 22374 15600
rect 22430 15544 22435 15600
rect 14181 15542 22435 15544
rect 22694 15602 22754 15678
rect 25129 15736 32555 15738
rect 25129 15680 25134 15736
rect 25190 15680 32494 15736
rect 32550 15680 32555 15736
rect 25129 15678 32555 15680
rect 25129 15675 25195 15678
rect 32489 15675 32555 15678
rect 35341 15738 35407 15741
rect 40125 15738 40191 15741
rect 35341 15736 40191 15738
rect 35341 15680 35346 15736
rect 35402 15680 40130 15736
rect 40186 15680 40191 15736
rect 35341 15678 40191 15680
rect 35341 15675 35407 15678
rect 40125 15675 40191 15678
rect 49049 15738 49115 15741
rect 50200 15738 51000 15768
rect 49049 15736 51000 15738
rect 49049 15680 49054 15736
rect 49110 15680 51000 15736
rect 49049 15678 51000 15680
rect 49049 15675 49115 15678
rect 50200 15648 51000 15678
rect 24485 15602 24551 15605
rect 26233 15602 26299 15605
rect 26969 15602 27035 15605
rect 48313 15602 48379 15605
rect 22694 15600 24551 15602
rect 22694 15544 24490 15600
rect 24546 15544 24551 15600
rect 22694 15542 24551 15544
rect 14181 15539 14247 15542
rect 22369 15539 22435 15542
rect 24485 15539 24551 15542
rect 25270 15600 48379 15602
rect 25270 15544 26238 15600
rect 26294 15544 26974 15600
rect 27030 15544 48318 15600
rect 48374 15544 48379 15600
rect 25270 15542 48379 15544
rect 0 15466 800 15496
rect 1301 15466 1367 15469
rect 0 15464 1367 15466
rect 0 15408 1306 15464
rect 1362 15408 1367 15464
rect 0 15406 1367 15408
rect 0 15376 800 15406
rect 1301 15403 1367 15406
rect 9397 15466 9463 15469
rect 22829 15466 22895 15469
rect 25270 15466 25330 15542
rect 26233 15539 26299 15542
rect 26969 15539 27035 15542
rect 48313 15539 48379 15542
rect 9397 15464 25330 15466
rect 9397 15408 9402 15464
rect 9458 15408 22834 15464
rect 22890 15408 25330 15464
rect 9397 15406 25330 15408
rect 25405 15466 25471 15469
rect 49233 15466 49299 15469
rect 25405 15464 49299 15466
rect 25405 15408 25410 15464
rect 25466 15408 49238 15464
rect 49294 15408 49299 15464
rect 25405 15406 49299 15408
rect 9397 15403 9463 15406
rect 22829 15403 22895 15406
rect 25405 15403 25471 15406
rect 49233 15403 49299 15406
rect 25957 15330 26023 15333
rect 26969 15330 27035 15333
rect 25957 15328 27035 15330
rect 25957 15272 25962 15328
rect 26018 15272 26974 15328
rect 27030 15272 27035 15328
rect 25957 15270 27035 15272
rect 25957 15267 26023 15270
rect 26969 15267 27035 15270
rect 31017 15330 31083 15333
rect 31753 15330 31819 15333
rect 31017 15328 31819 15330
rect 31017 15272 31022 15328
rect 31078 15272 31758 15328
rect 31814 15272 31819 15328
rect 31017 15270 31819 15272
rect 31017 15267 31083 15270
rect 31753 15267 31819 15270
rect 38561 15330 38627 15333
rect 40861 15330 40927 15333
rect 38561 15328 40927 15330
rect 38561 15272 38566 15328
rect 38622 15272 40866 15328
rect 40922 15272 40927 15328
rect 38561 15270 40927 15272
rect 38561 15267 38627 15270
rect 40861 15267 40927 15270
rect 49325 15330 49391 15333
rect 50200 15330 51000 15360
rect 49325 15328 51000 15330
rect 49325 15272 49330 15328
rect 49386 15272 51000 15328
rect 49325 15270 51000 15272
rect 49325 15267 49391 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 50200 15240 51000 15270
rect 47946 15199 48262 15200
rect 11973 15194 12039 15197
rect 15929 15194 15995 15197
rect 11973 15192 15995 15194
rect 11973 15136 11978 15192
rect 12034 15136 15934 15192
rect 15990 15136 15995 15192
rect 11973 15134 15995 15136
rect 11973 15131 12039 15134
rect 15929 15131 15995 15134
rect 19517 15194 19583 15197
rect 23289 15194 23355 15197
rect 19517 15192 23355 15194
rect 19517 15136 19522 15192
rect 19578 15136 23294 15192
rect 23350 15136 23355 15192
rect 19517 15134 23355 15136
rect 19517 15131 19583 15134
rect 23289 15131 23355 15134
rect 33225 15194 33291 15197
rect 34053 15194 34119 15197
rect 34973 15194 35039 15197
rect 33225 15192 35039 15194
rect 33225 15136 33230 15192
rect 33286 15136 34058 15192
rect 34114 15136 34978 15192
rect 35034 15136 35039 15192
rect 33225 15134 35039 15136
rect 33225 15131 33291 15134
rect 34053 15131 34119 15134
rect 34973 15131 35039 15134
rect 0 15058 800 15088
rect 1301 15058 1367 15061
rect 0 15056 1367 15058
rect 0 15000 1306 15056
rect 1362 15000 1367 15056
rect 0 14998 1367 15000
rect 0 14968 800 14998
rect 1301 14995 1367 14998
rect 12065 15058 12131 15061
rect 27061 15058 27127 15061
rect 12065 15056 27127 15058
rect 12065 15000 12070 15056
rect 12126 15000 27066 15056
rect 27122 15000 27127 15056
rect 12065 14998 27127 15000
rect 12065 14995 12131 14998
rect 27061 14995 27127 14998
rect 27245 15058 27311 15061
rect 48497 15058 48563 15061
rect 27245 15056 48563 15058
rect 27245 15000 27250 15056
rect 27306 15000 48502 15056
rect 48558 15000 48563 15056
rect 27245 14998 48563 15000
rect 27245 14995 27311 14998
rect 48497 14995 48563 14998
rect 10961 14922 11027 14925
rect 14641 14922 14707 14925
rect 16757 14922 16823 14925
rect 10961 14920 14474 14922
rect 10961 14864 10966 14920
rect 11022 14864 14474 14920
rect 10961 14862 14474 14864
rect 10961 14859 11027 14862
rect 14414 14786 14474 14862
rect 14641 14920 16823 14922
rect 14641 14864 14646 14920
rect 14702 14864 16762 14920
rect 16818 14864 16823 14920
rect 14641 14862 16823 14864
rect 14641 14859 14707 14862
rect 16757 14859 16823 14862
rect 21633 14922 21699 14925
rect 48313 14922 48379 14925
rect 21633 14920 48379 14922
rect 21633 14864 21638 14920
rect 21694 14864 48318 14920
rect 48374 14864 48379 14920
rect 21633 14862 48379 14864
rect 21633 14859 21699 14862
rect 48313 14859 48379 14862
rect 49049 14922 49115 14925
rect 50200 14922 51000 14952
rect 49049 14920 51000 14922
rect 49049 14864 49054 14920
rect 49110 14864 51000 14920
rect 49049 14862 51000 14864
rect 49049 14859 49115 14862
rect 50200 14832 51000 14862
rect 18873 14786 18939 14789
rect 14414 14784 18939 14786
rect 14414 14728 18878 14784
rect 18934 14728 18939 14784
rect 14414 14726 18939 14728
rect 18873 14723 18939 14726
rect 25221 14786 25287 14789
rect 30741 14786 30807 14789
rect 25221 14784 30807 14786
rect 25221 14728 25226 14784
rect 25282 14728 30746 14784
rect 30802 14728 30807 14784
rect 25221 14726 30807 14728
rect 25221 14723 25287 14726
rect 30741 14723 30807 14726
rect 33685 14786 33751 14789
rect 34145 14786 34211 14789
rect 33685 14784 34211 14786
rect 33685 14728 33690 14784
rect 33746 14728 34150 14784
rect 34206 14728 34211 14784
rect 33685 14726 34211 14728
rect 33685 14723 33751 14726
rect 34145 14723 34211 14726
rect 37549 14786 37615 14789
rect 39849 14786 39915 14789
rect 37549 14784 39915 14786
rect 37549 14728 37554 14784
rect 37610 14728 39854 14784
rect 39910 14728 39915 14784
rect 37549 14726 39915 14728
rect 37549 14723 37615 14726
rect 39849 14723 39915 14726
rect 2946 14720 3262 14721
rect 0 14650 800 14680
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 1301 14650 1367 14653
rect 0 14648 1367 14650
rect 0 14592 1306 14648
rect 1362 14592 1367 14648
rect 0 14590 1367 14592
rect 0 14560 800 14590
rect 1301 14587 1367 14590
rect 14273 14514 14339 14517
rect 17677 14514 17743 14517
rect 14273 14512 17743 14514
rect 14273 14456 14278 14512
rect 14334 14456 17682 14512
rect 17738 14456 17743 14512
rect 14273 14454 17743 14456
rect 14273 14451 14339 14454
rect 17677 14451 17743 14454
rect 18597 14514 18663 14517
rect 33225 14514 33291 14517
rect 33358 14514 33364 14516
rect 18597 14512 33364 14514
rect 18597 14456 18602 14512
rect 18658 14456 33230 14512
rect 33286 14456 33364 14512
rect 18597 14454 33364 14456
rect 18597 14451 18663 14454
rect 33225 14451 33291 14454
rect 33358 14452 33364 14454
rect 33428 14452 33434 14516
rect 33501 14514 33567 14517
rect 39481 14514 39547 14517
rect 33501 14512 39547 14514
rect 33501 14456 33506 14512
rect 33562 14456 39486 14512
rect 39542 14456 39547 14512
rect 33501 14454 39547 14456
rect 33501 14451 33567 14454
rect 39481 14451 39547 14454
rect 49049 14514 49115 14517
rect 50200 14514 51000 14544
rect 49049 14512 51000 14514
rect 49049 14456 49054 14512
rect 49110 14456 51000 14512
rect 49049 14454 51000 14456
rect 49049 14451 49115 14454
rect 50200 14424 51000 14454
rect 13445 14378 13511 14381
rect 15285 14378 15351 14381
rect 13445 14376 15351 14378
rect 13445 14320 13450 14376
rect 13506 14320 15290 14376
rect 15346 14320 15351 14376
rect 13445 14318 15351 14320
rect 13445 14315 13511 14318
rect 15285 14315 15351 14318
rect 16205 14378 16271 14381
rect 16849 14378 16915 14381
rect 19057 14378 19123 14381
rect 49233 14378 49299 14381
rect 16205 14376 19123 14378
rect 16205 14320 16210 14376
rect 16266 14320 16854 14376
rect 16910 14320 19062 14376
rect 19118 14320 19123 14376
rect 16205 14318 19123 14320
rect 16205 14315 16271 14318
rect 16849 14315 16915 14318
rect 19057 14315 19123 14318
rect 22694 14376 49299 14378
rect 22694 14320 49238 14376
rect 49294 14320 49299 14376
rect 22694 14318 49299 14320
rect 0 14242 800 14272
rect 933 14242 999 14245
rect 0 14240 999 14242
rect 0 14184 938 14240
rect 994 14184 999 14240
rect 0 14182 999 14184
rect 0 14152 800 14182
rect 933 14179 999 14182
rect 10685 14242 10751 14245
rect 14917 14242 14983 14245
rect 15142 14242 15148 14244
rect 10685 14240 15148 14242
rect 10685 14184 10690 14240
rect 10746 14184 14922 14240
rect 14978 14184 15148 14240
rect 10685 14182 15148 14184
rect 10685 14179 10751 14182
rect 14917 14179 14983 14182
rect 15142 14180 15148 14182
rect 15212 14180 15218 14244
rect 17217 14242 17283 14245
rect 17769 14242 17835 14245
rect 17217 14240 17835 14242
rect 17217 14184 17222 14240
rect 17278 14184 17774 14240
rect 17830 14184 17835 14240
rect 17217 14182 17835 14184
rect 17217 14179 17283 14182
rect 17769 14179 17835 14182
rect 22461 14242 22527 14245
rect 22694 14242 22754 14318
rect 49233 14315 49299 14318
rect 29269 14244 29335 14245
rect 29269 14242 29316 14244
rect 22461 14240 22754 14242
rect 22461 14184 22466 14240
rect 22522 14184 22754 14240
rect 22461 14182 22754 14184
rect 29224 14240 29316 14242
rect 29224 14184 29274 14240
rect 29224 14182 29316 14184
rect 22461 14179 22527 14182
rect 29269 14180 29316 14182
rect 29380 14180 29386 14244
rect 31661 14242 31727 14245
rect 32213 14242 32279 14245
rect 32949 14242 33015 14245
rect 31661 14240 33015 14242
rect 31661 14184 31666 14240
rect 31722 14184 32218 14240
rect 32274 14184 32954 14240
rect 33010 14184 33015 14240
rect 31661 14182 33015 14184
rect 29269 14179 29335 14180
rect 31661 14179 31727 14182
rect 32213 14179 32279 14182
rect 32949 14179 33015 14182
rect 33317 14242 33383 14245
rect 34053 14242 34119 14245
rect 33317 14240 34119 14242
rect 33317 14184 33322 14240
rect 33378 14184 34058 14240
rect 34114 14184 34119 14240
rect 33317 14182 34119 14184
rect 33317 14179 33383 14182
rect 34053 14179 34119 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 9857 14106 9923 14109
rect 16573 14106 16639 14109
rect 9857 14104 16639 14106
rect 9857 14048 9862 14104
rect 9918 14048 16578 14104
rect 16634 14048 16639 14104
rect 9857 14046 16639 14048
rect 9857 14043 9923 14046
rect 16573 14043 16639 14046
rect 18873 14106 18939 14109
rect 25405 14106 25471 14109
rect 18873 14104 25471 14106
rect 18873 14048 18878 14104
rect 18934 14048 25410 14104
rect 25466 14048 25471 14104
rect 18873 14046 25471 14048
rect 18873 14043 18939 14046
rect 25405 14043 25471 14046
rect 49141 14106 49207 14109
rect 50200 14106 51000 14136
rect 49141 14104 51000 14106
rect 49141 14048 49146 14104
rect 49202 14048 51000 14104
rect 49141 14046 51000 14048
rect 49141 14043 49207 14046
rect 50200 14016 51000 14046
rect 10317 13970 10383 13973
rect 16113 13970 16179 13973
rect 10317 13968 16179 13970
rect 10317 13912 10322 13968
rect 10378 13912 16118 13968
rect 16174 13912 16179 13968
rect 10317 13910 16179 13912
rect 10317 13907 10383 13910
rect 16113 13907 16179 13910
rect 16389 13970 16455 13973
rect 17585 13970 17651 13973
rect 30189 13970 30255 13973
rect 37273 13970 37339 13973
rect 40953 13970 41019 13973
rect 16389 13968 30255 13970
rect 16389 13912 16394 13968
rect 16450 13912 17590 13968
rect 17646 13912 30194 13968
rect 30250 13912 30255 13968
rect 16389 13910 30255 13912
rect 16389 13907 16455 13910
rect 17585 13907 17651 13910
rect 30189 13907 30255 13910
rect 31710 13910 37106 13970
rect 0 13834 800 13864
rect 2773 13834 2839 13837
rect 0 13832 2839 13834
rect 0 13776 2778 13832
rect 2834 13776 2839 13832
rect 0 13774 2839 13776
rect 0 13744 800 13774
rect 2773 13771 2839 13774
rect 10225 13834 10291 13837
rect 12617 13834 12683 13837
rect 17401 13834 17467 13837
rect 18781 13834 18847 13837
rect 31109 13834 31175 13837
rect 31710 13834 31770 13910
rect 37046 13834 37106 13910
rect 37273 13968 41019 13970
rect 37273 13912 37278 13968
rect 37334 13912 40958 13968
rect 41014 13912 41019 13968
rect 37273 13910 41019 13912
rect 37273 13907 37339 13910
rect 40953 13907 41019 13910
rect 37917 13834 37983 13837
rect 41321 13834 41387 13837
rect 10225 13832 12683 13834
rect 10225 13776 10230 13832
rect 10286 13776 12622 13832
rect 12678 13776 12683 13832
rect 10225 13774 12683 13776
rect 10225 13771 10291 13774
rect 12617 13771 12683 13774
rect 12758 13774 13554 13834
rect 9949 13698 10015 13701
rect 12758 13698 12818 13774
rect 9949 13696 12818 13698
rect 9949 13640 9954 13696
rect 10010 13640 12818 13696
rect 9949 13638 12818 13640
rect 13494 13698 13554 13774
rect 17401 13832 31770 13834
rect 17401 13776 17406 13832
rect 17462 13776 18786 13832
rect 18842 13776 31114 13832
rect 31170 13776 31770 13832
rect 17401 13774 31770 13776
rect 32814 13774 33426 13834
rect 37046 13832 41387 13834
rect 37046 13776 37922 13832
rect 37978 13776 41326 13832
rect 41382 13776 41387 13832
rect 37046 13774 41387 13776
rect 17401 13771 17467 13774
rect 18781 13771 18847 13774
rect 31109 13771 31175 13774
rect 19149 13698 19215 13701
rect 13494 13696 19215 13698
rect 13494 13640 19154 13696
rect 19210 13640 19215 13696
rect 13494 13638 19215 13640
rect 9949 13635 10015 13638
rect 19149 13635 19215 13638
rect 28717 13698 28783 13701
rect 32814 13698 32874 13774
rect 28717 13696 32874 13698
rect 28717 13640 28722 13696
rect 28778 13640 32874 13696
rect 28717 13638 32874 13640
rect 33366 13698 33426 13774
rect 37917 13771 37983 13774
rect 41321 13771 41387 13774
rect 42750 13774 43546 13834
rect 39849 13698 39915 13701
rect 33366 13696 39915 13698
rect 33366 13640 39854 13696
rect 39910 13640 39915 13696
rect 33366 13638 39915 13640
rect 28717 13635 28783 13638
rect 39849 13635 39915 13638
rect 40033 13698 40099 13701
rect 42750 13698 42810 13774
rect 40033 13696 42810 13698
rect 40033 13640 40038 13696
rect 40094 13640 42810 13696
rect 40033 13638 42810 13640
rect 43486 13698 43546 13774
rect 45277 13698 45343 13701
rect 43486 13696 45343 13698
rect 43486 13640 45282 13696
rect 45338 13640 45343 13696
rect 43486 13638 45343 13640
rect 40033 13635 40099 13638
rect 45277 13635 45343 13638
rect 48221 13698 48287 13701
rect 50200 13698 51000 13728
rect 48221 13696 51000 13698
rect 48221 13640 48226 13696
rect 48282 13640 51000 13696
rect 48221 13638 51000 13640
rect 48221 13635 48287 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 50200 13608 51000 13638
rect 42946 13567 43262 13568
rect 15101 13562 15167 13565
rect 17309 13562 17375 13565
rect 40677 13562 40743 13565
rect 15101 13560 17375 13562
rect 15101 13504 15106 13560
rect 15162 13504 17314 13560
rect 17370 13504 17375 13560
rect 15101 13502 17375 13504
rect 15101 13499 15167 13502
rect 17309 13499 17375 13502
rect 33366 13560 40743 13562
rect 33366 13504 40682 13560
rect 40738 13504 40743 13560
rect 33366 13502 40743 13504
rect 0 13426 800 13456
rect 1761 13426 1827 13429
rect 14457 13426 14523 13429
rect 0 13366 1594 13426
rect 0 13336 800 13366
rect 1534 13290 1594 13366
rect 1761 13424 14523 13426
rect 1761 13368 1766 13424
rect 1822 13368 14462 13424
rect 14518 13368 14523 13424
rect 1761 13366 14523 13368
rect 1761 13363 1827 13366
rect 14457 13363 14523 13366
rect 15009 13426 15075 13429
rect 23105 13426 23171 13429
rect 15009 13424 23171 13426
rect 15009 13368 15014 13424
rect 15070 13368 23110 13424
rect 23166 13368 23171 13424
rect 15009 13366 23171 13368
rect 15009 13363 15075 13366
rect 23105 13363 23171 13366
rect 32581 13426 32647 13429
rect 33366 13426 33426 13502
rect 40677 13499 40743 13502
rect 32581 13424 33426 13426
rect 32581 13368 32586 13424
rect 32642 13368 33426 13424
rect 32581 13366 33426 13368
rect 34421 13426 34487 13429
rect 45553 13426 45619 13429
rect 34421 13424 45619 13426
rect 34421 13368 34426 13424
rect 34482 13368 45558 13424
rect 45614 13368 45619 13424
rect 34421 13366 45619 13368
rect 32581 13363 32647 13366
rect 34421 13363 34487 13366
rect 45553 13363 45619 13366
rect 3509 13290 3575 13293
rect 1534 13288 3575 13290
rect 1534 13232 3514 13288
rect 3570 13232 3575 13288
rect 1534 13230 3575 13232
rect 3509 13227 3575 13230
rect 9949 13290 10015 13293
rect 14365 13290 14431 13293
rect 24577 13290 24643 13293
rect 9949 13288 24643 13290
rect 9949 13232 9954 13288
rect 10010 13232 14370 13288
rect 14426 13232 24582 13288
rect 24638 13232 24643 13288
rect 9949 13230 24643 13232
rect 9949 13227 10015 13230
rect 14365 13227 14431 13230
rect 24577 13227 24643 13230
rect 31477 13290 31543 13293
rect 38745 13290 38811 13293
rect 31477 13288 38811 13290
rect 31477 13232 31482 13288
rect 31538 13232 38750 13288
rect 38806 13232 38811 13288
rect 31477 13230 38811 13232
rect 31477 13227 31543 13230
rect 38745 13227 38811 13230
rect 49141 13290 49207 13293
rect 50200 13290 51000 13320
rect 49141 13288 51000 13290
rect 49141 13232 49146 13288
rect 49202 13232 51000 13288
rect 49141 13230 51000 13232
rect 49141 13227 49207 13230
rect 50200 13200 51000 13230
rect 10317 13154 10383 13157
rect 14825 13154 14891 13157
rect 15377 13154 15443 13157
rect 10317 13152 15443 13154
rect 10317 13096 10322 13152
rect 10378 13096 14830 13152
rect 14886 13096 15382 13152
rect 15438 13096 15443 13152
rect 10317 13094 15443 13096
rect 10317 13091 10383 13094
rect 14825 13091 14891 13094
rect 15377 13091 15443 13094
rect 15653 13154 15719 13157
rect 17125 13154 17191 13157
rect 21265 13156 21331 13157
rect 21214 13154 21220 13156
rect 15653 13152 17191 13154
rect 15653 13096 15658 13152
rect 15714 13096 17130 13152
rect 17186 13096 17191 13152
rect 15653 13094 17191 13096
rect 21174 13094 21220 13154
rect 21284 13152 21331 13156
rect 21326 13096 21331 13152
rect 15653 13091 15719 13094
rect 17125 13091 17191 13094
rect 21214 13092 21220 13094
rect 21284 13092 21331 13096
rect 21265 13091 21331 13092
rect 21633 13154 21699 13157
rect 27613 13154 27679 13157
rect 21633 13152 27679 13154
rect 21633 13096 21638 13152
rect 21694 13096 27618 13152
rect 27674 13096 27679 13152
rect 21633 13094 27679 13096
rect 21633 13091 21699 13094
rect 27613 13091 27679 13094
rect 7946 13088 8262 13089
rect 0 13018 800 13048
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 1209 13018 1275 13021
rect 0 13016 1275 13018
rect 0 12960 1214 13016
rect 1270 12960 1275 13016
rect 0 12958 1275 12960
rect 0 12928 800 12958
rect 1209 12955 1275 12958
rect 16021 12882 16087 12885
rect 24485 12882 24551 12885
rect 16021 12880 24551 12882
rect 16021 12824 16026 12880
rect 16082 12824 24490 12880
rect 24546 12824 24551 12880
rect 16021 12822 24551 12824
rect 16021 12819 16087 12822
rect 24485 12819 24551 12822
rect 26141 12882 26207 12885
rect 30005 12882 30071 12885
rect 26141 12880 30071 12882
rect 26141 12824 26146 12880
rect 26202 12824 30010 12880
rect 30066 12824 30071 12880
rect 26141 12822 30071 12824
rect 26141 12819 26207 12822
rect 30005 12819 30071 12822
rect 31845 12882 31911 12885
rect 39297 12882 39363 12885
rect 31845 12880 39363 12882
rect 31845 12824 31850 12880
rect 31906 12824 39302 12880
rect 39358 12824 39363 12880
rect 31845 12822 39363 12824
rect 31845 12819 31911 12822
rect 39297 12819 39363 12822
rect 49141 12882 49207 12885
rect 50200 12882 51000 12912
rect 49141 12880 51000 12882
rect 49141 12824 49146 12880
rect 49202 12824 51000 12880
rect 49141 12822 51000 12824
rect 49141 12819 49207 12822
rect 50200 12792 51000 12822
rect 9213 12746 9279 12749
rect 20621 12746 20687 12749
rect 9213 12744 20687 12746
rect 9213 12688 9218 12744
rect 9274 12688 20626 12744
rect 20682 12688 20687 12744
rect 9213 12686 20687 12688
rect 9213 12683 9279 12686
rect 20621 12683 20687 12686
rect 31569 12746 31635 12749
rect 34697 12746 34763 12749
rect 31569 12744 34763 12746
rect 31569 12688 31574 12744
rect 31630 12688 34702 12744
rect 34758 12688 34763 12744
rect 31569 12686 34763 12688
rect 31569 12683 31635 12686
rect 34697 12683 34763 12686
rect 36486 12684 36492 12748
rect 36556 12746 36562 12748
rect 40033 12746 40099 12749
rect 36556 12744 40099 12746
rect 36556 12688 40038 12744
rect 40094 12688 40099 12744
rect 36556 12686 40099 12688
rect 36556 12684 36562 12686
rect 40033 12683 40099 12686
rect 0 12610 800 12640
rect 1301 12610 1367 12613
rect 0 12608 1367 12610
rect 0 12552 1306 12608
rect 1362 12552 1367 12608
rect 0 12550 1367 12552
rect 0 12520 800 12550
rect 1301 12547 1367 12550
rect 16113 12610 16179 12613
rect 20253 12610 20319 12613
rect 21541 12610 21607 12613
rect 16113 12608 21607 12610
rect 16113 12552 16118 12608
rect 16174 12552 20258 12608
rect 20314 12552 21546 12608
rect 21602 12552 21607 12608
rect 16113 12550 21607 12552
rect 16113 12547 16179 12550
rect 20253 12547 20319 12550
rect 21541 12547 21607 12550
rect 34145 12610 34211 12613
rect 38745 12610 38811 12613
rect 34145 12608 38811 12610
rect 34145 12552 34150 12608
rect 34206 12552 38750 12608
rect 38806 12552 38811 12608
rect 34145 12550 38811 12552
rect 34145 12547 34211 12550
rect 38745 12547 38811 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 36445 12474 36511 12477
rect 38561 12474 38627 12477
rect 36445 12472 38627 12474
rect 36445 12416 36450 12472
rect 36506 12416 38566 12472
rect 38622 12416 38627 12472
rect 36445 12414 38627 12416
rect 36445 12411 36511 12414
rect 38561 12411 38627 12414
rect 49141 12474 49207 12477
rect 50200 12474 51000 12504
rect 49141 12472 51000 12474
rect 49141 12416 49146 12472
rect 49202 12416 51000 12472
rect 49141 12414 51000 12416
rect 49141 12411 49207 12414
rect 50200 12384 51000 12414
rect 26233 12338 26299 12341
rect 29453 12338 29519 12341
rect 26233 12336 29519 12338
rect 26233 12280 26238 12336
rect 26294 12280 29458 12336
rect 29514 12280 29519 12336
rect 26233 12278 29519 12280
rect 26233 12275 26299 12278
rect 29453 12275 29519 12278
rect 31017 12338 31083 12341
rect 37549 12338 37615 12341
rect 31017 12336 37615 12338
rect 31017 12280 31022 12336
rect 31078 12280 37554 12336
rect 37610 12280 37615 12336
rect 31017 12278 37615 12280
rect 31017 12275 31083 12278
rect 37549 12275 37615 12278
rect 0 12202 800 12232
rect 1209 12202 1275 12205
rect 0 12200 1275 12202
rect 0 12144 1214 12200
rect 1270 12144 1275 12200
rect 0 12142 1275 12144
rect 0 12112 800 12142
rect 1209 12139 1275 12142
rect 13905 12202 13971 12205
rect 16021 12202 16087 12205
rect 13905 12200 16087 12202
rect 13905 12144 13910 12200
rect 13966 12144 16026 12200
rect 16082 12144 16087 12200
rect 13905 12142 16087 12144
rect 13905 12139 13971 12142
rect 16021 12139 16087 12142
rect 17217 12202 17283 12205
rect 23749 12202 23815 12205
rect 17217 12200 23815 12202
rect 17217 12144 17222 12200
rect 17278 12144 23754 12200
rect 23810 12144 23815 12200
rect 17217 12142 23815 12144
rect 17217 12139 17283 12142
rect 23749 12139 23815 12142
rect 31753 12202 31819 12205
rect 48681 12202 48747 12205
rect 31753 12200 48747 12202
rect 31753 12144 31758 12200
rect 31814 12144 48686 12200
rect 48742 12144 48747 12200
rect 31753 12142 48747 12144
rect 31753 12139 31819 12142
rect 48681 12139 48747 12142
rect 13905 12066 13971 12069
rect 17125 12066 17191 12069
rect 13905 12064 17191 12066
rect 13905 12008 13910 12064
rect 13966 12008 17130 12064
rect 17186 12008 17191 12064
rect 13905 12006 17191 12008
rect 13905 12003 13971 12006
rect 17125 12003 17191 12006
rect 30925 12066 30991 12069
rect 34421 12066 34487 12069
rect 30925 12064 34487 12066
rect 30925 12008 30930 12064
rect 30986 12008 34426 12064
rect 34482 12008 34487 12064
rect 30925 12006 34487 12008
rect 30925 12003 30991 12006
rect 34421 12003 34487 12006
rect 49141 12066 49207 12069
rect 50200 12066 51000 12096
rect 49141 12064 51000 12066
rect 49141 12008 49146 12064
rect 49202 12008 51000 12064
rect 49141 12006 51000 12008
rect 49141 12003 49207 12006
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 50200 11976 51000 12006
rect 47946 11935 48262 11936
rect 17217 11930 17283 11933
rect 15150 11928 17283 11930
rect 15150 11872 17222 11928
rect 17278 11872 17283 11928
rect 15150 11870 17283 11872
rect 0 11794 800 11824
rect 1301 11794 1367 11797
rect 0 11792 1367 11794
rect 0 11736 1306 11792
rect 1362 11736 1367 11792
rect 0 11734 1367 11736
rect 0 11704 800 11734
rect 1301 11731 1367 11734
rect 12893 11794 12959 11797
rect 13445 11794 13511 11797
rect 15150 11794 15210 11870
rect 17217 11867 17283 11870
rect 19885 11930 19951 11933
rect 22369 11930 22435 11933
rect 19885 11928 22435 11930
rect 19885 11872 19890 11928
rect 19946 11872 22374 11928
rect 22430 11872 22435 11928
rect 19885 11870 22435 11872
rect 19885 11867 19951 11870
rect 22369 11867 22435 11870
rect 29177 11930 29243 11933
rect 29913 11930 29979 11933
rect 29177 11928 29979 11930
rect 29177 11872 29182 11928
rect 29238 11872 29918 11928
rect 29974 11872 29979 11928
rect 29177 11870 29979 11872
rect 29177 11867 29243 11870
rect 29913 11867 29979 11870
rect 32765 11930 32831 11933
rect 34789 11930 34855 11933
rect 32765 11928 34855 11930
rect 32765 11872 32770 11928
rect 32826 11872 34794 11928
rect 34850 11872 34855 11928
rect 32765 11870 34855 11872
rect 32765 11867 32831 11870
rect 34789 11867 34855 11870
rect 38326 11868 38332 11932
rect 38396 11930 38402 11932
rect 38396 11870 45570 11930
rect 38396 11868 38402 11870
rect 12893 11792 15210 11794
rect 12893 11736 12898 11792
rect 12954 11736 13450 11792
rect 13506 11736 15210 11792
rect 12893 11734 15210 11736
rect 12893 11731 12959 11734
rect 13445 11731 13511 11734
rect 15326 11732 15332 11796
rect 15396 11794 15402 11796
rect 15469 11794 15535 11797
rect 15396 11792 15535 11794
rect 15396 11736 15474 11792
rect 15530 11736 15535 11792
rect 15396 11734 15535 11736
rect 15396 11732 15402 11734
rect 15469 11731 15535 11734
rect 28809 11794 28875 11797
rect 38929 11794 38995 11797
rect 28809 11792 38995 11794
rect 28809 11736 28814 11792
rect 28870 11736 38934 11792
rect 38990 11736 38995 11792
rect 28809 11734 38995 11736
rect 45510 11794 45570 11870
rect 48957 11794 49023 11797
rect 45510 11792 49023 11794
rect 45510 11736 48962 11792
rect 49018 11736 49023 11792
rect 45510 11734 49023 11736
rect 28809 11731 28875 11734
rect 38929 11731 38995 11734
rect 48957 11731 49023 11734
rect 11789 11658 11855 11661
rect 16941 11658 17007 11661
rect 11789 11656 17007 11658
rect 11789 11600 11794 11656
rect 11850 11600 16946 11656
rect 17002 11600 17007 11656
rect 11789 11598 17007 11600
rect 11789 11595 11855 11598
rect 16941 11595 17007 11598
rect 20989 11658 21055 11661
rect 27429 11658 27495 11661
rect 28993 11658 29059 11661
rect 20989 11656 29059 11658
rect 20989 11600 20994 11656
rect 21050 11600 27434 11656
rect 27490 11600 28998 11656
rect 29054 11600 29059 11656
rect 20989 11598 29059 11600
rect 20989 11595 21055 11598
rect 27429 11595 27495 11598
rect 28993 11595 29059 11598
rect 32029 11658 32095 11661
rect 40125 11658 40191 11661
rect 32029 11656 40191 11658
rect 32029 11600 32034 11656
rect 32090 11600 40130 11656
rect 40186 11600 40191 11656
rect 32029 11598 40191 11600
rect 32029 11595 32095 11598
rect 40125 11595 40191 11598
rect 49141 11658 49207 11661
rect 50200 11658 51000 11688
rect 49141 11656 51000 11658
rect 49141 11600 49146 11656
rect 49202 11600 51000 11656
rect 49141 11598 51000 11600
rect 49141 11595 49207 11598
rect 50200 11568 51000 11598
rect 12065 11522 12131 11525
rect 12433 11522 12499 11525
rect 12065 11520 12499 11522
rect 12065 11464 12070 11520
rect 12126 11464 12438 11520
rect 12494 11464 12499 11520
rect 12065 11462 12499 11464
rect 12065 11459 12131 11462
rect 12433 11459 12499 11462
rect 14825 11522 14891 11525
rect 18597 11522 18663 11525
rect 14825 11520 18663 11522
rect 14825 11464 14830 11520
rect 14886 11464 18602 11520
rect 18658 11464 18663 11520
rect 14825 11462 18663 11464
rect 14825 11459 14891 11462
rect 18597 11459 18663 11462
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 1301 11386 1367 11389
rect 40033 11386 40099 11389
rect 40309 11386 40375 11389
rect 0 11384 1367 11386
rect 0 11328 1306 11384
rect 1362 11328 1367 11384
rect 0 11326 1367 11328
rect 0 11296 800 11326
rect 1301 11323 1367 11326
rect 34470 11384 40375 11386
rect 34470 11328 40038 11384
rect 40094 11328 40314 11384
rect 40370 11328 40375 11384
rect 34470 11326 40375 11328
rect 28993 11250 29059 11253
rect 34470 11250 34530 11326
rect 40033 11323 40099 11326
rect 40309 11323 40375 11326
rect 28993 11248 34530 11250
rect 28993 11192 28998 11248
rect 29054 11192 34530 11248
rect 28993 11190 34530 11192
rect 34697 11250 34763 11253
rect 40125 11250 40191 11253
rect 34697 11248 40191 11250
rect 34697 11192 34702 11248
rect 34758 11192 40130 11248
rect 40186 11192 40191 11248
rect 34697 11190 40191 11192
rect 28993 11187 29059 11190
rect 34697 11187 34763 11190
rect 40125 11187 40191 11190
rect 49233 11250 49299 11253
rect 50200 11250 51000 11280
rect 49233 11248 51000 11250
rect 49233 11192 49238 11248
rect 49294 11192 51000 11248
rect 49233 11190 51000 11192
rect 49233 11187 49299 11190
rect 50200 11160 51000 11190
rect 1761 11114 1827 11117
rect 14641 11114 14707 11117
rect 1761 11112 14707 11114
rect 1761 11056 1766 11112
rect 1822 11056 14646 11112
rect 14702 11056 14707 11112
rect 1761 11054 14707 11056
rect 1761 11051 1827 11054
rect 14641 11051 14707 11054
rect 15101 11114 15167 11117
rect 18505 11114 18571 11117
rect 15101 11112 18571 11114
rect 15101 11056 15106 11112
rect 15162 11056 18510 11112
rect 18566 11056 18571 11112
rect 15101 11054 18571 11056
rect 15101 11051 15167 11054
rect 18505 11051 18571 11054
rect 23289 11114 23355 11117
rect 23749 11114 23815 11117
rect 28625 11114 28691 11117
rect 28942 11114 28948 11116
rect 23289 11112 28948 11114
rect 23289 11056 23294 11112
rect 23350 11056 23754 11112
rect 23810 11056 28630 11112
rect 28686 11056 28948 11112
rect 23289 11054 28948 11056
rect 23289 11051 23355 11054
rect 23749 11051 23815 11054
rect 28625 11051 28691 11054
rect 28942 11052 28948 11054
rect 29012 11052 29018 11116
rect 31569 11114 31635 11117
rect 33961 11114 34027 11117
rect 31569 11112 34027 11114
rect 31569 11056 31574 11112
rect 31630 11056 33966 11112
rect 34022 11056 34027 11112
rect 31569 11054 34027 11056
rect 31569 11051 31635 11054
rect 33961 11051 34027 11054
rect 35249 11114 35315 11117
rect 40769 11114 40835 11117
rect 35249 11112 40835 11114
rect 35249 11056 35254 11112
rect 35310 11056 40774 11112
rect 40830 11056 40835 11112
rect 35249 11054 40835 11056
rect 35249 11051 35315 11054
rect 40769 11051 40835 11054
rect 0 10978 800 11008
rect 1577 10978 1643 10981
rect 0 10976 1643 10978
rect 0 10920 1582 10976
rect 1638 10920 1643 10976
rect 0 10918 1643 10920
rect 0 10888 800 10918
rect 1577 10915 1643 10918
rect 34329 10978 34395 10981
rect 37733 10978 37799 10981
rect 34329 10976 37799 10978
rect 34329 10920 34334 10976
rect 34390 10920 37738 10976
rect 37794 10920 37799 10976
rect 34329 10918 37799 10920
rect 34329 10915 34395 10918
rect 37733 10915 37799 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 19885 10842 19951 10845
rect 27337 10842 27403 10845
rect 35382 10842 35388 10844
rect 19885 10840 27403 10842
rect 19885 10784 19890 10840
rect 19946 10784 27342 10840
rect 27398 10784 27403 10840
rect 19885 10782 27403 10784
rect 19885 10779 19951 10782
rect 27337 10779 27403 10782
rect 28398 10782 35388 10842
rect 13721 10706 13787 10709
rect 20713 10706 20779 10709
rect 13721 10704 20779 10706
rect 13721 10648 13726 10704
rect 13782 10648 20718 10704
rect 20774 10648 20779 10704
rect 13721 10646 20779 10648
rect 13721 10643 13787 10646
rect 20713 10643 20779 10646
rect 22185 10706 22251 10709
rect 28398 10706 28458 10782
rect 35382 10780 35388 10782
rect 35452 10780 35458 10844
rect 49141 10842 49207 10845
rect 50200 10842 51000 10872
rect 49141 10840 51000 10842
rect 49141 10784 49146 10840
rect 49202 10784 51000 10840
rect 49141 10782 51000 10784
rect 49141 10779 49207 10782
rect 50200 10752 51000 10782
rect 40217 10706 40283 10709
rect 22185 10704 28458 10706
rect 22185 10648 22190 10704
rect 22246 10648 28458 10704
rect 22185 10646 28458 10648
rect 28582 10704 40283 10706
rect 28582 10648 40222 10704
rect 40278 10648 40283 10704
rect 28582 10646 40283 10648
rect 22185 10643 22251 10646
rect 0 10570 800 10600
rect 1301 10570 1367 10573
rect 0 10568 1367 10570
rect 0 10512 1306 10568
rect 1362 10512 1367 10568
rect 0 10510 1367 10512
rect 0 10480 800 10510
rect 1301 10507 1367 10510
rect 2497 10570 2563 10573
rect 15653 10570 15719 10573
rect 2497 10568 15719 10570
rect 2497 10512 2502 10568
rect 2558 10512 15658 10568
rect 15714 10512 15719 10568
rect 2497 10510 15719 10512
rect 2497 10507 2563 10510
rect 15653 10507 15719 10510
rect 25405 10570 25471 10573
rect 28582 10570 28642 10646
rect 40217 10643 40283 10646
rect 25405 10568 28642 10570
rect 25405 10512 25410 10568
rect 25466 10512 28642 10568
rect 25405 10510 28642 10512
rect 30557 10570 30623 10573
rect 48773 10570 48839 10573
rect 30557 10568 48839 10570
rect 30557 10512 30562 10568
rect 30618 10512 48778 10568
rect 48834 10512 48839 10568
rect 30557 10510 48839 10512
rect 25405 10507 25471 10510
rect 30557 10507 30623 10510
rect 48773 10507 48839 10510
rect 49325 10434 49391 10437
rect 50200 10434 51000 10464
rect 49325 10432 51000 10434
rect 49325 10376 49330 10432
rect 49386 10376 51000 10432
rect 49325 10374 51000 10376
rect 49325 10371 49391 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 50200 10344 51000 10374
rect 42946 10303 43262 10304
rect 15009 10298 15075 10301
rect 15837 10298 15903 10301
rect 19885 10298 19951 10301
rect 15009 10296 19951 10298
rect 15009 10240 15014 10296
rect 15070 10240 15842 10296
rect 15898 10240 19890 10296
rect 19946 10240 19951 10296
rect 15009 10238 19951 10240
rect 15009 10235 15075 10238
rect 15837 10235 15903 10238
rect 19885 10235 19951 10238
rect 0 10162 800 10192
rect 1209 10162 1275 10165
rect 0 10160 1275 10162
rect 0 10104 1214 10160
rect 1270 10104 1275 10160
rect 0 10102 1275 10104
rect 0 10072 800 10102
rect 1209 10099 1275 10102
rect 16481 10162 16547 10165
rect 27061 10162 27127 10165
rect 33685 10164 33751 10165
rect 33685 10162 33732 10164
rect 16481 10160 27127 10162
rect 16481 10104 16486 10160
rect 16542 10104 27066 10160
rect 27122 10104 27127 10160
rect 16481 10102 27127 10104
rect 33640 10160 33732 10162
rect 33796 10162 33802 10164
rect 34421 10162 34487 10165
rect 39481 10162 39547 10165
rect 33796 10160 39547 10162
rect 33640 10104 33690 10160
rect 33796 10104 34426 10160
rect 34482 10104 39486 10160
rect 39542 10104 39547 10160
rect 33640 10102 33732 10104
rect 16481 10099 16547 10102
rect 27061 10099 27127 10102
rect 33685 10100 33732 10102
rect 33796 10102 39547 10104
rect 33796 10100 33802 10102
rect 33685 10099 33751 10100
rect 34421 10099 34487 10102
rect 39481 10099 39547 10102
rect 11329 10026 11395 10029
rect 18597 10026 18663 10029
rect 11329 10024 18663 10026
rect 11329 9968 11334 10024
rect 11390 9968 18602 10024
rect 18658 9968 18663 10024
rect 11329 9966 18663 9968
rect 11329 9963 11395 9966
rect 18597 9963 18663 9966
rect 30557 10026 30623 10029
rect 38285 10026 38351 10029
rect 30557 10024 38351 10026
rect 30557 9968 30562 10024
rect 30618 9968 38290 10024
rect 38346 9968 38351 10024
rect 30557 9966 38351 9968
rect 30557 9963 30623 9966
rect 38285 9963 38351 9966
rect 49233 10026 49299 10029
rect 50200 10026 51000 10056
rect 49233 10024 51000 10026
rect 49233 9968 49238 10024
rect 49294 9968 51000 10024
rect 49233 9966 51000 9968
rect 49233 9963 49299 9966
rect 50200 9936 51000 9966
rect 7946 9824 8262 9825
rect 0 9754 800 9784
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 1301 9754 1367 9757
rect 0 9752 1367 9754
rect 0 9696 1306 9752
rect 1362 9696 1367 9752
rect 0 9694 1367 9696
rect 0 9664 800 9694
rect 1301 9691 1367 9694
rect 15142 9556 15148 9620
rect 15212 9618 15218 9620
rect 26049 9618 26115 9621
rect 36261 9618 36327 9621
rect 15212 9616 36327 9618
rect 15212 9560 26054 9616
rect 26110 9560 36266 9616
rect 36322 9560 36327 9616
rect 15212 9558 36327 9560
rect 15212 9556 15218 9558
rect 26049 9555 26115 9558
rect 36261 9555 36327 9558
rect 47301 9618 47367 9621
rect 50200 9618 51000 9648
rect 47301 9616 51000 9618
rect 47301 9560 47306 9616
rect 47362 9560 51000 9616
rect 47301 9558 51000 9560
rect 47301 9555 47367 9558
rect 50200 9528 51000 9558
rect 1853 9482 1919 9485
rect 23381 9482 23447 9485
rect 1853 9480 23447 9482
rect 1853 9424 1858 9480
rect 1914 9424 23386 9480
rect 23442 9424 23447 9480
rect 1853 9422 23447 9424
rect 1853 9419 1919 9422
rect 23381 9419 23447 9422
rect 32673 9482 32739 9485
rect 35525 9482 35591 9485
rect 32673 9480 35591 9482
rect 32673 9424 32678 9480
rect 32734 9424 35530 9480
rect 35586 9424 35591 9480
rect 32673 9422 35591 9424
rect 32673 9419 32739 9422
rect 35525 9419 35591 9422
rect 0 9346 800 9376
rect 1301 9346 1367 9349
rect 0 9344 1367 9346
rect 0 9288 1306 9344
rect 1362 9288 1367 9344
rect 0 9286 1367 9288
rect 0 9256 800 9286
rect 1301 9283 1367 9286
rect 15101 9346 15167 9349
rect 15326 9346 15332 9348
rect 15101 9344 15332 9346
rect 15101 9288 15106 9344
rect 15162 9288 15332 9344
rect 15101 9286 15332 9288
rect 15101 9283 15167 9286
rect 15326 9284 15332 9286
rect 15396 9284 15402 9348
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 49141 9210 49207 9213
rect 50200 9210 51000 9240
rect 49141 9208 51000 9210
rect 49141 9152 49146 9208
rect 49202 9152 51000 9208
rect 49141 9150 51000 9152
rect 49141 9147 49207 9150
rect 50200 9120 51000 9150
rect 22461 9074 22527 9077
rect 26141 9074 26207 9077
rect 22461 9072 26207 9074
rect 22461 9016 22466 9072
rect 22522 9016 26146 9072
rect 26202 9016 26207 9072
rect 22461 9014 26207 9016
rect 22461 9011 22527 9014
rect 26141 9011 26207 9014
rect 0 8938 800 8968
rect 1301 8938 1367 8941
rect 0 8936 1367 8938
rect 0 8880 1306 8936
rect 1362 8880 1367 8936
rect 0 8878 1367 8880
rect 0 8848 800 8878
rect 1301 8875 1367 8878
rect 2497 8938 2563 8941
rect 20529 8938 20595 8941
rect 2497 8936 20595 8938
rect 2497 8880 2502 8936
rect 2558 8880 20534 8936
rect 20590 8880 20595 8936
rect 2497 8878 20595 8880
rect 2497 8875 2563 8878
rect 20529 8875 20595 8878
rect 23473 8938 23539 8941
rect 33409 8938 33475 8941
rect 33961 8938 34027 8941
rect 23473 8936 34027 8938
rect 23473 8880 23478 8936
rect 23534 8880 33414 8936
rect 33470 8880 33966 8936
rect 34022 8880 34027 8936
rect 23473 8878 34027 8880
rect 23473 8875 23539 8878
rect 33409 8875 33475 8878
rect 33961 8875 34027 8878
rect 49233 8802 49299 8805
rect 50200 8802 51000 8832
rect 49233 8800 51000 8802
rect 49233 8744 49238 8800
rect 49294 8744 51000 8800
rect 49233 8742 51000 8744
rect 49233 8739 49299 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 50200 8712 51000 8742
rect 47946 8671 48262 8672
rect 0 8530 800 8560
rect 1209 8530 1275 8533
rect 0 8528 1275 8530
rect 0 8472 1214 8528
rect 1270 8472 1275 8528
rect 0 8470 1275 8472
rect 0 8440 800 8470
rect 1209 8467 1275 8470
rect 21541 8392 21607 8397
rect 21541 8336 21546 8392
rect 21602 8336 21607 8392
rect 21541 8331 21607 8336
rect 49325 8394 49391 8397
rect 50200 8394 51000 8424
rect 49325 8392 51000 8394
rect 49325 8336 49330 8392
rect 49386 8336 51000 8392
rect 49325 8334 51000 8336
rect 49325 8331 49391 8334
rect 16573 8258 16639 8261
rect 21544 8258 21604 8331
rect 50200 8304 51000 8334
rect 16573 8256 21604 8258
rect 16573 8200 16578 8256
rect 16634 8200 21604 8256
rect 16573 8198 21604 8200
rect 16573 8195 16639 8198
rect 2946 8192 3262 8193
rect 0 8122 800 8152
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 1393 8122 1459 8125
rect 0 8120 1459 8122
rect 0 8064 1398 8120
rect 1454 8064 1459 8120
rect 0 8062 1459 8064
rect 0 8032 800 8062
rect 1393 8059 1459 8062
rect 46841 7986 46907 7989
rect 50200 7986 51000 8016
rect 46841 7984 51000 7986
rect 46841 7928 46846 7984
rect 46902 7928 51000 7984
rect 46841 7926 51000 7928
rect 46841 7923 46907 7926
rect 50200 7896 51000 7926
rect 0 7714 800 7744
rect 1301 7714 1367 7717
rect 0 7712 1367 7714
rect 0 7656 1306 7712
rect 1362 7656 1367 7712
rect 0 7654 1367 7656
rect 0 7624 800 7654
rect 1301 7651 1367 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 28942 7516 28948 7580
rect 29012 7578 29018 7580
rect 37365 7578 37431 7581
rect 29012 7576 37431 7578
rect 29012 7520 37370 7576
rect 37426 7520 37431 7576
rect 29012 7518 37431 7520
rect 29012 7516 29018 7518
rect 37365 7515 37431 7518
rect 49141 7578 49207 7581
rect 50200 7578 51000 7608
rect 49141 7576 51000 7578
rect 49141 7520 49146 7576
rect 49202 7520 51000 7576
rect 49141 7518 51000 7520
rect 49141 7515 49207 7518
rect 50200 7488 51000 7518
rect 0 7306 800 7336
rect 1301 7306 1367 7309
rect 0 7304 1367 7306
rect 0 7248 1306 7304
rect 1362 7248 1367 7304
rect 0 7246 1367 7248
rect 0 7216 800 7246
rect 1301 7243 1367 7246
rect 49325 7170 49391 7173
rect 50200 7170 51000 7200
rect 49325 7168 51000 7170
rect 49325 7112 49330 7168
rect 49386 7112 51000 7168
rect 49325 7110 51000 7112
rect 49325 7107 49391 7110
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 50200 7080 51000 7110
rect 42946 7039 43262 7040
rect 0 6898 800 6928
rect 1209 6898 1275 6901
rect 0 6896 1275 6898
rect 0 6840 1214 6896
rect 1270 6840 1275 6896
rect 0 6838 1275 6840
rect 0 6808 800 6838
rect 1209 6835 1275 6838
rect 49233 6762 49299 6765
rect 50200 6762 51000 6792
rect 49233 6760 51000 6762
rect 49233 6704 49238 6760
rect 49294 6704 51000 6760
rect 49233 6702 51000 6704
rect 49233 6699 49299 6702
rect 50200 6672 51000 6702
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 1301 6490 1367 6493
rect 0 6488 1367 6490
rect 0 6432 1306 6488
rect 1362 6432 1367 6488
rect 0 6430 1367 6432
rect 0 6400 800 6430
rect 1301 6427 1367 6430
rect 48865 6354 48931 6357
rect 50200 6354 51000 6384
rect 48865 6352 51000 6354
rect 48865 6296 48870 6352
rect 48926 6296 51000 6352
rect 48865 6294 51000 6296
rect 48865 6291 48931 6294
rect 50200 6264 51000 6294
rect 0 6082 800 6112
rect 1301 6082 1367 6085
rect 0 6080 1367 6082
rect 0 6024 1306 6080
rect 1362 6024 1367 6080
rect 0 6022 1367 6024
rect 0 5992 800 6022
rect 1301 6019 1367 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 49141 5946 49207 5949
rect 50200 5946 51000 5976
rect 49141 5944 51000 5946
rect 49141 5888 49146 5944
rect 49202 5888 51000 5944
rect 49141 5886 51000 5888
rect 49141 5883 49207 5886
rect 50200 5856 51000 5886
rect 0 5674 800 5704
rect 1301 5674 1367 5677
rect 0 5672 1367 5674
rect 0 5616 1306 5672
rect 1362 5616 1367 5672
rect 0 5614 1367 5616
rect 0 5584 800 5614
rect 1301 5611 1367 5614
rect 29310 5612 29316 5676
rect 29380 5674 29386 5676
rect 34237 5674 34303 5677
rect 29380 5672 34303 5674
rect 29380 5616 34242 5672
rect 34298 5616 34303 5672
rect 29380 5614 34303 5616
rect 29380 5612 29386 5614
rect 34237 5611 34303 5614
rect 49417 5538 49483 5541
rect 50200 5538 51000 5568
rect 49417 5536 51000 5538
rect 49417 5480 49422 5536
rect 49478 5480 51000 5536
rect 49417 5478 51000 5480
rect 49417 5475 49483 5478
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 50200 5448 51000 5478
rect 47946 5407 48262 5408
rect 0 5266 800 5296
rect 2773 5266 2839 5269
rect 0 5264 2839 5266
rect 0 5208 2778 5264
rect 2834 5208 2839 5264
rect 0 5206 2839 5208
rect 0 5176 800 5206
rect 2773 5203 2839 5206
rect 8845 5130 8911 5133
rect 21214 5130 21220 5132
rect 8845 5128 21220 5130
rect 8845 5072 8850 5128
rect 8906 5072 21220 5128
rect 8845 5070 21220 5072
rect 8845 5067 8911 5070
rect 21214 5068 21220 5070
rect 21284 5130 21290 5132
rect 26233 5130 26299 5133
rect 21284 5128 26299 5130
rect 21284 5072 26238 5128
rect 26294 5072 26299 5128
rect 21284 5070 26299 5072
rect 21284 5068 21290 5070
rect 26233 5067 26299 5070
rect 49325 5130 49391 5133
rect 50200 5130 51000 5160
rect 49325 5128 51000 5130
rect 49325 5072 49330 5128
rect 49386 5072 51000 5128
rect 49325 5070 51000 5072
rect 49325 5067 49391 5070
rect 50200 5040 51000 5070
rect 2946 4928 3262 4929
rect 0 4858 800 4888
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 48313 4722 48379 4725
rect 50200 4722 51000 4752
rect 48313 4720 51000 4722
rect 48313 4664 48318 4720
rect 48374 4664 51000 4720
rect 48313 4662 51000 4664
rect 48313 4659 48379 4662
rect 50200 4632 51000 4662
rect 0 4450 800 4480
rect 1301 4450 1367 4453
rect 0 4448 1367 4450
rect 0 4392 1306 4448
rect 1362 4392 1367 4448
rect 0 4390 1367 4392
rect 0 4360 800 4390
rect 1301 4387 1367 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 49141 4314 49207 4317
rect 50200 4314 51000 4344
rect 49141 4312 51000 4314
rect 49141 4256 49146 4312
rect 49202 4256 51000 4312
rect 49141 4254 51000 4256
rect 49141 4251 49207 4254
rect 50200 4224 51000 4254
rect 0 4042 800 4072
rect 1393 4042 1459 4045
rect 0 4040 1459 4042
rect 0 3984 1398 4040
rect 1454 3984 1459 4040
rect 0 3982 1459 3984
rect 0 3952 800 3982
rect 1393 3979 1459 3982
rect 49233 3906 49299 3909
rect 50200 3906 51000 3936
rect 49233 3904 51000 3906
rect 49233 3848 49238 3904
rect 49294 3848 51000 3904
rect 49233 3846 51000 3848
rect 49233 3843 49299 3846
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 50200 3816 51000 3846
rect 42946 3775 43262 3776
rect 0 3634 800 3664
rect 1301 3634 1367 3637
rect 0 3632 1367 3634
rect 0 3576 1306 3632
rect 1362 3576 1367 3632
rect 0 3574 1367 3576
rect 0 3544 800 3574
rect 1301 3571 1367 3574
rect 49141 3498 49207 3501
rect 50200 3498 51000 3528
rect 49141 3496 51000 3498
rect 49141 3440 49146 3496
rect 49202 3440 51000 3496
rect 49141 3438 51000 3440
rect 49141 3435 49207 3438
rect 50200 3408 51000 3438
rect 7946 3296 8262 3297
rect 0 3226 800 3256
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 1301 3226 1367 3229
rect 0 3224 1367 3226
rect 0 3168 1306 3224
rect 1362 3168 1367 3224
rect 0 3166 1367 3168
rect 0 3136 800 3166
rect 1301 3163 1367 3166
rect 48681 3090 48747 3093
rect 50200 3090 51000 3120
rect 48681 3088 51000 3090
rect 48681 3032 48686 3088
rect 48742 3032 51000 3088
rect 48681 3030 51000 3032
rect 48681 3027 48747 3030
rect 50200 3000 51000 3030
rect 0 2818 800 2848
rect 1301 2818 1367 2821
rect 0 2816 1367 2818
rect 0 2760 1306 2816
rect 1362 2760 1367 2816
rect 0 2758 1367 2760
rect 0 2728 800 2758
rect 1301 2755 1367 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 46841 2682 46907 2685
rect 50200 2682 51000 2712
rect 46841 2680 51000 2682
rect 46841 2624 46846 2680
rect 46902 2624 51000 2680
rect 46841 2622 51000 2624
rect 46841 2619 46907 2622
rect 50200 2592 51000 2622
rect 0 2410 800 2440
rect 1301 2410 1367 2413
rect 0 2408 1367 2410
rect 0 2352 1306 2408
rect 1362 2352 1367 2408
rect 0 2350 1367 2352
rect 0 2320 800 2350
rect 1301 2347 1367 2350
rect 48497 2274 48563 2277
rect 50200 2274 51000 2304
rect 48497 2272 51000 2274
rect 48497 2216 48502 2272
rect 48558 2216 51000 2272
rect 48497 2214 51000 2216
rect 48497 2211 48563 2214
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 50200 2184 51000 2214
rect 47946 2143 48262 2144
rect 0 2002 800 2032
rect 1209 2002 1275 2005
rect 0 2000 1275 2002
rect 0 1944 1214 2000
rect 1270 1944 1275 2000
rect 0 1942 1275 1944
rect 0 1912 800 1942
rect 1209 1939 1275 1942
rect 46749 1866 46815 1869
rect 50200 1866 51000 1896
rect 46749 1864 51000 1866
rect 46749 1808 46754 1864
rect 46810 1808 51000 1864
rect 46749 1806 51000 1808
rect 46749 1803 46815 1806
rect 50200 1776 51000 1806
rect 0 1594 800 1624
rect 1301 1594 1367 1597
rect 0 1592 1367 1594
rect 0 1536 1306 1592
rect 1362 1536 1367 1592
rect 0 1534 1367 1536
rect 0 1504 800 1534
rect 1301 1531 1367 1534
rect 46657 1458 46723 1461
rect 50200 1458 51000 1488
rect 46657 1456 51000 1458
rect 46657 1400 46662 1456
rect 46718 1400 51000 1456
rect 46657 1398 51000 1400
rect 46657 1395 46723 1398
rect 50200 1368 51000 1398
<< via3 >>
rect 33548 26556 33612 26620
rect 45692 26284 45756 26348
rect 34284 26012 34348 26076
rect 19932 25604 19996 25668
rect 44220 25468 44284 25532
rect 30052 24652 30116 24716
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 36492 22748 36556 22812
rect 19932 22672 19996 22676
rect 19932 22616 19946 22672
rect 19946 22616 19996 22672
rect 19932 22612 19996 22616
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 34284 21660 34348 21724
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 44220 21660 44284 21724
rect 45692 21524 45756 21588
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 7788 20980 7852 21044
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 30052 19892 30116 19956
rect 31156 19892 31220 19956
rect 28948 19756 29012 19820
rect 34468 19756 34532 19820
rect 32812 19620 32876 19684
rect 35388 19680 35452 19684
rect 35388 19624 35402 19680
rect 35402 19624 35452 19680
rect 35388 19620 35452 19624
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 33364 19212 33428 19276
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 7788 18804 7852 18868
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 33732 18396 33796 18460
rect 38332 18260 38396 18324
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 33548 18124 33612 18188
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 34468 17852 34532 17916
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 28948 17308 29012 17372
rect 31156 17308 31220 17372
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 15332 16220 15396 16284
rect 16436 16220 16500 16284
rect 32812 16144 32876 16148
rect 32812 16088 32862 16144
rect 32862 16088 32876 16144
rect 32812 16084 32876 16088
rect 16436 15812 16500 15876
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 33364 14452 33428 14516
rect 15148 14180 15212 14244
rect 29316 14240 29380 14244
rect 29316 14184 29330 14240
rect 29330 14184 29380 14240
rect 29316 14180 29380 14184
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 21220 13152 21284 13156
rect 21220 13096 21270 13152
rect 21270 13096 21284 13152
rect 21220 13092 21284 13096
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 36492 12684 36556 12748
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 38332 11868 38396 11932
rect 15332 11732 15396 11796
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 28948 11052 29012 11116
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 35388 10780 35452 10844
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 33732 10160 33796 10164
rect 33732 10104 33746 10160
rect 33746 10104 33796 10160
rect 33732 10100 33796 10104
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 15148 9556 15212 9620
rect 15332 9284 15396 9348
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 28948 7516 29012 7580
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 29316 5612 29380 5676
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 21220 5068 21284 5132
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 33547 26620 33613 26621
rect 33547 26556 33548 26620
rect 33612 26556 33613 26620
rect 33547 26555 33613 26556
rect 19931 25668 19997 25669
rect 19931 25604 19932 25668
rect 19996 25604 19997 25668
rect 19931 25603 19997 25604
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7787 21044 7853 21045
rect 7787 20980 7788 21044
rect 7852 20980 7853 21044
rect 7787 20979 7853 20980
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 7790 18869 7850 20979
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7787 18868 7853 18869
rect 7787 18804 7788 18868
rect 7852 18804 7853 18868
rect 7787 18803 7853 18804
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 17944 23968 18264 24528
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 19934 22677 19994 25603
rect 30051 24716 30117 24717
rect 30051 24652 30052 24716
rect 30116 24652 30117 24716
rect 30051 24651 30117 24652
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 19931 22676 19997 22677
rect 19931 22612 19932 22676
rect 19996 22612 19997 22676
rect 19931 22611 19997 22612
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 15331 16284 15397 16285
rect 15331 16220 15332 16284
rect 15396 16220 15397 16284
rect 15331 16219 15397 16220
rect 16435 16284 16501 16285
rect 16435 16220 16436 16284
rect 16500 16220 16501 16284
rect 16435 16219 16501 16220
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 15147 14244 15213 14245
rect 15147 14180 15148 14244
rect 15212 14180 15213 14244
rect 15147 14179 15213 14180
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 15150 9621 15210 14179
rect 15334 11797 15394 16219
rect 16438 15877 16498 16219
rect 16435 15876 16501 15877
rect 16435 15812 16436 15876
rect 16500 15812 16501 15876
rect 16435 15811 16501 15812
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 21219 13156 21285 13157
rect 21219 13092 21220 13156
rect 21284 13092 21285 13156
rect 21219 13091 21285 13092
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 15331 11796 15397 11797
rect 15331 11732 15332 11796
rect 15396 11732 15397 11796
rect 15331 11731 15397 11732
rect 15147 9620 15213 9621
rect 15147 9556 15148 9620
rect 15212 9556 15213 9620
rect 15147 9555 15213 9556
rect 15334 9349 15394 11731
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 15331 9348 15397 9349
rect 15331 9284 15332 9348
rect 15396 9284 15397 9348
rect 15331 9283 15397 9284
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 21222 5133 21282 13091
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 21219 5132 21285 5133
rect 21219 5068 21220 5132
rect 21284 5068 21285 5132
rect 21219 5067 21285 5068
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 27944 23968 28264 24528
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 30054 19957 30114 24651
rect 32944 24512 33264 24528
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 30051 19956 30117 19957
rect 30051 19892 30052 19956
rect 30116 19892 30117 19956
rect 30051 19891 30117 19892
rect 31155 19956 31221 19957
rect 31155 19892 31156 19956
rect 31220 19892 31221 19956
rect 31155 19891 31221 19892
rect 28947 19820 29013 19821
rect 28947 19756 28948 19820
rect 29012 19756 29013 19820
rect 28947 19755 29013 19756
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27944 18528 28264 19552
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27944 17440 28264 18464
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 28950 17373 29010 19755
rect 31158 17373 31218 19891
rect 32811 19684 32877 19685
rect 32811 19620 32812 19684
rect 32876 19620 32877 19684
rect 32811 19619 32877 19620
rect 28947 17372 29013 17373
rect 28947 17308 28948 17372
rect 29012 17308 29013 17372
rect 28947 17307 29013 17308
rect 31155 17372 31221 17373
rect 31155 17308 31156 17372
rect 31220 17308 31221 17372
rect 31155 17307 31221 17308
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 32814 16149 32874 19619
rect 32944 19072 33264 20096
rect 33363 19276 33429 19277
rect 33363 19212 33364 19276
rect 33428 19212 33429 19276
rect 33363 19211 33429 19212
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32811 16148 32877 16149
rect 32811 16084 32812 16148
rect 32876 16084 32877 16148
rect 32811 16083 32877 16084
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27944 14176 28264 15200
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 29315 14244 29381 14245
rect 29315 14180 29316 14244
rect 29380 14180 29381 14244
rect 29315 14179 29381 14180
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 28947 11116 29013 11117
rect 28947 11052 28948 11116
rect 29012 11052 29013 11116
rect 28947 11051 29013 11052
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 28950 7581 29010 11051
rect 28947 7580 29013 7581
rect 28947 7516 28948 7580
rect 29012 7516 29013 7580
rect 28947 7515 29013 7516
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 29318 5677 29378 14179
rect 32944 13632 33264 14656
rect 33366 14517 33426 19211
rect 33550 18189 33610 26555
rect 45691 26348 45757 26349
rect 45691 26284 45692 26348
rect 45756 26284 45757 26348
rect 45691 26283 45757 26284
rect 34283 26076 34349 26077
rect 34283 26012 34284 26076
rect 34348 26012 34349 26076
rect 34283 26011 34349 26012
rect 34286 21725 34346 26011
rect 44219 25532 44285 25533
rect 44219 25468 44220 25532
rect 44284 25468 44285 25532
rect 44219 25467 44285 25468
rect 37944 23968 38264 24528
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 36491 22812 36557 22813
rect 36491 22748 36492 22812
rect 36556 22748 36557 22812
rect 36491 22747 36557 22748
rect 34283 21724 34349 21725
rect 34283 21660 34284 21724
rect 34348 21660 34349 21724
rect 34283 21659 34349 21660
rect 34467 19820 34533 19821
rect 34467 19756 34468 19820
rect 34532 19756 34533 19820
rect 34467 19755 34533 19756
rect 33731 18460 33797 18461
rect 33731 18396 33732 18460
rect 33796 18396 33797 18460
rect 33731 18395 33797 18396
rect 33547 18188 33613 18189
rect 33547 18124 33548 18188
rect 33612 18124 33613 18188
rect 33547 18123 33613 18124
rect 33363 14516 33429 14517
rect 33363 14452 33364 14516
rect 33428 14452 33429 14516
rect 33363 14451 33429 14452
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32944 10368 33264 11392
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 33734 10165 33794 18395
rect 34470 17917 34530 19755
rect 35387 19684 35453 19685
rect 35387 19620 35388 19684
rect 35452 19620 35453 19684
rect 35387 19619 35453 19620
rect 34467 17916 34533 17917
rect 34467 17852 34468 17916
rect 34532 17852 34533 17916
rect 34467 17851 34533 17852
rect 35390 10845 35450 19619
rect 36494 12749 36554 22747
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 42944 24512 43264 24528
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 44222 21725 44282 25467
rect 44219 21724 44285 21725
rect 44219 21660 44220 21724
rect 44284 21660 44285 21724
rect 44219 21659 44285 21660
rect 45694 21589 45754 26283
rect 47944 23968 48264 24528
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 45691 21588 45757 21589
rect 45691 21524 45692 21588
rect 45756 21524 45757 21588
rect 45691 21523 45757 21524
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 38331 18324 38397 18325
rect 38331 18260 38332 18324
rect 38396 18260 38397 18324
rect 38331 18259 38397 18260
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 36491 12748 36557 12749
rect 36491 12684 36492 12748
rect 36556 12684 36557 12748
rect 36491 12683 36557 12684
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 38334 11933 38394 18259
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 38331 11932 38397 11933
rect 38331 11868 38332 11932
rect 38396 11868 38397 11932
rect 38331 11867 38397 11868
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 35387 10844 35453 10845
rect 35387 10780 35388 10844
rect 35452 10780 35453 10844
rect 35387 10779 35453 10780
rect 33731 10164 33797 10165
rect 33731 10100 33732 10164
rect 33796 10100 33797 10164
rect 33731 10099 33797 10100
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 29315 5676 29381 5677
rect 29315 5612 29316 5676
rect 29380 5612 29381 5676
rect 29315 5611 29381 5612
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_2  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14260 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1679235063
transform 1 0 11040 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1679235063
transform 1 0 9476 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1679235063
transform 1 0 6440 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1679235063
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1679235063
transform 1 0 10856 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1679235063
transform 1 0 13432 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1679235063
transform 1 0 8096 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1679235063
transform 1 0 10488 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1679235063
transform 1 0 9292 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1679235063
transform 1 0 11684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1679235063
transform 1 0 9200 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1679235063
transform 1 0 16008 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1679235063
transform 1 0 16008 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1679235063
transform 1 0 11684 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1679235063
transform 1 0 7636 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1679235063
transform 1 0 10120 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1679235063
transform 1 0 11960 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1679235063
transform 1 0 16008 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1679235063
transform 1 0 5704 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1679235063
transform 1 0 9752 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1679235063
transform 1 0 9016 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _126_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 7636 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1679235063
transform 1 0 7728 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1679235063
transform 1 0 5244 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1679235063
transform 1 0 8280 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1679235063
transform 1 0 6164 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1679235063
transform 1 0 3956 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1679235063
transform 1 0 5244 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1679235063
transform 1 0 2024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1679235063
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1679235063
transform 1 0 37260 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1679235063
transform 1 0 37996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1679235063
transform 1 0 43608 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1679235063
transform 1 0 38456 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1679235063
transform 1 0 37720 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1679235063
transform 1 0 37444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1679235063
transform 1 0 43884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1679235063
transform 1 0 38456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1679235063
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1679235063
transform 1 0 37904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1679235063
transform 1 0 44712 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1679235063
transform 1 0 38640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1679235063
transform 1 0 40204 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1679235063
transform 1 0 39192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1679235063
transform 1 0 44068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1679235063
transform 1 0 40020 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1679235063
transform 1 0 38180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1679235063
transform 1 0 39652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1679235063
transform 1 0 44252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1679235063
transform 1 0 40756 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1679235063
transform 1 0 40020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1679235063
transform 1 0 40020 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1679235063
transform 1 0 44988 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1679235063
transform 1 0 45540 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1679235063
transform 1 0 41032 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1679235063
transform 1 0 45908 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1679235063
transform 1 0 46000 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1679235063
transform 1 0 45632 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1679235063
transform 1 0 44896 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1679235063
transform 1 0 6716 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1679235063
transform 1 0 5428 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1679235063
transform 1 0 5244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _167_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 4140 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _168_
timestamp 1679235063
transform 1 0 3404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1679235063
transform 1 0 4784 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1679235063
transform 1 0 3956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _171_
timestamp 1679235063
transform 1 0 5796 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1679235063
transform 1 0 6532 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _173_
timestamp 1679235063
transform 1 0 6532 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1679235063
transform 1 0 24656 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp 1679235063
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1679235063
transform 1 0 8556 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1679235063
transform 1 0 10948 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _178_
timestamp 1679235063
transform 1 0 13616 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _179_
timestamp 1679235063
transform 1 0 11776 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _180_
timestamp 1679235063
transform 1 0 14444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _181_
timestamp 1679235063
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1679235063
transform 1 0 8280 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _183_
timestamp 1679235063
transform 1 0 3956 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1679235063
transform 1 0 19504 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1679235063
transform 1 0 22540 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1679235063
transform 1 0 19688 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _187_
timestamp 1679235063
transform 1 0 21160 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1679235063
transform 1 0 14536 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1679235063
transform 1 0 23736 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1679235063
transform 1 0 19688 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1679235063
transform 1 0 29716 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _192_
timestamp 1679235063
transform 1 0 27140 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1679235063
transform 1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _194_
timestamp 1679235063
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1679235063
transform 1 0 17572 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1679235063
transform 1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1679235063
transform 1 0 20240 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9016 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1679235063
transform 1 0 19596 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1679235063
transform 1 0 8188 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1679235063
transform 1 0 17940 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1679235063
transform 1 0 27784 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1679235063
transform 1 0 30728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1679235063
transform 1 0 9016 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1679235063
transform 1 0 16744 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1679235063
transform 1 0 17664 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1679235063
transform 1 0 10764 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1679235063
transform 1 0 9844 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1679235063
transform 1 0 9108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1679235063
transform 1 0 9476 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1679235063
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1679235063
transform 1 0 9108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1679235063
transform 1 0 12512 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1679235063
transform 1 0 9752 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1679235063
transform 1 0 9292 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1679235063
transform 1 0 9936 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1679235063
transform 1 0 11592 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1679235063
transform 1 0 13064 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1679235063
transform 1 0 6716 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1679235063
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1679235063
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1679235063
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1679235063
transform 1 0 5888 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1679235063
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1679235063
transform 1 0 5336 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1679235063
transform 1 0 5888 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1679235063
transform 1 0 1656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1679235063
transform 1 0 36892 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1679235063
transform 1 0 36892 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A
timestamp 1679235063
transform 1 0 38548 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A
timestamp 1679235063
transform 1 0 39008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1679235063
transform 1 0 37352 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1679235063
transform 1 0 37996 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1679235063
transform 1 0 39008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1679235063
transform 1 0 37352 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1679235063
transform 1 0 37536 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1679235063
transform 1 0 39192 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1679235063
transform 1 0 40756 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1679235063
transform 1 0 39836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1679235063
transform 1 0 40572 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1679235063
transform 1 0 38732 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1679235063
transform 1 0 39468 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1679235063
transform 1 0 40572 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1679235063
transform 1 0 40204 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1679235063
transform 1 0 40756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1679235063
transform 1 0 41768 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__A
timestamp 1679235063
transform 1 0 5612 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A
timestamp 1679235063
transform 1 0 20792 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1679235063
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__A
timestamp 1679235063
transform 1 0 3312 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1679235063
transform 1 0 18768 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__187__A
timestamp 1679235063
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A
timestamp 1679235063
transform 1 0 23000 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 1679235063
transform 1 0 11592 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A
timestamp 1679235063
transform 1 0 19320 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19412 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 15180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 17848 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 18676 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20332 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 14996 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 15640 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16376 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 9476 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 9660 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 9936 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 10396 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10120 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11592 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11040 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 6624 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12328 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 15088 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 20608 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 10028 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 17756 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 25208 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 9476 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 12696 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 11592 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 12696 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 9200 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 16468 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 8556 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 18768 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 16836 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 10488 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 12972 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__S
timestamp 1679235063
transform 1 0 17940 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 12052 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 10120 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 11592 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 16376 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 17940 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 17480 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 14996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 10580 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 26588 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 31188 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1679235063
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1679235063
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1679235063
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1679235063
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1679235063
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1679235063
transform 1 0 20424 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1679235063
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1679235063
transform 1 0 25208 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1679235063
transform 1 0 22816 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1679235063
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1679235063
transform 1 0 31740 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1679235063
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1679235063
transform 1 0 36892 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1679235063
transform 1 0 32292 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1679235063
transform 1 0 32752 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1679235063
transform 1 0 38456 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1679235063
transform 1 0 37444 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold95_A
timestamp 1679235063
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold109_A
timestamp 1679235063
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1679235063
transform 1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1679235063
transform 1 0 47748 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1679235063
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1679235063
transform 1 0 3036 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1679235063
transform 1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1679235063
transform 1 0 2760 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1679235063
transform 1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1679235063
transform 1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1679235063
transform 1 0 2300 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1679235063
transform 1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1679235063
transform 1 0 2852 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1679235063
transform 1 0 3036 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1679235063
transform 1 0 2300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1679235063
transform 1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1679235063
transform 1 0 2116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1679235063
transform 1 0 2852 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1679235063
transform 1 0 3036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1679235063
transform 1 0 2300 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1679235063
transform 1 0 2760 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1679235063
transform 1 0 2852 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1679235063
transform 1 0 2116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1679235063
transform 1 0 3312 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1679235063
transform 1 0 2668 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1679235063
transform 1 0 3956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1679235063
transform 1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1679235063
transform 1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1679235063
transform 1 0 2116 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1679235063
transform 1 0 2852 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1679235063
transform 1 0 3036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1679235063
transform 1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1679235063
transform 1 0 2116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1679235063
transform 1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1679235063
transform 1 0 48668 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1679235063
transform 1 0 48484 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1679235063
transform 1 0 48668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1679235063
transform 1 0 48668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1679235063
transform 1 0 48484 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1679235063
transform 1 0 47840 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1679235063
transform 1 0 47656 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1679235063
transform 1 0 47840 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1679235063
transform 1 0 47656 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1679235063
transform 1 0 47748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1679235063
transform 1 0 47932 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1679235063
transform 1 0 48024 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1679235063
transform 1 0 48024 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1679235063
transform 1 0 47104 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1679235063
transform 1 0 49036 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1679235063
transform 1 0 48300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1679235063
transform 1 0 48024 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1679235063
transform 1 0 46644 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1679235063
transform 1 0 47932 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1679235063
transform 1 0 47932 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1679235063
transform 1 0 47288 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1679235063
transform 1 0 46920 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1679235063
transform 1 0 48484 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1679235063
transform 1 0 48668 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1679235063
transform 1 0 48760 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1679235063
transform 1 0 48668 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1679235063
transform 1 0 48484 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1679235063
transform 1 0 48668 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1679235063
transform 1 0 48668 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1679235063
transform 1 0 48484 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1679235063
transform 1 0 3496 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1679235063
transform 1 0 46920 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1679235063
transform 1 0 49220 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1679235063
transform 1 0 43240 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1679235063
transform 1 0 47104 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1679235063
transform 1 0 47012 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1679235063
transform 1 0 45816 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1679235063
transform 1 0 42780 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1679235063
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1679235063
transform 1 0 45632 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1679235063
transform 1 0 44528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1679235063
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1679235063
transform 1 0 47288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1679235063
transform 1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1679235063
transform 1 0 43792 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1679235063
transform 1 0 47564 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1679235063
transform 1 0 46000 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1679235063
transform 1 0 44160 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1679235063
transform 1 0 44344 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1679235063
transform 1 0 44712 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1679235063
transform 1 0 47748 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1679235063
transform 1 0 47564 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1679235063
transform 1 0 5152 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1679235063
transform 1 0 27876 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1679235063
transform 1 0 7544 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1679235063
transform 1 0 47196 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1679235063
transform 1 0 6440 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1679235063
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1679235063
transform 1 0 9384 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1679235063
transform 1 0 47012 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1679235063
transform 1 0 29164 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1679235063
transform 1 0 31280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1679235063
transform 1 0 33396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1679235063
transform 1 0 35512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1679235063
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1679235063
transform 1 0 47196 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1679235063
transform 1 0 47196 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1679235063
transform 1 0 47932 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1679235063
transform 1 0 47472 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1679235063
transform 1 0 47748 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1679235063
transform 1 0 48116 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1679235063
transform 1 0 47932 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1679235063
transform 1 0 47748 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1679235063
transform 1 0 46460 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 27048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 26588 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 25024 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23276 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 20332 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 17940 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21344 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21160 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 23920 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 20792 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23368 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24104 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 20700 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 20148 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 14260 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19412 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 13616 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23184 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25576 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 23460 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 29164 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 31740 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 32108 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 26496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 30912 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 26680 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 19596 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21896 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 28612 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 30728 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 34316 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 37260 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 37076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 37812 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 39376 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 41584 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 39192 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 39560 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 37812 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 36064 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 35880 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 34684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 35052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 36064 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 30728 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 33304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 33120 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 29164 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 30636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 32200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 34868 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 34500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 33948 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 31740 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 30176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 29072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 47564 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 35696 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 35512 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 36892 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 36892 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 38456 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 39376 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 39560 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 37628 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 36892 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 37076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 42136 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 43792 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 41768 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 41952 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 43056 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 42044 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 40020 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 37628 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 39468 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 42596 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 42596 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 43148 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 41952 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 41860 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 41676 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 41952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 41492 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 41768 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 42044 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 36892 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 27692 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25944 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 26588 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25576 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 26588 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 28980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23368 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 23552 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20424 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19872 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20792 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 22632 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23828 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21344 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 9844 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13156 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13892 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14260 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8280 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 9752 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 9292 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 9108 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 9200 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 10120 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 31740 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 30360 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 26496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 30176 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 22172 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 21988 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 18860 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 28980 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 24564 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 19412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 28980 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 26496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 25484 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 29348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 29164 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 25484 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 25300 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 14168 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 14720 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31740 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23092 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 18584 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 20240 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 19320 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 28888 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 29072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 24472 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 23552 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 21896 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 26312 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 24104 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23368 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 22632 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 22448 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 19136 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l2_in_1__S
timestamp 1679235063
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 34224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 27692 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 25116 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_37.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 34316 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_37.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 32108 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_37.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 23736 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_45.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 33304 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_45.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 30268 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 7360 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 24288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 19320 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 30452 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 40940 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 40756 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 37260 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 28888 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 27508 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 29072 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 35328 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 36892 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 30912 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 39836 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 37628 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 34224 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 35236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 34132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 36892 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 34684 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 34316 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 34316 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 30360 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 34224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 27140 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 29348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 33764 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 28152 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 28888 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 34500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 25944 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 25760 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 34500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 36708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 34316 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 31280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 31740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 27968 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31096 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 29808 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 27968 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 39560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 39192 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 39376 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 47012 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 44528 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 20332 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 22080 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 21896 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 31648 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 41032 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 44712 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 30728 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 34040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 37444 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 44344 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 34316 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 42872 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 42872 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 43056 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 36892 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 37444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 44620 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 44712 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 43608 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 37628 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 37444 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 36708 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 37260 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 42780 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 42504 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 42688 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 40020 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 43240 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 43424 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 36892 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 42136 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 42320 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 41768 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 42044 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 42412 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 34500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 29624 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 29072 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 24472 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23092 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 6532 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 28796 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 19044 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 28980 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 29164 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 24012 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_28.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21988 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 24380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_30.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20608 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_32.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_34.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18768 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 27140 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 27324 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 20976 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_40.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13708 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_42.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15272 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_42.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16468 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 10396 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_48.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14444 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14168 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_50.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16836 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17020 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_58.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14168 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_58.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18952 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 18032 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16836 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16744 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 16836 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14352 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 13616 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 14260 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14260 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10856 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 10672 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 11132 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12328 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13340 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 10764 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 8648 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14444 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 16836 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 16836 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 20700 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_
timestamp 1679235063
transform 1 0 15548 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15180 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 17848 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_
timestamp 1679235063
transform 1 0 17940 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_
timestamp 1679235063
transform 1 0 18308 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__246 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19044 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_
timestamp 1679235063
transform 1 0 18216 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20332 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12696 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_
timestamp 1679235063
transform 1 0 19596 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_
timestamp 1679235063
transform 1 0 15640 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_
timestamp 1679235063
transform 1 0 16744 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11776 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_
timestamp 1679235063
transform 1 0 17572 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_
timestamp 1679235063
transform 1 0 12972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_
timestamp 1679235063
transform 1 0 15732 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__247
timestamp 1679235063
transform 1 0 19412 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 13156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_
timestamp 1679235063
transform 1 0 15364 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_
timestamp 1679235063
transform 1 0 15364 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18124 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 7728 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 8004 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 18124 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_
timestamp 1679235063
transform 1 0 14444 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_
timestamp 1679235063
transform 1 0 19412 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9476 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_
timestamp 1679235063
transform 1 0 12972 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_
timestamp 1679235063
transform 1 0 11684 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__248
timestamp 1679235063
transform 1 0 10212 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_
timestamp 1679235063
transform 1 0 11960 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_
timestamp 1679235063
transform 1 0 12420 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14352 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_
timestamp 1679235063
transform 1 0 15548 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_
timestamp 1679235063
transform 1 0 18308 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_
timestamp 1679235063
transform 1 0 15088 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13156 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_
timestamp 1679235063
transform 1 0 15364 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_
timestamp 1679235063
transform 1 0 14536 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__249
timestamp 1679235063
transform 1 0 9844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_
timestamp 1679235063
transform 1 0 16376 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 11960 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_
timestamp 1679235063
transform 1 0 12972 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_
timestamp 1679235063
transform 1 0 11132 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16468 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 27140 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20884 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 22724 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14536 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 25208 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 23644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 22448 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 21160 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 24288 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 23460 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 19596 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24564 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 24564 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 22172 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 27600 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 18308 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 29072 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 27140 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17940 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1679235063
transform 1 0 19412 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1679235063
transform 1 0 22540 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1679235063
transform 1 0 22540 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1679235063
transform 1 0 17940 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1679235063
transform 1 0 17940 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1679235063
transform 1 0 22448 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1679235063
transform 1 0 22632 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1679235063
transform 1 0 29716 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1679235063
transform 1 0 29624 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1679235063
transform 1 0 34500 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1679235063
transform 1 0 34868 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1679235063
transform 1 0 29808 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1679235063
transform 1 0 30728 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1679235063
transform 1 0 34592 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1679235063
transform 1 0 34868 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17
timestamp 1679235063
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24
timestamp 1679235063
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1679235063
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1679235063
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1679235063
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1679235063
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_96
timestamp 1679235063
transform 1 0 9936 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100
timestamp 1679235063
transform 1 0 10304 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp 1679235063
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132
timestamp 1679235063
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1679235063
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_159 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 15732 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_165 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16284 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1679235063
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1679235063
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1679235063
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1679235063
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_205
timestamp 1679235063
transform 1 0 19964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_211
timestamp 1679235063
transform 1 0 20516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1679235063
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_225
timestamp 1679235063
transform 1 0 21804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_231
timestamp 1679235063
transform 1 0 22356 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_239
timestamp 1679235063
transform 1 0 23092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1679235063
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1679235063
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_275
timestamp 1679235063
transform 1 0 26404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1679235063
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_281
timestamp 1679235063
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_287
timestamp 1679235063
transform 1 0 27508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_295
timestamp 1679235063
transform 1 0 28244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_299
timestamp 1679235063
transform 1 0 28612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_303
timestamp 1679235063
transform 1 0 28980 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1679235063
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1679235063
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_321
timestamp 1679235063
transform 1 0 30636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_326
timestamp 1679235063
transform 1 0 31096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1679235063
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_337
timestamp 1679235063
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_345
timestamp 1679235063
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_349
timestamp 1679235063
transform 1 0 33212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_353
timestamp 1679235063
transform 1 0 33580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1679235063
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_365
timestamp 1679235063
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_372
timestamp 1679235063
transform 1 0 35328 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_376
timestamp 1679235063
transform 1 0 35696 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_388
timestamp 1679235063
transform 1 0 36800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1679235063
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1679235063
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1679235063
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_421
timestamp 1679235063
transform 1 0 39836 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_429
timestamp 1679235063
transform 1 0 40572 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1679235063
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1679235063
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1679235063
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1679235063
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_477
timestamp 1679235063
transform 1 0 44988 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_485
timestamp 1679235063
transform 1 0 45724 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1679235063
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_505
timestamp 1679235063
transform 1 0 47564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1679235063
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1679235063
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_9
timestamp 1679235063
transform 1 0 1932 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_19
timestamp 1679235063
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_31
timestamp 1679235063
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_43
timestamp 1679235063
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1679235063
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1679235063
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1679235063
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1679235063
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1679235063
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1679235063
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1679235063
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1679235063
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1679235063
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_137
timestamp 1679235063
transform 1 0 13708 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_145
timestamp 1679235063
transform 1 0 14444 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1679235063
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1679235063
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_187
timestamp 1679235063
transform 1 0 18308 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_196
timestamp 1679235063
transform 1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_200
timestamp 1679235063
transform 1 0 19504 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1679235063
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1679235063
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_233
timestamp 1679235063
transform 1 0 22540 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_256
timestamp 1679235063
transform 1 0 24656 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_268
timestamp 1679235063
transform 1 0 25760 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_281
timestamp 1679235063
transform 1 0 26956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_289
timestamp 1679235063
transform 1 0 27692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_299
timestamp 1679235063
transform 1 0 28612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_303
timestamp 1679235063
transform 1 0 28980 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_325
timestamp 1679235063
transform 1 0 31004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1679235063
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1679235063
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1679235063
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1679235063
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1679235063
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1679235063
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1679235063
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1679235063
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1679235063
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1679235063
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1679235063
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1679235063
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1679235063
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1679235063
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1679235063
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_461
timestamp 1679235063
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_465
timestamp 1679235063
transform 1 0 43884 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_482
timestamp 1679235063
transform 1 0 45448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1679235063
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_505
timestamp 1679235063
transform 1 0 47564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1679235063
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1679235063
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1679235063
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1679235063
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1679235063
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1679235063
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1679235063
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1679235063
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1679235063
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1679235063
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1679235063
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1679235063
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1679235063
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1679235063
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1679235063
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1679235063
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1679235063
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1679235063
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_165
timestamp 1679235063
transform 1 0 16284 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_170
timestamp 1679235063
transform 1 0 16744 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_178
timestamp 1679235063
transform 1 0 17480 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_182
timestamp 1679235063
transform 1 0 17848 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1679235063
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1679235063
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_207
timestamp 1679235063
transform 1 0 20148 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_215
timestamp 1679235063
transform 1 0 20884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_239
timestamp 1679235063
transform 1 0 23092 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1679235063
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1679235063
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_276
timestamp 1679235063
transform 1 0 26496 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_288
timestamp 1679235063
transform 1 0 27600 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_300
timestamp 1679235063
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1679235063
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1679235063
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1679235063
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1679235063
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1679235063
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1679235063
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1679235063
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_377
timestamp 1679235063
transform 1 0 35788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_387
timestamp 1679235063
transform 1 0 36708 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_391
timestamp 1679235063
transform 1 0 37076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_403
timestamp 1679235063
transform 1 0 38180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_415
timestamp 1679235063
transform 1 0 39284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1679235063
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1679235063
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1679235063
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1679235063
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1679235063
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1679235063
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1679235063
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1679235063
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_505
timestamp 1679235063
transform 1 0 47564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1679235063
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1679235063
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_9
timestamp 1679235063
transform 1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_17
timestamp 1679235063
transform 1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_23
timestamp 1679235063
transform 1 0 3220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_35
timestamp 1679235063
transform 1 0 4324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1679235063
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1679235063
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1679235063
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1679235063
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1679235063
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1679235063
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1679235063
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1679235063
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1679235063
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1679235063
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1679235063
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1679235063
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1679235063
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1679235063
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1679235063
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_181
timestamp 1679235063
transform 1 0 17756 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_208
timestamp 1679235063
transform 1 0 20240 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1679235063
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1679235063
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_247
timestamp 1679235063
transform 1 0 23828 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_251
timestamp 1679235063
transform 1 0 24196 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1679235063
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1679235063
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1679235063
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_304
timestamp 1679235063
transform 1 0 29072 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_316
timestamp 1679235063
transform 1 0 30176 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_328
timestamp 1679235063
transform 1 0 31280 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1679235063
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1679235063
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1679235063
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1679235063
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1679235063
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1679235063
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1679235063
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1679235063
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1679235063
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1679235063
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1679235063
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1679235063
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1679235063
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1679235063
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1679235063
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_485
timestamp 1679235063
transform 1 0 45724 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1679235063
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_505
timestamp 1679235063
transform 1 0 47564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1679235063
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1679235063
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_9
timestamp 1679235063
transform 1 0 1932 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1679235063
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1679235063
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1679235063
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1679235063
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1679235063
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1679235063
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1679235063
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1679235063
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1679235063
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1679235063
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1679235063
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1679235063
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1679235063
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1679235063
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1679235063
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1679235063
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1679235063
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1679235063
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1679235063
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1679235063
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1679235063
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1679235063
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_221
timestamp 1679235063
transform 1 0 21436 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_232
timestamp 1679235063
transform 1 0 22448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_239
timestamp 1679235063
transform 1 0 23092 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_248
timestamp 1679235063
transform 1 0 23920 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_253
timestamp 1679235063
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_261
timestamp 1679235063
transform 1 0 25116 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_283
timestamp 1679235063
transform 1 0 27140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_295
timestamp 1679235063
transform 1 0 28244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1679235063
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1679235063
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1679235063
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1679235063
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1679235063
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1679235063
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1679235063
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1679235063
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1679235063
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_391
timestamp 1679235063
transform 1 0 37076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_397
timestamp 1679235063
transform 1 0 37628 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1679235063
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_409
timestamp 1679235063
transform 1 0 38732 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_417
timestamp 1679235063
transform 1 0 39468 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1679235063
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1679235063
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1679235063
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1679235063
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1679235063
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1679235063
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1679235063
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1679235063
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_501
timestamp 1679235063
transform 1 0 47196 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1679235063
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1679235063
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1679235063
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1679235063
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1679235063
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1679235063
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1679235063
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1679235063
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1679235063
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1679235063
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1679235063
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1679235063
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1679235063
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1679235063
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1679235063
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1679235063
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1679235063
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1679235063
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1679235063
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1679235063
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1679235063
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1679235063
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1679235063
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1679235063
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1679235063
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1679235063
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1679235063
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1679235063
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1679235063
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1679235063
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1679235063
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1679235063
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1679235063
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1679235063
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1679235063
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1679235063
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1679235063
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1679235063
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1679235063
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1679235063
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1679235063
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1679235063
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1679235063
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_393
timestamp 1679235063
transform 1 0 37260 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_396
timestamp 1679235063
transform 1 0 37536 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_402
timestamp 1679235063
transform 1 0 38088 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_410
timestamp 1679235063
transform 1 0 38824 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_414
timestamp 1679235063
transform 1 0 39192 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_426
timestamp 1679235063
transform 1 0 40296 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_438
timestamp 1679235063
transform 1 0 41400 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_446
timestamp 1679235063
transform 1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1679235063
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1679235063
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1679235063
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_485
timestamp 1679235063
transform 1 0 45724 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1679235063
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_505
timestamp 1679235063
transform 1 0 47564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1679235063
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1679235063
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1679235063
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_17
timestamp 1679235063
transform 1 0 2668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1679235063
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1679235063
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1679235063
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1679235063
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1679235063
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1679235063
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1679235063
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1679235063
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1679235063
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1679235063
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1679235063
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1679235063
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1679235063
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1679235063
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1679235063
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1679235063
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1679235063
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1679235063
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1679235063
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1679235063
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1679235063
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1679235063
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1679235063
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1679235063
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1679235063
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1679235063
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1679235063
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1679235063
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1679235063
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1679235063
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1679235063
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1679235063
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1679235063
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1679235063
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1679235063
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1679235063
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1679235063
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1679235063
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1679235063
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1679235063
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1679235063
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1679235063
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1679235063
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1679235063
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1679235063
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1679235063
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1679235063
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_457
timestamp 1679235063
transform 1 0 43148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_461
timestamp 1679235063
transform 1 0 43516 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_466
timestamp 1679235063
transform 1 0 43976 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_474
timestamp 1679235063
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1679235063
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1679235063
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_501
timestamp 1679235063
transform 1 0 47196 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1679235063
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1679235063
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_9
timestamp 1679235063
transform 1 0 1932 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1679235063
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1679235063
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1679235063
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1679235063
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1679235063
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1679235063
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1679235063
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1679235063
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1679235063
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1679235063
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1679235063
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1679235063
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1679235063
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1679235063
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1679235063
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1679235063
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1679235063
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1679235063
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_181
timestamp 1679235063
transform 1 0 17756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_188
timestamp 1679235063
transform 1 0 18400 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_193
timestamp 1679235063
transform 1 0 18860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_205
timestamp 1679235063
transform 1 0 19964 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_212
timestamp 1679235063
transform 1 0 20608 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1679235063
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1679235063
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1679235063
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1679235063
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1679235063
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1679235063
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1679235063
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1679235063
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1679235063
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1679235063
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1679235063
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1679235063
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1679235063
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1679235063
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1679235063
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1679235063
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1679235063
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1679235063
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1679235063
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_399
timestamp 1679235063
transform 1 0 37812 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_403
timestamp 1679235063
transform 1 0 38180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_415
timestamp 1679235063
transform 1 0 39284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_427
timestamp 1679235063
transform 1 0 40388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_439
timestamp 1679235063
transform 1 0 41492 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1679235063
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1679235063
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_461
timestamp 1679235063
transform 1 0 43516 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_469
timestamp 1679235063
transform 1 0 44252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_481
timestamp 1679235063
transform 1 0 45356 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_493
timestamp 1679235063
transform 1 0 46460 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_501
timestamp 1679235063
transform 1 0 47196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_505
timestamp 1679235063
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1679235063
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1679235063
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_9
timestamp 1679235063
transform 1 0 1932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_16
timestamp 1679235063
transform 1 0 2576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1679235063
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1679235063
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1679235063
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1679235063
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1679235063
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1679235063
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1679235063
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1679235063
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1679235063
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1679235063
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1679235063
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1679235063
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1679235063
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1679235063
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1679235063
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_165
timestamp 1679235063
transform 1 0 16284 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_168
timestamp 1679235063
transform 1 0 16560 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_180
timestamp 1679235063
transform 1 0 17664 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_183
timestamp 1679235063
transform 1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1679235063
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1679235063
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_202
timestamp 1679235063
transform 1 0 19688 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_206
timestamp 1679235063
transform 1 0 20056 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_217
timestamp 1679235063
transform 1 0 21068 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_221
timestamp 1679235063
transform 1 0 21436 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_230
timestamp 1679235063
transform 1 0 22264 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_242
timestamp 1679235063
transform 1 0 23368 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1679235063
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1679235063
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1679235063
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1679235063
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1679235063
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1679235063
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1679235063
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_309
timestamp 1679235063
transform 1 0 29532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_317
timestamp 1679235063
transform 1 0 30268 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_326
timestamp 1679235063
transform 1 0 31096 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_330
timestamp 1679235063
transform 1 0 31464 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_342
timestamp 1679235063
transform 1 0 32568 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_354
timestamp 1679235063
transform 1 0 33672 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp 1679235063
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1679235063
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1679235063
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1679235063
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1679235063
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1679235063
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1679235063
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1679235063
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1679235063
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1679235063
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1679235063
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1679235063
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1679235063
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1679235063
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_505
timestamp 1679235063
transform 1 0 47564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1679235063
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1679235063
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_9
timestamp 1679235063
transform 1 0 1932 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_13
timestamp 1679235063
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_25
timestamp 1679235063
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_37
timestamp 1679235063
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1679235063
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1679235063
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1679235063
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1679235063
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1679235063
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1679235063
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1679235063
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1679235063
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1679235063
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1679235063
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1679235063
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_149
timestamp 1679235063
transform 1 0 14812 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_157
timestamp 1679235063
transform 1 0 15548 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_160
timestamp 1679235063
transform 1 0 15824 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1679235063
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1679235063
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_179
timestamp 1679235063
transform 1 0 17572 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_184
timestamp 1679235063
transform 1 0 18032 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_195
timestamp 1679235063
transform 1 0 19044 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_207
timestamp 1679235063
transform 1 0 20148 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_211
timestamp 1679235063
transform 1 0 20516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1679235063
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1679235063
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_235
timestamp 1679235063
transform 1 0 22724 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_247
timestamp 1679235063
transform 1 0 23828 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_259
timestamp 1679235063
transform 1 0 24932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_271
timestamp 1679235063
transform 1 0 26036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1679235063
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1679235063
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1679235063
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_305
timestamp 1679235063
transform 1 0 29164 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_309
timestamp 1679235063
transform 1 0 29532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_313
timestamp 1679235063
transform 1 0 29900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_325
timestamp 1679235063
transform 1 0 31004 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_332
timestamp 1679235063
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1679235063
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_347
timestamp 1679235063
transform 1 0 33028 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_359
timestamp 1679235063
transform 1 0 34132 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_371
timestamp 1679235063
transform 1 0 35236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_383
timestamp 1679235063
transform 1 0 36340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1679235063
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_393
timestamp 1679235063
transform 1 0 37260 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_396
timestamp 1679235063
transform 1 0 37536 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_402
timestamp 1679235063
transform 1 0 38088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_410
timestamp 1679235063
transform 1 0 38824 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_414
timestamp 1679235063
transform 1 0 39192 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_426
timestamp 1679235063
transform 1 0 40296 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_438
timestamp 1679235063
transform 1 0 41400 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_446
timestamp 1679235063
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1679235063
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1679235063
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_473
timestamp 1679235063
transform 1 0 44620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_478
timestamp 1679235063
transform 1 0 45080 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_490
timestamp 1679235063
transform 1 0 46184 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_502
timestamp 1679235063
transform 1 0 47288 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1679235063
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1679235063
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1679235063
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_9
timestamp 1679235063
transform 1 0 1932 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1679235063
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1679235063
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1679235063
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1679235063
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1679235063
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1679235063
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1679235063
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1679235063
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1679235063
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1679235063
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1679235063
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1679235063
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1679235063
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1679235063
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_141
timestamp 1679235063
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_149
timestamp 1679235063
transform 1 0 14812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_153
timestamp 1679235063
transform 1 0 15180 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_164
timestamp 1679235063
transform 1 0 16192 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_169
timestamp 1679235063
transform 1 0 16652 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_179
timestamp 1679235063
transform 1 0 17572 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_192
timestamp 1679235063
transform 1 0 18768 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1679235063
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_208
timestamp 1679235063
transform 1 0 20240 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_218
timestamp 1679235063
transform 1 0 21160 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_240
timestamp 1679235063
transform 1 0 23184 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_246
timestamp 1679235063
transform 1 0 23736 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1679235063
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_263
timestamp 1679235063
transform 1 0 25300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_275
timestamp 1679235063
transform 1 0 26404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_287
timestamp 1679235063
transform 1 0 27508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_291
timestamp 1679235063
transform 1 0 27876 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_294
timestamp 1679235063
transform 1 0 28152 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_302
timestamp 1679235063
transform 1 0 28888 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1679235063
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1679235063
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_319
timestamp 1679235063
transform 1 0 30452 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_323
timestamp 1679235063
transform 1 0 30820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_334
timestamp 1679235063
transform 1 0 31832 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_346
timestamp 1679235063
transform 1 0 32936 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_353
timestamp 1679235063
transform 1 0 33580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_361
timestamp 1679235063
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1679235063
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1679235063
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_389
timestamp 1679235063
transform 1 0 36892 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_395
timestamp 1679235063
transform 1 0 37444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_398
timestamp 1679235063
transform 1 0 37720 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_404
timestamp 1679235063
transform 1 0 38272 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_412
timestamp 1679235063
transform 1 0 39008 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_416
timestamp 1679235063
transform 1 0 39376 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1679235063
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1679235063
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1679235063
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1679235063
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1679235063
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1679235063
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1679235063
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1679235063
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_501
timestamp 1679235063
transform 1 0 47196 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1679235063
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1679235063
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1679235063
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1679235063
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1679235063
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1679235063
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1679235063
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1679235063
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1679235063
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1679235063
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1679235063
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1679235063
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1679235063
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1679235063
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1679235063
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_139
timestamp 1679235063
transform 1 0 13892 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_149
timestamp 1679235063
transform 1 0 14812 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_153
timestamp 1679235063
transform 1 0 15180 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_164
timestamp 1679235063
transform 1 0 16192 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1679235063
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp 1679235063
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_198
timestamp 1679235063
transform 1 0 19320 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1679235063
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_229
timestamp 1679235063
transform 1 0 22172 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_251
timestamp 1679235063
transform 1 0 24196 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_255
timestamp 1679235063
transform 1 0 24564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_266
timestamp 1679235063
transform 1 0 25576 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_272
timestamp 1679235063
transform 1 0 26128 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_281
timestamp 1679235063
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_297
timestamp 1679235063
transform 1 0 28428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_321
timestamp 1679235063
transform 1 0 30636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1679235063
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1679235063
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_359
timestamp 1679235063
transform 1 0 34132 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_365
timestamp 1679235063
transform 1 0 34684 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_376
timestamp 1679235063
transform 1 0 35696 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_388
timestamp 1679235063
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1679235063
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_398
timestamp 1679235063
transform 1 0 37720 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_410
timestamp 1679235063
transform 1 0 38824 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_414
timestamp 1679235063
transform 1 0 39192 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_422
timestamp 1679235063
transform 1 0 39928 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_429
timestamp 1679235063
transform 1 0 40572 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_433
timestamp 1679235063
transform 1 0 40940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_445
timestamp 1679235063
transform 1 0 42044 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1679235063
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_461
timestamp 1679235063
transform 1 0 43516 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_471
timestamp 1679235063
transform 1 0 44436 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_483
timestamp 1679235063
transform 1 0 45540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_502
timestamp 1679235063
transform 1 0 47288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_505
timestamp 1679235063
transform 1 0 47564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1679235063
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1679235063
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_9
timestamp 1679235063
transform 1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_17
timestamp 1679235063
transform 1 0 2668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1679235063
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1679235063
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1679235063
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1679235063
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1679235063
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1679235063
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1679235063
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1679235063
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1679235063
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1679235063
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1679235063
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_121
timestamp 1679235063
transform 1 0 12236 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1679235063
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1679235063
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_163
timestamp 1679235063
transform 1 0 16100 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_170
timestamp 1679235063
transform 1 0 16744 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1679235063
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1679235063
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1679235063
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_232
timestamp 1679235063
transform 1 0 22448 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_236
timestamp 1679235063
transform 1 0 22816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_248
timestamp 1679235063
transform 1 0 23920 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_253
timestamp 1679235063
transform 1 0 24380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_259
timestamp 1679235063
transform 1 0 24932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_271
timestamp 1679235063
transform 1 0 26036 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_278
timestamp 1679235063
transform 1 0 26680 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_290
timestamp 1679235063
transform 1 0 27784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_303
timestamp 1679235063
transform 1 0 28980 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1679235063
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1679235063
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_314
timestamp 1679235063
transform 1 0 29992 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_320
timestamp 1679235063
transform 1 0 30544 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_342
timestamp 1679235063
transform 1 0 32568 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_355
timestamp 1679235063
transform 1 0 33764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_361
timestamp 1679235063
transform 1 0 34316 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1679235063
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_376
timestamp 1679235063
transform 1 0 35696 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_382
timestamp 1679235063
transform 1 0 36248 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_389
timestamp 1679235063
transform 1 0 36892 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_400
timestamp 1679235063
transform 1 0 37904 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_412
timestamp 1679235063
transform 1 0 39008 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_418
timestamp 1679235063
transform 1 0 39560 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_423
timestamp 1679235063
transform 1 0 40020 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_435
timestamp 1679235063
transform 1 0 41124 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_447
timestamp 1679235063
transform 1 0 42228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_459
timestamp 1679235063
transform 1 0 43332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_471
timestamp 1679235063
transform 1 0 44436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1679235063
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1679235063
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1679235063
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_501
timestamp 1679235063
transform 1 0 47196 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1679235063
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1679235063
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_9
timestamp 1679235063
transform 1 0 1932 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1679235063
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1679235063
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1679235063
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1679235063
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1679235063
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1679235063
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1679235063
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1679235063
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1679235063
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1679235063
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1679235063
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 1679235063
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_121
timestamp 1679235063
transform 1 0 12236 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_132
timestamp 1679235063
transform 1 0 13248 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_156
timestamp 1679235063
transform 1 0 15456 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_161
timestamp 1679235063
transform 1 0 15916 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1679235063
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1679235063
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1679235063
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_218
timestamp 1679235063
transform 1 0 21160 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1679235063
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_236
timestamp 1679235063
transform 1 0 22816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_241
timestamp 1679235063
transform 1 0 23276 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_264
timestamp 1679235063
transform 1 0 25392 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1679235063
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_285
timestamp 1679235063
transform 1 0 27324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_307
timestamp 1679235063
transform 1 0 29348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_331
timestamp 1679235063
transform 1 0 31556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1679235063
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_337
timestamp 1679235063
transform 1 0 32108 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_340
timestamp 1679235063
transform 1 0 32384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_351
timestamp 1679235063
transform 1 0 33396 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_355
timestamp 1679235063
transform 1 0 33764 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_376
timestamp 1679235063
transform 1 0 35696 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_388
timestamp 1679235063
transform 1 0 36800 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_395
timestamp 1679235063
transform 1 0 37444 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_401
timestamp 1679235063
transform 1 0 37996 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_413
timestamp 1679235063
transform 1 0 39100 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_425
timestamp 1679235063
transform 1 0 40204 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_437
timestamp 1679235063
transform 1 0 41308 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_445
timestamp 1679235063
transform 1 0 42044 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1679235063
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1679235063
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1679235063
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1679235063
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1679235063
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1679235063
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_505
timestamp 1679235063
transform 1 0 47564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1679235063
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1679235063
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1679235063
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1679235063
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1679235063
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1679235063
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1679235063
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1679235063
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1679235063
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1679235063
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1679235063
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1679235063
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_109
timestamp 1679235063
transform 1 0 11132 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_125
timestamp 1679235063
transform 1 0 12604 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1679235063
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1679235063
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_166
timestamp 1679235063
transform 1 0 16376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_190
timestamp 1679235063
transform 1 0 18584 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_199
timestamp 1679235063
transform 1 0 19412 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_204
timestamp 1679235063
transform 1 0 19872 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_208
timestamp 1679235063
transform 1 0 20240 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_229
timestamp 1679235063
transform 1 0 22172 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_244
timestamp 1679235063
transform 1 0 23552 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1679235063
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1679235063
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_275
timestamp 1679235063
transform 1 0 26404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_279
timestamp 1679235063
transform 1 0 26772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_301
timestamp 1679235063
transform 1 0 28796 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_305
timestamp 1679235063
transform 1 0 29164 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1679235063
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_314
timestamp 1679235063
transform 1 0 29992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_338
timestamp 1679235063
transform 1 0 32200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_345
timestamp 1679235063
transform 1 0 32844 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_349
timestamp 1679235063
transform 1 0 33212 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_359
timestamp 1679235063
transform 1 0 34132 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1679235063
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1679235063
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_387
timestamp 1679235063
transform 1 0 36708 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_399
timestamp 1679235063
transform 1 0 37812 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_407
timestamp 1679235063
transform 1 0 38548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_411
timestamp 1679235063
transform 1 0 38916 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1679235063
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_421
timestamp 1679235063
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_427
timestamp 1679235063
transform 1 0 40388 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_431
timestamp 1679235063
transform 1 0 40756 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_443
timestamp 1679235063
transform 1 0 41860 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_455
timestamp 1679235063
transform 1 0 42964 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_467
timestamp 1679235063
transform 1 0 44068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_473
timestamp 1679235063
transform 1 0 44620 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1679235063
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_505
timestamp 1679235063
transform 1 0 47564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1679235063
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1679235063
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_9
timestamp 1679235063
transform 1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_17
timestamp 1679235063
transform 1 0 2668 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 1679235063
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1679235063
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1679235063
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1679235063
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1679235063
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1679235063
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1679235063
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1679235063
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_105
timestamp 1679235063
transform 1 0 10764 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_109
timestamp 1679235063
transform 1 0 11132 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1679235063
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_116
timestamp 1679235063
transform 1 0 11776 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_127
timestamp 1679235063
transform 1 0 12788 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_140
timestamp 1679235063
transform 1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1679235063
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1679235063
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_169
timestamp 1679235063
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1679235063
transform 1 0 17756 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_185
timestamp 1679235063
transform 1 0 18124 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1679235063
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1679235063
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1679235063
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1679235063
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_247
timestamp 1679235063
transform 1 0 23828 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_260
timestamp 1679235063
transform 1 0 25024 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_268
timestamp 1679235063
transform 1 0 25760 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1679235063
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1679235063
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_292
timestamp 1679235063
transform 1 0 27968 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_305
timestamp 1679235063
transform 1 0 29164 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_309
timestamp 1679235063
transform 1 0 29532 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_320
timestamp 1679235063
transform 1 0 30544 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_333
timestamp 1679235063
transform 1 0 31740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1679235063
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_348
timestamp 1679235063
transform 1 0 33120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_352
timestamp 1679235063
transform 1 0 33488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_376
timestamp 1679235063
transform 1 0 35696 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_389
timestamp 1679235063
transform 1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1679235063
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_403
timestamp 1679235063
transform 1 0 38180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_415
timestamp 1679235063
transform 1 0 39284 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_423
timestamp 1679235063
transform 1 0 40020 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_427
timestamp 1679235063
transform 1 0 40388 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_431
timestamp 1679235063
transform 1 0 40756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_443
timestamp 1679235063
transform 1 0 41860 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1679235063
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1679235063
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1679235063
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1679235063
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1679235063
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1679235063
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1679235063
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_505
timestamp 1679235063
transform 1 0 47564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1679235063
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1679235063
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_9
timestamp 1679235063
transform 1 0 1932 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1679235063
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1679235063
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1679235063
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1679235063
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1679235063
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1679235063
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1679235063
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1679235063
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1679235063
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_97
timestamp 1679235063
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_107
timestamp 1679235063
transform 1 0 10948 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_129
timestamp 1679235063
transform 1 0 12972 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_136
timestamp 1679235063
transform 1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1679235063
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_144
timestamp 1679235063
transform 1 0 14352 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_155
timestamp 1679235063
transform 1 0 15364 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_168
timestamp 1679235063
transform 1 0 16560 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_181
timestamp 1679235063
transform 1 0 17756 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1679235063
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_197
timestamp 1679235063
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_200
timestamp 1679235063
transform 1 0 19504 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_205
timestamp 1679235063
transform 1 0 19964 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_229
timestamp 1679235063
transform 1 0 22172 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_236
timestamp 1679235063
transform 1 0 22816 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_240
timestamp 1679235063
transform 1 0 23184 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1679235063
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1679235063
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_275
timestamp 1679235063
transform 1 0 26404 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_279
timestamp 1679235063
transform 1 0 26772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_300
timestamp 1679235063
transform 1 0 28704 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1679235063
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_322
timestamp 1679235063
transform 1 0 30728 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_346
timestamp 1679235063
transform 1 0 32936 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_350
timestamp 1679235063
transform 1 0 33304 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_361
timestamp 1679235063
transform 1 0 34316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_373
timestamp 1679235063
transform 1 0 35420 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_399
timestamp 1679235063
transform 1 0 37812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_411
timestamp 1679235063
transform 1 0 38916 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_418
timestamp 1679235063
transform 1 0 39560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_421
timestamp 1679235063
transform 1 0 39836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_427
timestamp 1679235063
transform 1 0 40388 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_435
timestamp 1679235063
transform 1 0 41124 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_442
timestamp 1679235063
transform 1 0 41768 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_454
timestamp 1679235063
transform 1 0 42872 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_466
timestamp 1679235063
transform 1 0 43976 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_474
timestamp 1679235063
transform 1 0 44712 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_477
timestamp 1679235063
transform 1 0 44988 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_487
timestamp 1679235063
transform 1 0 45908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_499
timestamp 1679235063
transform 1 0 47012 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_507
timestamp 1679235063
transform 1 0 47748 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1679235063
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1679235063
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1679235063
transform 1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_16
timestamp 1679235063
transform 1 0 2576 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_20
timestamp 1679235063
transform 1 0 2944 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_32
timestamp 1679235063
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_44
timestamp 1679235063
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1679235063
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1679235063
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1679235063
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_93
timestamp 1679235063
transform 1 0 9660 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_100
timestamp 1679235063
transform 1 0 10304 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1679235063
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1679235063
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1679235063
transform 1 0 11960 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_145
timestamp 1679235063
transform 1 0 14444 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_150
timestamp 1679235063
transform 1 0 14904 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_161
timestamp 1679235063
transform 1 0 15916 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1679235063
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_191
timestamp 1679235063
transform 1 0 18676 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_197
timestamp 1679235063
transform 1 0 19228 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_208
timestamp 1679235063
transform 1 0 20240 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_212
timestamp 1679235063
transform 1 0 20608 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1679235063
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_231
timestamp 1679235063
transform 1 0 22356 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1679235063
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_268
timestamp 1679235063
transform 1 0 25760 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_272
timestamp 1679235063
transform 1 0 26128 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1679235063
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1679235063
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_292
timestamp 1679235063
transform 1 0 27968 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_296
timestamp 1679235063
transform 1 0 28336 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_319
timestamp 1679235063
transform 1 0 30452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_332
timestamp 1679235063
transform 1 0 31648 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1679235063
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_348
timestamp 1679235063
transform 1 0 33120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_361
timestamp 1679235063
transform 1 0 34316 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_367
timestamp 1679235063
transform 1 0 34868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1679235063
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1679235063
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_404
timestamp 1679235063
transform 1 0 38272 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_417
timestamp 1679235063
transform 1 0 39468 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_429
timestamp 1679235063
transform 1 0 40572 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_433
timestamp 1679235063
transform 1 0 40940 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_445
timestamp 1679235063
transform 1 0 42044 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1679235063
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1679235063
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_473
timestamp 1679235063
transform 1 0 44620 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_481
timestamp 1679235063
transform 1 0 45356 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_493
timestamp 1679235063
transform 1 0 46460 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_501
timestamp 1679235063
transform 1 0 47196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_505
timestamp 1679235063
transform 1 0 47564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1679235063
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1679235063
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_15
timestamp 1679235063
transform 1 0 2484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_21
timestamp 1679235063
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1679235063
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1679235063
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1679235063
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1679235063
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1679235063
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1679235063
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1679235063
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1679235063
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1679235063
transform 1 0 9384 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_100
timestamp 1679235063
transform 1 0 10304 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_124
timestamp 1679235063
transform 1 0 12512 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_128
timestamp 1679235063
transform 1 0 12880 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1679235063
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_141
timestamp 1679235063
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_165
timestamp 1679235063
transform 1 0 16284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_169
timestamp 1679235063
transform 1 0 16652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1679235063
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1679235063
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1679235063
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1679235063
transform 1 0 20424 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_214
timestamp 1679235063
transform 1 0 20792 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_224
timestamp 1679235063
transform 1 0 21712 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_237
timestamp 1679235063
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1679235063
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1679235063
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_275
timestamp 1679235063
transform 1 0 26404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_279
timestamp 1679235063
transform 1 0 26772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_290
timestamp 1679235063
transform 1 0 27784 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_294
timestamp 1679235063
transform 1 0 28152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1679235063
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1679235063
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_331
timestamp 1679235063
transform 1 0 31556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_335
timestamp 1679235063
transform 1 0 31924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_358
timestamp 1679235063
transform 1 0 34040 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1679235063
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_387
timestamp 1679235063
transform 1 0 36708 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_400
timestamp 1679235063
transform 1 0 37904 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_412
timestamp 1679235063
transform 1 0 39008 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1679235063
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_427
timestamp 1679235063
transform 1 0 40388 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_434
timestamp 1679235063
transform 1 0 41032 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_441
timestamp 1679235063
transform 1 0 41676 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_453
timestamp 1679235063
transform 1 0 42780 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_465
timestamp 1679235063
transform 1 0 43884 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_473
timestamp 1679235063
transform 1 0 44620 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_477
timestamp 1679235063
transform 1 0 44988 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_485
timestamp 1679235063
transform 1 0 45724 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_490
timestamp 1679235063
transform 1 0 46184 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_502
timestamp 1679235063
transform 1 0 47288 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_508
timestamp 1679235063
transform 1 0 47840 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1679235063
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1679235063
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_15
timestamp 1679235063
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_22
timestamp 1679235063
transform 1 0 3128 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_26
timestamp 1679235063
transform 1 0 3496 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_38
timestamp 1679235063
transform 1 0 4600 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1679235063
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1679235063
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1679235063
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1679235063
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_93
timestamp 1679235063
transform 1 0 9660 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_99
timestamp 1679235063
transform 1 0 10212 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1679235063
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1679235063
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_124
timestamp 1679235063
transform 1 0 12512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_128
timestamp 1679235063
transform 1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_150
timestamp 1679235063
transform 1 0 14904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1679235063
transform 1 0 15364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1679235063
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1679235063
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_192
timestamp 1679235063
transform 1 0 18768 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_205
timestamp 1679235063
transform 1 0 19964 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_210
timestamp 1679235063
transform 1 0 20424 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_221
timestamp 1679235063
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1679235063
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_230
timestamp 1679235063
transform 1 0 22264 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_234
timestamp 1679235063
transform 1 0 22632 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_244
timestamp 1679235063
transform 1 0 23552 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_268
timestamp 1679235063
transform 1 0 25760 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_275
timestamp 1679235063
transform 1 0 26404 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1679235063
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_306
timestamp 1679235063
transform 1 0 29256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_321
timestamp 1679235063
transform 1 0 30636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1679235063
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1679235063
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_359
timestamp 1679235063
transform 1 0 34132 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_374
timestamp 1679235063
transform 1 0 35512 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_387
timestamp 1679235063
transform 1 0 36708 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1679235063
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1679235063
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_418
timestamp 1679235063
transform 1 0 39560 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_430
timestamp 1679235063
transform 1 0 40664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_438
timestamp 1679235063
transform 1 0 41400 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_444
timestamp 1679235063
transform 1 0 41952 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1679235063
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1679235063
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1679235063
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_485
timestamp 1679235063
transform 1 0 45724 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_491
timestamp 1679235063
transform 1 0 46276 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1679235063
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_505
timestamp 1679235063
transform 1 0 47564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1679235063
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1679235063
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1679235063
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1679235063
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1679235063
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1679235063
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1679235063
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1679235063
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1679235063
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1679235063
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1679235063
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_97
timestamp 1679235063
transform 1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_102
timestamp 1679235063
transform 1 0 10488 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_127
timestamp 1679235063
transform 1 0 12788 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_133
timestamp 1679235063
transform 1 0 13340 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1679235063
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1679235063
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_147
timestamp 1679235063
transform 1 0 14628 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1679235063
transform 1 0 14996 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1679235063
transform 1 0 16008 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_175
timestamp 1679235063
transform 1 0 17204 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_188
timestamp 1679235063
transform 1 0 18400 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_197
timestamp 1679235063
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_209
timestamp 1679235063
transform 1 0 20332 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_222
timestamp 1679235063
transform 1 0 21528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_235
timestamp 1679235063
transform 1 0 22724 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_248
timestamp 1679235063
transform 1 0 23920 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_253
timestamp 1679235063
transform 1 0 24380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_256
timestamp 1679235063
transform 1 0 24656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_267
timestamp 1679235063
transform 1 0 25668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_279
timestamp 1679235063
transform 1 0 26772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_291
timestamp 1679235063
transform 1 0 27876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_295
timestamp 1679235063
transform 1 0 28244 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_304
timestamp 1679235063
transform 1 0 29072 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1679235063
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_320
timestamp 1679235063
transform 1 0 30544 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_324
timestamp 1679235063
transform 1 0 30912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_348
timestamp 1679235063
transform 1 0 33120 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_361
timestamp 1679235063
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1679235063
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_378
timestamp 1679235063
transform 1 0 35880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_382
timestamp 1679235063
transform 1 0 36248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_404
timestamp 1679235063
transform 1 0 38272 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_416
timestamp 1679235063
transform 1 0 39376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_421
timestamp 1679235063
transform 1 0 39836 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_431
timestamp 1679235063
transform 1 0 40756 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_443
timestamp 1679235063
transform 1 0 41860 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_455
timestamp 1679235063
transform 1 0 42964 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_467
timestamp 1679235063
transform 1 0 44068 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1679235063
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1679235063
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1679235063
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_501
timestamp 1679235063
transform 1 0 47196 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1679235063
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1679235063
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1679235063
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_29
timestamp 1679235063
transform 1 0 3772 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1679235063
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1679235063
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1679235063
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1679235063
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1679235063
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_81
timestamp 1679235063
transform 1 0 8556 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_89
timestamp 1679235063
transform 1 0 9292 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_93
timestamp 1679235063
transform 1 0 9660 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_98
timestamp 1679235063
transform 1 0 10120 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1679235063
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1679235063
transform 1 0 11500 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_116
timestamp 1679235063
transform 1 0 11776 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_127
timestamp 1679235063
transform 1 0 12788 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_131
timestamp 1679235063
transform 1 0 13156 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_154
timestamp 1679235063
transform 1 0 15272 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1679235063
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_173
timestamp 1679235063
transform 1 0 17020 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_178
timestamp 1679235063
transform 1 0 17480 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_191
timestamp 1679235063
transform 1 0 18676 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1679235063
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1679235063
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1679235063
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_247
timestamp 1679235063
transform 1 0 23828 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_254
timestamp 1679235063
transform 1 0 24472 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1679235063
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1679235063
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_303
timestamp 1679235063
transform 1 0 28980 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_327
timestamp 1679235063
transform 1 0 31188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1679235063
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1679235063
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_359
timestamp 1679235063
transform 1 0 34132 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_372
timestamp 1679235063
transform 1 0 35328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_385
timestamp 1679235063
transform 1 0 36524 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1679235063
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1679235063
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_404
timestamp 1679235063
transform 1 0 38272 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_417
timestamp 1679235063
transform 1 0 39468 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_429
timestamp 1679235063
transform 1 0 40572 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_435
timestamp 1679235063
transform 1 0 41124 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_440
timestamp 1679235063
transform 1 0 41584 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_444
timestamp 1679235063
transform 1 0 41952 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1679235063
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1679235063
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_473
timestamp 1679235063
transform 1 0 44620 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_480
timestamp 1679235063
transform 1 0 45264 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_487
timestamp 1679235063
transform 1 0 45908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_499
timestamp 1679235063
transform 1 0 47012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1679235063
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_505
timestamp 1679235063
transform 1 0 47564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_509
timestamp 1679235063
transform 1 0 47932 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_512
timestamp 1679235063
transform 1 0 48208 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_517
timestamp 1679235063
transform 1 0 48668 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1679235063
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1679235063
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1679235063
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1679235063
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1679235063
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1679235063
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1679235063
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1679235063
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1679235063
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1679235063
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_89
timestamp 1679235063
transform 1 0 9292 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_95
timestamp 1679235063
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_103
timestamp 1679235063
transform 1 0 10580 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_107
timestamp 1679235063
transform 1 0 10948 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_112
timestamp 1679235063
transform 1 0 11408 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_125
timestamp 1679235063
transform 1 0 12604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1679235063
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1679235063
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1679235063
transform 1 0 15272 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_167
timestamp 1679235063
transform 1 0 16468 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_180
timestamp 1679235063
transform 1 0 17664 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_184
timestamp 1679235063
transform 1 0 18032 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1679235063
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_199
timestamp 1679235063
transform 1 0 19412 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_210
timestamp 1679235063
transform 1 0 20424 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_214
timestamp 1679235063
transform 1 0 20792 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_240
timestamp 1679235063
transform 1 0 23184 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1679235063
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_263
timestamp 1679235063
transform 1 0 25300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_287
timestamp 1679235063
transform 1 0 27508 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_300
timestamp 1679235063
transform 1 0 28704 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1679235063
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_320
timestamp 1679235063
transform 1 0 30544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_333
timestamp 1679235063
transform 1 0 31740 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_346
timestamp 1679235063
transform 1 0 32936 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_359
timestamp 1679235063
transform 1 0 34132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1679235063
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1679235063
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_387
timestamp 1679235063
transform 1 0 36708 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_411
timestamp 1679235063
transform 1 0 38916 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1679235063
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_421
timestamp 1679235063
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_431
timestamp 1679235063
transform 1 0 40756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_443
timestamp 1679235063
transform 1 0 41860 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_447
timestamp 1679235063
transform 1 0 42228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_459
timestamp 1679235063
transform 1 0 43332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_471
timestamp 1679235063
transform 1 0 44436 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1679235063
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1679235063
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1679235063
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1679235063
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_513
timestamp 1679235063
transform 1 0 48300 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_519
timestamp 1679235063
transform 1 0 48852 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1679235063
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1679235063
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_21
timestamp 1679235063
transform 1 0 3036 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_33
timestamp 1679235063
transform 1 0 4140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_45
timestamp 1679235063
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1679235063
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1679235063
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1679235063
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_81
timestamp 1679235063
transform 1 0 8556 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_89
timestamp 1679235063
transform 1 0 9292 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_100
timestamp 1679235063
transform 1 0 10304 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_104
timestamp 1679235063
transform 1 0 10672 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1679235063
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_113
timestamp 1679235063
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_125
timestamp 1679235063
transform 1 0 12604 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_149
timestamp 1679235063
transform 1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_156
timestamp 1679235063
transform 1 0 15456 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1679235063
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1679235063
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_180
timestamp 1679235063
transform 1 0 17664 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_185
timestamp 1679235063
transform 1 0 18124 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_196
timestamp 1679235063
transform 1 0 19136 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_209
timestamp 1679235063
transform 1 0 20332 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1679235063
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_225
timestamp 1679235063
transform 1 0 21804 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_228
timestamp 1679235063
transform 1 0 22080 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_233
timestamp 1679235063
transform 1 0 22540 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_246
timestamp 1679235063
transform 1 0 23736 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_259
timestamp 1679235063
transform 1 0 24932 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_267
timestamp 1679235063
transform 1 0 25668 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1679235063
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_291
timestamp 1679235063
transform 1 0 27876 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_313
timestamp 1679235063
transform 1 0 29900 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_326
timestamp 1679235063
transform 1 0 31096 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_330
timestamp 1679235063
transform 1 0 31464 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1679235063
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1679235063
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_348
timestamp 1679235063
transform 1 0 33120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_361
timestamp 1679235063
transform 1 0 34316 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_374
timestamp 1679235063
transform 1 0 35512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_387
timestamp 1679235063
transform 1 0 36708 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1679235063
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1679235063
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_415
timestamp 1679235063
transform 1 0 39284 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_428
timestamp 1679235063
transform 1 0 40480 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_440
timestamp 1679235063
transform 1 0 41584 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 1679235063
transform 1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_449
timestamp 1679235063
transform 1 0 42412 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_454
timestamp 1679235063
transform 1 0 42872 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_466
timestamp 1679235063
transform 1 0 43976 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_478
timestamp 1679235063
transform 1 0 45080 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_490
timestamp 1679235063
transform 1 0 46184 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_502
timestamp 1679235063
transform 1 0 47288 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1679235063
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_519
timestamp 1679235063
transform 1 0 48852 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1679235063
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1679235063
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1679235063
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1679235063
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1679235063
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1679235063
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1679235063
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_57
timestamp 1679235063
transform 1 0 6348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_62
timestamp 1679235063
transform 1 0 6808 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_74
timestamp 1679235063
transform 1 0 7912 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_80
timestamp 1679235063
transform 1 0 8464 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1679235063
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_87
timestamp 1679235063
transform 1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1679235063
transform 1 0 9660 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_98
timestamp 1679235063
transform 1 0 10120 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_103
timestamp 1679235063
transform 1 0 10580 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_125
timestamp 1679235063
transform 1 0 12604 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1679235063
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1679235063
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_151
timestamp 1679235063
transform 1 0 14996 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_164
timestamp 1679235063
transform 1 0 16192 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_169
timestamp 1679235063
transform 1 0 16652 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_180
timestamp 1679235063
transform 1 0 17664 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_184
timestamp 1679235063
transform 1 0 18032 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1679235063
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_201
timestamp 1679235063
transform 1 0 19596 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1679235063
transform 1 0 20608 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_216
timestamp 1679235063
transform 1 0 20976 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_227
timestamp 1679235063
transform 1 0 21988 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_234
timestamp 1679235063
transform 1 0 22632 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_247
timestamp 1679235063
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1679235063
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_253
timestamp 1679235063
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_265
timestamp 1679235063
transform 1 0 25484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_278
timestamp 1679235063
transform 1 0 26680 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_284
timestamp 1679235063
transform 1 0 27232 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_295
timestamp 1679235063
transform 1 0 28244 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1679235063
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_309
timestamp 1679235063
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_315
timestamp 1679235063
transform 1 0 30084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_339
timestamp 1679235063
transform 1 0 32292 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_352
timestamp 1679235063
transform 1 0 33488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_359
timestamp 1679235063
transform 1 0 34132 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1679235063
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1679235063
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_387
timestamp 1679235063
transform 1 0 36708 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_395
timestamp 1679235063
transform 1 0 37444 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_418
timestamp 1679235063
transform 1 0 39560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_421
timestamp 1679235063
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_443
timestamp 1679235063
transform 1 0 41860 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_455
timestamp 1679235063
transform 1 0 42964 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_467
timestamp 1679235063
transform 1 0 44068 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1679235063
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1679235063
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1679235063
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1679235063
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_513
timestamp 1679235063
transform 1 0 48300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_517
timestamp 1679235063
transform 1 0 48668 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_520
timestamp 1679235063
transform 1 0 48944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1679235063
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1679235063
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1679235063
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1679235063
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1679235063
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1679235063
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1679235063
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_69
timestamp 1679235063
transform 1 0 7452 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_84
timestamp 1679235063
transform 1 0 8832 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_92
timestamp 1679235063
transform 1 0 9568 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_100
timestamp 1679235063
transform 1 0 10304 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_106
timestamp 1679235063
transform 1 0 10856 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1679235063
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_116
timestamp 1679235063
transform 1 0 11776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_127
timestamp 1679235063
transform 1 0 12788 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_140
timestamp 1679235063
transform 1 0 13984 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1679235063
transform 1 0 15180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1679235063
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1679235063
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_175
timestamp 1679235063
transform 1 0 17204 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_191
timestamp 1679235063
transform 1 0 18676 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_216
timestamp 1679235063
transform 1 0 20976 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_220
timestamp 1679235063
transform 1 0 21344 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1679235063
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_235
timestamp 1679235063
transform 1 0 22724 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_248
timestamp 1679235063
transform 1 0 23920 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_252
timestamp 1679235063
transform 1 0 24288 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_275
timestamp 1679235063
transform 1 0 26404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1679235063
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1679235063
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_292
timestamp 1679235063
transform 1 0 27968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_316
timestamp 1679235063
transform 1 0 30176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_329
timestamp 1679235063
transform 1 0 31372 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1679235063
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1679235063
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_348
timestamp 1679235063
transform 1 0 33120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_361
timestamp 1679235063
transform 1 0 34316 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_367
timestamp 1679235063
transform 1 0 34868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1679235063
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_401
timestamp 1679235063
transform 1 0 37996 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_423
timestamp 1679235063
transform 1 0 40020 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_427
timestamp 1679235063
transform 1 0 40388 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_437
timestamp 1679235063
transform 1 0 41308 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_445
timestamp 1679235063
transform 1 0 42044 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_449
timestamp 1679235063
transform 1 0 42412 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_459
timestamp 1679235063
transform 1 0 43332 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_471
timestamp 1679235063
transform 1 0 44436 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_483
timestamp 1679235063
transform 1 0 45540 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_495
timestamp 1679235063
transform 1 0 46644 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1679235063
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1679235063
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_519
timestamp 1679235063
transform 1 0 48852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1679235063
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1679235063
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1679235063
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1679235063
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1679235063
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_34
timestamp 1679235063
transform 1 0 4232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_41
timestamp 1679235063
transform 1 0 4876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_48
timestamp 1679235063
transform 1 0 5520 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_56
timestamp 1679235063
transform 1 0 6256 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_62
timestamp 1679235063
transform 1 0 6808 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_70
timestamp 1679235063
transform 1 0 7544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1679235063
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_87
timestamp 1679235063
transform 1 0 9108 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_93
timestamp 1679235063
transform 1 0 9660 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_105
timestamp 1679235063
transform 1 0 10764 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_118
timestamp 1679235063
transform 1 0 11960 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_125
timestamp 1679235063
transform 1 0 12604 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1679235063
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_143
timestamp 1679235063
transform 1 0 14260 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1679235063
transform 1 0 15272 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_158
timestamp 1679235063
transform 1 0 15640 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_167
timestamp 1679235063
transform 1 0 16468 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_179
timestamp 1679235063
transform 1 0 17572 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1679235063
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1679235063
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_208
timestamp 1679235063
transform 1 0 20240 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_212
timestamp 1679235063
transform 1 0 20608 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1679235063
transform 1 0 20884 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_237
timestamp 1679235063
transform 1 0 22908 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1679235063
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1679235063
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_258
timestamp 1679235063
transform 1 0 24840 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_264
timestamp 1679235063
transform 1 0 25392 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_286
timestamp 1679235063
transform 1 0 27416 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_290
timestamp 1679235063
transform 1 0 27784 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_294
timestamp 1679235063
transform 1 0 28152 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1679235063
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1679235063
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_320
timestamp 1679235063
transform 1 0 30544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_328
timestamp 1679235063
transform 1 0 31280 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_351
timestamp 1679235063
transform 1 0 33396 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_358
timestamp 1679235063
transform 1 0 34040 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1679235063
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_378
timestamp 1679235063
transform 1 0 35880 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_391
timestamp 1679235063
transform 1 0 37076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_395
timestamp 1679235063
transform 1 0 37444 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1679235063
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_421
timestamp 1679235063
transform 1 0 39836 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_431
timestamp 1679235063
transform 1 0 40756 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_443
timestamp 1679235063
transform 1 0 41860 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_455
timestamp 1679235063
transform 1 0 42964 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_467
timestamp 1679235063
transform 1 0 44068 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1679235063
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1679235063
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1679235063
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1679235063
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_513
timestamp 1679235063
transform 1 0 48300 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_519
timestamp 1679235063
transform 1 0 48852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1679235063
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1679235063
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_21
timestamp 1679235063
transform 1 0 3036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_29
timestamp 1679235063
transform 1 0 3772 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_34
timestamp 1679235063
transform 1 0 4232 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_43
timestamp 1679235063
transform 1 0 5060 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_50
timestamp 1679235063
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1679235063
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_69
timestamp 1679235063
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_76
timestamp 1679235063
transform 1 0 8096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_83
timestamp 1679235063
transform 1 0 8740 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_90
timestamp 1679235063
transform 1 0 9384 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_97
timestamp 1679235063
transform 1 0 10028 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1679235063
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1679235063
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_119
timestamp 1679235063
transform 1 0 12052 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_124
timestamp 1679235063
transform 1 0 12512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_135
timestamp 1679235063
transform 1 0 13524 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_143
timestamp 1679235063
transform 1 0 14260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_153
timestamp 1679235063
transform 1 0 15180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1679235063
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_171
timestamp 1679235063
transform 1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_194
timestamp 1679235063
transform 1 0 18952 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_218
timestamp 1679235063
transform 1 0 21160 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1679235063
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_230
timestamp 1679235063
transform 1 0 22264 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_254
timestamp 1679235063
transform 1 0 24472 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_267
timestamp 1679235063
transform 1 0 25668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_274
timestamp 1679235063
transform 1 0 26312 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_283
timestamp 1679235063
transform 1 0 27140 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_294
timestamp 1679235063
transform 1 0 28152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_298
timestamp 1679235063
transform 1 0 28520 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_308
timestamp 1679235063
transform 1 0 29440 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_314
timestamp 1679235063
transform 1 0 29992 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_325
timestamp 1679235063
transform 1 0 31004 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_332
timestamp 1679235063
transform 1 0 31648 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1679235063
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_359
timestamp 1679235063
transform 1 0 34132 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_363
timestamp 1679235063
transform 1 0 34500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_375
timestamp 1679235063
transform 1 0 35604 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_388
timestamp 1679235063
transform 1 0 36800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1679235063
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_404
timestamp 1679235063
transform 1 0 38272 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_408
timestamp 1679235063
transform 1 0 38640 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_430
timestamp 1679235063
transform 1 0 40664 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_442
timestamp 1679235063
transform 1 0 41768 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_446
timestamp 1679235063
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1679235063
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1679235063
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1679235063
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1679235063
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1679235063
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1679235063
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1679235063
transform 1 0 47564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_513
timestamp 1679235063
transform 1 0 48300 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_517
timestamp 1679235063
transform 1 0 48668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1679235063
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1679235063
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1679235063
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1679235063
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_29
timestamp 1679235063
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_43
timestamp 1679235063
transform 1 0 5060 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1679235063
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1679235063
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_75
timestamp 1679235063
transform 1 0 8004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1679235063
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_85
timestamp 1679235063
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_91
timestamp 1679235063
transform 1 0 9476 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_104
timestamp 1679235063
transform 1 0 10672 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_128
timestamp 1679235063
transform 1 0 12880 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_132
timestamp 1679235063
transform 1 0 13248 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1679235063
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1679235063
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_163
timestamp 1679235063
transform 1 0 16100 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_168
timestamp 1679235063
transform 1 0 16560 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_179
timestamp 1679235063
transform 1 0 17572 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1679235063
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1679235063
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_202
timestamp 1679235063
transform 1 0 19688 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_206
timestamp 1679235063
transform 1 0 20056 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_227
timestamp 1679235063
transform 1 0 21988 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_231
timestamp 1679235063
transform 1 0 22356 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_243
timestamp 1679235063
transform 1 0 23460 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1679235063
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1679235063
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_264
timestamp 1679235063
transform 1 0 25392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_277
timestamp 1679235063
transform 1 0 26588 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_281
timestamp 1679235063
transform 1 0 26956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_302
timestamp 1679235063
transform 1 0 28888 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_309
timestamp 1679235063
transform 1 0 29532 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_323
timestamp 1679235063
transform 1 0 30820 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_327
timestamp 1679235063
transform 1 0 31188 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_337
timestamp 1679235063
transform 1 0 32108 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_341
timestamp 1679235063
transform 1 0 32476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_353
timestamp 1679235063
transform 1 0 33580 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_357
timestamp 1679235063
transform 1 0 33948 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1679235063
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1679235063
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_370
timestamp 1679235063
transform 1 0 35144 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_374
timestamp 1679235063
transform 1 0 35512 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_397
timestamp 1679235063
transform 1 0 37628 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_410
timestamp 1679235063
transform 1 0 38824 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_417
timestamp 1679235063
transform 1 0 39468 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_425
timestamp 1679235063
transform 1 0 40204 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_437
timestamp 1679235063
transform 1 0 41308 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_449
timestamp 1679235063
transform 1 0 42412 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_455
timestamp 1679235063
transform 1 0 42964 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_467
timestamp 1679235063
transform 1 0 44068 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1679235063
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1679235063
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1679235063
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1679235063
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_513
timestamp 1679235063
transform 1 0 48300 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_519
timestamp 1679235063
transform 1 0 48852 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1679235063
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1679235063
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_21
timestamp 1679235063
transform 1 0 3036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_29
timestamp 1679235063
transform 1 0 3772 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_40
timestamp 1679235063
transform 1 0 4784 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_47
timestamp 1679235063
transform 1 0 5428 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1679235063
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_57
timestamp 1679235063
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1679235063
transform 1 0 6808 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_67
timestamp 1679235063
transform 1 0 7268 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_75
timestamp 1679235063
transform 1 0 8004 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_80
timestamp 1679235063
transform 1 0 8464 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_103
timestamp 1679235063
transform 1 0 10580 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1679235063
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 1679235063
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_116
timestamp 1679235063
transform 1 0 11776 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_121
timestamp 1679235063
transform 1 0 12236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_145
timestamp 1679235063
transform 1 0 14444 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_158
timestamp 1679235063
transform 1 0 15640 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1679235063
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_175
timestamp 1679235063
transform 1 0 17204 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_186
timestamp 1679235063
transform 1 0 18216 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_194
timestamp 1679235063
transform 1 0 18952 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_199
timestamp 1679235063
transform 1 0 19412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1679235063
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1679235063
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_230
timestamp 1679235063
transform 1 0 22264 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_245
timestamp 1679235063
transform 1 0 23644 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_252
timestamp 1679235063
transform 1 0 24288 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_265
timestamp 1679235063
transform 1 0 25484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1679235063
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1679235063
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_292
timestamp 1679235063
transform 1 0 27968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_305
timestamp 1679235063
transform 1 0 29164 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_309
timestamp 1679235063
transform 1 0 29532 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_320
timestamp 1679235063
transform 1 0 30544 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_333
timestamp 1679235063
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1679235063
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_348
timestamp 1679235063
transform 1 0 33120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_352
timestamp 1679235063
transform 1 0 33488 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_373
timestamp 1679235063
transform 1 0 35420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_377
timestamp 1679235063
transform 1 0 35788 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_387
timestamp 1679235063
transform 1 0 36708 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1679235063
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_399
timestamp 1679235063
transform 1 0 37812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_421
timestamp 1679235063
transform 1 0 39836 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_425
timestamp 1679235063
transform 1 0 40204 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_436
timestamp 1679235063
transform 1 0 41216 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_443
timestamp 1679235063
transform 1 0 41860 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1679235063
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_449
timestamp 1679235063
transform 1 0 42412 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_459
timestamp 1679235063
transform 1 0 43332 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_471
timestamp 1679235063
transform 1 0 44436 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_483
timestamp 1679235063
transform 1 0 45540 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_495
timestamp 1679235063
transform 1 0 46644 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1679235063
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1679235063
transform 1 0 47564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_513
timestamp 1679235063
transform 1 0 48300 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_519
timestamp 1679235063
transform 1 0 48852 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1679235063
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1679235063
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1679235063
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1679235063
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1679235063
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_47
timestamp 1679235063
transform 1 0 5428 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_51
timestamp 1679235063
transform 1 0 5796 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_58
timestamp 1679235063
transform 1 0 6440 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_65
timestamp 1679235063
transform 1 0 7084 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_72
timestamp 1679235063
transform 1 0 7728 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_80
timestamp 1679235063
transform 1 0 8464 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1679235063
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_91
timestamp 1679235063
transform 1 0 9476 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_98
timestamp 1679235063
transform 1 0 10120 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_122
timestamp 1679235063
transform 1 0 12328 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_128
timestamp 1679235063
transform 1 0 12880 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1679235063
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1679235063
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_163
timestamp 1679235063
transform 1 0 16100 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_176
timestamp 1679235063
transform 1 0 17296 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_189
timestamp 1679235063
transform 1 0 18492 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_212
timestamp 1679235063
transform 1 0 20608 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_216
timestamp 1679235063
transform 1 0 20976 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_226
timestamp 1679235063
transform 1 0 21896 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1679235063
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1679235063
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_264
timestamp 1679235063
transform 1 0 25392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_268
timestamp 1679235063
transform 1 0 25760 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_289
timestamp 1679235063
transform 1 0 27692 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_301
timestamp 1679235063
transform 1 0 28796 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1679235063
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1679235063
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_320
timestamp 1679235063
transform 1 0 30544 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_333
timestamp 1679235063
transform 1 0 31740 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_346
timestamp 1679235063
transform 1 0 32936 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_359
timestamp 1679235063
transform 1 0 34132 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1679235063
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_365
timestamp 1679235063
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_370
timestamp 1679235063
transform 1 0 35144 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_374
timestamp 1679235063
transform 1 0 35512 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_395
timestamp 1679235063
transform 1 0 37444 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_399
timestamp 1679235063
transform 1 0 37812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_410
timestamp 1679235063
transform 1 0 38824 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_417
timestamp 1679235063
transform 1 0 39468 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_421
timestamp 1679235063
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_443
timestamp 1679235063
transform 1 0 41860 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_455
timestamp 1679235063
transform 1 0 42964 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_459
timestamp 1679235063
transform 1 0 43332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_471
timestamp 1679235063
transform 1 0 44436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1679235063
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1679235063
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1679235063
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1679235063
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_513
timestamp 1679235063
transform 1 0 48300 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_517
timestamp 1679235063
transform 1 0 48668 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1679235063
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1679235063
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1679235063
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1679235063
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_49
timestamp 1679235063
transform 1 0 5612 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_63
timestamp 1679235063
transform 1 0 6900 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_68
timestamp 1679235063
transform 1 0 7360 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_76
timestamp 1679235063
transform 1 0 8096 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_80
timestamp 1679235063
transform 1 0 8464 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_84
timestamp 1679235063
transform 1 0 8832 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_91
timestamp 1679235063
transform 1 0 9476 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_98
timestamp 1679235063
transform 1 0 10120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1679235063
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1679235063
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_119
timestamp 1679235063
transform 1 0 12052 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_132
timestamp 1679235063
transform 1 0 13248 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_140
timestamp 1679235063
transform 1 0 13984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1679235063
transform 1 0 14352 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_154
timestamp 1679235063
transform 1 0 15272 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1679235063
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1679235063
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_180
timestamp 1679235063
transform 1 0 17664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_207
timestamp 1679235063
transform 1 0 20148 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_211
timestamp 1679235063
transform 1 0 20516 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1679235063
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1679235063
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_236
timestamp 1679235063
transform 1 0 22816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_241
timestamp 1679235063
transform 1 0 23276 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_263
timestamp 1679235063
transform 1 0 25300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_267
timestamp 1679235063
transform 1 0 25668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1679235063
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_281
timestamp 1679235063
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_293
timestamp 1679235063
transform 1 0 28060 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_306
timestamp 1679235063
transform 1 0 29256 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_318
timestamp 1679235063
transform 1 0 30360 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1679235063
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1679235063
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_348
timestamp 1679235063
transform 1 0 33120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_361
timestamp 1679235063
transform 1 0 34316 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_374
timestamp 1679235063
transform 1 0 35512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_387
timestamp 1679235063
transform 1 0 36708 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1679235063
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_397
timestamp 1679235063
transform 1 0 37628 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_420
timestamp 1679235063
transform 1 0 39744 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_433
timestamp 1679235063
transform 1 0 40940 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_445
timestamp 1679235063
transform 1 0 42044 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_455
timestamp 1679235063
transform 1 0 42964 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_467
timestamp 1679235063
transform 1 0 44068 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_479
timestamp 1679235063
transform 1 0 45172 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_491
timestamp 1679235063
transform 1 0 46276 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1679235063
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_505
timestamp 1679235063
transform 1 0 47564 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_519
timestamp 1679235063
transform 1 0 48852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1679235063
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1679235063
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1679235063
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1679235063
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1679235063
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_47
timestamp 1679235063
transform 1 0 5428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_67
timestamp 1679235063
transform 1 0 7268 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_74
timestamp 1679235063
transform 1 0 7912 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1679235063
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_85
timestamp 1679235063
transform 1 0 8924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_91
timestamp 1679235063
transform 1 0 9476 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_96
timestamp 1679235063
transform 1 0 9936 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_102
timestamp 1679235063
transform 1 0 10488 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1679235063
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1679235063
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_147
timestamp 1679235063
transform 1 0 14628 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_157
timestamp 1679235063
transform 1 0 15548 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_169
timestamp 1679235063
transform 1 0 16652 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_193
timestamp 1679235063
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_197
timestamp 1679235063
transform 1 0 19228 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_200
timestamp 1679235063
transform 1 0 19504 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_206
timestamp 1679235063
transform 1 0 20056 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_230
timestamp 1679235063
transform 1 0 22264 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_238
timestamp 1679235063
transform 1 0 23000 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1679235063
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_257
timestamp 1679235063
transform 1 0 24748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_262
timestamp 1679235063
transform 1 0 25208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_275
timestamp 1679235063
transform 1 0 26404 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_288
timestamp 1679235063
transform 1 0 27600 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_301
timestamp 1679235063
transform 1 0 28796 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1679235063
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1679235063
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_320
timestamp 1679235063
transform 1 0 30544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_333
timestamp 1679235063
transform 1 0 31740 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_346
timestamp 1679235063
transform 1 0 32936 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_350
timestamp 1679235063
transform 1 0 33304 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_360
timestamp 1679235063
transform 1 0 34224 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1679235063
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_376
timestamp 1679235063
transform 1 0 35696 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_389
timestamp 1679235063
transform 1 0 36892 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_402
timestamp 1679235063
transform 1 0 38088 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_415
timestamp 1679235063
transform 1 0 39284 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1679235063
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1679235063
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_432
timestamp 1679235063
transform 1 0 40848 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_444
timestamp 1679235063
transform 1 0 41952 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_460
timestamp 1679235063
transform 1 0 43424 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_472
timestamp 1679235063
transform 1 0 44528 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1679235063
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_489
timestamp 1679235063
transform 1 0 46092 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_497
timestamp 1679235063
transform 1 0 46828 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_503
timestamp 1679235063
transform 1 0 47380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_512
timestamp 1679235063
transform 1 0 48208 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_517
timestamp 1679235063
transform 1 0 48668 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1679235063
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1679235063
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_21
timestamp 1679235063
transform 1 0 3036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_41
timestamp 1679235063
transform 1 0 4876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_49
timestamp 1679235063
transform 1 0 5612 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1679235063
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_75
timestamp 1679235063
transform 1 0 8004 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_82
timestamp 1679235063
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_90
timestamp 1679235063
transform 1 0 9384 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_98
timestamp 1679235063
transform 1 0 10120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1679235063
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_113
timestamp 1679235063
transform 1 0 11500 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_116
timestamp 1679235063
transform 1 0 11776 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_122
timestamp 1679235063
transform 1 0 12328 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_134
timestamp 1679235063
transform 1 0 13432 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_158
timestamp 1679235063
transform 1 0 15640 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1679235063
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_169
timestamp 1679235063
transform 1 0 16652 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_181
timestamp 1679235063
transform 1 0 17756 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_187
timestamp 1679235063
transform 1 0 18308 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_209
timestamp 1679235063
transform 1 0 20332 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1679235063
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_225
timestamp 1679235063
transform 1 0 21804 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_228
timestamp 1679235063
transform 1 0 22080 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_239
timestamp 1679235063
transform 1 0 23092 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_245
timestamp 1679235063
transform 1 0 23644 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_267
timestamp 1679235063
transform 1 0 25668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_274
timestamp 1679235063
transform 1 0 26312 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_281
timestamp 1679235063
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_304
timestamp 1679235063
transform 1 0 29072 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_317
timestamp 1679235063
transform 1 0 30268 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_330
timestamp 1679235063
transform 1 0 31464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1679235063
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_359
timestamp 1679235063
transform 1 0 34132 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_365
timestamp 1679235063
transform 1 0 34684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_376
timestamp 1679235063
transform 1 0 35696 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1679235063
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_395
timestamp 1679235063
transform 1 0 37444 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_418
timestamp 1679235063
transform 1 0 39560 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_431
timestamp 1679235063
transform 1 0 40756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_443
timestamp 1679235063
transform 1 0 41860 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1679235063
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_449
timestamp 1679235063
transform 1 0 42412 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_454
timestamp 1679235063
transform 1 0 42872 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_466
timestamp 1679235063
transform 1 0 43976 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_476
timestamp 1679235063
transform 1 0 44896 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_488
timestamp 1679235063
transform 1 0 46000 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_492
timestamp 1679235063
transform 1 0 46368 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_497
timestamp 1679235063
transform 1 0 46828 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_505
timestamp 1679235063
transform 1 0 47564 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_512
timestamp 1679235063
transform 1 0 48208 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_517
timestamp 1679235063
transform 1 0 48668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1679235063
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1679235063
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1679235063
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1679235063
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1679235063
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1679235063
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_67
timestamp 1679235063
transform 1 0 7268 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_74
timestamp 1679235063
transform 1 0 7912 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1679235063
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_91
timestamp 1679235063
transform 1 0 9476 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_101
timestamp 1679235063
transform 1 0 10396 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_113
timestamp 1679235063
transform 1 0 11500 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_125
timestamp 1679235063
transform 1 0 12604 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1679235063
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_145
timestamp 1679235063
transform 1 0 14444 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_167
timestamp 1679235063
transform 1 0 16468 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_171
timestamp 1679235063
transform 1 0 16836 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_181
timestamp 1679235063
transform 1 0 17756 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1679235063
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_197
timestamp 1679235063
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_204
timestamp 1679235063
transform 1 0 19872 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_228
timestamp 1679235063
transform 1 0 22080 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_232
timestamp 1679235063
transform 1 0 22448 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_237
timestamp 1679235063
transform 1 0 22908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1679235063
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1679235063
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_263
timestamp 1679235063
transform 1 0 25300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_276
timestamp 1679235063
transform 1 0 26496 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_289
timestamp 1679235063
transform 1 0 27692 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_293
timestamp 1679235063
transform 1 0 28060 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1679235063
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1679235063
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_314
timestamp 1679235063
transform 1 0 29992 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_320
timestamp 1679235063
transform 1 0 30544 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_331
timestamp 1679235063
transform 1 0 31556 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_339
timestamp 1679235063
transform 1 0 32292 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1679235063
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1679235063
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_387
timestamp 1679235063
transform 1 0 36708 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_395
timestamp 1679235063
transform 1 0 37444 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_417
timestamp 1679235063
transform 1 0 39468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_421
timestamp 1679235063
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_432
timestamp 1679235063
transform 1 0 40848 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_445
timestamp 1679235063
transform 1 0 42044 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_459
timestamp 1679235063
transform 1 0 43332 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_466
timestamp 1679235063
transform 1 0 43976 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_473
timestamp 1679235063
transform 1 0 44620 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_477
timestamp 1679235063
transform 1 0 44988 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_482
timestamp 1679235063
transform 1 0 45448 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_490
timestamp 1679235063
transform 1 0 46184 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_495
timestamp 1679235063
transform 1 0 46644 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_502
timestamp 1679235063
transform 1 0 47288 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_506
timestamp 1679235063
transform 1 0 47656 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_510
timestamp 1679235063
transform 1 0 48024 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_517
timestamp 1679235063
transform 1 0 48668 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_525
timestamp 1679235063
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1679235063
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1679235063
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_41
timestamp 1679235063
transform 1 0 4876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_48
timestamp 1679235063
transform 1 0 5520 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1679235063
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1679235063
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_75
timestamp 1679235063
transform 1 0 8004 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_95
timestamp 1679235063
transform 1 0 9844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_100
timestamp 1679235063
transform 1 0 10304 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1679235063
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1679235063
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_119
timestamp 1679235063
transform 1 0 12052 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_123
timestamp 1679235063
transform 1 0 12420 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_132
timestamp 1679235063
transform 1 0 13248 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_144
timestamp 1679235063
transform 1 0 14352 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_157
timestamp 1679235063
transform 1 0 15548 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_161
timestamp 1679235063
transform 1 0 15916 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1679235063
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1679235063
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_180
timestamp 1679235063
transform 1 0 17664 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_204
timestamp 1679235063
transform 1 0 19872 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_211
timestamp 1679235063
transform 1 0 20516 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1679235063
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_225
timestamp 1679235063
transform 1 0 21804 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_230
timestamp 1679235063
transform 1 0 22264 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_253
timestamp 1679235063
transform 1 0 24380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_266
timestamp 1679235063
transform 1 0 25576 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1679235063
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1679235063
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_292
timestamp 1679235063
transform 1 0 27968 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_305
timestamp 1679235063
transform 1 0 29164 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_318
timestamp 1679235063
transform 1 0 30360 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_331
timestamp 1679235063
transform 1 0 31556 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1679235063
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1679235063
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_342
timestamp 1679235063
transform 1 0 32568 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_346
timestamp 1679235063
transform 1 0 32936 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_358
timestamp 1679235063
transform 1 0 34040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_371
timestamp 1679235063
transform 1 0 35236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_375
timestamp 1679235063
transform 1 0 35604 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_385
timestamp 1679235063
transform 1 0 36524 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1679235063
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_399
timestamp 1679235063
transform 1 0 37812 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_421
timestamp 1679235063
transform 1 0 39836 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_434
timestamp 1679235063
transform 1 0 41032 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1679235063
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_449
timestamp 1679235063
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_459
timestamp 1679235063
transform 1 0 43332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_466
timestamp 1679235063
transform 1 0 43976 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_473
timestamp 1679235063
transform 1 0 44620 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_480
timestamp 1679235063
transform 1 0 45264 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_487
timestamp 1679235063
transform 1 0 45908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_494
timestamp 1679235063
transform 1 0 46552 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_501
timestamp 1679235063
transform 1 0 47196 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_511
timestamp 1679235063
transform 1 0 48116 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_517
timestamp 1679235063
transform 1 0 48668 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1679235063
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1679235063
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1679235063
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1679235063
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1679235063
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_47
timestamp 1679235063
transform 1 0 5428 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_67
timestamp 1679235063
transform 1 0 7268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_72
timestamp 1679235063
transform 1 0 7728 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1679235063
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1679235063
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_103
timestamp 1679235063
transform 1 0 10580 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_111
timestamp 1679235063
transform 1 0 11316 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_116
timestamp 1679235063
transform 1 0 11776 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_134
timestamp 1679235063
transform 1 0 13432 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_143
timestamp 1679235063
transform 1 0 14260 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_149
timestamp 1679235063
transform 1 0 14812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_173
timestamp 1679235063
transform 1 0 17020 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_177
timestamp 1679235063
transform 1 0 17388 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1679235063
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_203
timestamp 1679235063
transform 1 0 19780 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_214
timestamp 1679235063
transform 1 0 20792 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_238
timestamp 1679235063
transform 1 0 23000 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1679235063
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1679235063
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1679235063
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_268
timestamp 1679235063
transform 1 0 25760 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_279
timestamp 1679235063
transform 1 0 26772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_292
timestamp 1679235063
transform 1 0 27968 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_305
timestamp 1679235063
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1679235063
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_319
timestamp 1679235063
transform 1 0 30452 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_343
timestamp 1679235063
transform 1 0 32660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_356
timestamp 1679235063
transform 1 0 33856 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1679235063
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_376
timestamp 1679235063
transform 1 0 35696 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_389
timestamp 1679235063
transform 1 0 36892 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_414
timestamp 1679235063
transform 1 0 39192 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_421
timestamp 1679235063
transform 1 0 39836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_432
timestamp 1679235063
transform 1 0 40848 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_445
timestamp 1679235063
transform 1 0 42044 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_452
timestamp 1679235063
transform 1 0 42688 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_456
timestamp 1679235063
transform 1 0 43056 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_468
timestamp 1679235063
transform 1 0 44160 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_477
timestamp 1679235063
transform 1 0 44988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_482
timestamp 1679235063
transform 1 0 45448 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_496
timestamp 1679235063
transform 1 0 46736 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_503
timestamp 1679235063
transform 1 0 47380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_511
timestamp 1679235063
transform 1 0 48116 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_517
timestamp 1679235063
transform 1 0 48668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1679235063
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1679235063
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_21
timestamp 1679235063
transform 1 0 3036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_25
timestamp 1679235063
transform 1 0 3404 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_28
timestamp 1679235063
transform 1 0 3680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1679235063
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1679235063
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1679235063
transform 1 0 6532 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_65
timestamp 1679235063
transform 1 0 7084 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_85
timestamp 1679235063
transform 1 0 8924 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_92
timestamp 1679235063
transform 1 0 9568 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1679235063
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1679235063
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_125
timestamp 1679235063
transform 1 0 12604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_129
timestamp 1679235063
transform 1 0 12972 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_146
timestamp 1679235063
transform 1 0 14536 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1679235063
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1679235063
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_191
timestamp 1679235063
transform 1 0 18676 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_198
timestamp 1679235063
transform 1 0 19320 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_221
timestamp 1679235063
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1679235063
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_248
timestamp 1679235063
transform 1 0 23920 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_256
timestamp 1679235063
transform 1 0 24656 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1679235063
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1679235063
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_287
timestamp 1679235063
transform 1 0 27508 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_291
timestamp 1679235063
transform 1 0 27876 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_313
timestamp 1679235063
transform 1 0 29900 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_326
timestamp 1679235063
transform 1 0 31096 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_330
timestamp 1679235063
transform 1 0 31464 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1679235063
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1679235063
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_348
timestamp 1679235063
transform 1 0 33120 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_352
timestamp 1679235063
transform 1 0 33488 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_374
timestamp 1679235063
transform 1 0 35512 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_378
timestamp 1679235063
transform 1 0 35880 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_389
timestamp 1679235063
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1679235063
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_415
timestamp 1679235063
transform 1 0 39284 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_428
timestamp 1679235063
transform 1 0 40480 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_440
timestamp 1679235063
transform 1 0 41584 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1679235063
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_454
timestamp 1679235063
transform 1 0 42872 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_468
timestamp 1679235063
transform 1 0 44160 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_482
timestamp 1679235063
transform 1 0 45448 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_496
timestamp 1679235063
transform 1 0 46736 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_511
timestamp 1679235063
transform 1 0 48116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_517
timestamp 1679235063
transform 1 0 48668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1679235063
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1679235063
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_21
timestamp 1679235063
transform 1 0 3036 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1679235063
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_41
timestamp 1679235063
transform 1 0 4876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_45
timestamp 1679235063
transform 1 0 5244 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1679235063
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1679235063
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1679235063
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_97
timestamp 1679235063
transform 1 0 10028 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_101
timestamp 1679235063
transform 1 0 10396 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_118
timestamp 1679235063
transform 1 0 11960 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1679235063
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_141
timestamp 1679235063
transform 1 0 14076 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_144
timestamp 1679235063
transform 1 0 14352 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_150
timestamp 1679235063
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1679235063
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1679235063
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_197
timestamp 1679235063
transform 1 0 19228 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_200
timestamp 1679235063
transform 1 0 19504 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_205
timestamp 1679235063
transform 1 0 19964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_229
timestamp 1679235063
transform 1 0 22172 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_242
timestamp 1679235063
transform 1 0 23368 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1679235063
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1679235063
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_263
timestamp 1679235063
transform 1 0 25300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_287
timestamp 1679235063
transform 1 0 27508 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_300
timestamp 1679235063
transform 1 0 28704 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1679235063
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_320
timestamp 1679235063
transform 1 0 30544 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_326
timestamp 1679235063
transform 1 0 31096 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_350
timestamp 1679235063
transform 1 0 33304 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_362
timestamp 1679235063
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_365
timestamp 1679235063
transform 1 0 34684 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_388
timestamp 1679235063
transform 1 0 36800 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_412
timestamp 1679235063
transform 1 0 39008 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1679235063
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_432
timestamp 1679235063
transform 1 0 40848 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_436
timestamp 1679235063
transform 1 0 41216 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_462
timestamp 1679235063
transform 1 0 43608 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_466
timestamp 1679235063
transform 1 0 43976 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_472
timestamp 1679235063
transform 1 0 44528 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_477
timestamp 1679235063
transform 1 0 44988 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_489
timestamp 1679235063
transform 1 0 46092 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_503
timestamp 1679235063
transform 1 0 47380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_511
timestamp 1679235063
transform 1 0 48116 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_517
timestamp 1679235063
transform 1 0 48668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1679235063
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_3
timestamp 1679235063
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_8
timestamp 1679235063
transform 1 0 1840 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1679235063
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1679235063
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1679235063
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_57
timestamp 1679235063
transform 1 0 6348 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_60
timestamp 1679235063
transform 1 0 6624 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1679235063
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1679235063
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1679235063
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1679235063
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_126
timestamp 1679235063
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1679235063
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1679235063
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_169
timestamp 1679235063
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_188
timestamp 1679235063
transform 1 0 18400 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_212
timestamp 1679235063
transform 1 0 20608 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_216
timestamp 1679235063
transform 1 0 20976 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1679235063
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1679235063
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_236
timestamp 1679235063
transform 1 0 22816 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_244
timestamp 1679235063
transform 1 0 23552 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_254
timestamp 1679235063
transform 1 0 24472 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1679235063
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1679235063
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_291
timestamp 1679235063
transform 1 0 27876 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_303
timestamp 1679235063
transform 1 0 28980 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_310
timestamp 1679235063
transform 1 0 29624 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1679235063
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1679235063
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_348
timestamp 1679235063
transform 1 0 33120 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_372
timestamp 1679235063
transform 1 0 35328 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_376
timestamp 1679235063
transform 1 0 35696 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_387
timestamp 1679235063
transform 1 0 36708 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1679235063
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1679235063
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_404
timestamp 1679235063
transform 1 0 38272 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_408
timestamp 1679235063
transform 1 0 38640 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_419
timestamp 1679235063
transform 1 0 39652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_431
timestamp 1679235063
transform 1 0 40756 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_445
timestamp 1679235063
transform 1 0 42044 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_449
timestamp 1679235063
transform 1 0 42412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_461
timestamp 1679235063
transform 1 0 43516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_475
timestamp 1679235063
transform 1 0 44804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_489
timestamp 1679235063
transform 1 0 46092 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_497
timestamp 1679235063
transform 1 0 46828 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1679235063
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_505
timestamp 1679235063
transform 1 0 47564 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_511
timestamp 1679235063
transform 1 0 48116 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_519
timestamp 1679235063
transform 1 0 48852 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1679235063
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1679235063
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1679235063
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1679235063
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1679235063
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1679235063
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1679235063
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1679235063
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1679235063
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1679235063
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1679235063
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1679235063
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1679235063
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1679235063
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1679235063
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1679235063
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1679235063
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1679235063
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1679235063
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_174
timestamp 1679235063
transform 1 0 17112 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1679235063
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1679235063
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1679235063
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1679235063
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_225
timestamp 1679235063
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_243
timestamp 1679235063
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1679235063
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_253
timestamp 1679235063
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_260
timestamp 1679235063
transform 1 0 25024 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_272
timestamp 1679235063
transform 1 0 26128 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_281
timestamp 1679235063
transform 1 0 26956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_292
timestamp 1679235063
transform 1 0 27968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_304
timestamp 1679235063
transform 1 0 29072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1679235063
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_315
timestamp 1679235063
transform 1 0 30084 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_321
timestamp 1679235063
transform 1 0 30636 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_331
timestamp 1679235063
transform 1 0 31556 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_335
timestamp 1679235063
transform 1 0 31924 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_339
timestamp 1679235063
transform 1 0 32292 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_349
timestamp 1679235063
transform 1 0 33212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1679235063
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1679235063
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_376
timestamp 1679235063
transform 1 0 35696 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_389
timestamp 1679235063
transform 1 0 36892 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_393
timestamp 1679235063
transform 1 0 37260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_404
timestamp 1679235063
transform 1 0 38272 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_416
timestamp 1679235063
transform 1 0 39376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1679235063
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_431
timestamp 1679235063
transform 1 0 40756 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_445
timestamp 1679235063
transform 1 0 42044 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_449
timestamp 1679235063
transform 1 0 42412 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_471
timestamp 1679235063
transform 1 0 44436 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1679235063
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1679235063
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_489
timestamp 1679235063
transform 1 0 46092 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_497
timestamp 1679235063
transform 1 0 46828 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_503
timestamp 1679235063
transform 1 0 47380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_505
timestamp 1679235063
transform 1 0 47564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_511
timestamp 1679235063
transform 1 0 48116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_525
timestamp 1679235063
transform 1 0 49404 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16836 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1679235063
transform 1 0 41216 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1679235063
transform 1 0 16836 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold4 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9660 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold5
timestamp 1679235063
transform 1 0 41308 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1679235063
transform 1 0 15916 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1679235063
transform 1 0 21528 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1679235063
transform 1 0 11868 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold9
timestamp 1679235063
transform 1 0 40020 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1679235063
transform 1 0 10856 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1679235063
transform 1 0 19412 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1679235063
transform 1 0 27876 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1679235063
transform 1 0 19412 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold14
timestamp 1679235063
transform 1 0 38640 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1679235063
transform 1 0 28060 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1679235063
transform 1 0 27140 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1679235063
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold18
timestamp 1679235063
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1679235063
transform 1 0 24840 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1679235063
transform 1 0 15732 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1679235063
transform 1 0 25392 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1679235063
transform 1 0 25024 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1679235063
transform 1 0 15640 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1679235063
transform 1 0 18216 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1679235063
transform 1 0 27048 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1679235063
transform 1 0 10488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1679235063
transform 1 0 13616 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1679235063
transform 1 0 39836 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1679235063
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold30
timestamp 1679235063
transform 1 0 12696 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1679235063
transform 1 0 41124 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1679235063
transform 1 0 38548 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1679235063
transform 1 0 24564 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1679235063
transform 1 0 25300 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1679235063
transform 1 0 10488 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1679235063
transform 1 0 25944 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1679235063
transform 1 0 27140 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1679235063
transform 1 0 13064 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1679235063
transform 1 0 20792 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1679235063
transform 1 0 24564 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold41
timestamp 1679235063
transform 1 0 16836 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1679235063
transform 1 0 30820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1679235063
transform 1 0 33672 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold44
timestamp 1679235063
transform 1 0 11868 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold45
timestamp 1679235063
transform 1 0 32292 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold46
timestamp 1679235063
transform 1 0 10764 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1679235063
transform 1 0 19228 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold48
timestamp 1679235063
transform 1 0 38272 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold49
timestamp 1679235063
transform 1 0 26036 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold50
timestamp 1679235063
transform 1 0 14536 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold51
timestamp 1679235063
transform 1 0 14812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold52
timestamp 1679235063
transform 1 0 40848 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold53
timestamp 1679235063
transform 1 0 32200 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold54
timestamp 1679235063
transform 1 0 40020 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold55
timestamp 1679235063
transform 1 0 42596 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold56
timestamp 1679235063
transform 1 0 41124 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold57
timestamp 1679235063
transform 1 0 23092 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold58
timestamp 1679235063
transform 1 0 30268 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold59
timestamp 1679235063
transform 1 0 38640 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold60
timestamp 1679235063
transform 1 0 42228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold61
timestamp 1679235063
transform 1 0 10488 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold62
timestamp 1679235063
transform 1 0 12512 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold63
timestamp 1679235063
transform 1 0 25944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold64
timestamp 1679235063
transform 1 0 41124 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold65
timestamp 1679235063
transform 1 0 14444 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold66
timestamp 1679235063
transform 1 0 41032 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold67
timestamp 1679235063
transform 1 0 14260 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold68
timestamp 1679235063
transform 1 0 7912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold69
timestamp 1679235063
transform 1 0 21988 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold70
timestamp 1679235063
transform 1 0 41676 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold71
timestamp 1679235063
transform 1 0 42596 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold72
timestamp 1679235063
transform 1 0 29716 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold73
timestamp 1679235063
transform 1 0 32476 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold74
timestamp 1679235063
transform 1 0 20332 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold75
timestamp 1679235063
transform 1 0 30360 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold76
timestamp 1679235063
transform 1 0 28520 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold77
timestamp 1679235063
transform 1 0 38180 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold78
timestamp 1679235063
transform 1 0 28336 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold79
timestamp 1679235063
transform 1 0 10488 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold80
timestamp 1679235063
transform 1 0 21988 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold81
timestamp 1679235063
transform 1 0 41400 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold82
timestamp 1679235063
transform 1 0 16836 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold83
timestamp 1679235063
transform 1 0 23736 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold84
timestamp 1679235063
transform 1 0 27692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold85
timestamp 1679235063
transform 1 0 40020 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold86
timestamp 1679235063
transform 1 0 39836 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold87
timestamp 1679235063
transform 1 0 24564 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold88
timestamp 1679235063
transform 1 0 29624 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold89
timestamp 1679235063
transform 1 0 29808 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold90
timestamp 1679235063
transform 1 0 36064 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold91
timestamp 1679235063
transform 1 0 14076 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold92
timestamp 1679235063
transform 1 0 9568 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold93
timestamp 1679235063
transform 1 0 37076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold94
timestamp 1679235063
transform 1 0 27232 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold95
timestamp 1679235063
transform 1 0 37444 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold96
timestamp 1679235063
transform 1 0 24564 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold97
timestamp 1679235063
transform 1 0 40848 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold98
timestamp 1679235063
transform 1 0 40020 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold99
timestamp 1679235063
transform 1 0 39928 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold100
timestamp 1679235063
transform 1 0 40020 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold101
timestamp 1679235063
transform 1 0 41124 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold102
timestamp 1679235063
transform 1 0 42228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold103
timestamp 1679235063
transform 1 0 10028 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold104
timestamp 1679235063
transform 1 0 29716 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold105
timestamp 1679235063
transform 1 0 42228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold106
timestamp 1679235063
transform 1 0 23368 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold107
timestamp 1679235063
transform 1 0 42596 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold108
timestamp 1679235063
transform 1 0 28244 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold109
timestamp 1679235063
transform 1 0 6808 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold110
timestamp 1679235063
transform 1 0 28336 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1679235063
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1679235063
transform 1 0 47104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1679235063
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input4 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1679235063
transform 1 0 1564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1679235063
transform 1 0 2300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1679235063
transform 1 0 1564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1679235063
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1679235063
transform 1 0 1564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1679235063
transform 1 0 1564 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1679235063
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1679235063
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1679235063
transform 1 0 1564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1679235063
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1679235063
transform 1 0 1564 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1679235063
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1679235063
transform 1 0 1564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1679235063
transform 1 0 1564 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1679235063
transform 1 0 2300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1679235063
transform 1 0 1564 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1679235063
transform 1 0 1564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1679235063
transform 1 0 2852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1679235063
transform 1 0 1564 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1679235063
transform 1 0 3404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1679235063
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1679235063
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1679235063
transform 1 0 1564 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input28
timestamp 1679235063
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1679235063
transform 1 0 1564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 1679235063
transform 1 0 1564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1679235063
transform 1 0 1564 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1679235063
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1679235063
transform 1 0 48392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1679235063
transform 1 0 49036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1679235063
transform 1 0 49036 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1679235063
transform 1 0 48392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1679235063
transform 1 0 49036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1679235063
transform 1 0 49036 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1679235063
transform 1 0 49036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1679235063
transform 1 0 48392 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1679235063
transform 1 0 49036 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1679235063
transform 1 0 49036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1679235063
transform 1 0 49036 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1679235063
transform 1 0 49036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1679235063
transform 1 0 48392 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1679235063
transform 1 0 49036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1679235063
transform 1 0 48300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1679235063
transform 1 0 48300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1679235063
transform 1 0 47748 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1679235063
transform 1 0 46368 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1679235063
transform 1 0 48300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1679235063
transform 1 0 48392 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1679235063
transform 1 0 47012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1679235063
transform 1 0 48484 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1679235063
transform 1 0 49036 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1679235063
transform 1 0 49036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1679235063
transform 1 0 49128 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1679235063
transform 1 0 49036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1679235063
transform 1 0 49036 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1679235063
transform 1 0 49036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1679235063
transform 1 0 48392 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1679235063
transform 1 0 49036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1679235063
transform 1 0 3864 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1679235063
transform 1 0 41124 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1679235063
transform 1 0 45172 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1679235063
transform 1 0 43240 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1679235063
transform 1 0 43240 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1679235063
transform 1 0 45172 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1679235063
transform 1 0 45632 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1679235063
transform 1 0 41584 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1679235063
transform 1 0 46276 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1679235063
transform 1 0 45172 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1679235063
transform 1 0 44528 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1679235063
transform 1 0 21988 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1679235063
transform 1 0 45816 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1679235063
transform 1 0 45172 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1679235063
transform 1 0 43700 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input78
timestamp 1679235063
transform 1 0 46460 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input79
timestamp 1679235063
transform 1 0 45816 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1679235063
transform 1 0 44344 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1679235063
transform 1 0 43700 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1679235063
transform 1 0 44988 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1679235063
transform 1 0 46920 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1679235063
transform 1 0 45172 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input85
timestamp 1679235063
transform 1 0 9108 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1679235063
transform 1 0 26036 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input87
timestamp 1679235063
transform 1 0 11684 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input88
timestamp 1679235063
transform 1 0 43884 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input89
timestamp 1679235063
transform 1 0 11776 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1679235063
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1679235063
transform 1 0 16836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input92
timestamp 1679235063
transform 1 0 41124 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1679235063
transform 1 0 28704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1679235063
transform 1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1679235063
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1679235063
transform 1 0 35052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input97
timestamp 1679235063
transform 1 0 37444 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_16  input98
timestamp 1679235063
transform 1 0 42596 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  input99
timestamp 1679235063
transform 1 0 46460 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input100
timestamp 1679235063
transform 1 0 47748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1679235063
transform 1 0 47748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input102
timestamp 1679235063
transform 1 0 49036 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1679235063
transform 1 0 48484 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input104
timestamp 1679235063
transform 1 0 48300 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input105
timestamp 1679235063
transform 1 0 44160 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1679235063
transform 1 0 46460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output107 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 40664 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1679235063
transform 1 0 3404 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1679235063
transform 1 0 1564 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1679235063
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1679235063
transform 1 0 1564 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1679235063
transform 1 0 1564 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1679235063
transform 1 0 1564 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1679235063
transform 1 0 1564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1679235063
transform 1 0 1564 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1679235063
transform 1 0 3404 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1679235063
transform 1 0 1564 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1679235063
transform 1 0 1564 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1679235063
transform 1 0 1564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1679235063
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1679235063
transform 1 0 3956 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1679235063
transform 1 0 3956 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1679235063
transform 1 0 5796 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1679235063
transform 1 0 5796 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1679235063
transform 1 0 6532 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1679235063
transform 1 0 3956 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1679235063
transform 1 0 5796 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1679235063
transform 1 0 6532 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1679235063
transform 1 0 8372 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1679235063
transform 1 0 9108 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1679235063
transform 1 0 1564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1679235063
transform 1 0 1564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1679235063
transform 1 0 1564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1679235063
transform 1 0 1564 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1679235063
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1679235063
transform 1 0 1564 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1679235063
transform 1 0 1564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1679235063
transform 1 0 1564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1679235063
transform 1 0 45816 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1679235063
transform 1 0 47932 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1679235063
transform 1 0 47932 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1679235063
transform 1 0 46092 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1679235063
transform 1 0 47932 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1679235063
transform 1 0 47932 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1679235063
transform 1 0 47932 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1679235063
transform 1 0 45816 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1679235063
transform 1 0 47932 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1679235063
transform 1 0 47932 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1679235063
transform 1 0 47932 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1679235063
transform 1 0 43976 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1679235063
transform 1 0 46092 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1679235063
transform 1 0 47932 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1679235063
transform 1 0 47932 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1679235063
transform 1 0 47932 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1679235063
transform 1 0 47932 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1679235063
transform 1 0 47932 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1679235063
transform 1 0 47932 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1679235063
transform 1 0 47932 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1679235063
transform 1 0 47932 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1679235063
transform 1 0 47932 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1679235063
transform 1 0 45816 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1679235063
transform 1 0 45816 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1679235063
transform 1 0 46092 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1679235063
transform 1 0 47932 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1679235063
transform 1 0 47932 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1679235063
transform 1 0 47932 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1679235063
transform 1 0 45816 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1679235063
transform 1 0 47932 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1679235063
transform 1 0 3956 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1679235063
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1679235063
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1679235063
transform 1 0 9752 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1679235063
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1679235063
transform 1 0 10488 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1679235063
transform 1 0 11960 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1679235063
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1679235063
transform 1 0 12328 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1679235063
transform 1 0 13064 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1679235063
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1679235063
transform 1 0 3404 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1679235063
transform 1 0 13064 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1679235063
transform 1 0 14904 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1679235063
transform 1 0 15272 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1679235063
transform 1 0 14904 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1679235063
transform 1 0 17480 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1679235063
transform 1 0 14904 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1679235063
transform 1 0 16928 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1679235063
transform 1 0 17480 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1679235063
transform 1 0 21988 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1679235063
transform 1 0 20056 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1679235063
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1679235063
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1679235063
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1679235063
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1679235063
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1679235063
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1679235063
transform 1 0 7452 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1679235063
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1679235063
transform 1 0 11776 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1679235063
transform 1 0 14260 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1679235063
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output202
timestamp 1679235063
transform 1 0 17480 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1679235063
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1679235063
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1679235063
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1679235063
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1679235063
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1679235063
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1679235063
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1679235063
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1679235063
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1679235063
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1679235063
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1679235063
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1679235063
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1679235063
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1679235063
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1679235063
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1679235063
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1679235063
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1679235063
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1679235063
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1679235063
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1679235063
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1679235063
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1679235063
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1679235063
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1679235063
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1679235063
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1679235063
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1679235063
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1679235063
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1679235063
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1679235063
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1679235063
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1679235063
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1679235063
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1679235063
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1679235063
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1679235063
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1679235063
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1679235063
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1679235063
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1679235063
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1679235063
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1679235063
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1679235063
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1679235063
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1679235063
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1679235063
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1679235063
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1679235063
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1679235063
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1679235063
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1679235063
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1679235063
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1679235063
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1679235063
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1679235063
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1679235063
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1679235063
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1679235063
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1679235063
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1679235063
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1679235063
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1679235063
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1679235063
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1679235063
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1679235063
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1679235063
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1679235063
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1679235063
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1679235063
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1679235063
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1679235063
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1679235063
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1679235063
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1679235063
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1679235063
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1679235063
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1679235063
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1679235063
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1679235063
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1679235063
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 27140 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24564 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 22632 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20424 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 17020 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18492 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20148 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 17112 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19044 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 19688 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21068 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21068 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 19320 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19596 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20240 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 18032 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19504 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20332 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 18768 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23828 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 23460 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 25852 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 27048 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 25576 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 27232 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 28060 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 24840 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 25668 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24840 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 21160 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22448 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 28336 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 30452 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 31464 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 32292 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 34868 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 35052 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 34868 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 36432 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 37444 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 34868 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 35144 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 35696 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 33856 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 34868 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 33764 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 32292 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 32200 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 31188 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 28060 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 29716 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 28520 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 26956 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 28796 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 30360 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 31096 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 32292 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 30728 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 29716 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 27508 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 26864 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 41492 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 30820 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 29992 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 31372 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 33672 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 33488 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 34960 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 34868 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 32292 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 32476 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 37444 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 37168 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 37260 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 37996 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 37628 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 37720 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 35788 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 33580 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 35604 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 37904 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 37996 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 40020 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 38824 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 37720 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 38180 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 40020 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 37720 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 37444 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 37076 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 32292 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 29348 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 25668 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24840 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23920 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24564 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23920 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24564 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24564 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23552 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22356 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21344 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19412 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19320 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20332 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20332 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13064 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12972 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14260 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12604 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11040 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10488 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11960 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13800 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14628 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 15180 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30728 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 27232 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_2_
timestamp 1679235063
transform 1 0 22724 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_1.mux_l1_in_3__250
timestamp 1679235063
transform 1 0 26128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_3_
timestamp 1679235063
transform 1 0 20884 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 25852 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l2_in_1_
timestamp 1679235063
transform 1 0 23092 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18584 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27140 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_3.mux_l2_in_1__203
timestamp 1679235063
transform 1 0 10948 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l2_in_1_
timestamp 1679235063
transform 1 0 17848 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25576 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24656 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21068 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l2_in_1_
timestamp 1679235063
transform 1 0 18124 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_5.mux_l2_in_1__206
timestamp 1679235063
transform 1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l3_in_0_
timestamp 1679235063
transform 1 0 17388 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8464 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27140 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24656 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_2_
timestamp 1679235063
transform 1 0 18124 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23000 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_7.mux_l2_in_1__208
timestamp 1679235063
transform 1 0 19044 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l2_in_1_
timestamp 1679235063
transform 1 0 19504 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19780 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27968 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_1_
timestamp 1679235063
transform 1 0 25852 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_2_
timestamp 1679235063
transform 1 0 20700 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_11.mux_l1_in_3__251
timestamp 1679235063
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_3_
timestamp 1679235063
transform 1 0 20700 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23184 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l2_in_1_
timestamp 1679235063
transform 1 0 19504 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27140 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24748 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_2_
timestamp 1679235063
transform 1 0 21160 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_13.mux_l2_in_1__252
timestamp 1679235063
transform 1 0 9200 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l2_in_1_
timestamp 1679235063
transform 1 0 19780 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l3_in_0_
timestamp 1679235063
transform 1 0 16928 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7084 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27876 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_2_
timestamp 1679235063
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22540 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l2_in_1_
timestamp 1679235063
transform 1 0 18124 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_21.mux_l2_in_1__253
timestamp 1679235063
transform 1 0 8372 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l3_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5152 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_0_
timestamp 1679235063
transform 1 0 29532 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_1_
timestamp 1679235063
transform 1 0 26772 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_2_
timestamp 1679235063
transform 1 0 24104 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l2_in_0_
timestamp 1679235063
transform 1 0 25668 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l2_in_1_
timestamp 1679235063
transform 1 0 25760 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_29.mux_l2_in_1__254
timestamp 1679235063
transform 1 0 23828 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l3_in_0_
timestamp 1679235063
transform 1 0 22264 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9844 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l1_in_0_
timestamp 1679235063
transform 1 0 32292 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l1_in_1_
timestamp 1679235063
transform 1 0 29716 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l2_in_0_
timestamp 1679235063
transform 1 0 28336 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_37.mux_l2_in_1__204
timestamp 1679235063
transform 1 0 22264 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l2_in_1_
timestamp 1679235063
transform 1 0 22908 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l3_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17204 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l1_in_0_
timestamp 1679235063
transform 1 0 32292 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l2_in_0_
timestamp 1679235063
transform 1 0 28336 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_45.mux_l2_in_1__205
timestamp 1679235063
transform 1 0 31556 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l2_in_1_
timestamp 1679235063
transform 1 0 28336 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l3_in_0_
timestamp 1679235063
transform 1 0 26864 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30268 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l2_in_0_
timestamp 1679235063
transform 1 0 25944 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l2_in_1_
timestamp 1679235063
transform 1 0 20700 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_53.mux_l2_in_1__207
timestamp 1679235063
transform 1 0 24012 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19964 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7636 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 29440 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 35696 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 27876 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 31280 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_0.mux_l2_in_1__209
timestamp 1679235063
transform 1 0 29808 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 30912 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 33488 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 39284 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 33212 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 32292 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 29716 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 34684 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_2.mux_l2_in_1__212
timestamp 1679235063
transform 1 0 34868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 33488 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 37996 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 42596 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 34408 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 36248 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_2_
timestamp 1679235063
transform 1 0 31004 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 35972 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_4.mux_l2_in_1__216
timestamp 1679235063
transform 1 0 33856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l2_in_1_
timestamp 1679235063
transform 1 0 37076 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l3_in_0_
timestamp 1679235063
transform 1 0 38640 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 41308 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 34868 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 32752 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_2_
timestamp 1679235063
transform 1 0 33488 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_6.mux_l1_in_3__219
timestamp 1679235063
transform 1 0 32568 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_3_
timestamp 1679235063
transform 1 0 32936 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 35880 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 38640 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 37444 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 41400 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 33396 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 32660 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_2_
timestamp 1679235063
transform 1 0 33304 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_3_
timestamp 1679235063
transform 1 0 31004 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_10.mux_l1_in_3__210
timestamp 1679235063
transform 1 0 31372 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 34500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l2_in_1_
timestamp 1679235063
transform 1 0 34868 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l3_in_0_
timestamp 1679235063
transform 1 0 36064 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 41492 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 32108 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_1_
timestamp 1679235063
transform 1 0 32292 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_2_
timestamp 1679235063
transform 1 0 27140 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 33304 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l2_in_1_
timestamp 1679235063
transform 1 0 30912 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_12.mux_l2_in_1__211
timestamp 1679235063
transform 1 0 29716 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l3_in_0_
timestamp 1679235063
transform 1 0 35880 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 40756 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30636 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_1_
timestamp 1679235063
transform 1 0 29716 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_2_
timestamp 1679235063
transform 1 0 27140 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 30544 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_20.mux_l2_in_1__213
timestamp 1679235063
transform 1 0 31556 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l2_in_1_
timestamp 1679235063
transform 1 0 28428 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l3_in_0_
timestamp 1679235063
transform 1 0 33488 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 39284 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 29716 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_1_
timestamp 1679235063
transform 1 0 30268 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_2_
timestamp 1679235063
transform 1 0 25760 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 29716 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l2_in_1_
timestamp 1679235063
transform 1 0 28336 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_28.mux_l2_in_1__214
timestamp 1679235063
transform 1 0 29624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l3_in_0_
timestamp 1679235063
transform 1 0 32568 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 37628 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30912 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l1_in_1_
timestamp 1679235063
transform 1 0 32108 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l2_in_0_
timestamp 1679235063
transform 1 0 33488 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_36.mux_l2_in_1__215
timestamp 1679235063
transform 1 0 33304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l2_in_1_
timestamp 1679235063
transform 1 0 31004 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l3_in_0_
timestamp 1679235063
transform 1 0 34868 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 38916 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 29716 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l1_in_1_
timestamp 1679235063
transform 1 0 28152 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_44.mux_l1_in_1__217
timestamp 1679235063
transform 1 0 28980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 32292 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 37444 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l1_in_0_
timestamp 1679235063
transform 1 0 28612 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l1_in_1_
timestamp 1679235063
transform 1 0 26956 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_52.mux_l1_in_1__218
timestamp 1679235063
transform 1 0 26404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l2_in_0_
timestamp 1679235063
transform 1 0 30820 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 36616 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 34868 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 38824 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 23276 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_0.mux_l1_in_3__220
timestamp 1679235063
transform 1 0 32292 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 28428 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 35880 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 28336 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 29716 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 42596 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 34868 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 40020 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 30912 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 37444 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_2.mux_l2_in_1__226
timestamp 1679235063
transform 1 0 42412 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 33028 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 32292 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 27876 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 36064 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 40020 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 35696 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l2_in_1_
timestamp 1679235063
transform 1 0 30912 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_4.mux_l2_in_1__236
timestamp 1679235063
transform 1 0 33764 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l3_in_0_
timestamp 1679235063
transform 1 0 30728 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 29348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 40204 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 41216 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_2_
timestamp 1679235063
transform 1 0 33488 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 39652 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 36064 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_6.mux_l2_in_1__244
timestamp 1679235063
transform 1 0 39192 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 33580 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 42596 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1679235063
transform 1 0 37444 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_1_
timestamp 1679235063
transform 1 0 41216 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_2_
timestamp 1679235063
transform 1 0 33304 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 40020 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l2_in_1_
timestamp 1679235063
transform 1 0 36064 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_8.mux_l2_in_1__245
timestamp 1679235063
transform 1 0 42596 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l3_in_0_
timestamp 1679235063
transform 1 0 36064 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 42412 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 34868 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 40112 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 36064 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_10.mux_l2_in_1__221
timestamp 1679235063
transform 1 0 31372 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l2_in_1_
timestamp 1679235063
transform 1 0 30176 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l3_in_0_
timestamp 1679235063
transform 1 0 32108 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 24932 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 40020 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 40388 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_12.mux_l2_in_1__222
timestamp 1679235063
transform 1 0 34868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l2_in_1_
timestamp 1679235063
transform 1 0 37444 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l3_in_0_
timestamp 1679235063
transform 1 0 37260 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 44344 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 39928 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 40480 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_14.mux_l2_in_1__223
timestamp 1679235063
transform 1 0 34132 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l2_in_1_
timestamp 1679235063
transform 1 0 34684 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l3_in_0_
timestamp 1679235063
transform 1 0 35880 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 39192 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1679235063
transform 1 0 38456 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 40480 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_16.mux_l2_in_1__224
timestamp 1679235063
transform 1 0 31556 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l2_in_1_
timestamp 1679235063
transform 1 0 37444 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l3_in_0_
timestamp 1679235063
transform 1 0 35880 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 37996 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 39652 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l2_in_1_
timestamp 1679235063
transform 1 0 32292 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_18.mux_l2_in_1__225
timestamp 1679235063
transform 1 0 29716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l3_in_0_
timestamp 1679235063
transform 1 0 32292 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 26036 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27324 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_20.mux_l1_in_1__227
timestamp 1679235063
transform 1 0 24196 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24840 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24840 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21988 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25852 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_22.mux_l1_in_1__228
timestamp 1679235063
transform 1 0 24564 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l1_in_1_
timestamp 1679235063
transform 1 0 23276 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23092 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27140 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l1_in_1_
timestamp 1679235063
transform 1 0 22080 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_24.mux_l1_in_1__229
timestamp 1679235063
transform 1 0 22540 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 22356 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27416 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24196 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_26.mux_l1_in_1__230
timestamp 1679235063
transform 1 0 24656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21896 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23092 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_28.mux_l2_in_0__231
timestamp 1679235063
transform 1 0 19688 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 12328 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21620 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_30.mux_l2_in_0__232
timestamp 1679235063
transform 1 0 11684 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16928 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11960 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16928 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_32.mux_l2_in_0__233
timestamp 1679235063
transform 1 0 16100 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9200 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19504 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19136 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_34.mux_l2_in_0__234
timestamp 1679235063
transform 1 0 19596 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9752 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25852 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l1_in_1_
timestamp 1679235063
transform 1 0 21988 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_36.mux_l1_in_1__235
timestamp 1679235063
transform 1 0 26404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20608 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9200 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_40.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_40.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11960 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_40.mux_l2_in_0__237
timestamp 1679235063
transform 1 0 13340 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6808 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_42.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_42.mux_l2_in_0__238
timestamp 1679235063
transform 1 0 7452 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_42.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14812 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4508 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12420 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_44.mux_l2_in_0__239
timestamp 1679235063
transform 1 0 5796 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6992 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11776 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_46.mux_l2_in_0__240
timestamp 1679235063
transform 1 0 7728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9844 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16468 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_48.mux_l2_in_0__241
timestamp 1679235063
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7084 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17664 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_50.mux_l2_in_0__242
timestamp 1679235063
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14720 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_58.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_58.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16928 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_58.mux_l2_in_0__243
timestamp 1679235063
transform 1 0 9200 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4600 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1679235063
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1679235063
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1679235063
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1679235063
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1679235063
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1679235063
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1679235063
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1679235063
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1679235063
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1679235063
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1679235063
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1679235063
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1679235063
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1679235063
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1679235063
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1679235063
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1679235063
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1679235063
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1679235063
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1679235063
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1679235063
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1679235063
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1679235063
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1679235063
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1679235063
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1679235063
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1679235063
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1679235063
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1679235063
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1679235063
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1679235063
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1679235063
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1679235063
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1679235063
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1679235063
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1679235063
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1679235063
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1679235063
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1679235063
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1679235063
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1679235063
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1679235063
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1679235063
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1679235063
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1679235063
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1679235063
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1679235063
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1679235063
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1679235063
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1679235063
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1679235063
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1679235063
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1679235063
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1679235063
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1679235063
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1679235063
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1679235063
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1679235063
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1679235063
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1679235063
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1679235063
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1679235063
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1679235063
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1679235063
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1679235063
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1679235063
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1679235063
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1679235063
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1679235063
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1679235063
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1679235063
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1679235063
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1679235063
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1679235063
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1679235063
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1679235063
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1679235063
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1679235063
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1679235063
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1679235063
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1679235063
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1679235063
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1679235063
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1679235063
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1679235063
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1679235063
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1679235063
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1679235063
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1679235063
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1679235063
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1679235063
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1679235063
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1679235063
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1679235063
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1679235063
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1679235063
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1679235063
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1679235063
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1679235063
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1679235063
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1679235063
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1679235063
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1679235063
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1679235063
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1679235063
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1679235063
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1679235063
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1679235063
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1679235063
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1679235063
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1679235063
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1679235063
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1679235063
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1679235063
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1679235063
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1679235063
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1679235063
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1679235063
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1679235063
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1679235063
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1679235063
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1679235063
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1679235063
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1679235063
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1679235063
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1679235063
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1679235063
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1679235063
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1679235063
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1679235063
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1679235063
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1679235063
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1679235063
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1679235063
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1679235063
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1679235063
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1679235063
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1679235063
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1679235063
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1679235063
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1679235063
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1679235063
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1679235063
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1679235063
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1679235063
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1679235063
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1679235063
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1679235063
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1679235063
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1679235063
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1679235063
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1679235063
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1679235063
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1679235063
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1679235063
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1679235063
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1679235063
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1679235063
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1679235063
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1679235063
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1679235063
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1679235063
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1679235063
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1679235063
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1679235063
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1679235063
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1679235063
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1679235063
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1679235063
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1679235063
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1679235063
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1679235063
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1679235063
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1679235063
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1679235063
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1679235063
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1679235063
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1679235063
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1679235063
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1679235063
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1679235063
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1679235063
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1679235063
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1679235063
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1679235063
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1679235063
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1679235063
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1679235063
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1679235063
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1679235063
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1679235063
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1679235063
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1679235063
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1679235063
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1679235063
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1679235063
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1679235063
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1679235063
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1679235063
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1679235063
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1679235063
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1679235063
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1679235063
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1679235063
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1679235063
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1679235063
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1679235063
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1679235063
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1679235063
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1679235063
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1679235063
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1679235063
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1679235063
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1679235063
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1679235063
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1679235063
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1679235063
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1679235063
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1679235063
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1679235063
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1679235063
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1679235063
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1679235063
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1679235063
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1679235063
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1679235063
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1679235063
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1679235063
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1679235063
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1679235063
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1679235063
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1679235063
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1679235063
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1679235063
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1679235063
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1679235063
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1679235063
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1679235063
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1679235063
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1679235063
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1679235063
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1679235063
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1679235063
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1679235063
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1679235063
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1679235063
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1679235063
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1679235063
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1679235063
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1679235063
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1679235063
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1679235063
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1679235063
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1679235063
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1679235063
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1679235063
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1679235063
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1679235063
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1679235063
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1679235063
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1679235063
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1679235063
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1679235063
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1679235063
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1679235063
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1679235063
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1679235063
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1679235063
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1679235063
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1679235063
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1679235063
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1679235063
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1679235063
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1679235063
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1679235063
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1679235063
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1679235063
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1679235063
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1679235063
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1679235063
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1679235063
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1679235063
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1679235063
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1679235063
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1679235063
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1679235063
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1679235063
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1679235063
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1679235063
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1679235063
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1679235063
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1679235063
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1679235063
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1679235063
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1679235063
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1679235063
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1679235063
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1679235063
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1679235063
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1679235063
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1679235063
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1679235063
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1679235063
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1679235063
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1679235063
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1679235063
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1679235063
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1679235063
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1679235063
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1679235063
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1679235063
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1679235063
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1679235063
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1679235063
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1679235063
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1679235063
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1679235063
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1679235063
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1679235063
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1679235063
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1679235063
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1679235063
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1679235063
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1679235063
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1679235063
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1679235063
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1679235063
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1679235063
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1679235063
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1679235063
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1679235063
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1679235063
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1679235063
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1679235063
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1679235063
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1679235063
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1679235063
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1679235063
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1679235063
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1679235063
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1679235063
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1679235063
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1679235063
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1679235063
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1679235063
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1679235063
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1679235063
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1679235063
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1679235063
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1679235063
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1679235063
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1679235063
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1679235063
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1679235063
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1679235063
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1679235063
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1679235063
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1679235063
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1679235063
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1679235063
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1679235063
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1679235063
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1679235063
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1679235063
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1679235063
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1679235063
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1679235063
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1679235063
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1679235063
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1679235063
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1679235063
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1679235063
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1679235063
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1679235063
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1679235063
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1679235063
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1679235063
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1679235063
transform 1 0 26864 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1679235063
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1679235063
transform 1 0 32016 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1679235063
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1679235063
transform 1 0 37168 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1679235063
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1679235063
transform 1 0 42320 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1679235063
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1679235063
transform 1 0 47472 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 49238 26200 49294 27000 0 FreeSans 224 90 0 0 ccff_head_1
port 3 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1582 26200 1638 27000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[20]
port 18 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[21]
port 19 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[22]
port 20 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[23]
port 21 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[24]
port 22 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[25]
port 23 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[26]
port 24 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[27]
port 25 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[28]
port 26 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[29]
port 27 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 28 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 29 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 30 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 31 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 32 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 33 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 34 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 35 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 36 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 37 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 38 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 39 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 40 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 41 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 42 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 43 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 44 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 45 nsew signal tristate
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 46 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 47 nsew signal tristate
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 chanx_left_out[20]
port 48 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 chanx_left_out[21]
port 49 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 chanx_left_out[22]
port 50 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_out[23]
port 51 nsew signal tristate
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 chanx_left_out[24]
port 52 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 chanx_left_out[25]
port 53 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 chanx_left_out[26]
port 54 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 chanx_left_out[27]
port 55 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_out[28]
port 56 nsew signal tristate
flabel metal3 s 0 25576 800 25696 0 FreeSans 480 0 0 0 chanx_left_out[29]
port 57 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal3 s 50200 13608 51000 13728 0 FreeSans 480 0 0 0 chanx_right_in_0[0]
port 66 nsew signal input
flabel metal3 s 50200 17688 51000 17808 0 FreeSans 480 0 0 0 chanx_right_in_0[10]
port 67 nsew signal input
flabel metal3 s 50200 18096 51000 18216 0 FreeSans 480 0 0 0 chanx_right_in_0[11]
port 68 nsew signal input
flabel metal3 s 50200 18504 51000 18624 0 FreeSans 480 0 0 0 chanx_right_in_0[12]
port 69 nsew signal input
flabel metal3 s 50200 18912 51000 19032 0 FreeSans 480 0 0 0 chanx_right_in_0[13]
port 70 nsew signal input
flabel metal3 s 50200 19320 51000 19440 0 FreeSans 480 0 0 0 chanx_right_in_0[14]
port 71 nsew signal input
flabel metal3 s 50200 19728 51000 19848 0 FreeSans 480 0 0 0 chanx_right_in_0[15]
port 72 nsew signal input
flabel metal3 s 50200 20136 51000 20256 0 FreeSans 480 0 0 0 chanx_right_in_0[16]
port 73 nsew signal input
flabel metal3 s 50200 20544 51000 20664 0 FreeSans 480 0 0 0 chanx_right_in_0[17]
port 74 nsew signal input
flabel metal3 s 50200 20952 51000 21072 0 FreeSans 480 0 0 0 chanx_right_in_0[18]
port 75 nsew signal input
flabel metal3 s 50200 21360 51000 21480 0 FreeSans 480 0 0 0 chanx_right_in_0[19]
port 76 nsew signal input
flabel metal3 s 50200 14016 51000 14136 0 FreeSans 480 0 0 0 chanx_right_in_0[1]
port 77 nsew signal input
flabel metal3 s 50200 21768 51000 21888 0 FreeSans 480 0 0 0 chanx_right_in_0[20]
port 78 nsew signal input
flabel metal3 s 50200 22176 51000 22296 0 FreeSans 480 0 0 0 chanx_right_in_0[21]
port 79 nsew signal input
flabel metal3 s 50200 22584 51000 22704 0 FreeSans 480 0 0 0 chanx_right_in_0[22]
port 80 nsew signal input
flabel metal3 s 50200 22992 51000 23112 0 FreeSans 480 0 0 0 chanx_right_in_0[23]
port 81 nsew signal input
flabel metal3 s 50200 23400 51000 23520 0 FreeSans 480 0 0 0 chanx_right_in_0[24]
port 82 nsew signal input
flabel metal3 s 50200 23808 51000 23928 0 FreeSans 480 0 0 0 chanx_right_in_0[25]
port 83 nsew signal input
flabel metal3 s 50200 24216 51000 24336 0 FreeSans 480 0 0 0 chanx_right_in_0[26]
port 84 nsew signal input
flabel metal3 s 50200 24624 51000 24744 0 FreeSans 480 0 0 0 chanx_right_in_0[27]
port 85 nsew signal input
flabel metal3 s 50200 25032 51000 25152 0 FreeSans 480 0 0 0 chanx_right_in_0[28]
port 86 nsew signal input
flabel metal3 s 50200 25440 51000 25560 0 FreeSans 480 0 0 0 chanx_right_in_0[29]
port 87 nsew signal input
flabel metal3 s 50200 14424 51000 14544 0 FreeSans 480 0 0 0 chanx_right_in_0[2]
port 88 nsew signal input
flabel metal3 s 50200 14832 51000 14952 0 FreeSans 480 0 0 0 chanx_right_in_0[3]
port 89 nsew signal input
flabel metal3 s 50200 15240 51000 15360 0 FreeSans 480 0 0 0 chanx_right_in_0[4]
port 90 nsew signal input
flabel metal3 s 50200 15648 51000 15768 0 FreeSans 480 0 0 0 chanx_right_in_0[5]
port 91 nsew signal input
flabel metal3 s 50200 16056 51000 16176 0 FreeSans 480 0 0 0 chanx_right_in_0[6]
port 92 nsew signal input
flabel metal3 s 50200 16464 51000 16584 0 FreeSans 480 0 0 0 chanx_right_in_0[7]
port 93 nsew signal input
flabel metal3 s 50200 16872 51000 16992 0 FreeSans 480 0 0 0 chanx_right_in_0[8]
port 94 nsew signal input
flabel metal3 s 50200 17280 51000 17400 0 FreeSans 480 0 0 0 chanx_right_in_0[9]
port 95 nsew signal input
flabel metal3 s 50200 1368 51000 1488 0 FreeSans 480 0 0 0 chanx_right_out_0[0]
port 96 nsew signal tristate
flabel metal3 s 50200 5448 51000 5568 0 FreeSans 480 0 0 0 chanx_right_out_0[10]
port 97 nsew signal tristate
flabel metal3 s 50200 5856 51000 5976 0 FreeSans 480 0 0 0 chanx_right_out_0[11]
port 98 nsew signal tristate
flabel metal3 s 50200 6264 51000 6384 0 FreeSans 480 0 0 0 chanx_right_out_0[12]
port 99 nsew signal tristate
flabel metal3 s 50200 6672 51000 6792 0 FreeSans 480 0 0 0 chanx_right_out_0[13]
port 100 nsew signal tristate
flabel metal3 s 50200 7080 51000 7200 0 FreeSans 480 0 0 0 chanx_right_out_0[14]
port 101 nsew signal tristate
flabel metal3 s 50200 7488 51000 7608 0 FreeSans 480 0 0 0 chanx_right_out_0[15]
port 102 nsew signal tristate
flabel metal3 s 50200 7896 51000 8016 0 FreeSans 480 0 0 0 chanx_right_out_0[16]
port 103 nsew signal tristate
flabel metal3 s 50200 8304 51000 8424 0 FreeSans 480 0 0 0 chanx_right_out_0[17]
port 104 nsew signal tristate
flabel metal3 s 50200 8712 51000 8832 0 FreeSans 480 0 0 0 chanx_right_out_0[18]
port 105 nsew signal tristate
flabel metal3 s 50200 9120 51000 9240 0 FreeSans 480 0 0 0 chanx_right_out_0[19]
port 106 nsew signal tristate
flabel metal3 s 50200 1776 51000 1896 0 FreeSans 480 0 0 0 chanx_right_out_0[1]
port 107 nsew signal tristate
flabel metal3 s 50200 9528 51000 9648 0 FreeSans 480 0 0 0 chanx_right_out_0[20]
port 108 nsew signal tristate
flabel metal3 s 50200 9936 51000 10056 0 FreeSans 480 0 0 0 chanx_right_out_0[21]
port 109 nsew signal tristate
flabel metal3 s 50200 10344 51000 10464 0 FreeSans 480 0 0 0 chanx_right_out_0[22]
port 110 nsew signal tristate
flabel metal3 s 50200 10752 51000 10872 0 FreeSans 480 0 0 0 chanx_right_out_0[23]
port 111 nsew signal tristate
flabel metal3 s 50200 11160 51000 11280 0 FreeSans 480 0 0 0 chanx_right_out_0[24]
port 112 nsew signal tristate
flabel metal3 s 50200 11568 51000 11688 0 FreeSans 480 0 0 0 chanx_right_out_0[25]
port 113 nsew signal tristate
flabel metal3 s 50200 11976 51000 12096 0 FreeSans 480 0 0 0 chanx_right_out_0[26]
port 114 nsew signal tristate
flabel metal3 s 50200 12384 51000 12504 0 FreeSans 480 0 0 0 chanx_right_out_0[27]
port 115 nsew signal tristate
flabel metal3 s 50200 12792 51000 12912 0 FreeSans 480 0 0 0 chanx_right_out_0[28]
port 116 nsew signal tristate
flabel metal3 s 50200 13200 51000 13320 0 FreeSans 480 0 0 0 chanx_right_out_0[29]
port 117 nsew signal tristate
flabel metal3 s 50200 2184 51000 2304 0 FreeSans 480 0 0 0 chanx_right_out_0[2]
port 118 nsew signal tristate
flabel metal3 s 50200 2592 51000 2712 0 FreeSans 480 0 0 0 chanx_right_out_0[3]
port 119 nsew signal tristate
flabel metal3 s 50200 3000 51000 3120 0 FreeSans 480 0 0 0 chanx_right_out_0[4]
port 120 nsew signal tristate
flabel metal3 s 50200 3408 51000 3528 0 FreeSans 480 0 0 0 chanx_right_out_0[5]
port 121 nsew signal tristate
flabel metal3 s 50200 3816 51000 3936 0 FreeSans 480 0 0 0 chanx_right_out_0[6]
port 122 nsew signal tristate
flabel metal3 s 50200 4224 51000 4344 0 FreeSans 480 0 0 0 chanx_right_out_0[7]
port 123 nsew signal tristate
flabel metal3 s 50200 4632 51000 4752 0 FreeSans 480 0 0 0 chanx_right_out_0[8]
port 124 nsew signal tristate
flabel metal3 s 50200 5040 51000 5160 0 FreeSans 480 0 0 0 chanx_right_out_0[9]
port 125 nsew signal tristate
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 126 nsew signal input
flabel metal2 s 27986 26200 28042 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 127 nsew signal input
flabel metal2 s 28630 26200 28686 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 128 nsew signal input
flabel metal2 s 29274 26200 29330 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 129 nsew signal input
flabel metal2 s 29918 26200 29974 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 130 nsew signal input
flabel metal2 s 30562 26200 30618 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 131 nsew signal input
flabel metal2 s 31206 26200 31262 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 132 nsew signal input
flabel metal2 s 31850 26200 31906 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 133 nsew signal input
flabel metal2 s 32494 26200 32550 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 134 nsew signal input
flabel metal2 s 33138 26200 33194 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 135 nsew signal input
flabel metal2 s 33782 26200 33838 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 136 nsew signal input
flabel metal2 s 22190 26200 22246 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 137 nsew signal input
flabel metal2 s 34426 26200 34482 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 138 nsew signal input
flabel metal2 s 35070 26200 35126 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 139 nsew signal input
flabel metal2 s 35714 26200 35770 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 140 nsew signal input
flabel metal2 s 36358 26200 36414 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 141 nsew signal input
flabel metal2 s 37002 26200 37058 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 142 nsew signal input
flabel metal2 s 37646 26200 37702 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 143 nsew signal input
flabel metal2 s 38290 26200 38346 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 144 nsew signal input
flabel metal2 s 38934 26200 38990 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 145 nsew signal input
flabel metal2 s 39578 26200 39634 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 146 nsew signal input
flabel metal2 s 40222 26200 40278 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 147 nsew signal input
flabel metal2 s 22834 26200 22890 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 148 nsew signal input
flabel metal2 s 23478 26200 23534 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 149 nsew signal input
flabel metal2 s 24122 26200 24178 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 150 nsew signal input
flabel metal2 s 24766 26200 24822 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 151 nsew signal input
flabel metal2 s 25410 26200 25466 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 152 nsew signal input
flabel metal2 s 26054 26200 26110 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 153 nsew signal input
flabel metal2 s 26698 26200 26754 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 154 nsew signal input
flabel metal2 s 27342 26200 27398 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 155 nsew signal input
flabel metal2 s 2226 26200 2282 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 156 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 157 nsew signal tristate
flabel metal2 s 9310 26200 9366 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 158 nsew signal tristate
flabel metal2 s 9954 26200 10010 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 159 nsew signal tristate
flabel metal2 s 10598 26200 10654 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 160 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 161 nsew signal tristate
flabel metal2 s 11886 26200 11942 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 162 nsew signal tristate
flabel metal2 s 12530 26200 12586 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 163 nsew signal tristate
flabel metal2 s 13174 26200 13230 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 164 nsew signal tristate
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 165 nsew signal tristate
flabel metal2 s 14462 26200 14518 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 166 nsew signal tristate
flabel metal2 s 2870 26200 2926 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 167 nsew signal tristate
flabel metal2 s 15106 26200 15162 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 168 nsew signal tristate
flabel metal2 s 15750 26200 15806 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 169 nsew signal tristate
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 170 nsew signal tristate
flabel metal2 s 17038 26200 17094 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 171 nsew signal tristate
flabel metal2 s 17682 26200 17738 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 172 nsew signal tristate
flabel metal2 s 18326 26200 18382 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 173 nsew signal tristate
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 174 nsew signal tristate
flabel metal2 s 19614 26200 19670 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 175 nsew signal tristate
flabel metal2 s 20258 26200 20314 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 176 nsew signal tristate
flabel metal2 s 20902 26200 20958 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 177 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 178 nsew signal tristate
flabel metal2 s 4158 26200 4214 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 179 nsew signal tristate
flabel metal2 s 4802 26200 4858 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 180 nsew signal tristate
flabel metal2 s 5446 26200 5502 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 181 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 182 nsew signal tristate
flabel metal2 s 6734 26200 6790 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 183 nsew signal tristate
flabel metal2 s 7378 26200 7434 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 184 nsew signal tristate
flabel metal2 s 8022 26200 8078 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 185 nsew signal tristate
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 42154 26200 42210 27000 0 FreeSans 224 90 0 0 prog_reset
port 200 nsew signal input
flabel metal2 s 42798 26200 42854 27000 0 FreeSans 224 90 0 0 reset
port 201 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 202 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 203 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 204 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 205 nsew signal input
flabel metal2 s 43442 26200 43498 27000 0 FreeSans 224 90 0 0 test_enable
port 206 nsew signal input
flabel metal2 s 45374 26200 45430 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 207 nsew signal input
flabel metal2 s 46018 26200 46074 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 208 nsew signal input
flabel metal2 s 46662 26200 46718 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 209 nsew signal input
flabel metal2 s 47306 26200 47362 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 210 nsew signal input
flabel metal2 s 47950 26200 48006 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 211 nsew signal input
flabel metal2 s 48594 26200 48650 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 212 nsew signal input
flabel metal2 s 44086 26200 44142 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 213 nsew signal input
flabel metal2 s 44730 26200 44786 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 214 nsew signal input
flabel metal2 s 1122 0 1178 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_inpad_0_
port 215 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_1__pin_inpad_0_
port 216 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_2__pin_inpad_0_
port 217 nsew signal tristate
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_3__pin_inpad_0_
port 218 nsew signal tristate
rlabel metal1 25484 23936 25484 23936 0 VGND
rlabel metal1 25484 24480 25484 24480 0 VPWR
rlabel metal2 22770 4556 22770 4556 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal2 21206 4862 21206 4862 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 19596 3026 19596 3026 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 17434 4114 17434 4114 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 20516 22066 20516 22066 0 cbx_1__0_.cbx_8__0_.ccff_head
rlabel metal2 18630 8092 18630 8092 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
rlabel metal1 20332 19414 20332 19414 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
rlabel metal1 18308 13838 18308 13838 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
rlabel metal1 17618 10234 17618 10234 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
rlabel metal2 16054 8364 16054 8364 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
rlabel metal2 16238 15606 16238 15606 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
rlabel metal1 13800 12274 13800 12274 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
rlabel metal1 13984 8466 13984 8466 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
rlabel metal1 13248 9486 13248 9486 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
rlabel metal2 16974 14144 16974 14144 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
rlabel metal1 11638 12274 11638 12274 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
rlabel metal2 12282 11356 12282 11356 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
rlabel metal1 16284 16014 16284 16014 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
rlabel metal2 13754 15742 13754 15742 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
rlabel metal1 13064 15538 13064 15538 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
rlabel metal2 15686 14790 15686 14790 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18262 7480 18262 7480 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 20010 6290 20010 6290 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 15916 13294 15916 13294 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18446 13974 18446 13974 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19504 14042 19504 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17020 12614 17020 12614 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15042 10778 15042 10778 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 17848 14042 17848 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 18722 7786 18722 7786 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 18492 7514 18492 7514 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 19918 7956 19918 7956 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 12236 14314 12236 14314 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15594 7854 15594 7854 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 18124 6290 18124 6290 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 12098 14382 12098 14382 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18262 13294 18262 13294 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 17986 13634 17986 13634 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13478 12342 13478 12342 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13110 10778 13110 10778 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 14122 10642 14122 10642 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 15916 8602 15916 8602 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 15778 9792 15778 9792 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 15364 7922 15364 7922 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 9430 15062 9430 15062 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12788 9622 12788 9622 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 15180 7378 15180 7378 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 9890 15538 9890 15538 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13478 14484 13478 14484 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13938 14314 13938 14314 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16422 9894 16422 9894 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10672 12954 10672 12954 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11086 12818 11086 12818 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 12926 10234 12926 10234 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 12052 10778 12052 10778 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 12742 9554 12742 9554 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 13340 16150 13340 16150 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11546 16048 11546 16048 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 15870 8874 15870 8874 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13984 16218 13984 16218 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15870 15708 15870 15708 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18400 14858 18400 14858 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 15042 11356 15042 11356 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12834 16218 12834 16218 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 12374 15844 12374 15844 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 14030 15334 14030 15334 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 16008 13498 16008 13498 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 11822 16218 11822 16218 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 19458 3162 19458 3162 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 22126 2550 22126 2550 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 25691 3706 25691 3706 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 23230 2618 23230 2618 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 23138 2550 23138 2550 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 24633 4522 24633 4522 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 27002 2618 27002 2618 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 23690 2550 23690 2550 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal1 24288 4182 24288 4182 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 27186 2176 27186 2176 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 24196 3570 24196 3570 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 9798 2414 9798 2414 0 ccff_head
rlabel metal1 48576 22202 48576 22202 0 ccff_head_1
rlabel metal2 41354 1622 41354 1622 0 ccff_tail
rlabel metal1 3128 22202 3128 22202 0 ccff_tail_0
rlabel metal2 3266 2244 3266 2244 0 chanx_left_in[0]
rlabel metal1 1472 5678 1472 5678 0 chanx_left_in[10]
rlabel metal1 1472 6290 1472 6290 0 chanx_left_in[11]
rlabel metal1 1932 6766 1932 6766 0 chanx_left_in[12]
rlabel metal1 1472 6698 1472 6698 0 chanx_left_in[13]
rlabel metal1 1472 7378 1472 7378 0 chanx_left_in[14]
rlabel metal1 1472 7854 1472 7854 0 chanx_left_in[15]
rlabel metal1 1518 8398 1518 8398 0 chanx_left_in[16]
rlabel metal1 1794 8942 1794 8942 0 chanx_left_in[17]
rlabel metal1 1518 8874 1518 8874 0 chanx_left_in[18]
rlabel metal1 1518 9554 1518 9554 0 chanx_left_in[19]
rlabel metal1 2024 2414 2024 2414 0 chanx_left_in[1]
rlabel metal1 1472 10030 1472 10030 0 chanx_left_in[20]
rlabel metal1 2346 10676 2346 10676 0 chanx_left_in[21]
rlabel metal1 1472 10642 1472 10642 0 chanx_left_in[22]
rlabel metal2 1610 11033 1610 11033 0 chanx_left_in[23]
rlabel metal1 2530 11696 2530 11696 0 chanx_left_in[24]
rlabel metal1 1472 12206 1472 12206 0 chanx_left_in[25]
rlabel metal1 1426 11730 1426 11730 0 chanx_left_in[26]
rlabel metal2 1334 12699 1334 12699 0 chanx_left_in[27]
rlabel metal1 1426 12750 1426 12750 0 chanx_left_in[28]
rlabel metal3 1564 13328 1564 13328 0 chanx_left_in[29]
rlabel metal1 1610 2448 1610 2448 0 chanx_left_in[2]
rlabel metal1 1472 3026 1472 3026 0 chanx_left_in[3]
rlabel metal1 1472 3502 1472 3502 0 chanx_left_in[4]
rlabel metal1 1840 4114 1840 4114 0 chanx_left_in[5]
rlabel metal1 1564 4182 1564 4182 0 chanx_left_in[6]
rlabel metal1 1472 4590 1472 4590 0 chanx_left_in[7]
rlabel metal1 1472 5134 1472 5134 0 chanx_left_in[8]
rlabel metal1 2576 5678 2576 5678 0 chanx_left_in[9]
rlabel metal2 2806 13583 2806 13583 0 chanx_left_out[0]
rlabel metal3 1694 17884 1694 17884 0 chanx_left_out[10]
rlabel metal2 2898 18819 2898 18819 0 chanx_left_out[11]
rlabel metal3 1004 18700 1004 18700 0 chanx_left_out[12]
rlabel metal3 1004 19108 1004 19108 0 chanx_left_out[13]
rlabel metal3 1694 19516 1694 19516 0 chanx_left_out[14]
rlabel metal3 1050 19924 1050 19924 0 chanx_left_out[15]
rlabel via2 3910 20349 3910 20349 0 chanx_left_out[16]
rlabel metal3 1004 20740 1004 20740 0 chanx_left_out[17]
rlabel metal1 2852 22542 2852 22542 0 chanx_left_out[18]
rlabel metal3 1694 21556 1694 21556 0 chanx_left_out[19]
rlabel metal3 820 14212 820 14212 0 chanx_left_out[1]
rlabel metal2 3818 22015 3818 22015 0 chanx_left_out[20]
rlabel metal3 1579 22372 1579 22372 0 chanx_left_out[21]
rlabel metal3 1924 22780 1924 22780 0 chanx_left_out[22]
rlabel metal3 2062 23188 2062 23188 0 chanx_left_out[23]
rlabel metal3 2062 23596 2062 23596 0 chanx_left_out[24]
rlabel metal3 2108 24004 2108 24004 0 chanx_left_out[25]
rlabel metal3 1740 24412 1740 24412 0 chanx_left_out[26]
rlabel metal3 2062 24820 2062 24820 0 chanx_left_out[27]
rlabel metal3 2154 25228 2154 25228 0 chanx_left_out[28]
rlabel metal3 1878 25636 1878 25636 0 chanx_left_out[29]
rlabel metal3 1004 14620 1004 14620 0 chanx_left_out[2]
rlabel metal3 1004 15028 1004 15028 0 chanx_left_out[3]
rlabel metal3 1004 15436 1004 15436 0 chanx_left_out[4]
rlabel metal3 1004 15844 1004 15844 0 chanx_left_out[5]
rlabel metal3 1004 16252 1004 16252 0 chanx_left_out[6]
rlabel metal3 1004 16660 1004 16660 0 chanx_left_out[7]
rlabel metal3 958 17068 958 17068 0 chanx_left_out[8]
rlabel metal2 2806 17833 2806 17833 0 chanx_left_out[9]
rlabel metal1 48438 13906 48438 13906 0 chanx_right_in_0[0]
rlabel metal2 49082 18003 49082 18003 0 chanx_right_in_0[10]
rlabel metal1 49128 18734 49128 18734 0 chanx_right_in_0[11]
rlabel metal2 48806 18479 48806 18479 0 chanx_right_in_0[12]
rlabel metal2 49174 19159 49174 19159 0 chanx_right_in_0[13]
rlabel metal1 49266 19754 49266 19754 0 chanx_right_in_0[14]
rlabel metal2 49082 20111 49082 20111 0 chanx_right_in_0[15]
rlabel metal2 48622 20315 48622 20315 0 chanx_right_in_0[16]
rlabel metal2 49082 20757 49082 20757 0 chanx_right_in_0[17]
rlabel metal1 48806 21522 48806 21522 0 chanx_right_in_0[18]
rlabel metal3 49734 21420 49734 21420 0 chanx_right_in_0[19]
rlabel metal2 49174 14025 49174 14025 0 chanx_right_in_0[1]
rlabel metal1 48668 19822 48668 19822 0 chanx_right_in_0[20]
rlabel metal1 48300 20502 48300 20502 0 chanx_right_in_0[21]
rlabel metal1 48714 21998 48714 21998 0 chanx_right_in_0[22]
rlabel via2 48346 23069 48346 23069 0 chanx_right_in_0[23]
rlabel metal1 47840 20910 47840 20910 0 chanx_right_in_0[24]
rlabel metal1 46506 20910 46506 20910 0 chanx_right_in_0[25]
rlabel metal1 47886 23290 47886 23290 0 chanx_right_in_0[26]
rlabel metal1 47702 21658 47702 21658 0 chanx_right_in_0[27]
rlabel metal1 47150 20910 47150 20910 0 chanx_right_in_0[28]
rlabel metal1 47104 20570 47104 20570 0 chanx_right_in_0[29]
rlabel metal2 49082 14433 49082 14433 0 chanx_right_in_0[2]
rlabel metal2 49082 14943 49082 14943 0 chanx_right_in_0[3]
rlabel metal2 49358 15385 49358 15385 0 chanx_right_in_0[4]
rlabel metal2 49082 15895 49082 15895 0 chanx_right_in_0[5]
rlabel metal1 49128 16558 49128 16558 0 chanx_right_in_0[6]
rlabel metal1 49220 17170 49220 17170 0 chanx_right_in_0[7]
rlabel metal2 48806 16847 48806 16847 0 chanx_right_in_0[8]
rlabel metal2 49082 17493 49082 17493 0 chanx_right_in_0[9]
rlabel metal2 46690 2737 46690 2737 0 chanx_right_out_0[0]
rlabel metal1 49312 4658 49312 4658 0 chanx_right_out_0[10]
rlabel metal2 49174 5593 49174 5593 0 chanx_right_out_0[11]
rlabel metal3 49596 6324 49596 6324 0 chanx_right_out_0[12]
rlabel metal1 49220 5746 49220 5746 0 chanx_right_out_0[13]
rlabel metal1 49266 6358 49266 6358 0 chanx_right_out_0[14]
rlabel metal3 49734 7548 49734 7548 0 chanx_right_out_0[15]
rlabel metal2 46874 8177 46874 8177 0 chanx_right_out_0[16]
rlabel metal1 49266 7446 49266 7446 0 chanx_right_out_0[17]
rlabel metal1 49220 7922 49220 7922 0 chanx_right_out_0[18]
rlabel metal2 49174 8857 49174 8857 0 chanx_right_out_0[19]
rlabel metal2 46782 2397 46782 2397 0 chanx_right_out_0[1]
rlabel metal3 48814 9588 48814 9588 0 chanx_right_out_0[20]
rlabel metal1 49220 9010 49220 9010 0 chanx_right_out_0[21]
rlabel metal1 49266 9622 49266 9622 0 chanx_right_out_0[22]
rlabel metal2 49174 10455 49174 10455 0 chanx_right_out_0[23]
rlabel metal1 49220 10710 49220 10710 0 chanx_right_out_0[24]
rlabel metal2 49174 11407 49174 11407 0 chanx_right_out_0[25]
rlabel metal2 49174 11917 49174 11917 0 chanx_right_out_0[26]
rlabel metal3 49734 12444 49734 12444 0 chanx_right_out_0[27]
rlabel via2 49174 12835 49174 12835 0 chanx_right_out_0[28]
rlabel metal3 49734 13260 49734 13260 0 chanx_right_out_0[29]
rlabel metal3 49412 2244 49412 2244 0 chanx_right_out_0[2]
rlabel metal2 46874 2805 46874 2805 0 chanx_right_out_0[3]
rlabel metal3 49504 3060 49504 3060 0 chanx_right_out_0[4]
rlabel metal2 49174 2975 49174 2975 0 chanx_right_out_0[5]
rlabel metal1 49220 3094 49220 3094 0 chanx_right_out_0[6]
rlabel metal2 49174 3927 49174 3927 0 chanx_right_out_0[7]
rlabel metal1 47610 5134 47610 5134 0 chanx_right_out_0[8]
rlabel metal1 49266 4114 49266 4114 0 chanx_right_out_0[9]
rlabel metal1 3956 22610 3956 22610 0 chany_top_in[0]
rlabel metal3 38548 23120 38548 23120 0 chany_top_in[10]
rlabel via1 28934 26299 28934 26299 0 chany_top_in[11]
rlabel metal1 43332 21998 43332 21998 0 chany_top_in[12]
rlabel metal2 30406 25840 30406 25840 0 chany_top_in[13]
rlabel metal3 38295 12716 38295 12716 0 chany_top_in[14]
rlabel via2 45862 21539 45862 21539 0 chany_top_in[15]
rlabel metal2 32154 25704 32154 25704 0 chany_top_in[16]
rlabel metal1 46230 21522 46230 21522 0 chany_top_in[17]
rlabel metal2 33442 26231 33442 26231 0 chany_top_in[18]
rlabel metal2 33810 26156 33810 26156 0 chany_top_in[19]
rlabel metal1 21942 17170 21942 17170 0 chany_top_in[1]
rlabel metal2 34454 26190 34454 26190 0 chany_top_in[20]
rlabel metal2 35466 24820 35466 24820 0 chany_top_in[21]
rlabel metal2 36018 25721 36018 25721 0 chany_top_in[22]
rlabel metal2 36754 25585 36754 25585 0 chany_top_in[23]
rlabel metal2 37030 26122 37030 26122 0 chany_top_in[24]
rlabel metal2 37674 25612 37674 25612 0 chany_top_in[25]
rlabel metal2 38502 24548 38502 24548 0 chany_top_in[26]
rlabel metal1 41354 22984 41354 22984 0 chany_top_in[27]
rlabel metal1 40434 22610 40434 22610 0 chany_top_in[28]
rlabel metal1 45540 21998 45540 21998 0 chany_top_in[29]
rlabel metal1 9200 23086 9200 23086 0 chany_top_in[2]
rlabel metal1 27094 21114 27094 21114 0 chany_top_in[3]
rlabel metal1 11776 22542 11776 22542 0 chany_top_in[4]
rlabel metal2 43930 24990 43930 24990 0 chany_top_in[5]
rlabel metal2 11822 24174 11822 24174 0 chany_top_in[6]
rlabel metal1 14122 22066 14122 22066 0 chany_top_in[7]
rlabel metal1 17112 24174 17112 24174 0 chany_top_in[8]
rlabel metal2 40066 25296 40066 25296 0 chany_top_in[9]
rlabel metal1 3404 22134 3404 22134 0 chany_top_out[0]
rlabel metal1 8464 24242 8464 24242 0 chany_top_out[10]
rlabel metal1 9246 23766 9246 23766 0 chany_top_out[11]
rlabel metal1 10120 22542 10120 22542 0 chany_top_out[12]
rlabel metal2 10718 25041 10718 25041 0 chany_top_out[13]
rlabel metal2 11270 24728 11270 24728 0 chany_top_out[14]
rlabel metal2 11914 24218 11914 24218 0 chany_top_out[15]
rlabel metal2 12558 25204 12558 25204 0 chany_top_out[16]
rlabel metal2 13386 24735 13386 24735 0 chany_top_out[17]
rlabel metal2 13846 24422 13846 24422 0 chany_top_out[18]
rlabel metal1 14030 24242 14030 24242 0 chany_top_out[19]
rlabel metal1 3588 22678 3588 22678 0 chany_top_out[1]
rlabel metal1 14536 23766 14536 23766 0 chany_top_out[20]
rlabel metal2 15870 24497 15870 24497 0 chany_top_out[21]
rlabel metal2 16422 24728 16422 24728 0 chany_top_out[22]
rlabel metal1 16606 23766 16606 23766 0 chany_top_out[23]
rlabel metal1 18308 21930 18308 21930 0 chany_top_out[24]
rlabel metal1 17250 24242 17250 24242 0 chany_top_out[25]
rlabel metal1 18584 23766 18584 23766 0 chany_top_out[26]
rlabel metal1 18998 24242 18998 24242 0 chany_top_out[27]
rlabel metal2 20286 25204 20286 25204 0 chany_top_out[28]
rlabel metal2 20930 25272 20930 25272 0 chany_top_out[29]
rlabel metal1 3404 24242 3404 24242 0 chany_top_out[2]
rlabel metal1 4094 23630 4094 23630 0 chany_top_out[3]
rlabel metal2 5106 24429 5106 24429 0 chany_top_out[4]
rlabel metal2 5474 24966 5474 24966 0 chany_top_out[5]
rlabel metal2 6118 24728 6118 24728 0 chany_top_out[6]
rlabel metal1 6164 24242 6164 24242 0 chany_top_out[7]
rlabel metal1 7820 22542 7820 22542 0 chany_top_out[8]
rlabel metal2 7866 23919 7866 23919 0 chany_top_out[9]
rlabel metal1 18170 16490 18170 16490 0 clknet_0_prog_clk
rlabel metal1 19366 9418 19366 9418 0 clknet_4_0_0_prog_clk
rlabel metal1 35098 12750 35098 12750 0 clknet_4_10_0_prog_clk
rlabel metal2 36478 13090 36478 13090 0 clknet_4_11_0_prog_clk
rlabel metal1 32338 17204 32338 17204 0 clknet_4_12_0_prog_clk
rlabel metal2 35650 19108 35650 19108 0 clknet_4_13_0_prog_clk
rlabel metal2 34914 14960 34914 14960 0 clknet_4_14_0_prog_clk
rlabel metal2 37766 19856 37766 19856 0 clknet_4_15_0_prog_clk
rlabel metal1 12374 11798 12374 11798 0 clknet_4_1_0_prog_clk
rlabel metal1 23322 2482 23322 2482 0 clknet_4_2_0_prog_clk
rlabel metal1 22034 13974 22034 13974 0 clknet_4_3_0_prog_clk
rlabel metal1 14720 17714 14720 17714 0 clknet_4_4_0_prog_clk
rlabel metal2 13846 19584 13846 19584 0 clknet_4_5_0_prog_clk
rlabel metal2 21114 15538 21114 15538 0 clknet_4_6_0_prog_clk
rlabel metal2 18814 23426 18814 23426 0 clknet_4_7_0_prog_clk
rlabel metal1 28842 8500 28842 8500 0 clknet_4_8_0_prog_clk
rlabel metal1 30360 12886 30360 12886 0 clknet_4_9_0_prog_clk
rlabel metal2 11730 1622 11730 1622 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 13846 1622 13846 1622 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 15962 1761 15962 1761 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 18078 823 18078 823 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 28796 2414 28796 2414 0 gfpga_pad_io_soc_in[0]
rlabel metal1 30912 2414 30912 2414 0 gfpga_pad_io_soc_in[1]
rlabel metal2 33166 1989 33166 1989 0 gfpga_pad_io_soc_in[2]
rlabel metal1 35144 2414 35144 2414 0 gfpga_pad_io_soc_in[3]
rlabel metal2 20194 2404 20194 2404 0 gfpga_pad_io_soc_out[0]
rlabel metal1 21896 2958 21896 2958 0 gfpga_pad_io_soc_out[1]
rlabel metal1 23736 3434 23736 3434 0 gfpga_pad_io_soc_out[2]
rlabel metal1 25576 2958 25576 2958 0 gfpga_pad_io_soc_out[3]
rlabel metal2 37122 1520 37122 1520 0 isol_n
rlabel metal1 10396 2618 10396 2618 0 net1
rlabel metal1 2990 8466 2990 8466 0 net10
rlabel metal2 17388 15062 17388 15062 0 net100
rlabel metal1 16330 17170 16330 17170 0 net101
rlabel metal1 35190 19686 35190 19686 0 net102
rlabel metal2 16974 18377 16974 18377 0 net103
rlabel metal1 18630 18734 18630 18734 0 net104
rlabel metal2 37214 21556 37214 21556 0 net105
rlabel metal1 40434 20332 40434 20332 0 net106
rlabel metal1 40710 2482 40710 2482 0 net107
rlabel metal1 7866 19958 7866 19958 0 net108
rlabel metal2 1794 13345 1794 13345 0 net109
rlabel metal2 2530 8857 2530 8857 0 net11
rlabel metal1 1794 18768 1794 18768 0 net110
rlabel metal1 1794 19380 1794 19380 0 net111
rlabel metal2 1794 19873 1794 19873 0 net112
rlabel metal1 1840 20434 1840 20434 0 net113
rlabel metal1 1794 20944 1794 20944 0 net114
rlabel metal2 3450 21318 3450 21318 0 net115
rlabel metal2 3634 20230 3634 20230 0 net116
rlabel metal2 1794 21794 1794 21794 0 net117
rlabel metal1 1840 22610 1840 22610 0 net118
rlabel metal1 2576 23086 2576 23086 0 net119
rlabel metal2 1794 8670 1794 8670 0 net12
rlabel metal1 1794 13940 1794 13940 0 net120
rlabel metal1 4094 21930 4094 21930 0 net121
rlabel metal1 4094 20876 4094 20876 0 net122
rlabel metal2 7682 21556 7682 21556 0 net123
rlabel metal1 6532 20910 6532 20910 0 net124
rlabel metal1 5336 16422 5336 16422 0 net125
rlabel metal1 4186 18734 4186 18734 0 net126
rlabel metal1 6118 18938 6118 18938 0 net127
rlabel metal2 4002 16320 4002 16320 0 net128
rlabel metal1 5566 20536 5566 20536 0 net129
rlabel via2 1886 9469 1886 9469 0 net13
rlabel metal1 5566 23596 5566 23596 0 net130
rlabel metal1 5796 14382 5796 14382 0 net131
rlabel metal2 6670 15164 6670 15164 0 net132
rlabel metal2 9706 15028 9706 15028 0 net133
rlabel metal2 5474 15300 5474 15300 0 net134
rlabel metal2 4094 16354 4094 16354 0 net135
rlabel metal1 1794 17204 1794 17204 0 net136
rlabel metal1 1794 17612 1794 17612 0 net137
rlabel metal2 1794 18020 1794 18020 0 net138
rlabel metal1 37950 3706 37950 3706 0 net139
rlabel metal1 4715 2550 4715 2550 0 net14
rlabel metal1 47518 4590 47518 4590 0 net140
rlabel metal1 47610 5202 47610 5202 0 net141
rlabel metal2 40618 7276 40618 7276 0 net142
rlabel metal1 47794 5678 47794 5678 0 net143
rlabel metal2 42734 7582 42734 7582 0 net144
rlabel metal1 47840 6766 47840 6766 0 net145
rlabel metal2 45862 9282 45862 9282 0 net146
rlabel metal2 46966 8772 46966 8772 0 net147
rlabel metal2 47058 9214 47058 9214 0 net148
rlabel metal2 46782 9214 46782 9214 0 net149
rlabel metal2 1886 10438 1886 10438 0 net15
rlabel metal2 39422 3740 39422 3740 0 net150
rlabel metal2 44206 10540 44206 10540 0 net151
rlabel metal2 47150 10132 47150 10132 0 net152
rlabel metal2 47242 10846 47242 10846 0 net153
rlabel metal2 46690 10812 46690 10812 0 net154
rlabel metal1 47472 10642 47472 10642 0 net155
rlabel metal1 47978 11186 47978 11186 0 net156
rlabel metal1 46966 11730 46966 11730 0 net157
rlabel metal1 47012 12614 47012 12614 0 net158
rlabel metal1 47932 12818 47932 12818 0 net159
rlabel metal2 2530 10489 2530 10489 0 net16
rlabel metal1 47288 13294 47288 13294 0 net160
rlabel metal2 44482 3434 44482 3434 0 net161
rlabel metal2 45862 4318 45862 4318 0 net162
rlabel metal2 40066 4284 40066 4284 0 net163
rlabel metal2 47242 3604 47242 3604 0 net164
rlabel metal2 47334 4454 47334 4454 0 net165
rlabel metal2 46966 4828 46966 4828 0 net166
rlabel metal1 42090 7208 42090 7208 0 net167
rlabel metal1 47564 4114 47564 4114 0 net168
rlabel metal1 6348 22406 6348 22406 0 net169
rlabel metal1 4347 10506 4347 10506 0 net17
rlabel metal2 7406 24225 7406 24225 0 net170
rlabel metal2 4002 23902 4002 23902 0 net171
rlabel metal1 9131 19482 9131 19482 0 net172
rlabel metal1 10028 23698 10028 23698 0 net173
rlabel metal1 10718 23052 10718 23052 0 net174
rlabel metal2 11822 21828 11822 21828 0 net175
rlabel metal1 10396 24174 10396 24174 0 net176
rlabel metal2 12466 23562 12466 23562 0 net177
rlabel metal1 9798 22542 9798 22542 0 net178
rlabel metal2 5290 23664 5290 23664 0 net179
rlabel metal2 1794 11169 1794 11169 0 net18
rlabel metal1 5290 17306 5290 17306 0 net180
rlabel metal1 19090 21046 19090 21046 0 net181
rlabel metal1 15134 22678 15134 22678 0 net182
rlabel metal1 19734 20026 19734 20026 0 net183
rlabel metal1 14950 23732 14950 23732 0 net184
rlabel metal1 16192 23018 16192 23018 0 net185
rlabel metal1 15134 24140 15134 24140 0 net186
rlabel metal2 19734 23562 19734 23562 0 net187
rlabel metal1 17756 24174 17756 24174 0 net188
rlabel metal1 22402 24174 22402 24174 0 net189
rlabel metal1 3358 11866 3358 11866 0 net19
rlabel metal1 20102 24106 20102 24106 0 net190
rlabel metal1 2300 24174 2300 24174 0 net191
rlabel metal1 3174 23698 3174 23698 0 net192
rlabel metal1 4370 22610 4370 22610 0 net193
rlabel metal2 4830 20502 4830 20502 0 net194
rlabel metal1 4922 23086 4922 23086 0 net195
rlabel metal1 4876 24174 4876 24174 0 net196
rlabel metal1 7222 22610 7222 22610 0 net197
rlabel metal1 7176 23086 7176 23086 0 net198
rlabel metal1 12282 2414 12282 2414 0 net199
rlabel metal1 46184 21862 46184 21862 0 net2
rlabel metal1 3588 12274 3588 12274 0 net20
rlabel metal1 14950 2414 14950 2414 0 net200
rlabel metal1 17066 2958 17066 2958 0 net201
rlabel metal1 17710 2346 17710 2346 0 net202
rlabel via2 17710 16099 17710 16099 0 net203
rlabel metal1 22816 14994 22816 14994 0 net204
rlabel metal1 29808 23018 29808 23018 0 net205
rlabel metal1 13938 13226 13938 13226 0 net206
rlabel metal1 23966 18326 23966 18326 0 net207
rlabel metal1 19780 13294 19780 13294 0 net208
rlabel metal1 31234 14382 31234 14382 0 net209
rlabel metal1 4347 11594 4347 11594 0 net21
rlabel metal2 31418 7990 31418 7990 0 net210
rlabel metal1 30544 10098 30544 10098 0 net211
rlabel metal1 34224 15130 34224 15130 0 net212
rlabel metal1 31004 14042 31004 14042 0 net213
rlabel metal2 29670 9078 29670 9078 0 net214
rlabel metal1 32384 7786 32384 7786 0 net215
rlabel metal2 37582 12580 37582 12580 0 net216
rlabel metal2 29026 8398 29026 8398 0 net217
rlabel metal1 26910 11866 26910 11866 0 net218
rlabel metal2 33350 9486 33350 9486 0 net219
rlabel metal2 5658 15062 5658 15062 0 net22
rlabel metal2 32062 20468 32062 20468 0 net220
rlabel metal1 31004 17170 31004 17170 0 net221
rlabel metal1 37168 17170 37168 17170 0 net222
rlabel metal1 34914 15130 34914 15130 0 net223
rlabel metal1 37812 14042 37812 14042 0 net224
rlabel metal1 29946 9010 29946 9010 0 net225
rlabel metal1 42412 22066 42412 22066 0 net226
rlabel metal2 25254 13634 25254 13634 0 net227
rlabel metal1 24012 11118 24012 11118 0 net228
rlabel metal1 22540 11186 22540 11186 0 net229
rlabel metal2 14490 18139 14490 18139 0 net23
rlabel metal1 24656 9010 24656 9010 0 net230
rlabel metal1 21022 10778 21022 10778 0 net231
rlabel metal2 12190 11424 12190 11424 0 net232
rlabel metal1 16376 9622 16376 9622 0 net233
rlabel metal1 19596 10098 19596 10098 0 net234
rlabel metal1 26450 9044 26450 9044 0 net235
rlabel metal1 33718 16558 33718 16558 0 net236
rlabel metal1 13064 11186 13064 11186 0 net237
rlabel metal2 15226 18496 15226 18496 0 net238
rlabel metal1 6118 18326 6118 18326 0 net239
rlabel metal2 20378 21029 20378 21029 0 net24
rlabel metal1 9016 17578 9016 17578 0 net240
rlabel metal1 6578 24310 6578 24310 0 net241
rlabel metal2 15134 21869 15134 21869 0 net242
rlabel metal2 16790 19533 16790 19533 0 net243
rlabel metal2 39238 17935 39238 17935 0 net244
rlabel metal1 40434 20468 40434 20468 0 net245
rlabel metal1 18906 8602 18906 8602 0 net246
rlabel metal1 17526 8398 17526 8398 0 net247
rlabel metal2 12098 13056 12098 13056 0 net248
rlabel metal1 16698 13226 16698 13226 0 net249
rlabel metal1 1794 2312 1794 2312 0 net25
rlabel metal2 21298 12444 21298 12444 0 net250
rlabel metal1 21574 11866 21574 11866 0 net251
rlabel via2 19642 18717 19642 18717 0 net252
rlabel via2 17986 20859 17986 20859 0 net253
rlabel metal1 25024 17578 25024 17578 0 net254
rlabel metal1 18722 17850 18722 17850 0 net255
rlabel metal2 40986 19533 40986 19533 0 net256
rlabel metal1 16928 7514 16928 7514 0 net257
rlabel metal1 15962 22576 15962 22576 0 net258
rlabel via2 38502 18819 38502 18819 0 net259
rlabel metal1 6532 2890 6532 2890 0 net26
rlabel metal1 17986 19278 17986 19278 0 net260
rlabel metal1 21804 6834 21804 6834 0 net261
rlabel metal1 14030 20366 14030 20366 0 net262
rlabel via2 40710 16507 40710 16507 0 net263
rlabel metal2 10810 19176 10810 19176 0 net264
rlabel metal2 22310 3876 22310 3876 0 net265
rlabel metal1 28980 2958 28980 2958 0 net266
rlabel metal1 19688 7514 19688 7514 0 net267
rlabel metal2 39330 13005 39330 13005 0 net268
rlabel metal1 28658 18938 28658 18938 0 net269
rlabel metal1 4738 3502 4738 3502 0 net27
rlabel metal1 26496 22542 26496 22542 0 net270
rlabel metal1 11316 14042 11316 14042 0 net271
rlabel metal1 18574 13702 18574 13702 0 net272
rlabel metal2 25530 9044 25530 9044 0 net273
rlabel metal1 16514 16762 16514 16762 0 net274
rlabel metal2 25990 23596 25990 23596 0 net275
rlabel metal1 25300 2822 25300 2822 0 net276
rlabel metal2 16330 19618 16330 19618 0 net277
rlabel metal1 18170 6834 18170 6834 0 net278
rlabel metal1 27600 12886 27600 12886 0 net279
rlabel metal1 4715 3978 4715 3978 0 net28
rlabel metal1 11720 20026 11720 20026 0 net280
rlabel metal1 18262 21454 18262 21454 0 net281
rlabel metal2 36018 11288 36018 11288 0 net282
rlabel metal1 16882 14042 16882 14042 0 net283
rlabel metal1 13662 20570 13662 20570 0 net284
rlabel metal1 37766 12920 37766 12920 0 net285
rlabel metal1 34086 10744 34086 10744 0 net286
rlabel metal2 25254 8228 25254 8228 0 net287
rlabel metal1 25438 9146 25438 9146 0 net288
rlabel metal2 11362 18496 11362 18496 0 net289
rlabel metal1 3680 3910 3680 3910 0 net29
rlabel metal1 25753 10234 25753 10234 0 net290
rlabel metal1 27416 13158 27416 13158 0 net291
rlabel metal1 14168 18666 14168 18666 0 net292
rlabel metal2 21482 7956 21482 7956 0 net293
rlabel metal1 23223 18938 23223 18938 0 net294
rlabel metal1 17342 8058 17342 8058 0 net295
rlabel metal2 31694 23596 31694 23596 0 net296
rlabel metal1 32844 20978 32844 20978 0 net297
rlabel metal1 12604 10234 12604 10234 0 net298
rlabel metal1 32936 7514 32936 7514 0 net299
rlabel metal2 9522 2448 9522 2448 0 net3
rlabel metal1 1794 4488 1794 4488 0 net30
rlabel metal1 14076 20842 14076 20842 0 net300
rlabel metal1 19780 6426 19780 6426 0 net301
rlabel metal2 38962 11917 38962 11917 0 net302
rlabel metal1 25944 13498 25944 13498 0 net303
rlabel metal1 13156 18190 13156 18190 0 net304
rlabel metal2 15502 20162 15502 20162 0 net305
rlabel metal2 40158 15419 40158 15419 0 net306
rlabel metal2 30682 8976 30682 8976 0 net307
rlabel via2 38778 13243 38778 13243 0 net308
rlabel metal2 43378 17578 43378 17578 0 net309
rlabel metal1 6348 5134 6348 5134 0 net31
rlabel metal2 39698 16133 39698 16133 0 net310
rlabel metal1 21666 7752 21666 7752 0 net311
rlabel metal1 30268 7446 30268 7446 0 net312
rlabel metal2 35282 23664 35282 23664 0 net313
rlabel metal2 40066 15130 40066 15130 0 net314
rlabel via2 11178 21437 11178 21437 0 net315
rlabel metal1 13294 21658 13294 21658 0 net316
rlabel metal1 26404 18802 26404 18802 0 net317
rlabel metal1 38778 14280 38778 14280 0 net318
rlabel metal1 17204 16150 17204 16150 0 net319
rlabel metal1 2530 5576 2530 5576 0 net32
rlabel metal1 40158 17000 40158 17000 0 net320
rlabel metal1 14766 15674 14766 15674 0 net321
rlabel metal1 16514 23188 16514 23188 0 net322
rlabel metal1 22494 7514 22494 7514 0 net323
rlabel metal2 42366 18326 42366 18326 0 net324
rlabel metal2 42366 15708 42366 15708 0 net325
rlabel metal2 30406 22372 30406 22372 0 net326
rlabel metal1 33948 22678 33948 22678 0 net327
rlabel metal1 20378 6834 20378 6834 0 net328
rlabel metal1 30544 6834 30544 6834 0 net329
rlabel metal2 48438 14552 48438 14552 0 net33
rlabel metal1 29992 15538 29992 15538 0 net330
rlabel metal1 38134 11254 38134 11254 0 net331
rlabel metal1 22494 22678 22494 22678 0 net332
rlabel metal1 11638 11526 11638 11526 0 net333
rlabel metal3 28106 12852 28106 12852 0 net334
rlabel metal1 38042 20536 38042 20536 0 net335
rlabel metal1 20838 16490 20838 16490 0 net336
rlabel metal2 21666 22984 21666 22984 0 net337
rlabel metal1 28014 8602 28014 8602 0 net338
rlabel metal1 38081 22202 38081 22202 0 net339
rlabel metal1 19826 11696 19826 11696 0 net34
rlabel metal2 36754 13668 36754 13668 0 net340
rlabel metal2 24242 13566 24242 13566 0 net341
rlabel metal1 28835 17850 28835 17850 0 net342
rlabel metal1 28658 14926 28658 14926 0 net343
rlabel metal1 33994 8398 33994 8398 0 net344
rlabel metal1 14674 8602 14674 8602 0 net345
rlabel metal1 11362 11186 11362 11186 0 net346
rlabel metal1 36478 10098 36478 10098 0 net347
rlabel metal1 25162 23800 25162 23800 0 net348
rlabel metal1 32568 12886 32568 12886 0 net349
rlabel metal1 19642 19958 19642 19958 0 net35
rlabel metal1 24564 19278 24564 19278 0 net350
rlabel metal1 37766 22712 37766 22712 0 net351
rlabel metal1 37490 22984 37490 22984 0 net352
rlabel metal3 36478 12580 36478 12580 0 net353
rlabel metal2 32614 13617 32614 13617 0 net354
rlabel metal4 34500 18836 34500 18836 0 net355
rlabel metal2 42182 16048 42182 16048 0 net356
rlabel metal1 10166 16490 10166 16490 0 net357
rlabel metal2 30406 8228 30406 8228 0 net358
rlabel metal2 38318 18105 38318 18105 0 net359
rlabel metal2 48438 18462 48438 18462 0 net36
rlabel metal1 21850 20842 21850 20842 0 net360
rlabel metal1 39698 21012 39698 21012 0 net361
rlabel metal2 20654 23256 20654 23256 0 net362
rlabel metal2 17250 23596 17250 23596 0 net363
rlabel metal1 29072 13498 29072 13498 0 net364
rlabel via2 16146 20451 16146 20451 0 net37
rlabel metal1 16606 18258 16606 18258 0 net38
rlabel metal2 18722 17255 18722 17255 0 net39
rlabel metal2 12834 12517 12834 12517 0 net4
rlabel metal2 40526 19363 40526 19363 0 net40
rlabel metal2 16054 14416 16054 14416 0 net41
rlabel metal2 21482 20672 21482 20672 0 net42
rlabel metal3 45540 11832 45540 11832 0 net43
rlabel via2 14398 13243 14398 13243 0 net44
rlabel metal1 48622 19958 48622 19958 0 net45
rlabel metal2 15962 16031 15962 16031 0 net46
rlabel metal2 18538 18224 18538 18224 0 net47
rlabel metal2 15778 20689 15778 20689 0 net48
rlabel metal1 47702 21114 47702 21114 0 net49
rlabel metal1 5934 6154 5934 6154 0 net5
rlabel metal2 40526 21488 40526 21488 0 net50
rlabel metal2 12466 19601 12466 19601 0 net51
rlabel metal1 48392 21114 48392 21114 0 net52
rlabel metal1 39238 23630 39238 23630 0 net53
rlabel metal2 19090 23103 19090 23103 0 net54
rlabel metal1 18722 10030 18722 10030 0 net55
rlabel metal1 21574 15130 21574 15130 0 net56
rlabel metal1 49082 15674 49082 15674 0 net57
rlabel via2 20286 12597 20286 12597 0 net58
rlabel metal2 18860 12852 18860 12852 0 net59
rlabel metal1 2392 6630 2392 6630 0 net6
rlabel metal2 13570 17969 13570 17969 0 net60
rlabel metal2 48438 17442 48438 17442 0 net61
rlabel metal4 16468 16048 16468 16048 0 net62
rlabel via2 4186 22525 4186 22525 0 net63
rlabel metal3 35788 19992 35788 19992 0 net64
rlabel metal1 35236 20570 35236 20570 0 net65
rlabel metal2 38962 25466 38962 25466 0 net66
rlabel metal1 28658 23018 28658 23018 0 net67
rlabel metal1 37260 20434 37260 20434 0 net68
rlabel metal2 45218 20621 45218 20621 0 net69
rlabel metal1 39008 7854 39008 7854 0 net7
rlabel metal2 35282 19771 35282 19771 0 net70
rlabel metal2 34822 21335 34822 21335 0 net71
rlabel metal2 33626 21403 33626 21403 0 net72
rlabel metal2 35834 24820 35834 24820 0 net73
rlabel metal2 22034 17340 22034 17340 0 net74
rlabel metal1 26174 19686 26174 19686 0 net75
rlabel metal2 31786 17425 31786 17425 0 net76
rlabel metal3 36524 19448 36524 19448 0 net77
rlabel metal1 34638 19754 34638 19754 0 net78
rlabel metal1 28014 23154 28014 23154 0 net79
rlabel metal2 18814 14365 18814 14365 0 net8
rlabel metal1 44666 21114 44666 21114 0 net80
rlabel metal1 42550 19992 42550 19992 0 net81
rlabel metal1 35512 20434 35512 20434 0 net82
rlabel metal2 45770 21097 45770 21097 0 net83
rlabel via2 33718 21437 33718 21437 0 net84
rlabel via2 9430 23171 9430 23171 0 net85
rlabel metal1 32752 16218 32752 16218 0 net86
rlabel metal2 12006 23613 12006 23613 0 net87
rlabel metal2 33258 17408 33258 17408 0 net88
rlabel via2 12098 23715 12098 23715 0 net89
rlabel metal1 1794 7752 1794 7752 0 net9
rlabel metal1 32982 18258 32982 18258 0 net90
rlabel metal1 27462 21862 27462 21862 0 net91
rlabel metal1 29210 17170 29210 17170 0 net92
rlabel metal2 27462 2448 27462 2448 0 net93
rlabel metal1 30774 2278 30774 2278 0 net94
rlabel metal1 32338 2618 32338 2618 0 net95
rlabel metal1 34362 2618 34362 2618 0 net96
rlabel metal1 23782 2414 23782 2414 0 net97
rlabel metal1 25109 2346 25109 2346 0 net98
rlabel via2 35374 19669 35374 19669 0 net99
rlabel metal2 34270 4879 34270 4879 0 prog_clk
rlabel metal1 44068 24106 44068 24106 0 prog_reset
rlabel metal2 43470 2098 43470 2098 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 45586 2200 45586 2200 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 47702 2166 47702 2166 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 49818 2064 49818 2064 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 29026 11254 29026 11254 0 sb_1__0_.mem_left_track_1.ccff_head
rlabel metal1 25162 17748 25162 17748 0 sb_1__0_.mem_left_track_1.ccff_tail
rlabel metal1 29578 20774 29578 20774 0 sb_1__0_.mem_left_track_1.mem_out\[0\]
rlabel metal2 19366 16218 19366 16218 0 sb_1__0_.mem_left_track_1.mem_out\[1\]
rlabel metal1 21252 14042 21252 14042 0 sb_1__0_.mem_left_track_11.ccff_head
rlabel metal1 20286 16966 20286 16966 0 sb_1__0_.mem_left_track_11.ccff_tail
rlabel metal2 21390 12512 21390 12512 0 sb_1__0_.mem_left_track_11.mem_out\[0\]
rlabel metal2 20102 16014 20102 16014 0 sb_1__0_.mem_left_track_11.mem_out\[1\]
rlabel metal1 17526 20944 17526 20944 0 sb_1__0_.mem_left_track_13.ccff_tail
rlabel metal1 21574 18054 21574 18054 0 sb_1__0_.mem_left_track_13.mem_out\[0\]
rlabel metal1 21344 21114 21344 21114 0 sb_1__0_.mem_left_track_13.mem_out\[1\]
rlabel metal1 17296 21590 17296 21590 0 sb_1__0_.mem_left_track_21.ccff_tail
rlabel metal1 21988 22542 21988 22542 0 sb_1__0_.mem_left_track_21.mem_out\[0\]
rlabel metal2 6854 23494 6854 23494 0 sb_1__0_.mem_left_track_21.mem_out\[1\]
rlabel metal1 25346 19210 25346 19210 0 sb_1__0_.mem_left_track_29.ccff_tail
rlabel metal2 24150 17612 24150 17612 0 sb_1__0_.mem_left_track_29.mem_out\[0\]
rlabel metal1 25990 17714 25990 17714 0 sb_1__0_.mem_left_track_29.mem_out\[1\]
rlabel metal1 17204 19278 17204 19278 0 sb_1__0_.mem_left_track_3.ccff_tail
rlabel metal1 27646 22066 27646 22066 0 sb_1__0_.mem_left_track_3.mem_out\[0\]
rlabel metal1 21160 19278 21160 19278 0 sb_1__0_.mem_left_track_3.mem_out\[1\]
rlabel metal1 26266 16422 26266 16422 0 sb_1__0_.mem_left_track_37.ccff_tail
rlabel metal1 32338 19244 32338 19244 0 sb_1__0_.mem_left_track_37.mem_out\[0\]
rlabel metal1 25852 16490 25852 16490 0 sb_1__0_.mem_left_track_37.mem_out\[1\]
rlabel metal1 27094 23494 27094 23494 0 sb_1__0_.mem_left_track_45.ccff_tail
rlabel metal1 32338 22508 32338 22508 0 sb_1__0_.mem_left_track_45.mem_out\[0\]
rlabel metal2 29946 22270 29946 22270 0 sb_1__0_.mem_left_track_45.mem_out\[1\]
rlabel metal1 17158 17306 17158 17306 0 sb_1__0_.mem_left_track_5.ccff_tail
rlabel metal1 20332 20230 20332 20230 0 sb_1__0_.mem_left_track_5.mem_out\[0\]
rlabel metal1 18400 15538 18400 15538 0 sb_1__0_.mem_left_track_5.mem_out\[1\]
rlabel metal2 27462 22848 27462 22848 0 sb_1__0_.mem_left_track_53.mem_out\[0\]
rlabel metal1 26542 22100 26542 22100 0 sb_1__0_.mem_left_track_53.mem_out\[1\]
rlabel metal1 21850 15912 21850 15912 0 sb_1__0_.mem_left_track_7.mem_out\[0\]
rlabel metal1 19964 13362 19964 13362 0 sb_1__0_.mem_left_track_7.mem_out\[1\]
rlabel metal1 17434 21862 17434 21862 0 sb_1__0_.mem_right_track_0.ccff_head
rlabel metal2 34178 16252 34178 16252 0 sb_1__0_.mem_right_track_0.ccff_tail
rlabel metal1 36294 13804 36294 13804 0 sb_1__0_.mem_right_track_0.mem_out\[0\]
rlabel metal1 30268 16218 30268 16218 0 sb_1__0_.mem_right_track_0.mem_out\[1\]
rlabel metal1 38134 11730 38134 11730 0 sb_1__0_.mem_right_track_10.ccff_head
rlabel metal1 37674 10574 37674 10574 0 sb_1__0_.mem_right_track_10.ccff_tail
rlabel metal1 33810 9520 33810 9520 0 sb_1__0_.mem_right_track_10.mem_out\[0\]
rlabel metal1 35098 13770 35098 13770 0 sb_1__0_.mem_right_track_10.mem_out\[1\]
rlabel metal1 38778 13328 38778 13328 0 sb_1__0_.mem_right_track_12.ccff_tail
rlabel metal1 32798 19890 32798 19890 0 sb_1__0_.mem_right_track_12.mem_out\[0\]
rlabel metal2 39054 12988 39054 12988 0 sb_1__0_.mem_right_track_12.mem_out\[1\]
rlabel metal1 36662 15368 36662 15368 0 sb_1__0_.mem_right_track_2.ccff_tail
rlabel metal2 32890 18020 32890 18020 0 sb_1__0_.mem_right_track_2.mem_out\[0\]
rlabel metal1 34546 17034 34546 17034 0 sb_1__0_.mem_right_track_2.mem_out\[1\]
rlabel metal1 34362 11662 34362 11662 0 sb_1__0_.mem_right_track_20.ccff_tail
rlabel metal2 32338 13056 32338 13056 0 sb_1__0_.mem_right_track_20.mem_out\[0\]
rlabel metal2 22034 15844 22034 15844 0 sb_1__0_.mem_right_track_20.mem_out\[1\]
rlabel metal2 32246 8670 32246 8670 0 sb_1__0_.mem_right_track_28.ccff_tail
rlabel metal1 30866 14994 30866 14994 0 sb_1__0_.mem_right_track_28.mem_out\[0\]
rlabel metal1 30268 13362 30268 13362 0 sb_1__0_.mem_right_track_28.mem_out\[1\]
rlabel metal2 34086 7854 34086 7854 0 sb_1__0_.mem_right_track_36.ccff_tail
rlabel metal1 32890 14450 32890 14450 0 sb_1__0_.mem_right_track_36.mem_out\[0\]
rlabel metal2 32936 12886 32936 12886 0 sb_1__0_.mem_right_track_36.mem_out\[1\]
rlabel metal1 39330 13804 39330 13804 0 sb_1__0_.mem_right_track_4.ccff_tail
rlabel metal1 35190 21454 35190 21454 0 sb_1__0_.mem_right_track_4.mem_out\[0\]
rlabel metal1 36616 14518 36616 14518 0 sb_1__0_.mem_right_track_4.mem_out\[1\]
rlabel metal1 32890 10540 32890 10540 0 sb_1__0_.mem_right_track_44.ccff_tail
rlabel metal1 30130 16626 30130 16626 0 sb_1__0_.mem_right_track_44.mem_out\[0\]
rlabel metal1 29486 17102 29486 17102 0 sb_1__0_.mem_right_track_52.mem_out\[0\]
rlabel metal1 33580 17714 33580 17714 0 sb_1__0_.mem_right_track_6.mem_out\[0\]
rlabel metal1 36616 14926 36616 14926 0 sb_1__0_.mem_right_track_6.mem_out\[1\]
rlabel metal1 30590 24174 30590 24174 0 sb_1__0_.mem_top_track_0.ccff_tail
rlabel metal1 39468 21998 39468 21998 0 sb_1__0_.mem_top_track_0.mem_out\[0\]
rlabel metal2 32614 22525 32614 22525 0 sb_1__0_.mem_top_track_0.mem_out\[1\]
rlabel metal1 39330 21114 39330 21114 0 sb_1__0_.mem_top_track_10.ccff_head
rlabel metal1 36294 18054 36294 18054 0 sb_1__0_.mem_top_track_10.ccff_tail
rlabel metal1 40802 19244 40802 19244 0 sb_1__0_.mem_top_track_10.mem_out\[0\]
rlabel metal2 33902 17578 33902 17578 0 sb_1__0_.mem_top_track_10.mem_out\[1\]
rlabel metal1 39238 18394 39238 18394 0 sb_1__0_.mem_top_track_12.ccff_tail
rlabel metal1 40388 19890 40388 19890 0 sb_1__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 39238 19142 39238 19142 0 sb_1__0_.mem_top_track_12.mem_out\[1\]
rlabel metal1 38272 16762 38272 16762 0 sb_1__0_.mem_top_track_14.ccff_tail
rlabel metal2 41078 19652 41078 19652 0 sb_1__0_.mem_top_track_14.mem_out\[0\]
rlabel metal2 40618 16796 40618 16796 0 sb_1__0_.mem_top_track_14.mem_out\[1\]
rlabel metal2 39514 15793 39514 15793 0 sb_1__0_.mem_top_track_16.ccff_tail
rlabel metal1 39790 15878 39790 15878 0 sb_1__0_.mem_top_track_16.mem_out\[0\]
rlabel metal2 41078 14858 41078 14858 0 sb_1__0_.mem_top_track_16.mem_out\[1\]
rlabel metal1 34316 13838 34316 13838 0 sb_1__0_.mem_top_track_18.ccff_tail
rlabel metal1 38778 14790 38778 14790 0 sb_1__0_.mem_top_track_18.mem_out\[0\]
rlabel metal1 38916 14246 38916 14246 0 sb_1__0_.mem_top_track_18.mem_out\[1\]
rlabel metal1 35420 23834 35420 23834 0 sb_1__0_.mem_top_track_2.ccff_tail
rlabel metal1 35696 24242 35696 24242 0 sb_1__0_.mem_top_track_2.mem_out\[0\]
rlabel metal1 35512 22474 35512 22474 0 sb_1__0_.mem_top_track_2.mem_out\[1\]
rlabel metal1 25806 13294 25806 13294 0 sb_1__0_.mem_top_track_20.ccff_tail
rlabel metal1 28382 13328 28382 13328 0 sb_1__0_.mem_top_track_20.mem_out\[0\]
rlabel metal1 24748 12954 24748 12954 0 sb_1__0_.mem_top_track_22.ccff_tail
rlabel metal1 24334 14382 24334 14382 0 sb_1__0_.mem_top_track_22.mem_out\[0\]
rlabel metal1 25668 11866 25668 11866 0 sb_1__0_.mem_top_track_24.ccff_tail
rlabel metal1 27554 15946 27554 15946 0 sb_1__0_.mem_top_track_24.mem_out\[0\]
rlabel metal1 22586 13328 22586 13328 0 sb_1__0_.mem_top_track_26.ccff_tail
rlabel metal1 27324 15538 27324 15538 0 sb_1__0_.mem_top_track_26.mem_out\[0\]
rlabel metal1 21390 10540 21390 10540 0 sb_1__0_.mem_top_track_28.ccff_tail
rlabel metal1 23828 9010 23828 9010 0 sb_1__0_.mem_top_track_28.mem_out\[0\]
rlabel metal1 21252 8602 21252 8602 0 sb_1__0_.mem_top_track_30.ccff_tail
rlabel metal2 20838 7718 20838 7718 0 sb_1__0_.mem_top_track_30.mem_out\[0\]
rlabel metal1 18860 9146 18860 9146 0 sb_1__0_.mem_top_track_32.ccff_tail
rlabel metal1 18676 6766 18676 6766 0 sb_1__0_.mem_top_track_32.mem_out\[0\]
rlabel metal1 20286 12750 20286 12750 0 sb_1__0_.mem_top_track_34.ccff_tail
rlabel metal1 21160 9350 21160 9350 0 sb_1__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 20562 7310 20562 7310 0 sb_1__0_.mem_top_track_36.ccff_tail
rlabel metal1 23092 9486 23092 9486 0 sb_1__0_.mem_top_track_36.mem_out\[0\]
rlabel metal1 34040 20570 34040 20570 0 sb_1__0_.mem_top_track_4.ccff_tail
rlabel metal1 35972 20978 35972 20978 0 sb_1__0_.mem_top_track_4.mem_out\[0\]
rlabel metal1 36524 21454 36524 21454 0 sb_1__0_.mem_top_track_4.mem_out\[1\]
rlabel metal1 12558 13770 12558 13770 0 sb_1__0_.mem_top_track_40.ccff_tail
rlabel metal1 10534 11662 10534 11662 0 sb_1__0_.mem_top_track_40.mem_out\[0\]
rlabel metal1 15410 18224 15410 18224 0 sb_1__0_.mem_top_track_42.ccff_tail
rlabel metal1 16100 14858 16100 14858 0 sb_1__0_.mem_top_track_42.mem_out\[0\]
rlabel metal1 13294 19278 13294 19278 0 sb_1__0_.mem_top_track_44.ccff_tail
rlabel metal1 15318 18938 15318 18938 0 sb_1__0_.mem_top_track_44.mem_out\[0\]
rlabel metal2 10534 19074 10534 19074 0 sb_1__0_.mem_top_track_46.ccff_tail
rlabel metal2 11730 18666 11730 18666 0 sb_1__0_.mem_top_track_46.mem_out\[0\]
rlabel metal1 13938 20978 13938 20978 0 sb_1__0_.mem_top_track_48.ccff_tail
rlabel metal1 13708 19686 13708 19686 0 sb_1__0_.mem_top_track_48.mem_out\[0\]
rlabel metal2 15318 21284 15318 21284 0 sb_1__0_.mem_top_track_50.ccff_tail
rlabel metal1 16790 18870 16790 18870 0 sb_1__0_.mem_top_track_50.mem_out\[0\]
rlabel metal2 18630 22984 18630 22984 0 sb_1__0_.mem_top_track_58.mem_out\[0\]
rlabel metal1 38870 23290 38870 23290 0 sb_1__0_.mem_top_track_6.ccff_tail
rlabel metal1 34224 20774 34224 20774 0 sb_1__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 37996 22542 37996 22542 0 sb_1__0_.mem_top_track_6.mem_out\[1\]
rlabel metal1 38226 21454 38226 21454 0 sb_1__0_.mem_top_track_8.mem_out\[0\]
rlabel metal1 39054 21318 39054 21318 0 sb_1__0_.mem_top_track_8.mem_out\[1\]
rlabel metal2 2162 24174 2162 24174 0 sb_1__0_.mux_left_track_1.out
rlabel metal1 26358 18156 26358 18156 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 26772 18394 26772 18394 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23184 12954 23184 12954 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23598 16150 23598 16150 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 25070 17884 25070 17884 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24104 16218 24104 16218 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 21206 18258 21206 18258 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7406 16218 7406 16218 0 sb_1__0_.mux_left_track_11.out
rlabel metal1 25852 19754 25852 19754 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24748 19482 24748 19482 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20378 13498 20378 13498 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20240 14994 20240 14994 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20332 16490 20332 16490 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 19688 15130 19688 15130 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal3 15916 16456 15916 16456 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7912 19346 7912 19346 0 sb_1__0_.mux_left_track_13.out
rlabel via2 27186 21675 27186 21675 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24794 21216 24794 21216 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21022 15674 21022 15674 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17434 21012 17434 21012 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18584 18938 18584 18938 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 7774 20468 7774 20468 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 5198 19822 5198 19822 0 sb_1__0_.mux_left_track_21.out
rlabel metal1 23046 23222 23046 23222 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24196 22202 24196 22202 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21896 19482 21896 19482 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18998 21658 18998 21658 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17710 21114 17710 21114 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 16882 21165 16882 21165 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 14858 14722 14858 14722 0 sb_1__0_.mux_left_track_29.out
rlabel metal2 26174 21080 26174 21080 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 26818 20434 26818 20434 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 25116 15130 25116 15130 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22770 20706 22770 20706 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 25254 17850 25254 17850 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 18354 19737 18354 19737 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9016 24038 9016 24038 0 sb_1__0_.mux_left_track_3.out
rlabel metal1 21252 19482 21252 19482 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24334 18938 24334 18938 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19044 19482 19044 19482 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17572 16218 17572 16218 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 9706 23868 9706 23868 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 15962 14059 15962 14059 0 sb_1__0_.mux_left_track_37.out
rlabel metal2 31786 18581 31786 18581 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 28750 18224 28750 18224 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23782 16660 23782 16660 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23230 15130 23230 15130 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19550 14535 19550 14535 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 8418 18003 8418 18003 0 sb_1__0_.mux_left_track_45.out
rlabel metal1 32062 22746 32062 22746 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27508 20842 27508 20842 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 27922 20910 27922 20910 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 8602 17697 8602 17697 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 6348 16966 6348 16966 0 sb_1__0_.mux_left_track_5.out
rlabel metal1 21827 18734 21827 18734 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21482 18496 21482 18496 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17894 18530 17894 18530 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18308 15674 18308 15674 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8694 17136 8694 17136 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 6762 15402 6762 15402 0 sb_1__0_.mux_left_track_53.out
rlabel metal1 29854 22202 29854 22202 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 25990 21896 25990 21896 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20746 21250 20746 21250 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20010 21505 20010 21505 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 14352 16082 14352 16082 0 sb_1__0_.mux_left_track_7.out
rlabel metal1 23690 15470 23690 15470 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23690 15402 23690 15402 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19550 13226 19550 13226 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23046 15368 23046 15368 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19734 13498 19734 13498 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 18630 15810 18630 15810 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 39330 14110 39330 14110 0 sb_1__0_.mux_right_track_0.out
rlabel metal1 30728 19822 30728 19822 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 35742 14824 35742 14824 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 30544 14314 30544 14314 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 33994 17000 33994 17000 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 33902 15334 33902 15334 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 39514 14433 39514 14433 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 41538 11220 41538 11220 0 sb_1__0_.mux_right_track_10.out
rlabel metal1 34960 13974 34960 13974 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34868 14042 34868 14042 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35098 9010 35098 9010 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33534 8840 33534 8840 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 35374 14042 35374 14042 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 35696 9146 35696 9146 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 38088 10506 38088 10506 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 40802 11934 40802 11934 0 sb_1__0_.mux_right_track_12.out
rlabel metal1 33718 14450 33718 14450 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33580 14382 33580 14382 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 29302 10778 29302 10778 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 35604 12886 35604 12886 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 30958 11271 30958 11271 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 37214 12614 37214 12614 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 45862 14348 45862 14348 0 sb_1__0_.mux_right_track_2.out
rlabel metal2 35190 20434 35190 20434 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33442 18054 33442 18054 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 30314 14586 30314 14586 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 38318 17714 38318 17714 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 34316 14790 34316 14790 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 40434 17578 40434 17578 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 43286 9962 43286 9962 0 sb_1__0_.mux_right_track_20.out
rlabel metal1 30866 16218 30866 16218 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 30958 17102 30958 17102 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 27186 11900 27186 11900 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33488 11662 33488 11662 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 30130 11832 30130 11832 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 39514 11220 39514 11220 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 39606 8670 39606 8670 0 sb_1__0_.mux_right_track_28.out
rlabel metal1 30130 13158 30130 13158 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 30130 14042 30130 14042 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 26634 9418 26634 9418 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32752 9554 32752 9554 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32361 9622 32361 9622 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 37858 8976 37858 8976 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 44850 8024 44850 8024 0 sb_1__0_.mux_right_track_36.out
rlabel metal2 33994 13532 33994 13532 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33396 13294 33396 13294 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34454 13158 34454 13158 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 35282 8262 35282 8262 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 39146 8500 39146 8500 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 41446 14144 41446 14144 0 sb_1__0_.mux_right_track_4.out
rlabel metal1 35972 17102 35972 17102 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36340 16762 36340 16762 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 37582 12291 37582 12291 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 38732 13838 38732 13838 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 37490 13838 37490 13838 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 39790 13872 39790 13872 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 42734 6358 42734 6358 0 sb_1__0_.mux_right_track_44.out
rlabel metal2 31464 13124 31464 13124 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 29072 9146 29072 9146 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37674 8432 37674 8432 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 40066 7378 40066 7378 0 sb_1__0_.mux_right_track_52.out
rlabel metal2 31280 11866 31280 11866 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 30774 11866 30774 11866 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel via1 31786 11509 31786 11509 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 43493 12342 43493 12342 0 sb_1__0_.mux_right_track_6.out
rlabel metal1 35972 14926 35972 14926 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 36294 16218 36294 16218 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34684 11254 34684 11254 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33764 9146 33764 9146 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 36662 14858 36662 14858 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 38272 11866 38272 11866 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 41630 11900 41630 11900 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 21942 22984 21942 22984 0 sb_1__0_.mux_top_track_0.out
rlabel metal1 35052 21862 35052 21862 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37582 23834 37582 23834 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28842 21012 28842 21012 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 28612 19482 28612 19482 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 36110 23494 36110 23494 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 29256 21114 29256 21114 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 29808 23290 29808 23290 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 14674 21403 14674 21403 0 sb_1__0_.mux_top_track_10.out
rlabel metal1 35742 19754 35742 19754 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38318 19482 38318 19482 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34270 18666 34270 18666 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 32062 17952 32062 17952 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 31947 18938 31947 18938 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 14214 21573 14214 21573 0 sb_1__0_.mux_top_track_12.out
rlabel metal1 40480 18394 40480 18394 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40434 18156 40434 18156 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37582 17306 37582 17306 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 37306 20179 37306 20179 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19412 18870 19412 18870 0 sb_1__0_.mux_top_track_14.out
rlabel metal1 40480 17714 40480 17714 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39560 17850 39560 17850 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34730 14926 34730 14926 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 38318 18734 38318 18734 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22770 20910 22770 20910 0 sb_1__0_.mux_top_track_16.out
rlabel metal1 39836 16218 39836 16218 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40204 15946 40204 15946 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37398 14042 37398 14042 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 34684 18394 34684 18394 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 20286 19346 20286 19346 0 sb_1__0_.mux_top_track_18.out
rlabel metal1 40020 14994 40020 14994 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34592 15062 34592 15062 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32522 11866 32522 11866 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 27554 17034 27554 17034 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 27692 16422 27692 16422 0 sb_1__0_.mux_top_track_2.out
rlabel metal1 36570 23766 36570 23766 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 40066 23392 40066 23392 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 33534 21046 33534 21046 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37076 23562 37076 23562 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32890 21862 32890 21862 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 28290 16558 28290 16558 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 4002 22661 4002 22661 0 sb_1__0_.mux_top_track_20.out
rlabel metal1 26358 17306 26358 17306 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24932 13498 24932 13498 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 24886 17782 24886 17782 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 9890 19839 9890 19839 0 sb_1__0_.mux_top_track_22.out
rlabel metal1 24748 13226 24748 13226 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 23276 12818 23276 12818 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14950 16796 14950 16796 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11776 24174 11776 24174 0 sb_1__0_.mux_top_track_24.out
rlabel metal1 24564 14450 24564 14450 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23690 12240 23690 12240 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22954 12410 22954 12410 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17710 17782 17710 17782 0 sb_1__0_.mux_top_track_26.out
rlabel metal1 22402 13430 22402 13430 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24242 10540 24242 10540 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21666 13498 21666 13498 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12190 16422 12190 16422 0 sb_1__0_.mux_top_track_28.out
rlabel metal1 22908 9146 22908 9146 0 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13110 16558 13110 16558 0 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12052 18122 12052 18122 0 sb_1__0_.mux_top_track_30.out
rlabel metal1 21252 9146 21252 9146 0 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 16974 11475 16974 11475 0 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10212 17850 10212 17850 0 sb_1__0_.mux_top_track_32.out
rlabel metal1 16514 10778 16514 10778 0 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14674 15980 14674 15980 0 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9292 17306 9292 17306 0 sb_1__0_.mux_top_track_34.out
rlabel metal1 19596 10778 19596 10778 0 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19182 13175 19182 13175 0 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5060 24106 5060 24106 0 sb_1__0_.mux_top_track_36.out
rlabel metal2 22678 13736 22678 13736 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21988 9554 21988 9554 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 20654 12699 20654 12699 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 29394 23970 29394 23970 0 sb_1__0_.mux_top_track_4.out
rlabel metal1 36156 20570 36156 20570 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 40066 21760 40066 21760 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 35742 21216 35742 21216 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 31050 18394 31050 18394 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 30682 21114 30682 21114 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 6578 17884 6578 17884 0 sb_1__0_.mux_top_track_40.out
rlabel metal1 12696 9146 12696 9146 0 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10764 13702 10764 13702 0 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6624 16558 6624 16558 0 sb_1__0_.mux_top_track_42.out
rlabel metal1 16836 15130 16836 15130 0 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13294 18360 13294 18360 0 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6440 17714 6440 17714 0 sb_1__0_.mux_top_track_44.out
rlabel metal2 15594 18224 15594 18224 0 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12466 19040 12466 19040 0 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4186 17102 4186 17102 0 sb_1__0_.mux_top_track_46.out
rlabel metal1 11086 15130 11086 15130 0 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8050 17204 8050 17204 0 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 5014 17340 5014 17340 0 sb_1__0_.mux_top_track_48.out
rlabel metal1 13616 20774 13616 20774 0 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10994 17510 10994 17510 0 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 3542 16966 3542 16966 0 sb_1__0_.mux_top_track_50.out
rlabel metal2 17710 19006 17710 19006 0 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 14766 21675 14766 21675 0 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6348 22610 6348 22610 0 sb_1__0_.mux_top_track_58.out
rlabel metal1 18308 24038 18308 24038 0 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15226 17119 15226 17119 0 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19918 22865 19918 22865 0 sb_1__0_.mux_top_track_6.out
rlabel metal1 40204 21658 40204 21658 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40664 22202 40664 22202 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34086 19482 34086 19482 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 39698 23562 39698 23562 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 35880 22746 35880 22746 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 38962 23783 38962 23783 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal3 38364 22984 38364 22984 0 sb_1__0_.mux_top_track_8.out
rlabel metal1 40250 20978 40250 20978 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40848 20842 40848 20842 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34960 18938 34960 18938 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 40204 21114 40204 21114 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 36156 21862 36156 21862 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 36110 23749 36110 23749 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 46736 20026 46736 20026 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
rlabel metal1 47610 19210 47610 19210 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
rlabel metal1 47426 23766 47426 23766 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
rlabel metal1 47564 22746 47564 22746 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
rlabel metal1 47978 19278 47978 19278 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
rlabel metal1 48346 22066 48346 22066 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
rlabel metal1 44206 23086 44206 23086 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
rlabel metal1 46690 20570 46690 20570 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
rlabel metal2 1150 2166 1150 2166 0 top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 3266 1095 3266 1095 0 top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 5382 2234 5382 2234 0 top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 7498 2336 7498 2336 0 top_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 27000
<< end >>
