magic
tech sky130A
magscale 1 2
timestamp 1656242709
<< obsli1 >>
rect 1104 2159 21896 20689
<< obsm1 >>
rect 14 1368 22056 20720
<< metal2 >>
rect 5722 22200 5778 23000
rect 17222 22200 17278 23000
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
<< obsm2 >>
rect 20 22144 5666 22200
rect 5834 22144 17166 22200
rect 17334 22144 22050 22200
rect 20 856 22050 22144
rect 20 734 2170 856
rect 2338 734 2538 856
rect 2706 734 2906 856
rect 3074 734 3274 856
rect 3442 734 3642 856
rect 3810 734 4010 856
rect 4178 734 4378 856
rect 4546 734 4746 856
rect 4914 734 5114 856
rect 5282 734 5482 856
rect 5650 734 5850 856
rect 6018 734 6218 856
rect 6386 734 6586 856
rect 6754 734 6954 856
rect 7122 734 7322 856
rect 7490 734 7690 856
rect 7858 734 8058 856
rect 8226 734 8426 856
rect 8594 734 8794 856
rect 8962 734 9162 856
rect 9330 734 9530 856
rect 9698 734 9898 856
rect 10066 734 10266 856
rect 10434 734 10634 856
rect 10802 734 11002 856
rect 11170 734 11370 856
rect 11538 734 11738 856
rect 11906 734 12106 856
rect 12274 734 12474 856
rect 12642 734 12842 856
rect 13010 734 13210 856
rect 13378 734 13578 856
rect 13746 734 13946 856
rect 14114 734 14314 856
rect 14482 734 14682 856
rect 14850 734 15050 856
rect 15218 734 15418 856
rect 15586 734 15786 856
rect 15954 734 16154 856
rect 16322 734 16522 856
rect 16690 734 16890 856
rect 17058 734 17258 856
rect 17426 734 17626 856
rect 17794 734 17994 856
rect 18162 734 18362 856
rect 18530 734 18730 856
rect 18898 734 19098 856
rect 19266 734 19466 856
rect 19634 734 19834 856
rect 20002 734 20202 856
rect 20370 734 20570 856
rect 20738 734 22050 856
<< metal3 >>
rect 0 21224 800 21344
rect 22200 21224 23000 21344
rect 0 20816 800 20936
rect 22200 20816 23000 20936
rect 0 20408 800 20528
rect 22200 20408 23000 20528
rect 0 20000 800 20120
rect 22200 20000 23000 20120
rect 0 19592 800 19712
rect 22200 19592 23000 19712
rect 0 19184 800 19304
rect 22200 19184 23000 19304
rect 0 18776 800 18896
rect 22200 18776 23000 18896
rect 0 18368 800 18488
rect 22200 18368 23000 18488
rect 0 17960 800 18080
rect 22200 17960 23000 18080
rect 0 17552 800 17672
rect 22200 17552 23000 17672
rect 0 17144 800 17264
rect 22200 17144 23000 17264
rect 0 16736 800 16856
rect 22200 16736 23000 16856
rect 0 16328 800 16448
rect 22200 16328 23000 16448
rect 0 15920 800 16040
rect 22200 15920 23000 16040
rect 0 15512 800 15632
rect 22200 15512 23000 15632
rect 0 15104 800 15224
rect 22200 15104 23000 15224
rect 0 14696 800 14816
rect 22200 14696 23000 14816
rect 0 14288 800 14408
rect 22200 14288 23000 14408
rect 0 13880 800 14000
rect 22200 13880 23000 14000
rect 0 13472 800 13592
rect 22200 13472 23000 13592
rect 0 13064 800 13184
rect 22200 13064 23000 13184
rect 0 12656 800 12776
rect 22200 12656 23000 12776
rect 0 12248 800 12368
rect 22200 12248 23000 12368
rect 0 11840 800 11960
rect 22200 11840 23000 11960
rect 0 11432 800 11552
rect 22200 11432 23000 11552
rect 0 11024 800 11144
rect 22200 11024 23000 11144
rect 0 10616 800 10736
rect 22200 10616 23000 10736
rect 0 10208 800 10328
rect 22200 10208 23000 10328
rect 0 9800 800 9920
rect 22200 9800 23000 9920
rect 0 9392 800 9512
rect 22200 9392 23000 9512
rect 0 8984 800 9104
rect 22200 8984 23000 9104
rect 0 8576 800 8696
rect 22200 8576 23000 8696
rect 0 8168 800 8288
rect 22200 8168 23000 8288
rect 0 7760 800 7880
rect 22200 7760 23000 7880
rect 0 7352 800 7472
rect 22200 7352 23000 7472
rect 0 6944 800 7064
rect 22200 6944 23000 7064
rect 0 6536 800 6656
rect 22200 6536 23000 6656
rect 0 6128 800 6248
rect 22200 6128 23000 6248
rect 0 5720 800 5840
rect 22200 5720 23000 5840
rect 0 5312 800 5432
rect 22200 5312 23000 5432
rect 0 4904 800 5024
rect 22200 4904 23000 5024
rect 0 4496 800 4616
rect 22200 4496 23000 4616
rect 0 4088 800 4208
rect 22200 4088 23000 4208
rect 0 3680 800 3800
rect 22200 3680 23000 3800
rect 0 3272 800 3392
rect 22200 3272 23000 3392
rect 0 2864 800 2984
rect 22200 2864 23000 2984
rect 0 2456 800 2576
rect 22200 2456 23000 2576
rect 0 2048 800 2168
rect 22200 2048 23000 2168
rect 0 1640 800 1760
rect 22200 1640 23000 1760
<< obsm3 >>
rect 880 21144 22120 21317
rect 800 21016 22202 21144
rect 880 20736 22120 21016
rect 800 20608 22202 20736
rect 880 20328 22120 20608
rect 800 20200 22202 20328
rect 880 19920 22120 20200
rect 800 19792 22202 19920
rect 880 19512 22120 19792
rect 800 19384 22202 19512
rect 880 19104 22120 19384
rect 800 18976 22202 19104
rect 880 18696 22120 18976
rect 800 18568 22202 18696
rect 880 18288 22120 18568
rect 800 18160 22202 18288
rect 880 17880 22120 18160
rect 800 17752 22202 17880
rect 880 17472 22120 17752
rect 800 17344 22202 17472
rect 880 17064 22120 17344
rect 800 16936 22202 17064
rect 880 16656 22120 16936
rect 800 16528 22202 16656
rect 880 16248 22120 16528
rect 800 16120 22202 16248
rect 880 15840 22120 16120
rect 800 15712 22202 15840
rect 880 15432 22120 15712
rect 800 15304 22202 15432
rect 880 15024 22120 15304
rect 800 14896 22202 15024
rect 880 14616 22120 14896
rect 800 14488 22202 14616
rect 880 14208 22120 14488
rect 800 14080 22202 14208
rect 880 13800 22120 14080
rect 800 13672 22202 13800
rect 880 13392 22120 13672
rect 800 13264 22202 13392
rect 880 12984 22120 13264
rect 800 12856 22202 12984
rect 880 12576 22120 12856
rect 800 12448 22202 12576
rect 880 12168 22120 12448
rect 800 12040 22202 12168
rect 880 11760 22120 12040
rect 800 11632 22202 11760
rect 880 11352 22120 11632
rect 800 11224 22202 11352
rect 880 10944 22120 11224
rect 800 10816 22202 10944
rect 880 10536 22120 10816
rect 800 10408 22202 10536
rect 880 10128 22120 10408
rect 800 10000 22202 10128
rect 880 9720 22120 10000
rect 800 9592 22202 9720
rect 880 9312 22120 9592
rect 800 9184 22202 9312
rect 880 8904 22120 9184
rect 800 8776 22202 8904
rect 880 8496 22120 8776
rect 800 8368 22202 8496
rect 880 8088 22120 8368
rect 800 7960 22202 8088
rect 880 7680 22120 7960
rect 800 7552 22202 7680
rect 880 7272 22120 7552
rect 800 7144 22202 7272
rect 880 6864 22120 7144
rect 800 6736 22202 6864
rect 880 6456 22120 6736
rect 800 6328 22202 6456
rect 880 6048 22120 6328
rect 800 5920 22202 6048
rect 880 5640 22120 5920
rect 800 5512 22202 5640
rect 880 5232 22120 5512
rect 800 5104 22202 5232
rect 880 4824 22120 5104
rect 800 4696 22202 4824
rect 880 4416 22120 4696
rect 800 4288 22202 4416
rect 880 4008 22120 4288
rect 800 3880 22202 4008
rect 880 3600 22120 3880
rect 800 3472 22202 3600
rect 880 3192 22120 3472
rect 800 3064 22202 3192
rect 880 2784 22120 3064
rect 800 2656 22202 2784
rect 880 2376 22120 2656
rect 800 2248 22202 2376
rect 880 1968 22120 2248
rect 800 1840 22202 1968
rect 880 1560 22120 1840
rect 800 1531 22202 1560
<< metal4 >>
rect 3543 2128 3863 20720
rect 6142 2128 6462 20720
rect 8741 2128 9061 20720
rect 11340 2128 11660 20720
rect 13939 2128 14259 20720
rect 16538 2128 16858 20720
rect 19137 2128 19457 20720
rect 21736 2128 22056 20720
<< obsm4 >>
rect 979 2048 3463 20501
rect 3943 2048 6062 20501
rect 6542 2048 8661 20501
rect 9141 2048 11260 20501
rect 11740 2048 13859 20501
rect 14339 2048 16458 20501
rect 16938 2048 19057 20501
rect 19537 2048 20549 20501
rect 979 1667 20549 2048
<< labels >>
rlabel metal2 s 19890 0 19946 800 6 SC_IN_BOT
port 1 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 SC_OUT_BOT
port 2 nsew signal output
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 21736 2128 22056 20720 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 4 nsew power bidirectional
rlabel metal2 s 2226 0 2282 800 6 bottom_left_grid_pin_42_
port 5 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 bottom_left_grid_pin_43_
port 6 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 bottom_left_grid_pin_44_
port 7 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 bottom_left_grid_pin_45_
port 8 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 bottom_left_grid_pin_46_
port 9 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 bottom_left_grid_pin_47_
port 10 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 bottom_left_grid_pin_48_
port 11 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 bottom_left_grid_pin_49_
port 12 nsew signal input
rlabel metal2 s 5722 22200 5778 23000 6 ccff_head
port 13 nsew signal input
rlabel metal2 s 17222 22200 17278 23000 6 ccff_tail
port 14 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 chanx_left_in[0]
port 15 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[10]
port 16 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[11]
port 17 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 chanx_left_in[12]
port 18 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 chanx_left_in[13]
port 19 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 chanx_left_in[14]
port 20 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 chanx_left_in[15]
port 21 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 chanx_left_in[16]
port 22 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[17]
port 23 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[18]
port 24 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[19]
port 25 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 chanx_left_in[1]
port 26 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[2]
port 27 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[3]
port 28 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 chanx_left_in[4]
port 29 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 chanx_left_in[5]
port 30 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 chanx_left_in[6]
port 31 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 chanx_left_in[7]
port 32 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 chanx_left_in[8]
port 33 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[9]
port 34 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 chanx_left_out[0]
port 35 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 chanx_left_out[10]
port 36 nsew signal output
rlabel metal3 s 0 17552 800 17672 6 chanx_left_out[11]
port 37 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[12]
port 38 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[13]
port 39 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[14]
port 40 nsew signal output
rlabel metal3 s 0 19184 800 19304 6 chanx_left_out[15]
port 41 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 chanx_left_out[16]
port 42 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 chanx_left_out[17]
port 43 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 chanx_left_out[18]
port 44 nsew signal output
rlabel metal3 s 0 20816 800 20936 6 chanx_left_out[19]
port 45 nsew signal output
rlabel metal3 s 0 13472 800 13592 6 chanx_left_out[1]
port 46 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 chanx_left_out[2]
port 47 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 chanx_left_out[3]
port 48 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 chanx_left_out[4]
port 49 nsew signal output
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[5]
port 50 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[6]
port 51 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 chanx_left_out[7]
port 52 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 chanx_left_out[8]
port 53 nsew signal output
rlabel metal3 s 0 16736 800 16856 6 chanx_left_out[9]
port 54 nsew signal output
rlabel metal3 s 22200 4904 23000 5024 6 chanx_right_in[0]
port 55 nsew signal input
rlabel metal3 s 22200 8984 23000 9104 6 chanx_right_in[10]
port 56 nsew signal input
rlabel metal3 s 22200 9392 23000 9512 6 chanx_right_in[11]
port 57 nsew signal input
rlabel metal3 s 22200 9800 23000 9920 6 chanx_right_in[12]
port 58 nsew signal input
rlabel metal3 s 22200 10208 23000 10328 6 chanx_right_in[13]
port 59 nsew signal input
rlabel metal3 s 22200 10616 23000 10736 6 chanx_right_in[14]
port 60 nsew signal input
rlabel metal3 s 22200 11024 23000 11144 6 chanx_right_in[15]
port 61 nsew signal input
rlabel metal3 s 22200 11432 23000 11552 6 chanx_right_in[16]
port 62 nsew signal input
rlabel metal3 s 22200 11840 23000 11960 6 chanx_right_in[17]
port 63 nsew signal input
rlabel metal3 s 22200 12248 23000 12368 6 chanx_right_in[18]
port 64 nsew signal input
rlabel metal3 s 22200 12656 23000 12776 6 chanx_right_in[19]
port 65 nsew signal input
rlabel metal3 s 22200 5312 23000 5432 6 chanx_right_in[1]
port 66 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 chanx_right_in[2]
port 67 nsew signal input
rlabel metal3 s 22200 6128 23000 6248 6 chanx_right_in[3]
port 68 nsew signal input
rlabel metal3 s 22200 6536 23000 6656 6 chanx_right_in[4]
port 69 nsew signal input
rlabel metal3 s 22200 6944 23000 7064 6 chanx_right_in[5]
port 70 nsew signal input
rlabel metal3 s 22200 7352 23000 7472 6 chanx_right_in[6]
port 71 nsew signal input
rlabel metal3 s 22200 7760 23000 7880 6 chanx_right_in[7]
port 72 nsew signal input
rlabel metal3 s 22200 8168 23000 8288 6 chanx_right_in[8]
port 73 nsew signal input
rlabel metal3 s 22200 8576 23000 8696 6 chanx_right_in[9]
port 74 nsew signal input
rlabel metal3 s 22200 13064 23000 13184 6 chanx_right_out[0]
port 75 nsew signal output
rlabel metal3 s 22200 17144 23000 17264 6 chanx_right_out[10]
port 76 nsew signal output
rlabel metal3 s 22200 17552 23000 17672 6 chanx_right_out[11]
port 77 nsew signal output
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[12]
port 78 nsew signal output
rlabel metal3 s 22200 18368 23000 18488 6 chanx_right_out[13]
port 79 nsew signal output
rlabel metal3 s 22200 18776 23000 18896 6 chanx_right_out[14]
port 80 nsew signal output
rlabel metal3 s 22200 19184 23000 19304 6 chanx_right_out[15]
port 81 nsew signal output
rlabel metal3 s 22200 19592 23000 19712 6 chanx_right_out[16]
port 82 nsew signal output
rlabel metal3 s 22200 20000 23000 20120 6 chanx_right_out[17]
port 83 nsew signal output
rlabel metal3 s 22200 20408 23000 20528 6 chanx_right_out[18]
port 84 nsew signal output
rlabel metal3 s 22200 20816 23000 20936 6 chanx_right_out[19]
port 85 nsew signal output
rlabel metal3 s 22200 13472 23000 13592 6 chanx_right_out[1]
port 86 nsew signal output
rlabel metal3 s 22200 13880 23000 14000 6 chanx_right_out[2]
port 87 nsew signal output
rlabel metal3 s 22200 14288 23000 14408 6 chanx_right_out[3]
port 88 nsew signal output
rlabel metal3 s 22200 14696 23000 14816 6 chanx_right_out[4]
port 89 nsew signal output
rlabel metal3 s 22200 15104 23000 15224 6 chanx_right_out[5]
port 90 nsew signal output
rlabel metal3 s 22200 15512 23000 15632 6 chanx_right_out[6]
port 91 nsew signal output
rlabel metal3 s 22200 15920 23000 16040 6 chanx_right_out[7]
port 92 nsew signal output
rlabel metal3 s 22200 16328 23000 16448 6 chanx_right_out[8]
port 93 nsew signal output
rlabel metal3 s 22200 16736 23000 16856 6 chanx_right_out[9]
port 94 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 chany_bottom_in[0]
port 95 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 chany_bottom_in[10]
port 96 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[11]
port 97 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[12]
port 98 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 chany_bottom_in[13]
port 99 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 chany_bottom_in[14]
port 100 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 chany_bottom_in[15]
port 101 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 chany_bottom_in[16]
port 102 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[17]
port 103 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 chany_bottom_in[18]
port 104 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 chany_bottom_in[19]
port 105 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 chany_bottom_in[1]
port 106 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 chany_bottom_in[2]
port 107 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 chany_bottom_in[3]
port 108 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 chany_bottom_in[4]
port 109 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 chany_bottom_in[5]
port 110 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 chany_bottom_in[6]
port 111 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 chany_bottom_in[7]
port 112 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[8]
port 113 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 chany_bottom_in[9]
port 114 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 chany_bottom_out[0]
port 115 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 chany_bottom_out[10]
port 116 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 chany_bottom_out[11]
port 117 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_out[12]
port 118 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 chany_bottom_out[13]
port 119 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_out[14]
port 120 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 chany_bottom_out[15]
port 121 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 chany_bottom_out[16]
port 122 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 chany_bottom_out[17]
port 123 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 chany_bottom_out[18]
port 124 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 chany_bottom_out[19]
port 125 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 chany_bottom_out[1]
port 126 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_out[2]
port 127 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 chany_bottom_out[3]
port 128 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 chany_bottom_out[4]
port 129 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 chany_bottom_out[5]
port 130 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_out[6]
port 131 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 chany_bottom_out[7]
port 132 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_out[8]
port 133 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 chany_bottom_out[9]
port 134 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 left_bottom_grid_pin_34_
port 135 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 left_bottom_grid_pin_35_
port 136 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_36_
port 137 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_37_
port 138 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 left_bottom_grid_pin_38_
port 139 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 left_bottom_grid_pin_39_
port 140 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 left_bottom_grid_pin_40_
port 141 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 left_bottom_grid_pin_41_
port 142 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 left_top_grid_pin_1_
port 143 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 prog_clk_0_S_in
port 144 nsew signal input
rlabel metal3 s 22200 1640 23000 1760 6 right_bottom_grid_pin_34_
port 145 nsew signal input
rlabel metal3 s 22200 2048 23000 2168 6 right_bottom_grid_pin_35_
port 146 nsew signal input
rlabel metal3 s 22200 2456 23000 2576 6 right_bottom_grid_pin_36_
port 147 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_37_
port 148 nsew signal input
rlabel metal3 s 22200 3272 23000 3392 6 right_bottom_grid_pin_38_
port 149 nsew signal input
rlabel metal3 s 22200 3680 23000 3800 6 right_bottom_grid_pin_39_
port 150 nsew signal input
rlabel metal3 s 22200 4088 23000 4208 6 right_bottom_grid_pin_40_
port 151 nsew signal input
rlabel metal3 s 22200 4496 23000 4616 6 right_bottom_grid_pin_41_
port 152 nsew signal input
rlabel metal3 s 22200 21224 23000 21344 6 right_top_grid_pin_1_
port 153 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1867384
string GDS_FILE /home/marwan/clear_signoff_final/openlane/sb_1__2_/runs/sb_1__2_/results/signoff/sb_1__2_.magic.gds
string GDS_START 94420
<< end >>

