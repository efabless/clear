magic
tech sky130A
magscale 1 2
timestamp 1680902895
<< viali >>
rect 26433 24361 26467 24395
rect 27261 24361 27295 24395
rect 29745 24361 29779 24395
rect 31493 24361 31527 24395
rect 38669 24361 38703 24395
rect 39313 24361 39347 24395
rect 41061 24361 41095 24395
rect 43729 24361 43763 24395
rect 44373 24361 44407 24395
rect 24593 24293 24627 24327
rect 25789 24293 25823 24327
rect 31677 24293 31711 24327
rect 32965 24293 32999 24327
rect 38209 24293 38243 24327
rect 46673 24293 46707 24327
rect 2973 24225 3007 24259
rect 5825 24225 5859 24259
rect 8217 24225 8251 24259
rect 10701 24225 10735 24259
rect 13277 24225 13311 24259
rect 15853 24225 15887 24259
rect 18429 24225 18463 24259
rect 20913 24225 20947 24259
rect 22477 24225 22511 24259
rect 25145 24225 25179 24259
rect 29193 24225 29227 24259
rect 34253 24225 34287 24259
rect 35081 24225 35115 24259
rect 36737 24225 36771 24259
rect 37565 24225 37599 24259
rect 40601 24225 40635 24259
rect 41429 24225 41463 24259
rect 48513 24225 48547 24259
rect 3433 24157 3467 24191
rect 3985 24157 4019 24191
rect 4629 24157 4663 24191
rect 6561 24157 6595 24191
rect 7389 24157 7423 24191
rect 9321 24157 9355 24191
rect 11161 24157 11195 24191
rect 11897 24157 11931 24191
rect 13737 24157 13771 24191
rect 14473 24157 14507 24191
rect 16313 24157 16347 24191
rect 18889 24157 18923 24191
rect 19625 24157 19659 24191
rect 21373 24157 21407 24191
rect 22017 24157 22051 24191
rect 23857 24157 23891 24191
rect 25973 24157 26007 24191
rect 27905 24157 27939 24191
rect 28549 24157 28583 24191
rect 29929 24157 29963 24191
rect 30389 24157 30423 24191
rect 31033 24157 31067 24191
rect 32505 24157 32539 24191
rect 33149 24157 33183 24191
rect 36553 24157 36587 24191
rect 38853 24157 38887 24191
rect 39497 24157 39531 24191
rect 40417 24157 40451 24191
rect 42073 24157 42107 24191
rect 42625 24157 42659 24191
rect 43269 24157 43303 24191
rect 43913 24157 43947 24191
rect 44557 24157 44591 24191
rect 46213 24157 46247 24191
rect 46857 24157 46891 24191
rect 47225 24157 47259 24191
rect 48053 24157 48087 24191
rect 48789 24157 48823 24191
rect 24961 24089 24995 24123
rect 26617 24089 26651 24123
rect 26801 24089 26835 24123
rect 27353 24089 27387 24123
rect 29009 24089 29043 24123
rect 33977 24089 34011 24123
rect 35173 24089 35207 24123
rect 36461 24089 36495 24123
rect 37841 24089 37875 24123
rect 40509 24089 40543 24123
rect 45385 24089 45419 24123
rect 4169 24021 4203 24055
rect 6745 24021 6779 24055
rect 9137 24021 9171 24055
rect 11713 24021 11747 24055
rect 14289 24021 14323 24055
rect 17049 24021 17083 24055
rect 19441 24021 19475 24055
rect 24041 24021 24075 24055
rect 25053 24021 25087 24055
rect 28089 24021 28123 24055
rect 28733 24021 28767 24055
rect 30573 24021 30607 24055
rect 31217 24021 31251 24055
rect 31953 24021 31987 24055
rect 32321 24021 32355 24055
rect 33609 24021 33643 24055
rect 34069 24021 34103 24055
rect 35265 24021 35299 24055
rect 35633 24021 35667 24055
rect 36093 24021 36127 24055
rect 37749 24021 37783 24055
rect 40049 24021 40083 24055
rect 45293 24021 45327 24055
rect 46029 24021 46063 24055
rect 47869 24021 47903 24055
rect 2329 23817 2363 23851
rect 21465 23817 21499 23851
rect 23765 23817 23799 23851
rect 28457 23817 28491 23851
rect 32321 23817 32355 23851
rect 32781 23817 32815 23851
rect 37473 23817 37507 23851
rect 37841 23817 37875 23851
rect 41981 23817 42015 23851
rect 42257 23817 42291 23851
rect 47593 23817 47627 23851
rect 49341 23817 49375 23851
rect 14289 23749 14323 23783
rect 20269 23749 20303 23783
rect 21005 23749 21039 23783
rect 24501 23749 24535 23783
rect 26341 23749 26375 23783
rect 31493 23749 31527 23783
rect 37933 23749 37967 23783
rect 41797 23749 41831 23783
rect 42533 23749 42567 23783
rect 46949 23749 46983 23783
rect 47777 23749 47811 23783
rect 2145 23681 2179 23715
rect 4077 23681 4111 23715
rect 4721 23681 4755 23715
rect 6837 23681 6871 23715
rect 7297 23681 7331 23715
rect 9321 23681 9355 23715
rect 11161 23681 11195 23715
rect 12357 23681 12391 23715
rect 13093 23681 13127 23715
rect 16313 23681 16347 23715
rect 18245 23681 18279 23715
rect 21281 23681 21315 23715
rect 22845 23681 22879 23715
rect 23673 23681 23707 23715
rect 27353 23681 27387 23715
rect 27813 23681 27847 23715
rect 28641 23681 28675 23715
rect 29101 23681 29135 23715
rect 29561 23681 29595 23715
rect 32689 23681 32723 23715
rect 36277 23681 36311 23715
rect 39221 23681 39255 23715
rect 40233 23681 40267 23715
rect 40969 23681 41003 23715
rect 42625 23681 42659 23715
rect 43085 23681 43119 23715
rect 44833 23681 44867 23715
rect 45937 23681 45971 23715
rect 46765 23681 46799 23715
rect 47409 23681 47443 23715
rect 48881 23681 48915 23715
rect 3709 23613 3743 23647
rect 5457 23613 5491 23647
rect 8861 23613 8895 23647
rect 10609 23613 10643 23647
rect 12633 23613 12667 23647
rect 15853 23613 15887 23647
rect 17877 23613 17911 23647
rect 20545 23613 20579 23647
rect 22569 23613 22603 23647
rect 23857 23613 23891 23647
rect 26617 23613 26651 23647
rect 31769 23613 31803 23647
rect 32965 23613 32999 23647
rect 35081 23613 35115 23647
rect 35357 23613 35391 23647
rect 36369 23613 36403 23647
rect 36461 23613 36495 23647
rect 38025 23613 38059 23647
rect 38577 23613 38611 23647
rect 39313 23613 39347 23647
rect 39497 23613 39531 23647
rect 40693 23613 40727 23647
rect 46397 23613 46431 23647
rect 49157 23613 49191 23647
rect 7481 23545 7515 23579
rect 35909 23545 35943 23579
rect 38853 23545 38887 23579
rect 40049 23545 40083 23579
rect 48237 23545 48271 23579
rect 6653 23477 6687 23511
rect 18797 23477 18831 23511
rect 23305 23477 23339 23511
rect 24409 23477 24443 23511
rect 24869 23477 24903 23511
rect 27169 23477 27203 23511
rect 27997 23477 28031 23511
rect 29285 23477 29319 23511
rect 30021 23477 30055 23511
rect 33609 23477 33643 23511
rect 36921 23477 36955 23511
rect 45293 23477 45327 23511
rect 46213 23477 46247 23511
rect 4721 23273 4755 23307
rect 20361 23273 20395 23307
rect 25237 23273 25271 23307
rect 27905 23273 27939 23307
rect 29101 23273 29135 23307
rect 30757 23273 30791 23307
rect 31125 23273 31159 23307
rect 34161 23273 34195 23307
rect 38779 23273 38813 23307
rect 44281 23273 44315 23307
rect 45201 23273 45235 23307
rect 46673 23273 46707 23307
rect 46949 23273 46983 23307
rect 9137 23205 9171 23239
rect 14197 23205 14231 23239
rect 19625 23205 19659 23239
rect 24593 23205 24627 23239
rect 29009 23205 29043 23239
rect 29745 23205 29779 23239
rect 34437 23205 34471 23239
rect 37289 23205 37323 23239
rect 40049 23205 40083 23239
rect 44741 23205 44775 23239
rect 6101 23137 6135 23171
rect 7849 23137 7883 23171
rect 10057 23137 10091 23171
rect 11253 23137 11287 23171
rect 13277 23137 13311 23171
rect 15761 23137 15795 23171
rect 22109 23137 22143 23171
rect 23949 23137 23983 23171
rect 25973 23137 26007 23171
rect 28457 23137 28491 23171
rect 30205 23137 30239 23171
rect 30297 23137 30331 23171
rect 33149 23137 33183 23171
rect 35081 23137 35115 23171
rect 39037 23137 39071 23171
rect 39497 23137 39531 23171
rect 40601 23137 40635 23171
rect 43545 23137 43579 23171
rect 45661 23137 45695 23171
rect 2973 23069 3007 23103
rect 4261 23069 4295 23103
rect 4905 23069 4939 23103
rect 5365 23069 5399 23103
rect 7205 23069 7239 23103
rect 9321 23069 9355 23103
rect 11897 23069 11931 23103
rect 13737 23069 13771 23103
rect 14841 23069 14875 23103
rect 16681 23069 16715 23103
rect 18889 23069 18923 23103
rect 22753 23069 22787 23103
rect 23673 23069 23707 23103
rect 25697 23069 25731 23103
rect 28365 23069 28399 23103
rect 29377 23069 29411 23103
rect 31401 23069 31435 23103
rect 33885 23069 33919 23103
rect 34713 23069 34747 23103
rect 41061 23069 41095 23103
rect 44373 23069 44407 23103
rect 45385 23069 45419 23103
rect 46305 23069 46339 23103
rect 47133 23069 47167 23103
rect 47869 23069 47903 23103
rect 48605 23069 48639 23103
rect 49341 23069 49375 23103
rect 1777 23001 1811 23035
rect 18613 23001 18647 23035
rect 19809 23001 19843 23035
rect 21833 23001 21867 23035
rect 22569 23001 22603 23035
rect 24777 23001 24811 23035
rect 31677 23001 31711 23035
rect 35357 23001 35391 23035
rect 40509 23001 40543 23035
rect 41521 23001 41555 23035
rect 43269 23001 43303 23035
rect 4077 22933 4111 22967
rect 14381 22933 14415 22967
rect 14657 22933 14691 22967
rect 17141 22933 17175 22967
rect 19349 22933 19383 22967
rect 23305 22933 23339 22967
rect 23765 22933 23799 22967
rect 25329 22933 25363 22967
rect 27445 22933 27479 22967
rect 28273 22933 28307 22967
rect 30113 22933 30147 22967
rect 33701 22933 33735 22967
rect 36829 22933 36863 22967
rect 39405 22933 39439 22967
rect 40417 22933 40451 22967
rect 43821 22933 43855 22967
rect 46121 22933 46155 22967
rect 47685 22933 47719 22967
rect 48421 22933 48455 22967
rect 49157 22933 49191 22967
rect 7205 22729 7239 22763
rect 18613 22729 18647 22763
rect 19165 22729 19199 22763
rect 21189 22729 21223 22763
rect 32321 22729 32355 22763
rect 32781 22729 32815 22763
rect 35449 22729 35483 22763
rect 37473 22729 37507 22763
rect 40509 22729 40543 22763
rect 46397 22729 46431 22763
rect 4813 22661 4847 22695
rect 9965 22661 9999 22695
rect 11897 22661 11931 22695
rect 12817 22661 12851 22695
rect 15117 22661 15151 22695
rect 17141 22661 17175 22695
rect 22293 22661 22327 22695
rect 24133 22661 24167 22695
rect 26341 22661 26375 22695
rect 27721 22661 27755 22695
rect 30665 22661 30699 22695
rect 30757 22661 30791 22695
rect 38945 22661 38979 22695
rect 40417 22661 40451 22695
rect 47593 22661 47627 22695
rect 2973 22593 3007 22627
rect 3985 22593 4019 22627
rect 6009 22593 6043 22627
rect 6653 22593 6687 22627
rect 7481 22593 7515 22627
rect 9321 22593 9355 22627
rect 11161 22593 11195 22627
rect 14013 22593 14047 22627
rect 16313 22593 16347 22627
rect 22017 22593 22051 22627
rect 24409 22593 24443 22627
rect 26617 22593 26651 22627
rect 27169 22593 27203 22627
rect 29837 22593 29871 22627
rect 31677 22593 31711 22627
rect 32689 22593 32723 22627
rect 33425 22593 33459 22627
rect 33701 22593 33735 22627
rect 36461 22593 36495 22627
rect 39221 22593 39255 22627
rect 39497 22593 39531 22627
rect 39773 22593 39807 22627
rect 41429 22593 41463 22627
rect 42073 22593 42107 22627
rect 44097 22593 44131 22627
rect 44741 22593 44775 22627
rect 45385 22593 45419 22627
rect 45661 22593 45695 22627
rect 47225 22593 47259 22627
rect 47777 22593 47811 22627
rect 48605 22593 48639 22627
rect 49341 22593 49375 22627
rect 2513 22525 2547 22559
rect 7941 22525 7975 22559
rect 9505 22525 9539 22559
rect 16865 22525 16899 22559
rect 18889 22525 18923 22559
rect 19448 22525 19482 22559
rect 19717 22525 19751 22559
rect 24869 22525 24903 22559
rect 28089 22525 28123 22559
rect 29561 22525 29595 22559
rect 30849 22525 30883 22559
rect 32873 22525 32907 22559
rect 33977 22525 34011 22559
rect 36553 22525 36587 22559
rect 36737 22525 36771 22559
rect 40601 22525 40635 22559
rect 42625 22525 42659 22559
rect 42901 22525 42935 22559
rect 46765 22525 46799 22559
rect 4169 22457 4203 22491
rect 6837 22457 6871 22491
rect 11713 22457 11747 22491
rect 14565 22457 14599 22491
rect 23765 22457 23799 22491
rect 27353 22457 27387 22491
rect 36093 22457 36127 22491
rect 41889 22457 41923 22491
rect 45201 22457 45235 22491
rect 46581 22457 46615 22491
rect 47961 22457 47995 22491
rect 12265 22389 12299 22423
rect 14381 22389 14415 22423
rect 21649 22389 21683 22423
rect 24501 22389 24535 22423
rect 30297 22389 30331 22423
rect 31493 22389 31527 22423
rect 35817 22389 35851 22423
rect 40049 22389 40083 22423
rect 41245 22389 41279 22423
rect 43913 22389 43947 22423
rect 44557 22389 44591 22423
rect 45845 22389 45879 22423
rect 47041 22389 47075 22423
rect 48421 22389 48455 22423
rect 49157 22389 49191 22423
rect 12357 22185 12391 22219
rect 25605 22185 25639 22219
rect 28365 22185 28399 22219
rect 30297 22185 30331 22219
rect 39497 22185 39531 22219
rect 40233 22185 40267 22219
rect 44741 22185 44775 22219
rect 47041 22185 47075 22219
rect 47225 22185 47259 22219
rect 14197 22117 14231 22151
rect 24593 22117 24627 22151
rect 47685 22117 47719 22151
rect 6009 22049 6043 22083
rect 9781 22049 9815 22083
rect 11897 22049 11931 22083
rect 13645 22049 13679 22083
rect 14473 22049 14507 22083
rect 15209 22049 15243 22083
rect 16957 22049 16991 22083
rect 17601 22049 17635 22083
rect 19901 22049 19935 22083
rect 22017 22049 22051 22083
rect 23213 22049 23247 22083
rect 25145 22049 25179 22083
rect 26525 22049 26559 22083
rect 27629 22049 27663 22083
rect 27721 22049 27755 22083
rect 28917 22049 28951 22083
rect 33517 22049 33551 22083
rect 33701 22049 33735 22083
rect 34989 22049 35023 22083
rect 36277 22049 36311 22083
rect 38853 22049 38887 22083
rect 39129 22049 39163 22083
rect 40877 22049 40911 22083
rect 41981 22049 42015 22083
rect 43545 22049 43579 22083
rect 44373 22049 44407 22083
rect 44649 22049 44683 22083
rect 46857 22049 46891 22083
rect 2973 21981 3007 22015
rect 5365 21981 5399 22015
rect 7205 21981 7239 22015
rect 7849 21981 7883 22015
rect 8585 21981 8619 22015
rect 9137 21981 9171 22015
rect 11621 21981 11655 22015
rect 12541 21981 12575 22015
rect 13369 21981 13403 22015
rect 13461 21981 13495 22015
rect 18797 21981 18831 22015
rect 19441 21981 19475 22015
rect 24041 21981 24075 22015
rect 25053 21981 25087 22015
rect 26433 21981 26467 22015
rect 27537 21981 27571 22015
rect 29929 21981 29963 22015
rect 30849 21981 30883 22015
rect 34069 21981 34103 22015
rect 34437 21981 34471 22015
rect 41889 21981 41923 22015
rect 42809 21981 42843 22015
rect 43269 21981 43303 22015
rect 47869 21981 47903 22015
rect 48513 21981 48547 22015
rect 1777 21913 1811 21947
rect 4169 21913 4203 21947
rect 7665 21913 7699 21947
rect 14657 21913 14691 21947
rect 16681 21913 16715 21947
rect 21189 21913 21223 21947
rect 21833 21913 21867 21947
rect 23029 21913 23063 21947
rect 24961 21913 24995 21947
rect 26341 21913 26375 21947
rect 28825 21913 28859 21947
rect 31125 21913 31159 21947
rect 35265 21913 35299 21947
rect 40693 21913 40727 21947
rect 47409 21913 47443 21947
rect 49065 21913 49099 21947
rect 49249 21913 49283 21947
rect 8401 21845 8435 21879
rect 13001 21845 13035 21879
rect 21465 21845 21499 21879
rect 21925 21845 21959 21879
rect 22661 21845 22695 21879
rect 23121 21845 23155 21879
rect 23857 21845 23891 21879
rect 25973 21845 26007 21879
rect 27169 21845 27203 21879
rect 28733 21845 28767 21879
rect 29745 21845 29779 21879
rect 30389 21845 30423 21879
rect 32597 21845 32631 21879
rect 33057 21845 33091 21879
rect 33425 21845 33459 21879
rect 34345 21845 34379 21879
rect 35173 21845 35207 21879
rect 35633 21845 35667 21879
rect 36369 21845 36403 21879
rect 36461 21845 36495 21879
rect 36829 21845 36863 21879
rect 37381 21845 37415 21879
rect 39681 21845 39715 21879
rect 39865 21845 39899 21879
rect 40601 21845 40635 21879
rect 41429 21845 41463 21879
rect 41797 21845 41831 21879
rect 42625 21845 42659 21879
rect 48421 21845 48455 21879
rect 10517 21641 10551 21675
rect 13921 21641 13955 21675
rect 17417 21641 17451 21675
rect 17877 21641 17911 21675
rect 24777 21641 24811 21675
rect 27169 21641 27203 21675
rect 27629 21641 27663 21675
rect 30021 21641 30055 21675
rect 32781 21641 32815 21675
rect 33977 21641 34011 21675
rect 36093 21641 36127 21675
rect 40141 21641 40175 21675
rect 40325 21641 40359 21675
rect 40509 21641 40543 21675
rect 40693 21641 40727 21675
rect 43361 21641 43395 21675
rect 43637 21641 43671 21675
rect 43913 21641 43947 21675
rect 3617 21573 3651 21607
rect 13093 21573 13127 21607
rect 14841 21573 14875 21607
rect 21189 21573 21223 21607
rect 22753 21573 22787 21607
rect 27537 21573 27571 21607
rect 31125 21573 31159 21607
rect 33609 21573 33643 21607
rect 34805 21573 34839 21607
rect 38301 21573 38335 21607
rect 42533 21573 42567 21607
rect 42717 21573 42751 21607
rect 42993 21573 43027 21607
rect 2973 21505 3007 21539
rect 4629 21505 4663 21539
rect 5733 21505 5767 21539
rect 6653 21505 6687 21539
rect 8493 21505 8527 21539
rect 10701 21505 10735 21539
rect 11161 21505 11195 21539
rect 12357 21505 12391 21539
rect 13277 21505 13311 21539
rect 14105 21505 14139 21539
rect 17785 21505 17819 21539
rect 21373 21505 21407 21539
rect 25145 21505 25179 21539
rect 26065 21505 26099 21539
rect 26617 21505 26651 21539
rect 28733 21505 28767 21539
rect 29929 21505 29963 21539
rect 31217 21505 31251 21539
rect 33517 21505 33551 21539
rect 34713 21505 34747 21539
rect 43269 21505 43303 21539
rect 47961 21505 47995 21539
rect 48605 21505 48639 21539
rect 49341 21505 49375 21539
rect 1777 21437 1811 21471
rect 7021 21437 7055 21471
rect 8861 21437 8895 21471
rect 11713 21437 11747 21471
rect 11897 21437 11931 21471
rect 12817 21437 12851 21471
rect 14565 21437 14599 21471
rect 16313 21437 16347 21471
rect 18061 21437 18095 21471
rect 18613 21437 18647 21471
rect 18889 21437 18923 21471
rect 22477 21437 22511 21471
rect 24225 21437 24259 21471
rect 25237 21437 25271 21471
rect 25421 21437 25455 21471
rect 27721 21437 27755 21471
rect 28825 21437 28859 21471
rect 28917 21437 28951 21471
rect 30113 21437 30147 21471
rect 31401 21437 31435 21471
rect 31769 21437 31803 21471
rect 33425 21437 33459 21471
rect 34529 21437 34563 21471
rect 36185 21437 36219 21471
rect 36277 21437 36311 21471
rect 36829 21437 36863 21471
rect 37289 21437 37323 21471
rect 37657 21437 37691 21471
rect 38014 21437 38048 21471
rect 41245 21437 41279 21471
rect 41521 21437 41555 21471
rect 5917 21369 5951 21403
rect 16773 21369 16807 21403
rect 17141 21369 17175 21403
rect 20361 21369 20395 21403
rect 26433 21369 26467 21403
rect 47777 21369 47811 21403
rect 48421 21369 48455 21403
rect 11345 21301 11379 21335
rect 12265 21301 12299 21335
rect 16957 21301 16991 21335
rect 20729 21301 20763 21335
rect 20913 21301 20947 21335
rect 22017 21301 22051 21335
rect 22201 21301 22235 21335
rect 25881 21301 25915 21335
rect 28365 21301 28399 21335
rect 29561 21301 29595 21335
rect 30757 21301 30791 21335
rect 35173 21301 35207 21335
rect 35725 21301 35759 21335
rect 36921 21301 36955 21335
rect 37565 21301 37599 21335
rect 39773 21301 39807 21335
rect 40877 21301 40911 21335
rect 42809 21301 42843 21335
rect 49157 21301 49191 21335
rect 9229 21097 9263 21131
rect 12449 21097 12483 21131
rect 14289 21097 14323 21131
rect 17141 21097 17175 21131
rect 24041 21097 24075 21131
rect 24225 21097 24259 21131
rect 26893 21097 26927 21131
rect 29745 21097 29779 21131
rect 30205 21097 30239 21131
rect 37657 21097 37691 21131
rect 40049 21097 40083 21131
rect 42441 21097 42475 21131
rect 42993 21097 43027 21131
rect 48053 21097 48087 21131
rect 48605 21097 48639 21131
rect 11805 21029 11839 21063
rect 19993 21029 20027 21063
rect 21189 21029 21223 21063
rect 23397 21029 23431 21063
rect 24777 21029 24811 21063
rect 25237 21029 25271 21063
rect 25421 21029 25455 21063
rect 30389 21029 30423 21063
rect 31953 21029 31987 21063
rect 34897 21029 34931 21063
rect 37381 21029 37415 21063
rect 49157 21029 49191 21063
rect 2513 20961 2547 20995
rect 4169 20961 4203 20995
rect 6009 20961 6043 20995
rect 10057 20961 10091 20995
rect 12725 20961 12759 20995
rect 20545 20961 20579 20995
rect 26341 20961 26375 20995
rect 27905 20961 27939 20995
rect 28549 20961 28583 20995
rect 31309 20961 31343 20995
rect 31493 20961 31527 20995
rect 32781 20961 32815 20995
rect 39405 20961 39439 20995
rect 40509 20961 40543 20995
rect 40601 20961 40635 20995
rect 41797 20961 41831 20995
rect 42625 20961 42659 20995
rect 42901 20961 42935 20995
rect 47961 20961 47995 20995
rect 2973 20893 3007 20927
rect 5365 20893 5399 20927
rect 7205 20893 7239 20927
rect 8033 20893 8067 20927
rect 8401 20893 8435 20927
rect 9413 20893 9447 20927
rect 11345 20889 11379 20923
rect 13737 20893 13771 20927
rect 16037 20893 16071 20927
rect 18889 20893 18923 20927
rect 20361 20893 20395 20927
rect 22937 20893 22971 20927
rect 24593 20893 24627 20927
rect 29929 20893 29963 20927
rect 32505 20893 32539 20927
rect 36645 20893 36679 20927
rect 41613 20893 41647 20927
rect 48421 20893 48455 20927
rect 49341 20893 49375 20927
rect 11989 20825 12023 20859
rect 12909 20825 12943 20859
rect 15761 20825 15795 20859
rect 16681 20825 16715 20859
rect 18613 20825 18647 20859
rect 20453 20825 20487 20859
rect 22661 20825 22695 20859
rect 23581 20825 23615 20859
rect 26065 20825 26099 20859
rect 27445 20825 27479 20859
rect 36369 20825 36403 20859
rect 37197 20825 37231 20859
rect 39129 20825 39163 20859
rect 40417 20825 40451 20859
rect 48789 20825 48823 20859
rect 7573 20757 7607 20791
rect 7849 20757 7883 20791
rect 10701 20757 10735 20791
rect 11161 20757 11195 20791
rect 13553 20757 13587 20791
rect 19349 20757 19383 20791
rect 19533 20757 19567 20791
rect 19625 20757 19659 20791
rect 25697 20757 25731 20791
rect 26157 20757 26191 20791
rect 26709 20757 26743 20791
rect 28641 20757 28675 20791
rect 28733 20757 28767 20791
rect 29101 20757 29135 20791
rect 30849 20757 30883 20791
rect 31217 20757 31251 20791
rect 34253 20757 34287 20791
rect 37013 20757 37047 20791
rect 41245 20757 41279 20791
rect 41705 20757 41739 20791
rect 42257 20757 42291 20791
rect 5457 20553 5491 20587
rect 9689 20553 9723 20587
rect 10333 20553 10367 20587
rect 11161 20553 11195 20587
rect 13737 20553 13771 20587
rect 14105 20553 14139 20587
rect 14933 20553 14967 20587
rect 15577 20553 15611 20587
rect 15945 20553 15979 20587
rect 16037 20553 16071 20587
rect 18797 20553 18831 20587
rect 19717 20553 19751 20587
rect 35265 20553 35299 20587
rect 40325 20553 40359 20587
rect 3617 20485 3651 20519
rect 12449 20485 12483 20519
rect 22385 20485 22419 20519
rect 29837 20485 29871 20519
rect 31033 20485 31067 20519
rect 31769 20485 31803 20519
rect 36553 20485 36587 20519
rect 40233 20485 40267 20519
rect 41797 20485 41831 20519
rect 2973 20417 3007 20451
rect 4813 20417 4847 20451
rect 5273 20417 5307 20451
rect 6561 20417 6595 20451
rect 9229 20417 9263 20451
rect 9873 20417 9907 20451
rect 10517 20417 10551 20451
rect 11713 20417 11747 20451
rect 11897 20417 11931 20451
rect 12633 20417 12667 20451
rect 14197 20417 14231 20451
rect 15117 20417 15151 20451
rect 17049 20417 17083 20451
rect 21465 20417 21499 20451
rect 23397 20417 23431 20451
rect 23857 20417 23891 20451
rect 26065 20417 26099 20451
rect 27261 20417 27295 20451
rect 29745 20417 29779 20451
rect 34897 20417 34931 20451
rect 35541 20417 35575 20451
rect 36461 20417 36495 20451
rect 39497 20417 39531 20451
rect 41613 20417 41647 20451
rect 48605 20417 48639 20451
rect 49341 20417 49375 20451
rect 2513 20349 2547 20383
rect 7021 20349 7055 20383
rect 14289 20349 14323 20383
rect 16221 20349 16255 20383
rect 17325 20349 17359 20383
rect 21189 20349 21223 20383
rect 22477 20349 22511 20383
rect 22569 20349 22603 20383
rect 24133 20349 24167 20383
rect 25605 20349 25639 20383
rect 27537 20349 27571 20383
rect 29009 20349 29043 20383
rect 29561 20349 29595 20383
rect 31125 20349 31159 20383
rect 31309 20349 31343 20383
rect 32321 20349 32355 20383
rect 33793 20349 33827 20383
rect 34069 20349 34103 20383
rect 34713 20349 34747 20383
rect 34805 20349 34839 20383
rect 36737 20349 36771 20383
rect 39221 20349 39255 20383
rect 40141 20349 40175 20383
rect 41153 20349 41187 20383
rect 19073 20281 19107 20315
rect 23213 20281 23247 20315
rect 26617 20281 26651 20315
rect 31953 20281 31987 20315
rect 36093 20281 36127 20315
rect 49157 20281 49191 20315
rect 9045 20213 9079 20247
rect 13093 20213 13127 20247
rect 13277 20213 13311 20247
rect 13461 20213 13495 20247
rect 16773 20213 16807 20247
rect 19349 20213 19383 20247
rect 22017 20213 22051 20247
rect 26249 20213 26283 20247
rect 30205 20213 30239 20247
rect 30665 20213 30699 20247
rect 35725 20213 35759 20247
rect 37289 20213 37323 20247
rect 37749 20213 37783 20247
rect 40693 20213 40727 20247
rect 48421 20213 48455 20247
rect 11345 20009 11379 20043
rect 14473 20009 14507 20043
rect 16865 20009 16899 20043
rect 25605 20009 25639 20043
rect 26801 20009 26835 20043
rect 29101 20009 29135 20043
rect 41061 20009 41095 20043
rect 48789 20009 48823 20043
rect 9965 19941 9999 19975
rect 10609 19941 10643 19975
rect 14933 19941 14967 19975
rect 15669 19941 15703 19975
rect 19625 19941 19659 19975
rect 22937 19941 22971 19975
rect 24041 19941 24075 19975
rect 36093 19941 36127 19975
rect 39589 19941 39623 19975
rect 41245 19941 41279 19975
rect 4261 19873 4295 19907
rect 6009 19873 6043 19907
rect 11989 19873 12023 19907
rect 16313 19873 16347 19907
rect 17417 19873 17451 19907
rect 18797 19873 18831 19907
rect 22293 19873 22327 19907
rect 23397 19873 23431 19907
rect 23581 19873 23615 19907
rect 24593 19873 24627 19907
rect 25329 19873 25363 19907
rect 26157 19873 26191 19907
rect 27353 19873 27387 19907
rect 28549 19873 28583 19907
rect 30389 19873 30423 19907
rect 31125 19873 31159 19907
rect 32689 19873 32723 19907
rect 33609 19873 33643 19907
rect 34437 19873 34471 19907
rect 35081 19873 35115 19907
rect 36645 19873 36679 19907
rect 37933 19873 37967 19907
rect 38117 19873 38151 19907
rect 39037 19873 39071 19907
rect 40141 19873 40175 19907
rect 40325 19873 40359 19907
rect 2973 19805 3007 19839
rect 5273 19805 5307 19839
rect 7205 19805 7239 19839
rect 7941 19805 7975 19839
rect 10149 19805 10183 19839
rect 10793 19805 10827 19839
rect 14289 19805 14323 19839
rect 15117 19805 15151 19839
rect 17325 19805 17359 19839
rect 30205 19805 30239 19839
rect 32505 19805 32539 19839
rect 33793 19805 33827 19839
rect 35173 19805 35207 19839
rect 35265 19805 35299 19839
rect 38209 19805 38243 19839
rect 38853 19805 38887 19839
rect 1777 19737 1811 19771
rect 11437 19737 11471 19771
rect 12265 19737 12299 19771
rect 16037 19737 16071 19771
rect 19809 19737 19843 19771
rect 22017 19737 22051 19771
rect 25973 19737 26007 19771
rect 28457 19737 28491 19771
rect 30113 19737 30147 19771
rect 32597 19737 32631 19771
rect 33701 19737 33735 19771
rect 36461 19737 36495 19771
rect 40417 19737 40451 19771
rect 48605 19737 48639 19771
rect 49249 19737 49283 19771
rect 7757 19669 7791 19703
rect 13737 19669 13771 19703
rect 16129 19669 16163 19703
rect 17233 19669 17267 19703
rect 18153 19669 18187 19703
rect 18521 19669 18555 19703
rect 18613 19669 18647 19703
rect 19349 19669 19383 19703
rect 20269 19669 20303 19703
rect 20545 19669 20579 19703
rect 22661 19669 22695 19703
rect 22845 19669 22879 19703
rect 23673 19669 23707 19703
rect 25145 19669 25179 19703
rect 26065 19669 26099 19703
rect 27169 19669 27203 19703
rect 27261 19669 27295 19703
rect 27997 19669 28031 19703
rect 28365 19669 28399 19703
rect 29285 19669 29319 19703
rect 29745 19669 29779 19703
rect 31217 19669 31251 19703
rect 31309 19669 31343 19703
rect 31677 19669 31711 19703
rect 32137 19669 32171 19703
rect 34161 19669 34195 19703
rect 35633 19669 35667 19703
rect 36553 19669 36587 19703
rect 37381 19669 37415 19703
rect 37565 19669 37599 19703
rect 38577 19669 38611 19703
rect 40785 19669 40819 19703
rect 49157 19669 49191 19703
rect 10977 19465 11011 19499
rect 16865 19465 16899 19499
rect 17325 19465 17359 19499
rect 20729 19465 20763 19499
rect 21189 19465 21223 19499
rect 26157 19465 26191 19499
rect 26249 19465 26283 19499
rect 28457 19465 28491 19499
rect 33057 19465 33091 19499
rect 34253 19465 34287 19499
rect 35449 19465 35483 19499
rect 37289 19465 37323 19499
rect 40141 19465 40175 19499
rect 40601 19465 40635 19499
rect 41337 19465 41371 19499
rect 3617 19397 3651 19431
rect 10517 19397 10551 19431
rect 14933 19397 14967 19431
rect 16221 19397 16255 19431
rect 22937 19397 22971 19431
rect 31493 19397 31527 19431
rect 32597 19397 32631 19431
rect 32689 19397 32723 19431
rect 33793 19397 33827 19431
rect 35081 19397 35115 19431
rect 36185 19397 36219 19431
rect 39405 19397 39439 19431
rect 40509 19397 40543 19431
rect 1777 19329 1811 19363
rect 2973 19329 3007 19363
rect 4813 19329 4847 19363
rect 5457 19329 5491 19363
rect 11161 19329 11195 19363
rect 11713 19329 11747 19363
rect 12173 19329 12207 19363
rect 14473 19329 14507 19363
rect 15485 19329 15519 19363
rect 17233 19329 17267 19363
rect 18061 19329 18095 19363
rect 21097 19329 21131 19363
rect 22201 19329 22235 19363
rect 25237 19329 25271 19363
rect 27629 19329 27663 19363
rect 28825 19329 28859 19363
rect 29745 19329 29779 19363
rect 30757 19329 30791 19363
rect 33885 19329 33919 19363
rect 34989 19329 35023 19363
rect 36277 19329 36311 19363
rect 37565 19329 37599 19363
rect 39681 19329 39715 19363
rect 48605 19329 48639 19363
rect 49249 19329 49283 19363
rect 5273 19261 5307 19295
rect 9873 19261 9907 19295
rect 11989 19261 12023 19295
rect 14197 19261 14231 19295
rect 15301 19261 15335 19295
rect 16037 19261 16071 19295
rect 17417 19261 17451 19295
rect 19809 19261 19843 19295
rect 20085 19261 20119 19295
rect 21373 19261 21407 19295
rect 24961 19261 24995 19295
rect 26433 19261 26467 19295
rect 27721 19261 27755 19295
rect 27905 19261 27939 19295
rect 28917 19261 28951 19295
rect 29009 19261 29043 19295
rect 32413 19261 32447 19295
rect 33701 19261 33735 19295
rect 34805 19261 34839 19295
rect 36001 19261 36035 19295
rect 40693 19261 40727 19295
rect 14841 19193 14875 19227
rect 49065 19193 49099 19227
rect 5917 19125 5951 19159
rect 12725 19125 12759 19159
rect 20453 19125 20487 19159
rect 23489 19125 23523 19159
rect 25789 19125 25823 19159
rect 27261 19125 27295 19159
rect 30205 19125 30239 19159
rect 30389 19125 30423 19159
rect 36645 19125 36679 19159
rect 36921 19125 36955 19159
rect 37933 19125 37967 19159
rect 41245 19125 41279 19159
rect 48789 19125 48823 19159
rect 9229 18921 9263 18955
rect 11897 18921 11931 18955
rect 12541 18921 12575 18955
rect 16037 18921 16071 18955
rect 16957 18921 16991 18955
rect 18153 18921 18187 18955
rect 19901 18921 19935 18955
rect 21097 18921 21131 18955
rect 28089 18921 28123 18955
rect 31493 18921 31527 18955
rect 33425 18921 33459 18955
rect 37381 18921 37415 18955
rect 42073 18921 42107 18955
rect 13737 18853 13771 18887
rect 27537 18853 27571 18887
rect 29009 18853 29043 18887
rect 30941 18853 30975 18887
rect 33885 18853 33919 18887
rect 38025 18853 38059 18887
rect 4169 18785 4203 18819
rect 10977 18785 11011 18819
rect 13093 18785 13127 18819
rect 14289 18785 14323 18819
rect 17509 18785 17543 18819
rect 18797 18785 18831 18819
rect 20361 18785 20395 18819
rect 20453 18785 20487 18819
rect 21649 18785 21683 18819
rect 25237 18785 25271 18819
rect 25789 18785 25823 18819
rect 27813 18785 27847 18819
rect 28457 18785 28491 18819
rect 29837 18785 29871 18819
rect 31953 18785 31987 18819
rect 32137 18785 32171 18819
rect 32873 18785 32907 18819
rect 32965 18785 32999 18819
rect 34161 18785 34195 18819
rect 35633 18785 35667 18819
rect 38577 18785 38611 18819
rect 41797 18785 41831 18819
rect 2973 18717 3007 18751
rect 5365 18717 5399 18751
rect 8309 18717 8343 18751
rect 12081 18717 12115 18751
rect 12909 18717 12943 18751
rect 18521 18717 18555 18751
rect 18613 18717 18647 18751
rect 21465 18717 21499 18751
rect 24041 18717 24075 18751
rect 29193 18717 29227 18751
rect 31861 18717 31895 18751
rect 35173 18717 35207 18751
rect 38393 18717 38427 18751
rect 48605 18717 48639 18751
rect 49341 18717 49375 18751
rect 1777 18649 1811 18683
rect 8125 18649 8159 18683
rect 10701 18649 10735 18683
rect 13001 18649 13035 18683
rect 14565 18649 14599 18683
rect 16313 18649 16347 18683
rect 17417 18649 17451 18683
rect 19349 18649 19383 18683
rect 20269 18649 20303 18683
rect 23765 18649 23799 18683
rect 26065 18649 26099 18683
rect 30113 18649 30147 18683
rect 30757 18649 30791 18683
rect 35909 18649 35943 18683
rect 39589 18649 39623 18683
rect 41521 18649 41555 18683
rect 11253 18581 11287 18615
rect 11529 18581 11563 18615
rect 13921 18581 13955 18615
rect 16681 18581 16715 18615
rect 17325 18581 17359 18615
rect 19625 18581 19659 18615
rect 21557 18581 21591 18615
rect 22293 18581 22327 18615
rect 24593 18581 24627 18615
rect 24961 18581 24995 18615
rect 25053 18581 25087 18615
rect 28181 18581 28215 18615
rect 28641 18581 28675 18615
rect 30021 18581 30055 18615
rect 30481 18581 30515 18615
rect 31125 18581 31159 18615
rect 33057 18581 33091 18615
rect 33701 18581 33735 18615
rect 34253 18581 34287 18615
rect 34529 18581 34563 18615
rect 37657 18581 37691 18615
rect 38485 18581 38519 18615
rect 40049 18581 40083 18615
rect 48421 18581 48455 18615
rect 49157 18581 49191 18615
rect 3617 18377 3651 18411
rect 10793 18377 10827 18411
rect 17969 18377 18003 18411
rect 18337 18377 18371 18411
rect 19073 18377 19107 18411
rect 22477 18377 22511 18411
rect 26249 18377 26283 18411
rect 27629 18377 27663 18411
rect 28733 18377 28767 18411
rect 30849 18377 30883 18411
rect 33057 18377 33091 18411
rect 36921 18377 36955 18411
rect 37473 18377 37507 18411
rect 40417 18377 40451 18411
rect 40877 18377 40911 18411
rect 48789 18377 48823 18411
rect 7665 18309 7699 18343
rect 13185 18309 13219 18343
rect 14289 18309 14323 18343
rect 14381 18309 14415 18343
rect 17417 18309 17451 18343
rect 19901 18309 19935 18343
rect 23305 18309 23339 18343
rect 24133 18309 24167 18343
rect 25145 18309 25179 18343
rect 28825 18309 28859 18343
rect 40141 18309 40175 18343
rect 2973 18241 3007 18275
rect 3433 18241 3467 18275
rect 4445 18241 4479 18275
rect 7849 18241 7883 18275
rect 9965 18241 9999 18275
rect 10885 18241 10919 18275
rect 13461 18241 13495 18275
rect 15117 18241 15151 18275
rect 16313 18241 16347 18275
rect 22569 18241 22603 18275
rect 25053 18241 25087 18275
rect 26341 18241 26375 18275
rect 27537 18241 27571 18275
rect 30389 18241 30423 18275
rect 30481 18241 30515 18275
rect 31309 18241 31343 18275
rect 32597 18241 32631 18275
rect 32689 18241 32723 18275
rect 36277 18241 36311 18275
rect 36369 18241 36403 18275
rect 39773 18241 39807 18275
rect 40785 18241 40819 18275
rect 48605 18241 48639 18275
rect 49341 18241 49375 18275
rect 1777 18173 1811 18207
rect 4169 18173 4203 18207
rect 10977 18173 11011 18207
rect 11713 18173 11747 18207
rect 14565 18173 14599 18207
rect 15669 18173 15703 18207
rect 18429 18173 18463 18207
rect 18613 18173 18647 18207
rect 19349 18173 19383 18207
rect 19625 18173 19659 18207
rect 22661 18173 22695 18207
rect 25237 18173 25271 18207
rect 26525 18173 26559 18207
rect 27721 18173 27755 18207
rect 28917 18173 28951 18207
rect 30205 18173 30239 18207
rect 32413 18173 32447 18207
rect 33609 18173 33643 18207
rect 33885 18173 33919 18207
rect 36553 18173 36587 18207
rect 37289 18173 37323 18207
rect 39497 18173 39531 18207
rect 40969 18173 41003 18207
rect 9781 18105 9815 18139
rect 13921 18105 13955 18139
rect 16129 18105 16163 18139
rect 17233 18105 17267 18139
rect 22109 18105 22143 18139
rect 24685 18105 24719 18139
rect 28365 18105 28399 18139
rect 35909 18105 35943 18139
rect 38025 18105 38059 18139
rect 10425 18037 10459 18071
rect 15025 18037 15059 18071
rect 16681 18037 16715 18071
rect 16957 18037 16991 18071
rect 21373 18037 21407 18071
rect 25881 18037 25915 18071
rect 27169 18037 27203 18071
rect 29745 18037 29779 18071
rect 35357 18037 35391 18071
rect 37657 18037 37691 18071
rect 49157 18037 49191 18071
rect 10149 17833 10183 17867
rect 10609 17833 10643 17867
rect 12909 17833 12943 17867
rect 14289 17833 14323 17867
rect 17509 17833 17543 17867
rect 19441 17833 19475 17867
rect 24593 17833 24627 17867
rect 33517 17833 33551 17867
rect 33885 17833 33919 17867
rect 40509 17833 40543 17867
rect 23305 17765 23339 17799
rect 25789 17765 25823 17799
rect 26341 17765 26375 17799
rect 29653 17765 29687 17799
rect 34253 17765 34287 17799
rect 38761 17765 38795 17799
rect 10333 17697 10367 17731
rect 12357 17697 12391 17731
rect 16037 17697 16071 17731
rect 16865 17697 16899 17731
rect 18797 17697 18831 17731
rect 20269 17697 20303 17731
rect 21741 17697 21775 17731
rect 22017 17697 22051 17731
rect 23949 17697 23983 17731
rect 25053 17697 25087 17731
rect 25145 17697 25179 17731
rect 31493 17697 31527 17731
rect 32965 17697 32999 17731
rect 33057 17697 33091 17731
rect 35817 17697 35851 17731
rect 38117 17697 38151 17731
rect 40969 17697 41003 17731
rect 41061 17697 41095 17731
rect 2973 17629 3007 17663
rect 13093 17629 13127 17663
rect 13737 17629 13771 17663
rect 17141 17629 17175 17663
rect 19625 17629 19659 17663
rect 25973 17629 26007 17663
rect 28825 17629 28859 17663
rect 31677 17629 31711 17663
rect 34069 17629 34103 17663
rect 37565 17629 37599 17663
rect 48605 17629 48639 17663
rect 49341 17629 49375 17663
rect 1777 17561 1811 17595
rect 12081 17561 12115 17595
rect 15761 17561 15795 17595
rect 17969 17561 18003 17595
rect 22293 17561 22327 17595
rect 22845 17561 22879 17595
rect 23673 17561 23707 17595
rect 28549 17561 28583 17595
rect 29377 17561 29411 17595
rect 29929 17561 29963 17595
rect 30757 17561 30791 17595
rect 37289 17561 37323 17595
rect 38393 17561 38427 17595
rect 40877 17561 40911 17595
rect 13553 17493 13587 17527
rect 16497 17493 16531 17527
rect 17049 17493 17083 17527
rect 23765 17493 23799 17527
rect 24961 17493 24995 17527
rect 26433 17493 26467 17527
rect 27077 17493 27111 17527
rect 29193 17493 29227 17527
rect 31585 17493 31619 17527
rect 32045 17493 32079 17527
rect 32413 17493 32447 17527
rect 33149 17493 33183 17527
rect 34529 17493 34563 17527
rect 35081 17493 35115 17527
rect 35449 17493 35483 17527
rect 38301 17493 38335 17527
rect 39037 17493 39071 17527
rect 39313 17493 39347 17527
rect 48697 17493 48731 17527
rect 49157 17493 49191 17527
rect 13829 17289 13863 17323
rect 14933 17289 14967 17323
rect 15577 17289 15611 17323
rect 19165 17289 19199 17323
rect 22661 17289 22695 17323
rect 24869 17289 24903 17323
rect 25329 17289 25363 17323
rect 27353 17289 27387 17323
rect 27721 17289 27755 17323
rect 29009 17289 29043 17323
rect 30205 17289 30239 17323
rect 37841 17289 37875 17323
rect 48421 17289 48455 17323
rect 11897 17221 11931 17255
rect 13001 17221 13035 17255
rect 13093 17221 13127 17255
rect 14289 17221 14323 17255
rect 15945 17221 15979 17255
rect 17969 17221 18003 17255
rect 18705 17221 18739 17255
rect 20637 17221 20671 17255
rect 25881 17221 25915 17255
rect 28917 17221 28951 17255
rect 30113 17221 30147 17255
rect 31309 17221 31343 17255
rect 35541 17221 35575 17255
rect 37013 17221 37047 17255
rect 40417 17221 40451 17255
rect 40969 17221 41003 17255
rect 49249 17221 49283 17255
rect 2973 17153 3007 17187
rect 9873 17153 9907 17187
rect 10793 17153 10827 17187
rect 11713 17153 11747 17187
rect 12449 17153 12483 17187
rect 15117 17153 15151 17187
rect 17049 17153 17083 17187
rect 20913 17153 20947 17187
rect 24409 17153 24443 17187
rect 25237 17153 25271 17187
rect 27813 17153 27847 17187
rect 31401 17153 31435 17187
rect 32321 17153 32355 17187
rect 36277 17153 36311 17187
rect 36369 17153 36403 17187
rect 37933 17153 37967 17187
rect 48605 17153 48639 17187
rect 1777 17085 1811 17119
rect 10517 17085 10551 17119
rect 10701 17085 10735 17119
rect 12817 17085 12851 17119
rect 16037 17085 16071 17119
rect 16129 17085 16163 17119
rect 21281 17085 21315 17119
rect 21649 17085 21683 17119
rect 22201 17085 22235 17119
rect 24133 17085 24167 17119
rect 25513 17085 25547 17119
rect 27905 17085 27939 17119
rect 28825 17085 28859 17119
rect 30021 17085 30055 17119
rect 31125 17085 31159 17119
rect 32597 17085 32631 17119
rect 34069 17085 34103 17119
rect 34805 17085 34839 17119
rect 36185 17085 36219 17119
rect 38025 17085 38059 17119
rect 40693 17085 40727 17119
rect 49065 17085 49099 17119
rect 9781 17017 9815 17051
rect 10057 17017 10091 17051
rect 11161 17017 11195 17051
rect 29377 17017 29411 17051
rect 37473 17017 37507 17051
rect 9505 16949 9539 16983
rect 13461 16949 13495 16983
rect 14197 16949 14231 16983
rect 16957 16949 16991 16983
rect 17417 16949 17451 16983
rect 21925 16949 21959 16983
rect 30573 16949 30607 16983
rect 31769 16949 31803 16983
rect 36737 16949 36771 16983
rect 38577 16949 38611 16983
rect 38945 16949 38979 16983
rect 18631 16745 18665 16779
rect 21005 16745 21039 16779
rect 24685 16745 24719 16779
rect 28825 16745 28859 16779
rect 36277 16745 36311 16779
rect 41061 16745 41095 16779
rect 41521 16745 41555 16779
rect 48789 16745 48823 16779
rect 10333 16677 10367 16711
rect 12541 16677 12575 16711
rect 27721 16677 27755 16711
rect 29193 16677 29227 16711
rect 34253 16677 34287 16711
rect 41245 16677 41279 16711
rect 7941 16609 7975 16643
rect 8033 16609 8067 16643
rect 11161 16609 11195 16643
rect 13185 16609 13219 16643
rect 14657 16609 14691 16643
rect 16129 16609 16163 16643
rect 16221 16609 16255 16643
rect 18889 16609 18923 16643
rect 22477 16609 22511 16643
rect 22753 16609 22787 16643
rect 23765 16609 23799 16643
rect 23949 16609 23983 16643
rect 25605 16609 25639 16643
rect 27077 16609 27111 16643
rect 27997 16609 28031 16643
rect 28549 16609 28583 16643
rect 29285 16609 29319 16643
rect 29929 16609 29963 16643
rect 31125 16609 31159 16643
rect 32229 16609 32263 16643
rect 34437 16609 34471 16643
rect 35081 16609 35115 16643
rect 36737 16609 36771 16643
rect 36829 16609 36863 16643
rect 39221 16609 39255 16643
rect 40233 16609 40267 16643
rect 2973 16541 3007 16575
rect 12357 16541 12391 16575
rect 20269 16541 20303 16575
rect 27353 16541 27387 16575
rect 28365 16541 28399 16575
rect 30021 16541 30055 16575
rect 35817 16541 35851 16575
rect 37289 16541 37323 16575
rect 39497 16541 39531 16575
rect 48605 16541 48639 16575
rect 49341 16541 49375 16575
rect 1777 16473 1811 16507
rect 8125 16473 8159 16507
rect 10057 16473 10091 16507
rect 10517 16473 10551 16507
rect 11437 16473 11471 16507
rect 24593 16473 24627 16507
rect 28273 16473 28307 16507
rect 30113 16473 30147 16507
rect 32505 16473 32539 16507
rect 40325 16473 40359 16507
rect 40417 16473 40451 16507
rect 8493 16405 8527 16439
rect 9045 16405 9079 16439
rect 11345 16405 11379 16439
rect 11805 16405 11839 16439
rect 13277 16405 13311 16439
rect 13369 16405 13403 16439
rect 13737 16405 13771 16439
rect 14197 16405 14231 16439
rect 14749 16405 14783 16439
rect 14841 16405 14875 16439
rect 15209 16405 15243 16439
rect 15669 16405 15703 16439
rect 16037 16405 16071 16439
rect 16681 16405 16715 16439
rect 17141 16405 17175 16439
rect 19441 16405 19475 16439
rect 20085 16405 20119 16439
rect 20637 16405 20671 16439
rect 23305 16405 23339 16439
rect 23673 16405 23707 16439
rect 30481 16405 30515 16439
rect 31217 16405 31251 16439
rect 31309 16405 31343 16439
rect 31677 16405 31711 16439
rect 33977 16405 34011 16439
rect 36645 16405 36679 16439
rect 37749 16405 37783 16439
rect 40785 16405 40819 16439
rect 49157 16405 49191 16439
rect 8309 16201 8343 16235
rect 9229 16201 9263 16235
rect 10977 16201 11011 16235
rect 11989 16201 12023 16235
rect 12449 16201 12483 16235
rect 13185 16201 13219 16235
rect 13645 16201 13679 16235
rect 14381 16201 14415 16235
rect 15945 16201 15979 16235
rect 17417 16201 17451 16235
rect 17785 16201 17819 16235
rect 18797 16201 18831 16235
rect 22845 16201 22879 16235
rect 23857 16201 23891 16235
rect 26709 16201 26743 16235
rect 27537 16201 27571 16235
rect 27629 16201 27663 16235
rect 30941 16201 30975 16235
rect 33793 16201 33827 16235
rect 40509 16201 40543 16235
rect 40969 16201 41003 16235
rect 41521 16201 41555 16235
rect 13553 16133 13587 16167
rect 19441 16133 19475 16167
rect 30849 16133 30883 16167
rect 33885 16133 33919 16167
rect 38485 16133 38519 16167
rect 2973 16065 3007 16099
rect 8217 16065 8251 16099
rect 9321 16065 9355 16099
rect 10425 16065 10459 16099
rect 11069 16065 11103 16099
rect 12357 16065 12391 16099
rect 14749 16065 14783 16099
rect 14841 16065 14875 16099
rect 19165 16065 19199 16099
rect 23489 16065 23523 16099
rect 26341 16065 26375 16099
rect 28365 16065 28399 16099
rect 32689 16065 32723 16099
rect 36921 16065 36955 16099
rect 38209 16065 38243 16099
rect 40877 16065 40911 16099
rect 48789 16065 48823 16099
rect 49341 16065 49375 16099
rect 1777 15997 1811 16031
rect 8125 15997 8159 16031
rect 12633 15997 12667 16031
rect 13829 15997 13863 16031
rect 14933 15997 14967 16031
rect 15761 15997 15795 16031
rect 15853 15997 15887 16031
rect 16773 15997 16807 16031
rect 17877 15997 17911 16031
rect 17969 15997 18003 16031
rect 20913 15997 20947 16031
rect 23305 15997 23339 16031
rect 23397 15997 23431 16031
rect 24593 15997 24627 16031
rect 26065 15997 26099 16031
rect 27721 15997 27755 16031
rect 28641 15997 28675 16031
rect 30665 15997 30699 16031
rect 32413 15997 32447 16031
rect 32597 15997 32631 16031
rect 33609 15997 33643 16031
rect 34713 15997 34747 16031
rect 35173 15997 35207 16031
rect 36645 15997 36679 16031
rect 37473 15997 37507 16031
rect 41061 15997 41095 16031
rect 8677 15929 8711 15963
rect 16313 15929 16347 15963
rect 31585 15929 31619 15963
rect 34529 15929 34563 15963
rect 49157 15929 49191 15963
rect 10517 15861 10551 15895
rect 11621 15861 11655 15895
rect 16957 15861 16991 15895
rect 17141 15861 17175 15895
rect 21373 15861 21407 15895
rect 27169 15861 27203 15895
rect 30113 15861 30147 15895
rect 31309 15861 31343 15895
rect 31861 15861 31895 15895
rect 33057 15861 33091 15895
rect 34253 15861 34287 15895
rect 39957 15861 39991 15895
rect 10793 15657 10827 15691
rect 16773 15657 16807 15691
rect 17877 15657 17911 15691
rect 22477 15657 22511 15691
rect 32229 15657 32263 15691
rect 34345 15657 34379 15691
rect 36645 15657 36679 15691
rect 37749 15657 37783 15691
rect 42073 15657 42107 15691
rect 49157 15657 49191 15691
rect 18061 15589 18095 15623
rect 18981 15589 19015 15623
rect 19901 15589 19935 15623
rect 27445 15589 27479 15623
rect 29285 15589 29319 15623
rect 41797 15589 41831 15623
rect 10517 15521 10551 15555
rect 12265 15521 12299 15555
rect 12541 15521 12575 15555
rect 13185 15521 13219 15555
rect 14933 15521 14967 15555
rect 16129 15521 16163 15555
rect 17325 15521 17359 15555
rect 19257 15521 19291 15555
rect 20361 15521 20395 15555
rect 20545 15521 20579 15555
rect 21741 15521 21775 15555
rect 23673 15521 23707 15555
rect 25237 15521 25271 15555
rect 26433 15521 26467 15555
rect 27997 15521 28031 15555
rect 28733 15521 28767 15555
rect 30481 15521 30515 15555
rect 32873 15521 32907 15555
rect 32965 15521 32999 15555
rect 34897 15521 34931 15555
rect 35173 15521 35207 15555
rect 39497 15521 39531 15555
rect 40049 15521 40083 15555
rect 40325 15521 40359 15555
rect 2973 15453 3007 15487
rect 13277 15453 13311 15487
rect 13369 15453 13403 15487
rect 14749 15453 14783 15487
rect 18613 15453 18647 15487
rect 21649 15453 21683 15487
rect 23581 15453 23615 15487
rect 27813 15453 27847 15487
rect 28457 15453 28491 15487
rect 48881 15453 48915 15487
rect 49341 15453 49375 15487
rect 1777 15385 1811 15419
rect 6377 15385 6411 15419
rect 6561 15385 6595 15419
rect 15945 15385 15979 15419
rect 21557 15385 21591 15419
rect 23489 15385 23523 15419
rect 25053 15385 25087 15419
rect 26341 15385 26375 15419
rect 27905 15385 27939 15419
rect 29193 15385 29227 15419
rect 30757 15385 30791 15419
rect 39221 15385 39255 15419
rect 9045 15317 9079 15351
rect 13737 15317 13771 15351
rect 14289 15317 14323 15351
rect 14657 15317 14691 15351
rect 15577 15317 15611 15351
rect 16037 15317 16071 15351
rect 17141 15317 17175 15351
rect 17233 15317 17267 15351
rect 18429 15317 18463 15351
rect 19533 15317 19567 15351
rect 20269 15317 20303 15351
rect 21189 15317 21223 15351
rect 22293 15317 22327 15351
rect 23121 15317 23155 15351
rect 24685 15317 24719 15351
rect 25145 15317 25179 15351
rect 25881 15317 25915 15351
rect 26249 15317 26283 15351
rect 26893 15317 26927 15351
rect 27169 15317 27203 15351
rect 29009 15317 29043 15351
rect 30021 15317 30055 15351
rect 33057 15317 33091 15351
rect 33425 15317 33459 15351
rect 33885 15317 33919 15351
rect 37105 15317 37139 15351
rect 9689 15113 9723 15147
rect 9781 15113 9815 15147
rect 10149 15113 10183 15147
rect 11897 15113 11931 15147
rect 15945 15113 15979 15147
rect 18337 15113 18371 15147
rect 18705 15113 18739 15147
rect 19533 15113 19567 15147
rect 22937 15113 22971 15147
rect 24133 15113 24167 15147
rect 24593 15113 24627 15147
rect 26341 15113 26375 15147
rect 27445 15113 27479 15147
rect 31401 15113 31435 15147
rect 32321 15113 32355 15147
rect 33885 15113 33919 15147
rect 35081 15113 35115 15147
rect 39221 15113 39255 15147
rect 40141 15113 40175 15147
rect 10885 15045 10919 15079
rect 11069 15045 11103 15079
rect 12909 15045 12943 15079
rect 14841 15045 14875 15079
rect 16037 15045 16071 15079
rect 19901 15045 19935 15079
rect 21097 15045 21131 15079
rect 21833 15045 21867 15079
rect 23397 15045 23431 15079
rect 27077 15045 27111 15079
rect 36185 15045 36219 15079
rect 36277 15045 36311 15079
rect 37749 15045 37783 15079
rect 40049 15045 40083 15079
rect 1777 14977 1811 15011
rect 2973 14977 3007 15011
rect 12265 14977 12299 15011
rect 15117 14977 15151 15011
rect 17233 14977 17267 15011
rect 19993 14977 20027 15011
rect 23305 14977 23339 15011
rect 24501 14977 24535 15011
rect 25329 14977 25363 15011
rect 25605 14977 25639 15011
rect 26249 14977 26283 15011
rect 27261 14977 27295 15011
rect 27997 14977 28031 15011
rect 30573 14977 30607 15011
rect 32689 14977 32723 15011
rect 32781 14977 32815 15011
rect 36921 14977 36955 15011
rect 37473 14977 37507 15011
rect 40877 14977 40911 15011
rect 48789 14977 48823 15011
rect 49341 14977 49375 15011
rect 9597 14909 9631 14943
rect 11621 14909 11655 14943
rect 12357 14909 12391 14943
rect 12449 14909 12483 14943
rect 16129 14909 16163 14943
rect 17325 14909 17359 14943
rect 17417 14909 17451 14943
rect 18061 14909 18095 14943
rect 18797 14909 18831 14943
rect 18889 14909 18923 14943
rect 20177 14909 20211 14943
rect 21189 14909 21223 14943
rect 21281 14909 21315 14943
rect 22017 14909 22051 14943
rect 23581 14909 23615 14943
rect 24685 14909 24719 14943
rect 26433 14909 26467 14943
rect 28273 14909 28307 14943
rect 29745 14909 29779 14943
rect 30665 14909 30699 14943
rect 30757 14909 30791 14943
rect 31861 14909 31895 14943
rect 32873 14909 32907 14943
rect 33701 14909 33735 14943
rect 33793 14909 33827 14943
rect 34897 14909 34931 14943
rect 34989 14909 35023 14943
rect 36093 14909 36127 14943
rect 40233 14909 40267 14943
rect 20729 14841 20763 14875
rect 27629 14841 27663 14875
rect 35449 14841 35483 14875
rect 36645 14841 36679 14875
rect 39681 14841 39715 14875
rect 49157 14841 49191 14875
rect 10609 14773 10643 14807
rect 13369 14773 13403 14807
rect 15577 14773 15611 14807
rect 16865 14773 16899 14807
rect 25145 14773 25179 14807
rect 25881 14773 25915 14807
rect 30205 14773 30239 14807
rect 34253 14773 34287 14807
rect 41061 14773 41095 14807
rect 11805 14569 11839 14603
rect 13001 14569 13035 14603
rect 14105 14569 14139 14603
rect 14473 14569 14507 14603
rect 17601 14569 17635 14603
rect 18153 14569 18187 14603
rect 25605 14569 25639 14603
rect 30481 14569 30515 14603
rect 36645 14569 36679 14603
rect 37105 14569 37139 14603
rect 39957 14569 39991 14603
rect 40049 14569 40083 14603
rect 10241 14501 10275 14535
rect 20729 14501 20763 14535
rect 22845 14501 22879 14535
rect 24685 14501 24719 14535
rect 31677 14501 31711 14535
rect 34069 14501 34103 14535
rect 1777 14433 1811 14467
rect 12449 14433 12483 14467
rect 13645 14433 13679 14467
rect 15025 14433 15059 14467
rect 16957 14433 16991 14467
rect 17509 14433 17543 14467
rect 18705 14433 18739 14467
rect 20085 14433 20119 14467
rect 21097 14433 21131 14467
rect 27905 14433 27939 14467
rect 29837 14433 29871 14467
rect 30021 14433 30055 14467
rect 31033 14433 31067 14467
rect 32229 14433 32263 14467
rect 33425 14433 33459 14467
rect 33609 14433 33643 14467
rect 34897 14433 34931 14467
rect 38853 14433 38887 14467
rect 2973 14365 3007 14399
rect 9505 14365 9539 14399
rect 10425 14365 10459 14399
rect 14933 14365 14967 14399
rect 16865 14365 16899 14399
rect 18613 14365 18647 14399
rect 19901 14365 19935 14399
rect 23213 14365 23247 14399
rect 23489 14365 23523 14399
rect 27353 14365 27387 14399
rect 28181 14365 28215 14399
rect 33701 14365 33735 14399
rect 39313 14365 39347 14399
rect 49065 14365 49099 14399
rect 49249 14365 49283 14399
rect 9689 14297 9723 14331
rect 11253 14297 11287 14331
rect 12173 14297 12207 14331
rect 13369 14297 13403 14331
rect 15945 14297 15979 14331
rect 16773 14297 16807 14331
rect 17877 14297 17911 14331
rect 21373 14297 21407 14331
rect 27077 14297 27111 14331
rect 31217 14297 31251 14331
rect 32413 14297 32447 14331
rect 32505 14297 32539 14331
rect 35173 14297 35207 14331
rect 38577 14297 38611 14331
rect 48605 14297 48639 14331
rect 11161 14229 11195 14263
rect 12265 14229 12299 14263
rect 13461 14229 13495 14263
rect 14841 14229 14875 14263
rect 16405 14229 16439 14263
rect 18521 14229 18555 14263
rect 19533 14229 19567 14263
rect 19993 14229 20027 14263
rect 20545 14229 20579 14263
rect 23857 14229 23891 14263
rect 24409 14229 24443 14263
rect 25145 14229 25179 14263
rect 28089 14229 28123 14263
rect 28549 14229 28583 14263
rect 29009 14229 29043 14263
rect 30113 14229 30147 14263
rect 31309 14229 31343 14263
rect 32873 14229 32907 14263
rect 34345 14229 34379 14263
rect 39497 14229 39531 14263
rect 48697 14229 48731 14263
rect 3617 14025 3651 14059
rect 9965 14025 9999 14059
rect 10425 14025 10459 14059
rect 11989 14025 12023 14059
rect 15577 14025 15611 14059
rect 15945 14025 15979 14059
rect 17141 14025 17175 14059
rect 17509 14025 17543 14059
rect 17601 14025 17635 14059
rect 18337 14025 18371 14059
rect 18705 14025 18739 14059
rect 19441 14025 19475 14059
rect 21465 14025 21499 14059
rect 24869 14025 24903 14059
rect 27629 14025 27663 14059
rect 29377 14025 29411 14059
rect 31769 14025 31803 14059
rect 36093 14025 36127 14059
rect 36461 14025 36495 14059
rect 37841 14025 37875 14059
rect 38209 14025 38243 14059
rect 45845 14025 45879 14059
rect 48421 14025 48455 14059
rect 49157 14025 49191 14059
rect 1777 13957 1811 13991
rect 10701 13957 10735 13991
rect 13277 13957 13311 13991
rect 15025 13957 15059 13991
rect 15301 13957 15335 13991
rect 16037 13957 16071 13991
rect 26341 13957 26375 13991
rect 34897 13957 34931 13991
rect 37749 13957 37783 13991
rect 38577 13957 38611 13991
rect 38945 13957 38979 13991
rect 45017 13957 45051 13991
rect 48145 13957 48179 13991
rect 49249 13957 49283 13991
rect 2973 13889 3007 13923
rect 3525 13889 3559 13923
rect 3985 13889 4019 13923
rect 11161 13889 11195 13923
rect 12081 13889 12115 13923
rect 16865 13889 16899 13923
rect 18797 13889 18831 13923
rect 28917 13889 28951 13923
rect 31125 13889 31159 13923
rect 34805 13889 34839 13923
rect 36921 13889 36955 13923
rect 45661 13889 45695 13923
rect 48605 13889 48639 13923
rect 11897 13821 11931 13855
rect 13001 13821 13035 13855
rect 14749 13821 14783 13855
rect 16221 13821 16255 13855
rect 17785 13821 17819 13855
rect 18889 13821 18923 13855
rect 19717 13821 19751 13855
rect 22017 13821 22051 13855
rect 23489 13821 23523 13855
rect 23765 13821 23799 13855
rect 24225 13821 24259 13855
rect 26617 13821 26651 13855
rect 30849 13821 30883 13855
rect 32321 13821 32355 13855
rect 34069 13821 34103 13855
rect 34621 13821 34655 13855
rect 35909 13821 35943 13855
rect 36001 13821 36035 13855
rect 37657 13821 37691 13855
rect 45201 13821 45235 13855
rect 12449 13753 12483 13787
rect 35265 13753 35299 13787
rect 19980 13685 20014 13719
rect 33811 13685 33845 13719
rect 36737 13685 36771 13719
rect 12541 13481 12575 13515
rect 13737 13481 13771 13515
rect 14933 13481 14967 13515
rect 18153 13481 18187 13515
rect 20453 13481 20487 13515
rect 20913 13481 20947 13515
rect 22109 13481 22143 13515
rect 24041 13481 24075 13515
rect 25605 13481 25639 13515
rect 26709 13481 26743 13515
rect 27445 13481 27479 13515
rect 27813 13481 27847 13515
rect 28181 13481 28215 13515
rect 29193 13481 29227 13515
rect 35633 13481 35667 13515
rect 38209 13481 38243 13515
rect 38577 13481 38611 13515
rect 39589 13481 39623 13515
rect 10517 13413 10551 13447
rect 14289 13413 14323 13447
rect 31125 13413 31159 13447
rect 33333 13413 33367 13447
rect 36093 13413 36127 13447
rect 1777 13345 1811 13379
rect 10793 13345 10827 13379
rect 13093 13345 13127 13379
rect 13921 13345 13955 13379
rect 15393 13345 15427 13379
rect 15485 13345 15519 13379
rect 16405 13345 16439 13379
rect 19901 13345 19935 13379
rect 21465 13345 21499 13379
rect 22753 13345 22787 13379
rect 23489 13345 23523 13379
rect 23581 13345 23615 13379
rect 25053 13345 25087 13379
rect 28641 13345 28675 13379
rect 29837 13345 29871 13379
rect 30021 13345 30055 13379
rect 33885 13345 33919 13379
rect 34345 13345 34379 13379
rect 35081 13345 35115 13379
rect 2973 13277 3007 13311
rect 14473 13277 14507 13311
rect 24501 13277 24535 13311
rect 25237 13277 25271 13311
rect 28825 13277 28859 13311
rect 30113 13277 30147 13311
rect 32873 13277 32907 13311
rect 36461 13277 36495 13311
rect 41337 13277 41371 13311
rect 47961 13277 47995 13311
rect 49157 13277 49191 13311
rect 11069 13209 11103 13243
rect 16681 13209 16715 13243
rect 18889 13209 18923 13243
rect 20085 13209 20119 13243
rect 21373 13209 21407 13243
rect 22477 13209 22511 13243
rect 26065 13209 26099 13243
rect 27721 13209 27755 13243
rect 32597 13209 32631 13243
rect 33701 13209 33735 13243
rect 35173 13209 35207 13243
rect 35265 13209 35299 13243
rect 36737 13209 36771 13243
rect 15577 13141 15611 13175
rect 15945 13141 15979 13175
rect 19349 13141 19383 13175
rect 19993 13141 20027 13175
rect 21281 13141 21315 13175
rect 22569 13141 22603 13175
rect 23673 13141 23707 13175
rect 25145 13141 25179 13175
rect 28733 13141 28767 13175
rect 30481 13141 30515 13175
rect 33793 13141 33827 13175
rect 35909 13141 35943 13175
rect 41521 13141 41555 13175
rect 3065 12937 3099 12971
rect 10977 12937 11011 12971
rect 11161 12937 11195 12971
rect 11989 12937 12023 12971
rect 12725 12937 12759 12971
rect 13093 12937 13127 12971
rect 15301 12937 15335 12971
rect 15853 12937 15887 12971
rect 19257 12937 19291 12971
rect 22937 12937 22971 12971
rect 23397 12937 23431 12971
rect 26065 12937 26099 12971
rect 26249 12937 26283 12971
rect 26709 12937 26743 12971
rect 31769 12937 31803 12971
rect 33425 12937 33459 12971
rect 36461 12937 36495 12971
rect 1685 12869 1719 12903
rect 2145 12869 2179 12903
rect 15945 12869 15979 12903
rect 18705 12869 18739 12903
rect 25329 12869 25363 12903
rect 29653 12869 29687 12903
rect 30297 12869 30331 12903
rect 32689 12869 32723 12903
rect 34805 12869 34839 12903
rect 35725 12869 35759 12903
rect 37105 12869 37139 12903
rect 2881 12801 2915 12835
rect 3341 12801 3375 12835
rect 12081 12801 12115 12835
rect 17877 12801 17911 12835
rect 19625 12801 19659 12835
rect 21097 12801 21131 12835
rect 23029 12801 23063 12835
rect 25605 12801 25639 12835
rect 26433 12801 26467 12835
rect 27169 12801 27203 12835
rect 29193 12801 29227 12835
rect 30021 12801 30055 12835
rect 34069 12801 34103 12835
rect 35817 12801 35851 12835
rect 36737 12801 36771 12835
rect 37473 12801 37507 12835
rect 40049 12801 40083 12835
rect 40509 12801 40543 12835
rect 45937 12801 45971 12835
rect 47961 12801 47995 12835
rect 49157 12801 49191 12835
rect 1869 12733 1903 12767
rect 11805 12733 11839 12767
rect 14565 12733 14599 12767
rect 14841 12733 14875 12767
rect 15761 12733 15795 12767
rect 17417 12733 17451 12767
rect 19717 12733 19751 12767
rect 19901 12733 19935 12767
rect 21189 12733 21223 12767
rect 21281 12733 21315 12767
rect 22017 12733 22051 12767
rect 22753 12733 22787 12767
rect 23857 12733 23891 12767
rect 28917 12733 28951 12767
rect 32413 12733 32447 12767
rect 32597 12733 32631 12767
rect 35633 12733 35667 12767
rect 37749 12733 37783 12767
rect 39497 12733 39531 12767
rect 16313 12665 16347 12699
rect 20729 12665 20763 12699
rect 33057 12665 33091 12699
rect 36185 12665 36219 12699
rect 40233 12665 40267 12699
rect 11253 12597 11287 12631
rect 12449 12597 12483 12631
rect 16773 12597 16807 12631
rect 16865 12597 16899 12631
rect 20453 12597 20487 12631
rect 25973 12597 26007 12631
rect 33517 12597 33551 12631
rect 33701 12597 33735 12631
rect 36921 12597 36955 12631
rect 46121 12597 46155 12631
rect 11253 12393 11287 12427
rect 14381 12393 14415 12427
rect 16405 12393 16439 12427
rect 21649 12393 21683 12427
rect 23305 12393 23339 12427
rect 27721 12393 27755 12427
rect 35160 12393 35194 12427
rect 36645 12393 36679 12427
rect 39313 12393 39347 12427
rect 26341 12325 26375 12359
rect 39037 12325 39071 12359
rect 40325 12325 40359 12359
rect 2421 12257 2455 12291
rect 2697 12257 2731 12291
rect 9505 12257 9539 12291
rect 11713 12257 11747 12291
rect 13737 12257 13771 12291
rect 16129 12257 16163 12291
rect 17417 12257 17451 12291
rect 19993 12257 20027 12291
rect 20637 12257 20671 12291
rect 21005 12257 21039 12291
rect 21189 12257 21223 12291
rect 22293 12257 22327 12291
rect 23765 12257 23799 12291
rect 23949 12257 23983 12291
rect 24869 12257 24903 12291
rect 27169 12257 27203 12291
rect 28365 12257 28399 12291
rect 29745 12257 29779 12291
rect 31769 12257 31803 12291
rect 33885 12257 33919 12291
rect 37197 12257 37231 12291
rect 38393 12257 38427 12291
rect 38577 12257 38611 12291
rect 49157 12257 49191 12291
rect 2145 12189 2179 12223
rect 17141 12189 17175 12223
rect 19809 12189 19843 12223
rect 21281 12189 21315 12223
rect 24593 12189 24627 12223
rect 27261 12189 27295 12223
rect 29193 12189 29227 12223
rect 32137 12189 32171 12223
rect 34897 12189 34931 12223
rect 37381 12189 37415 12223
rect 40785 12189 40819 12223
rect 41429 12189 41463 12223
rect 45937 12189 45971 12223
rect 47961 12189 47995 12223
rect 9781 12121 9815 12155
rect 11989 12121 12023 12155
rect 15853 12121 15887 12155
rect 18153 12121 18187 12155
rect 18889 12121 18923 12155
rect 22477 12121 22511 12155
rect 23673 12121 23707 12155
rect 26709 12121 26743 12155
rect 30021 12121 30055 12155
rect 32413 12121 32447 12155
rect 39497 12121 39531 12155
rect 40141 12121 40175 12155
rect 16773 12053 16807 12087
rect 17233 12053 17267 12087
rect 19441 12053 19475 12087
rect 19901 12053 19935 12087
rect 22385 12053 22419 12087
rect 22845 12053 22879 12087
rect 27353 12053 27387 12087
rect 31493 12053 31527 12087
rect 34161 12053 34195 12087
rect 34345 12053 34379 12087
rect 37473 12053 37507 12087
rect 37841 12053 37875 12087
rect 38669 12053 38703 12087
rect 40969 12053 41003 12087
rect 41613 12053 41647 12087
rect 46121 12053 46155 12087
rect 11529 11849 11563 11883
rect 11989 11849 12023 11883
rect 14197 11849 14231 11883
rect 14289 11849 14323 11883
rect 19257 11849 19291 11883
rect 20269 11849 20303 11883
rect 20729 11849 20763 11883
rect 21189 11849 21223 11883
rect 21833 11849 21867 11883
rect 22109 11849 22143 11883
rect 26617 11849 26651 11883
rect 27537 11849 27571 11883
rect 27905 11849 27939 11883
rect 31493 11849 31527 11883
rect 32597 11849 32631 11883
rect 32689 11849 32723 11883
rect 33885 11849 33919 11883
rect 34713 11849 34747 11883
rect 37749 11849 37783 11883
rect 38669 11849 38703 11883
rect 40417 11849 40451 11883
rect 19073 11781 19107 11815
rect 19809 11781 19843 11815
rect 21097 11781 21131 11815
rect 30021 11781 30055 11815
rect 31769 11781 31803 11815
rect 39129 11781 39163 11815
rect 45109 11781 45143 11815
rect 49157 11781 49191 11815
rect 1593 11713 1627 11747
rect 2329 11713 2363 11747
rect 12725 11713 12759 11747
rect 12817 11713 12851 11747
rect 15485 11713 15519 11747
rect 16405 11713 16439 11747
rect 19901 11713 19935 11747
rect 22569 11713 22603 11747
rect 23397 11713 23431 11747
rect 23949 11713 23983 11747
rect 26157 11713 26191 11747
rect 31125 11713 31159 11747
rect 33793 11713 33827 11747
rect 37841 11713 37875 11747
rect 39037 11713 39071 11747
rect 39957 11713 39991 11747
rect 40601 11713 40635 11747
rect 47961 11713 47995 11747
rect 2789 11645 2823 11679
rect 12909 11645 12943 11679
rect 13645 11645 13679 11679
rect 14013 11645 14047 11679
rect 15577 11645 15611 11679
rect 15669 11645 15703 11679
rect 18337 11645 18371 11679
rect 18613 11645 18647 11679
rect 19625 11645 19659 11679
rect 21373 11645 21407 11679
rect 24225 11645 24259 11679
rect 27261 11645 27295 11679
rect 27445 11645 27479 11679
rect 28549 11645 28583 11679
rect 30297 11645 30331 11679
rect 30849 11645 30883 11679
rect 31033 11645 31067 11679
rect 32505 11645 32539 11679
rect 33609 11645 33643 11679
rect 35173 11645 35207 11679
rect 35449 11645 35483 11679
rect 37565 11645 37599 11679
rect 39221 11645 39255 11679
rect 1777 11577 1811 11611
rect 14657 11577 14691 11611
rect 16865 11577 16899 11611
rect 33057 11577 33091 11611
rect 34253 11577 34287 11611
rect 36921 11577 36955 11611
rect 40141 11577 40175 11611
rect 45293 11577 45327 11611
rect 2513 11509 2547 11543
rect 12357 11509 12391 11543
rect 13369 11509 13403 11543
rect 15117 11509 15151 11543
rect 16313 11509 16347 11543
rect 22293 11509 22327 11543
rect 25697 11509 25731 11543
rect 34621 11509 34655 11543
rect 38209 11509 38243 11543
rect 2145 11305 2179 11339
rect 14381 11305 14415 11339
rect 16773 11305 16807 11339
rect 17969 11305 18003 11339
rect 19073 11305 19107 11339
rect 19349 11305 19383 11339
rect 23305 11305 23339 11339
rect 26341 11305 26375 11339
rect 29009 11305 29043 11339
rect 34713 11305 34747 11339
rect 38761 11305 38795 11339
rect 39589 11305 39623 11339
rect 1777 11237 1811 11271
rect 19533 11237 19567 11271
rect 28641 11237 28675 11271
rect 30481 11237 30515 11271
rect 38393 11237 38427 11271
rect 40969 11237 41003 11271
rect 10977 11169 11011 11203
rect 12449 11169 12483 11203
rect 14841 11169 14875 11203
rect 15025 11169 15059 11203
rect 15761 11169 15795 11203
rect 15853 11169 15887 11203
rect 17417 11169 17451 11203
rect 18613 11169 18647 11203
rect 19993 11169 20027 11203
rect 20453 11169 20487 11203
rect 21925 11169 21959 11203
rect 23949 11169 23983 11203
rect 24869 11169 24903 11203
rect 27169 11169 27203 11203
rect 29929 11169 29963 11203
rect 32873 11169 32907 11203
rect 37749 11169 37783 11203
rect 49157 11169 49191 11203
rect 1593 11101 1627 11135
rect 2329 11101 2363 11135
rect 12725 11101 12759 11135
rect 17233 11101 17267 11135
rect 22201 11101 22235 11135
rect 24593 11101 24627 11135
rect 26893 11101 26927 11135
rect 31125 11101 31159 11135
rect 33333 11101 33367 11135
rect 38209 11101 38243 11135
rect 40141 11101 40175 11135
rect 40785 11101 40819 11135
rect 45661 11101 45695 11135
rect 47961 11101 47995 11135
rect 13001 11033 13035 11067
rect 13277 11033 13311 11067
rect 13737 11033 13771 11067
rect 15945 11033 15979 11067
rect 17141 11033 17175 11067
rect 23673 11033 23707 11067
rect 31401 11033 31435 11067
rect 34069 11033 34103 11067
rect 35725 11033 35759 11067
rect 37473 11033 37507 11067
rect 40325 11033 40359 11067
rect 45845 11033 45879 11067
rect 14749 10965 14783 10999
rect 16313 10965 16347 10999
rect 18337 10965 18371 10999
rect 18429 10965 18463 10999
rect 22661 10965 22695 10999
rect 23765 10965 23799 10999
rect 29193 10965 29227 10999
rect 29285 10965 29319 10999
rect 30021 10965 30055 10999
rect 30113 10965 30147 10999
rect 30757 10965 30791 10999
rect 2513 10761 2547 10795
rect 12449 10761 12483 10795
rect 13185 10761 13219 10795
rect 14381 10761 14415 10795
rect 15577 10761 15611 10795
rect 15945 10761 15979 10795
rect 17141 10761 17175 10795
rect 19533 10761 19567 10795
rect 21097 10761 21131 10795
rect 24225 10761 24259 10795
rect 25881 10761 25915 10795
rect 26433 10761 26467 10795
rect 26801 10761 26835 10795
rect 28549 10761 28583 10795
rect 31401 10761 31435 10795
rect 33057 10761 33091 10795
rect 36829 10761 36863 10795
rect 37289 10761 37323 10795
rect 37473 10761 37507 10795
rect 17509 10693 17543 10727
rect 19993 10693 20027 10727
rect 21189 10693 21223 10727
rect 27445 10693 27479 10727
rect 28825 10693 28859 10727
rect 35357 10693 35391 10727
rect 49157 10693 49191 10727
rect 1593 10625 1627 10659
rect 2329 10625 2363 10659
rect 2881 10625 2915 10659
rect 13553 10625 13587 10659
rect 14749 10625 14783 10659
rect 14841 10625 14875 10659
rect 16865 10625 16899 10659
rect 18705 10625 18739 10659
rect 19901 10625 19935 10659
rect 24593 10625 24627 10659
rect 25421 10625 25455 10659
rect 26065 10625 26099 10659
rect 27537 10625 27571 10659
rect 30573 10625 30607 10659
rect 32689 10625 32723 10659
rect 33333 10625 33367 10659
rect 35633 10625 35667 10659
rect 36461 10625 36495 10659
rect 39773 10625 39807 10659
rect 40233 10625 40267 10659
rect 47961 10625 47995 10659
rect 3065 10557 3099 10591
rect 12725 10557 12759 10591
rect 13645 10557 13679 10591
rect 13829 10557 13863 10591
rect 14933 10557 14967 10591
rect 16037 10557 16071 10591
rect 16129 10557 16163 10591
rect 17601 10557 17635 10591
rect 17693 10557 17727 10591
rect 18797 10557 18831 10591
rect 18889 10557 18923 10591
rect 20177 10557 20211 10591
rect 21373 10557 21407 10591
rect 22017 10557 22051 10591
rect 22293 10557 22327 10591
rect 24685 10557 24719 10591
rect 24869 10557 24903 10591
rect 27353 10557 27387 10591
rect 29561 10557 29595 10591
rect 30389 10557 30423 10591
rect 30481 10557 30515 10591
rect 32413 10557 32447 10591
rect 32597 10557 32631 10591
rect 33885 10557 33919 10591
rect 36185 10557 36219 10591
rect 36369 10557 36403 10591
rect 1777 10489 1811 10523
rect 23765 10489 23799 10523
rect 26249 10489 26283 10523
rect 27905 10489 27939 10523
rect 39957 10489 39991 10523
rect 12265 10421 12299 10455
rect 12817 10421 12851 10455
rect 18337 10421 18371 10455
rect 20729 10421 20763 10455
rect 30941 10421 30975 10455
rect 31953 10421 31987 10455
rect 13461 10217 13495 10251
rect 18153 10217 18187 10251
rect 20269 10217 20303 10251
rect 23765 10217 23799 10251
rect 24593 10217 24627 10251
rect 26709 10217 26743 10251
rect 28733 10217 28767 10251
rect 30389 10217 30423 10251
rect 36645 10217 36679 10251
rect 36921 10217 36955 10251
rect 13921 10149 13955 10183
rect 16589 10149 16623 10183
rect 23949 10149 23983 10183
rect 2145 10081 2179 10115
rect 12909 10081 12943 10115
rect 13001 10081 13035 10115
rect 16405 10081 16439 10115
rect 17417 10081 17451 10115
rect 17601 10081 17635 10115
rect 18613 10081 18647 10115
rect 18797 10081 18831 10115
rect 19717 10081 19751 10115
rect 21741 10081 21775 10115
rect 26065 10081 26099 10115
rect 26341 10081 26375 10115
rect 26985 10081 27019 10115
rect 29377 10081 29411 10115
rect 29929 10081 29963 10115
rect 32137 10081 32171 10115
rect 32781 10081 32815 10115
rect 35173 10081 35207 10115
rect 38485 10081 38519 10115
rect 49157 10081 49191 10115
rect 2421 10013 2455 10047
rect 16037 10013 16071 10047
rect 22017 10013 22051 10047
rect 23305 10013 23339 10047
rect 32873 10013 32907 10047
rect 34897 10013 34931 10047
rect 38301 10013 38335 10047
rect 38761 10013 38795 10047
rect 40141 10013 40175 10047
rect 40601 10013 40635 10047
rect 44373 10013 44407 10047
rect 46121 10013 46155 10047
rect 47961 10013 47995 10047
rect 15761 9945 15795 9979
rect 22477 9945 22511 9979
rect 27261 9945 27295 9979
rect 29101 9945 29135 9979
rect 31861 9945 31895 9979
rect 33793 9945 33827 9979
rect 40325 9945 40359 9979
rect 44557 9945 44591 9979
rect 47317 9945 47351 9979
rect 12449 9877 12483 9911
rect 13093 9877 13127 9911
rect 14289 9877 14323 9911
rect 16957 9877 16991 9911
rect 17325 9877 17359 9911
rect 18521 9877 18555 9911
rect 24133 9877 24167 9911
rect 32965 9877 32999 9911
rect 33333 9877 33367 9911
rect 2145 9673 2179 9707
rect 21097 9673 21131 9707
rect 22293 9673 22327 9707
rect 32965 9673 32999 9707
rect 35633 9673 35667 9707
rect 36093 9673 36127 9707
rect 13369 9605 13403 9639
rect 15853 9605 15887 9639
rect 16037 9605 16071 9639
rect 16313 9605 16347 9639
rect 19625 9605 19659 9639
rect 21373 9605 21407 9639
rect 29009 9605 29043 9639
rect 31861 9605 31895 9639
rect 49157 9605 49191 9639
rect 1593 9537 1627 9571
rect 2329 9537 2363 9571
rect 12541 9537 12575 9571
rect 22661 9537 22695 9571
rect 22753 9537 22787 9571
rect 25237 9537 25271 9571
rect 26065 9537 26099 9571
rect 32873 9537 32907 9571
rect 33885 9537 33919 9571
rect 47961 9537 47995 9571
rect 12265 9469 12299 9503
rect 12449 9469 12483 9503
rect 15117 9469 15151 9503
rect 15393 9469 15427 9503
rect 16865 9469 16899 9503
rect 18613 9469 18647 9503
rect 18889 9469 18923 9503
rect 19349 9469 19383 9503
rect 22937 9469 22971 9503
rect 24961 9469 24995 9503
rect 25881 9469 25915 9503
rect 25973 9469 26007 9503
rect 29285 9469 29319 9503
rect 29745 9469 29779 9503
rect 30021 9469 30055 9503
rect 31493 9469 31527 9503
rect 32689 9469 32723 9503
rect 34161 9469 34195 9503
rect 35909 9469 35943 9503
rect 1777 9401 1811 9435
rect 12909 9401 12943 9435
rect 21649 9401 21683 9435
rect 26433 9401 26467 9435
rect 27537 9401 27571 9435
rect 15669 9333 15703 9367
rect 16405 9333 16439 9367
rect 21833 9333 21867 9367
rect 23489 9333 23523 9367
rect 32229 9333 32263 9367
rect 33333 9333 33367 9367
rect 17889 9129 17923 9163
rect 19441 9129 19475 9163
rect 22293 9129 22327 9163
rect 24409 9129 24443 9163
rect 28917 9129 28951 9163
rect 34069 9129 34103 9163
rect 36737 9129 36771 9163
rect 1869 9061 1903 9095
rect 14473 9061 14507 9095
rect 30757 9061 30791 9095
rect 34345 9061 34379 9095
rect 37841 9061 37875 9095
rect 2881 8993 2915 9027
rect 15301 8993 15335 9027
rect 15485 8993 15519 9027
rect 18153 8993 18187 9027
rect 20913 8993 20947 9027
rect 23765 8993 23799 9027
rect 28365 8993 28399 9027
rect 32229 8993 32263 9027
rect 32505 8993 32539 9027
rect 33425 8993 33459 9027
rect 34989 8993 35023 9027
rect 39865 8993 39899 9027
rect 49157 8993 49191 9027
rect 2329 8925 2363 8959
rect 3065 8925 3099 8959
rect 14289 8925 14323 8959
rect 15577 8925 15611 8959
rect 18705 8925 18739 8959
rect 21189 8925 21223 8959
rect 24041 8925 24075 8959
rect 25605 8925 25639 8959
rect 35173 8925 35207 8959
rect 36553 8925 36587 8959
rect 37657 8925 37691 8959
rect 39313 8925 39347 8959
rect 39497 8925 39531 8959
rect 47961 8925 47995 8959
rect 1685 8857 1719 8891
rect 28549 8857 28583 8891
rect 29745 8857 29779 8891
rect 2513 8789 2547 8823
rect 14933 8789 14967 8823
rect 15945 8789 15979 8823
rect 16405 8789 16439 8823
rect 21833 8789 21867 8823
rect 24593 8789 24627 8823
rect 24777 8789 24811 8823
rect 25329 8789 25363 8823
rect 25697 8789 25731 8823
rect 27813 8789 27847 8823
rect 28457 8789 28491 8823
rect 30297 8789 30331 8823
rect 32873 8789 32907 8823
rect 33057 8789 33091 8823
rect 33609 8789 33643 8823
rect 33701 8789 33735 8823
rect 35265 8789 35299 8823
rect 35633 8789 35667 8823
rect 18613 8585 18647 8619
rect 19717 8585 19751 8619
rect 22017 8585 22051 8619
rect 24041 8585 24075 8619
rect 31769 8585 31803 8619
rect 34069 8585 34103 8619
rect 37657 8585 37691 8619
rect 13921 8517 13955 8551
rect 17141 8517 17175 8551
rect 21189 8517 21223 8551
rect 29101 8517 29135 8551
rect 31309 8517 31343 8551
rect 34805 8517 34839 8551
rect 40325 8517 40359 8551
rect 40785 8517 40819 8551
rect 44189 8517 44223 8551
rect 49157 8517 49191 8551
rect 2145 8449 2179 8483
rect 16865 8449 16899 8483
rect 23765 8449 23799 8483
rect 31401 8449 31435 8483
rect 32321 8449 32355 8483
rect 37473 8449 37507 8483
rect 38945 8449 38979 8483
rect 40509 8449 40543 8483
rect 45845 8449 45879 8483
rect 47961 8449 47995 8483
rect 2421 8381 2455 8415
rect 13645 8381 13679 8415
rect 15393 8381 15427 8415
rect 19073 8381 19107 8415
rect 21465 8381 21499 8415
rect 23489 8381 23523 8415
rect 28825 8381 28859 8415
rect 31217 8381 31251 8415
rect 32597 8381 32631 8415
rect 44373 8381 44407 8415
rect 46857 8381 46891 8415
rect 15761 8313 15795 8347
rect 16221 8313 16255 8347
rect 30573 8313 30607 8347
rect 34345 8313 34379 8347
rect 34621 8313 34655 8347
rect 39129 8313 39163 8347
rect 2145 8041 2179 8075
rect 18981 8041 19015 8075
rect 19441 8041 19475 8075
rect 22017 8041 22051 8075
rect 30389 8041 30423 8075
rect 31769 8041 31803 8075
rect 15761 7973 15795 8007
rect 33057 7973 33091 8007
rect 16773 7905 16807 7939
rect 16957 7905 16991 7939
rect 18061 7905 18095 7939
rect 20913 7905 20947 7939
rect 22569 7905 22603 7939
rect 29929 7905 29963 7939
rect 31217 7905 31251 7939
rect 32505 7905 32539 7939
rect 33425 7905 33459 7939
rect 49157 7905 49191 7939
rect 1593 7837 1627 7871
rect 2329 7837 2363 7871
rect 15577 7837 15611 7871
rect 17049 7837 17083 7871
rect 18153 7837 18187 7871
rect 21189 7837 21223 7871
rect 22385 7837 22419 7871
rect 31309 7837 31343 7871
rect 32689 7837 32723 7871
rect 38761 7837 38795 7871
rect 39221 7837 39255 7871
rect 47961 7837 47995 7871
rect 18245 7769 18279 7803
rect 30481 7769 30515 7803
rect 37565 7769 37599 7803
rect 38025 7769 38059 7803
rect 38945 7769 38979 7803
rect 1777 7701 1811 7735
rect 17417 7701 17451 7735
rect 18613 7701 18647 7735
rect 21465 7701 21499 7735
rect 21649 7701 21683 7735
rect 22477 7701 22511 7735
rect 23029 7701 23063 7735
rect 30665 7701 30699 7735
rect 31401 7701 31435 7735
rect 32597 7701 32631 7735
rect 38117 7701 38151 7735
rect 22017 7497 22051 7531
rect 22477 7497 22511 7531
rect 23029 7497 23063 7531
rect 31125 7497 31159 7531
rect 32321 7497 32355 7531
rect 39037 7497 39071 7531
rect 18337 7429 18371 7463
rect 18797 7429 18831 7463
rect 19073 7429 19107 7463
rect 31953 7429 31987 7463
rect 38577 7429 38611 7463
rect 49157 7429 49191 7463
rect 1593 7361 1627 7395
rect 2145 7361 2179 7395
rect 22385 7361 22419 7395
rect 37841 7361 37875 7395
rect 44925 7361 44959 7395
rect 47961 7361 47995 7395
rect 22569 7293 22603 7327
rect 1777 7225 1811 7259
rect 37381 7225 37415 7259
rect 38761 7225 38795 7259
rect 45109 7225 45143 7259
rect 21189 7157 21223 7191
rect 21373 7157 21407 7191
rect 21649 7157 21683 7191
rect 32873 7157 32907 7191
rect 37933 7157 37967 7191
rect 21833 6817 21867 6851
rect 49157 6817 49191 6851
rect 2329 6749 2363 6783
rect 2789 6749 2823 6783
rect 17693 6749 17727 6783
rect 19625 6749 19659 6783
rect 46121 6749 46155 6783
rect 47961 6749 47995 6783
rect 1685 6681 1719 6715
rect 47317 6681 47351 6715
rect 1777 6613 1811 6647
rect 2513 6613 2547 6647
rect 17877 6613 17911 6647
rect 19809 6613 19843 6647
rect 2145 6409 2179 6443
rect 37565 6341 37599 6375
rect 38025 6341 38059 6375
rect 44005 6341 44039 6375
rect 49157 6341 49191 6375
rect 1593 6273 1627 6307
rect 2329 6273 2363 6307
rect 18061 6273 18095 6307
rect 47961 6273 47995 6307
rect 18245 6205 18279 6239
rect 1777 6137 1811 6171
rect 44189 6137 44223 6171
rect 18705 6069 18739 6103
rect 37657 6069 37691 6103
rect 2513 5797 2547 5831
rect 3065 5729 3099 5763
rect 49157 5729 49191 5763
rect 1593 5661 1627 5695
rect 2329 5661 2363 5695
rect 2881 5661 2915 5695
rect 43729 5661 43763 5695
rect 47961 5661 47995 5695
rect 43913 5593 43947 5627
rect 1777 5525 1811 5559
rect 37381 5253 37415 5287
rect 37749 5253 37783 5287
rect 38485 5253 38519 5287
rect 38945 5253 38979 5287
rect 49157 5253 49191 5287
rect 2145 5185 2179 5219
rect 18889 5185 18923 5219
rect 45845 5185 45879 5219
rect 47961 5185 47995 5219
rect 2421 5117 2455 5151
rect 19073 5117 19107 5151
rect 46857 5117 46891 5151
rect 38669 5049 38703 5083
rect 19533 4981 19567 5015
rect 37841 4981 37875 5015
rect 2145 4777 2179 4811
rect 1777 4709 1811 4743
rect 22569 4709 22603 4743
rect 46489 4709 46523 4743
rect 20453 4641 20487 4675
rect 21925 4641 21959 4675
rect 26801 4641 26835 4675
rect 36829 4641 36863 4675
rect 47225 4641 47259 4675
rect 49157 4641 49191 4675
rect 1593 4573 1627 4607
rect 2329 4573 2363 4607
rect 20637 4573 20671 4607
rect 22109 4573 22143 4607
rect 23096 4573 23130 4607
rect 26985 4573 27019 4607
rect 37289 4573 37323 4607
rect 47961 4573 47995 4607
rect 25145 4505 25179 4539
rect 38025 4505 38059 4539
rect 38485 4505 38519 4539
rect 46673 4505 46707 4539
rect 47409 4505 47443 4539
rect 21097 4437 21131 4471
rect 23167 4437 23201 4471
rect 37381 4437 37415 4471
rect 38117 4437 38151 4471
rect 46213 4437 46247 4471
rect 2513 4233 2547 4267
rect 1685 4165 1719 4199
rect 25881 4165 25915 4199
rect 2329 4097 2363 4131
rect 22360 4096 22394 4130
rect 22972 4097 23006 4131
rect 23075 4097 23109 4131
rect 23616 4097 23650 4131
rect 26065 4097 26099 4131
rect 45845 4097 45879 4131
rect 47961 4097 47995 4131
rect 49157 4097 49191 4131
rect 3065 4029 3099 4063
rect 24869 4029 24903 4063
rect 27169 4029 27203 4063
rect 28825 4029 28859 4063
rect 29009 4029 29043 4063
rect 46673 4029 46707 4063
rect 1869 3961 1903 3995
rect 23719 3961 23753 3995
rect 2881 3893 2915 3927
rect 22431 3893 22465 3927
rect 47685 3893 47719 3927
rect 23029 3689 23063 3723
rect 23581 3689 23615 3723
rect 23949 3689 23983 3723
rect 45385 3621 45419 3655
rect 2145 3553 2179 3587
rect 26249 3553 26283 3587
rect 26433 3553 26467 3587
rect 49157 3553 49191 3587
rect 2421 3485 2455 3519
rect 16589 3485 16623 3519
rect 21005 3485 21039 3519
rect 23305 3485 23339 3519
rect 24041 3485 24075 3519
rect 46121 3485 46155 3519
rect 47961 3485 47995 3519
rect 16405 3417 16439 3451
rect 21281 3417 21315 3451
rect 24593 3417 24627 3451
rect 36461 3417 36495 3451
rect 36645 3417 36679 3451
rect 45109 3417 45143 3451
rect 45569 3417 45603 3451
rect 47317 3417 47351 3451
rect 22753 3349 22787 3383
rect 36921 3349 36955 3383
rect 2145 3145 2179 3179
rect 9873 3145 9907 3179
rect 16313 3145 16347 3179
rect 19993 3145 20027 3179
rect 21465 3145 21499 3179
rect 28365 3145 28399 3179
rect 16773 3077 16807 3111
rect 49157 3077 49191 3111
rect 1593 3009 1627 3043
rect 2513 3009 2547 3043
rect 9689 3009 9723 3043
rect 12357 3009 12391 3043
rect 14565 3009 14599 3043
rect 17601 3009 17635 3043
rect 19533 3009 19567 3043
rect 20177 3009 20211 3043
rect 20637 3009 20671 3043
rect 21281 3009 21315 3043
rect 22661 3009 22695 3043
rect 23029 3009 23063 3043
rect 23765 3009 23799 3043
rect 26433 3009 26467 3043
rect 27997 3009 28031 3043
rect 28917 3009 28951 3043
rect 44005 3009 44039 3043
rect 45845 3009 45879 3043
rect 47961 3009 47995 3043
rect 13001 2941 13035 2975
rect 14841 2941 14875 2975
rect 18337 2941 18371 2975
rect 24225 2941 24259 2975
rect 24501 2941 24535 2975
rect 25973 2941 26007 2975
rect 29193 2941 29227 2975
rect 31033 2941 31067 2975
rect 45201 2941 45235 2975
rect 46857 2941 46891 2975
rect 1777 2873 1811 2907
rect 20821 2873 20855 2907
rect 22201 2873 22235 2907
rect 27537 2873 27571 2907
rect 2329 2805 2363 2839
rect 2789 2805 2823 2839
rect 17417 2805 17451 2839
rect 22385 2805 22419 2839
rect 23305 2805 23339 2839
rect 23489 2805 23523 2839
rect 26617 2805 26651 2839
rect 27905 2805 27939 2839
rect 30665 2805 30699 2839
rect 2513 2601 2547 2635
rect 24041 2601 24075 2635
rect 26341 2601 26375 2635
rect 29009 2601 29043 2635
rect 35081 2601 35115 2635
rect 1777 2533 1811 2567
rect 3249 2533 3283 2567
rect 10333 2533 10367 2567
rect 30849 2533 30883 2567
rect 32965 2533 32999 2567
rect 20545 2465 20579 2499
rect 22845 2465 22879 2499
rect 25053 2465 25087 2499
rect 27629 2465 27663 2499
rect 37749 2465 37783 2499
rect 41429 2465 41463 2499
rect 43821 2465 43855 2499
rect 49157 2465 49191 2499
rect 1593 2397 1627 2431
rect 3065 2397 3099 2431
rect 3525 2397 3559 2431
rect 9689 2397 9723 2431
rect 13185 2397 13219 2431
rect 15669 2397 15703 2431
rect 18245 2397 18279 2431
rect 18889 2397 18923 2431
rect 19441 2397 19475 2431
rect 20085 2397 20119 2431
rect 22385 2397 22419 2431
rect 24593 2397 24627 2431
rect 27169 2397 27203 2431
rect 29193 2397 29227 2431
rect 29561 2397 29595 2431
rect 31033 2397 31067 2431
rect 31309 2397 31343 2431
rect 33149 2397 33183 2431
rect 33425 2397 33459 2431
rect 35265 2397 35299 2431
rect 35541 2397 35575 2431
rect 37473 2397 37507 2431
rect 40693 2397 40727 2431
rect 43545 2397 43579 2431
rect 45845 2397 45879 2431
rect 47961 2397 47995 2431
rect 2421 2329 2455 2363
rect 11989 2329 12023 2363
rect 14473 2329 14507 2363
rect 17049 2329 17083 2363
rect 47041 2329 47075 2363
rect 9413 2261 9447 2295
rect 18705 2261 18739 2295
rect 19625 2261 19659 2295
rect 37105 2261 37139 2295
rect 43269 2261 43303 2295
<< metal1 >>
rect 30558 25236 30564 25288
rect 30616 25276 30622 25288
rect 37918 25276 37924 25288
rect 30616 25248 37924 25276
rect 30616 25236 30622 25248
rect 37918 25236 37924 25248
rect 37976 25236 37982 25288
rect 3418 24828 3424 24880
rect 3476 24868 3482 24880
rect 9766 24868 9772 24880
rect 3476 24840 9772 24868
rect 3476 24828 3482 24840
rect 9766 24828 9772 24840
rect 9824 24828 9830 24880
rect 33318 24868 33324 24880
rect 32968 24840 33324 24868
rect 3602 24760 3608 24812
rect 3660 24800 3666 24812
rect 5902 24800 5908 24812
rect 3660 24772 5908 24800
rect 3660 24760 3666 24772
rect 5902 24760 5908 24772
rect 5960 24760 5966 24812
rect 17218 24760 17224 24812
rect 17276 24800 17282 24812
rect 24026 24800 24032 24812
rect 17276 24772 24032 24800
rect 17276 24760 17282 24772
rect 24026 24760 24032 24772
rect 24084 24760 24090 24812
rect 24762 24760 24768 24812
rect 24820 24800 24826 24812
rect 30374 24800 30380 24812
rect 24820 24772 30380 24800
rect 24820 24760 24826 24772
rect 30374 24760 30380 24772
rect 30432 24760 30438 24812
rect 18874 24692 18880 24744
rect 18932 24732 18938 24744
rect 27246 24732 27252 24744
rect 18932 24704 27252 24732
rect 18932 24692 18938 24704
rect 27246 24692 27252 24704
rect 27304 24692 27310 24744
rect 29914 24692 29920 24744
rect 29972 24732 29978 24744
rect 32968 24732 32996 24840
rect 33318 24828 33324 24840
rect 33376 24828 33382 24880
rect 39574 24828 39580 24880
rect 39632 24868 39638 24880
rect 45278 24868 45284 24880
rect 39632 24840 45284 24868
rect 39632 24828 39638 24840
rect 45278 24828 45284 24840
rect 45336 24828 45342 24880
rect 38930 24760 38936 24812
rect 38988 24800 38994 24812
rect 42058 24800 42064 24812
rect 38988 24772 42064 24800
rect 38988 24760 38994 24772
rect 42058 24760 42064 24772
rect 42116 24760 42122 24812
rect 34606 24732 34612 24744
rect 29972 24704 32996 24732
rect 33060 24704 34612 24732
rect 29972 24692 29978 24704
rect 22554 24624 22560 24676
rect 22612 24664 22618 24676
rect 26326 24664 26332 24676
rect 22612 24636 26332 24664
rect 22612 24624 22618 24636
rect 26326 24624 26332 24636
rect 26384 24624 26390 24676
rect 26418 24624 26424 24676
rect 26476 24664 26482 24676
rect 33060 24664 33088 24704
rect 34606 24692 34612 24704
rect 34664 24692 34670 24744
rect 34882 24692 34888 24744
rect 34940 24732 34946 24744
rect 40310 24732 40316 24744
rect 34940 24704 40316 24732
rect 34940 24692 34946 24704
rect 40310 24692 40316 24704
rect 40368 24692 40374 24744
rect 26476 24636 33088 24664
rect 26476 24624 26482 24636
rect 33134 24624 33140 24676
rect 33192 24664 33198 24676
rect 39942 24664 39948 24676
rect 33192 24636 39948 24664
rect 33192 24624 33198 24636
rect 39942 24624 39948 24636
rect 40000 24624 40006 24676
rect 40218 24624 40224 24676
rect 40276 24664 40282 24676
rect 43990 24664 43996 24676
rect 40276 24636 43996 24664
rect 40276 24624 40282 24636
rect 43990 24624 43996 24636
rect 44048 24624 44054 24676
rect 20530 24556 20536 24608
rect 20588 24596 20594 24608
rect 29730 24596 29736 24608
rect 20588 24568 29736 24596
rect 20588 24556 20594 24568
rect 29730 24556 29736 24568
rect 29788 24556 29794 24608
rect 29822 24556 29828 24608
rect 29880 24596 29886 24608
rect 31570 24596 31576 24608
rect 29880 24568 31576 24596
rect 29880 24556 29886 24568
rect 31570 24556 31576 24568
rect 31628 24556 31634 24608
rect 31846 24556 31852 24608
rect 31904 24596 31910 24608
rect 39482 24596 39488 24608
rect 31904 24568 39488 24596
rect 31904 24556 31910 24568
rect 39482 24556 39488 24568
rect 39540 24556 39546 24608
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 9582 24392 9588 24404
rect 6886 24364 9588 24392
rect 2961 24259 3019 24265
rect 2961 24225 2973 24259
rect 3007 24256 3019 24259
rect 3510 24256 3516 24268
rect 3007 24228 3516 24256
rect 3007 24225 3019 24228
rect 2961 24219 3019 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 5813 24259 5871 24265
rect 5813 24225 5825 24259
rect 5859 24256 5871 24259
rect 6730 24256 6736 24268
rect 5859 24228 6736 24256
rect 5859 24225 5871 24228
rect 5813 24219 5871 24225
rect 6730 24216 6736 24228
rect 6788 24216 6794 24268
rect 3421 24191 3479 24197
rect 3421 24157 3433 24191
rect 3467 24188 3479 24191
rect 3878 24188 3884 24200
rect 3467 24160 3884 24188
rect 3467 24157 3479 24160
rect 3421 24151 3479 24157
rect 3878 24148 3884 24160
rect 3936 24148 3942 24200
rect 3973 24191 4031 24197
rect 3973 24157 3985 24191
rect 4019 24157 4031 24191
rect 3973 24151 4031 24157
rect 3988 24120 4016 24151
rect 4614 24148 4620 24200
rect 4672 24148 4678 24200
rect 6549 24191 6607 24197
rect 6549 24157 6561 24191
rect 6595 24188 6607 24191
rect 6886 24188 6914 24364
rect 9582 24352 9588 24364
rect 9640 24352 9646 24404
rect 12342 24352 12348 24404
rect 12400 24392 12406 24404
rect 17218 24392 17224 24404
rect 12400 24364 17224 24392
rect 12400 24352 12406 24364
rect 17218 24352 17224 24364
rect 17276 24352 17282 24404
rect 18598 24352 18604 24404
rect 18656 24392 18662 24404
rect 18656 24364 25176 24392
rect 18656 24352 18662 24364
rect 11882 24324 11888 24336
rect 10704 24296 11888 24324
rect 8205 24259 8263 24265
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 8662 24256 8668 24268
rect 8251 24228 8668 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 8662 24216 8668 24228
rect 8720 24216 8726 24268
rect 10704 24265 10732 24296
rect 11882 24284 11888 24296
rect 11940 24284 11946 24336
rect 15470 24324 15476 24336
rect 12406 24296 15476 24324
rect 10689 24259 10747 24265
rect 10689 24225 10701 24259
rect 10735 24225 10747 24259
rect 12406 24256 12434 24296
rect 15470 24284 15476 24296
rect 15528 24284 15534 24336
rect 16022 24284 16028 24336
rect 16080 24324 16086 24336
rect 19610 24324 19616 24336
rect 16080 24296 17816 24324
rect 16080 24284 16086 24296
rect 10689 24219 10747 24225
rect 11072 24228 12434 24256
rect 13265 24259 13323 24265
rect 6595 24160 6914 24188
rect 6595 24157 6607 24160
rect 6549 24151 6607 24157
rect 7190 24148 7196 24200
rect 7248 24188 7254 24200
rect 7377 24191 7435 24197
rect 7377 24188 7389 24191
rect 7248 24160 7389 24188
rect 7248 24148 7254 24160
rect 7377 24157 7389 24160
rect 7423 24188 7435 24191
rect 7926 24188 7932 24200
rect 7423 24160 7932 24188
rect 7423 24157 7435 24160
rect 7377 24151 7435 24157
rect 7926 24148 7932 24160
rect 7984 24148 7990 24200
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24188 9367 24191
rect 11072 24188 11100 24228
rect 13265 24225 13277 24259
rect 13311 24256 13323 24259
rect 13814 24256 13820 24268
rect 13311 24228 13820 24256
rect 13311 24225 13323 24228
rect 13265 24219 13323 24225
rect 13814 24216 13820 24228
rect 13872 24216 13878 24268
rect 15841 24259 15899 24265
rect 15841 24225 15853 24259
rect 15887 24256 15899 24259
rect 17678 24256 17684 24268
rect 15887 24228 17684 24256
rect 15887 24225 15899 24228
rect 15841 24219 15899 24225
rect 17678 24216 17684 24228
rect 17736 24216 17742 24268
rect 9355 24160 11100 24188
rect 11149 24191 11207 24197
rect 9355 24157 9367 24160
rect 9309 24151 9367 24157
rect 11149 24157 11161 24191
rect 11195 24157 11207 24191
rect 11149 24151 11207 24157
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24188 11943 24191
rect 13725 24191 13783 24197
rect 11931 24160 13676 24188
rect 11931 24157 11943 24160
rect 11885 24151 11943 24157
rect 10134 24120 10140 24132
rect 3988 24092 10140 24120
rect 10134 24080 10140 24092
rect 10192 24080 10198 24132
rect 11164 24120 11192 24151
rect 12618 24120 12624 24132
rect 11164 24092 12624 24120
rect 12618 24080 12624 24092
rect 12676 24080 12682 24132
rect 13648 24120 13676 24160
rect 13725 24157 13737 24191
rect 13771 24188 13783 24191
rect 14274 24188 14280 24200
rect 13771 24160 14280 24188
rect 13771 24157 13783 24160
rect 13725 24151 13783 24157
rect 14274 24148 14280 24160
rect 14332 24148 14338 24200
rect 14458 24148 14464 24200
rect 14516 24148 14522 24200
rect 16301 24191 16359 24197
rect 16301 24157 16313 24191
rect 16347 24157 16359 24191
rect 17788 24188 17816 24296
rect 18432 24296 19616 24324
rect 18432 24265 18460 24296
rect 19610 24284 19616 24296
rect 19668 24284 19674 24336
rect 20254 24284 20260 24336
rect 20312 24324 20318 24336
rect 24581 24327 24639 24333
rect 20312 24296 22508 24324
rect 20312 24284 20318 24296
rect 18417 24259 18475 24265
rect 18417 24225 18429 24259
rect 18463 24225 18475 24259
rect 18417 24219 18475 24225
rect 18524 24228 20760 24256
rect 18524 24188 18552 24228
rect 17788 24160 18552 24188
rect 16301 24151 16359 24157
rect 14918 24120 14924 24132
rect 13648 24092 14924 24120
rect 14918 24080 14924 24092
rect 14976 24080 14982 24132
rect 16316 24120 16344 24151
rect 18874 24148 18880 24200
rect 18932 24148 18938 24200
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24188 19671 24191
rect 20530 24188 20536 24200
rect 19659 24160 20536 24188
rect 19659 24157 19671 24160
rect 19613 24151 19671 24157
rect 20530 24148 20536 24160
rect 20588 24148 20594 24200
rect 20622 24120 20628 24132
rect 16316 24092 20628 24120
rect 20622 24080 20628 24092
rect 20680 24080 20686 24132
rect 20732 24120 20760 24228
rect 20898 24216 20904 24268
rect 20956 24216 20962 24268
rect 22370 24256 22376 24268
rect 21376 24228 22376 24256
rect 21376 24197 21404 24228
rect 22370 24216 22376 24228
rect 22428 24216 22434 24268
rect 22480 24265 22508 24296
rect 24581 24293 24593 24327
rect 24627 24293 24639 24327
rect 24581 24287 24639 24293
rect 22465 24259 22523 24265
rect 22465 24225 22477 24259
rect 22511 24225 22523 24259
rect 24596 24256 24624 24287
rect 25148 24265 25176 24364
rect 26418 24352 26424 24404
rect 26476 24352 26482 24404
rect 27246 24352 27252 24404
rect 27304 24352 27310 24404
rect 29730 24352 29736 24404
rect 29788 24352 29794 24404
rect 30374 24352 30380 24404
rect 30432 24392 30438 24404
rect 31481 24395 31539 24401
rect 31481 24392 31493 24395
rect 30432 24364 31493 24392
rect 30432 24352 30438 24364
rect 31481 24361 31493 24364
rect 31527 24361 31539 24395
rect 31481 24355 31539 24361
rect 37292 24364 37964 24392
rect 25774 24284 25780 24336
rect 25832 24284 25838 24336
rect 22465 24219 22523 24225
rect 22848 24228 24624 24256
rect 25133 24259 25191 24265
rect 21361 24191 21419 24197
rect 21361 24157 21373 24191
rect 21407 24157 21419 24191
rect 21361 24151 21419 24157
rect 21450 24148 21456 24200
rect 21508 24188 21514 24200
rect 22005 24191 22063 24197
rect 22005 24188 22017 24191
rect 21508 24160 22017 24188
rect 21508 24148 21514 24160
rect 22005 24157 22017 24160
rect 22051 24157 22063 24191
rect 22005 24151 22063 24157
rect 22848 24120 22876 24228
rect 25133 24225 25145 24259
rect 25179 24225 25191 24259
rect 26436 24256 26464 24352
rect 28626 24284 28632 24336
rect 28684 24324 28690 24336
rect 31665 24327 31723 24333
rect 31665 24324 31677 24327
rect 28684 24296 31677 24324
rect 28684 24284 28690 24296
rect 25133 24219 25191 24225
rect 25976 24228 26464 24256
rect 23845 24191 23903 24197
rect 23845 24157 23857 24191
rect 23891 24188 23903 24191
rect 25406 24188 25412 24200
rect 23891 24160 25412 24188
rect 23891 24157 23903 24160
rect 23845 24151 23903 24157
rect 25406 24148 25412 24160
rect 25464 24148 25470 24200
rect 25976 24197 26004 24228
rect 27338 24216 27344 24268
rect 27396 24256 27402 24268
rect 29181 24259 29239 24265
rect 29181 24256 29193 24259
rect 27396 24228 29193 24256
rect 27396 24216 27402 24228
rect 25961 24191 26019 24197
rect 25961 24157 25973 24191
rect 26007 24157 26019 24191
rect 25961 24151 26019 24157
rect 26234 24148 26240 24200
rect 26292 24188 26298 24200
rect 28552 24197 28580 24228
rect 29181 24225 29193 24228
rect 29227 24225 29239 24259
rect 29181 24219 29239 24225
rect 27893 24191 27951 24197
rect 27893 24188 27905 24191
rect 26292 24160 27905 24188
rect 26292 24148 26298 24160
rect 27893 24157 27905 24160
rect 27939 24157 27951 24191
rect 27893 24151 27951 24157
rect 28537 24191 28595 24197
rect 28537 24157 28549 24191
rect 28583 24157 28595 24191
rect 28537 24151 28595 24157
rect 29917 24191 29975 24197
rect 29917 24157 29929 24191
rect 29963 24157 29975 24191
rect 29917 24151 29975 24157
rect 20732 24092 22876 24120
rect 24949 24123 25007 24129
rect 24949 24089 24961 24123
rect 24995 24120 25007 24123
rect 25314 24120 25320 24132
rect 24995 24092 25320 24120
rect 24995 24089 25007 24092
rect 24949 24083 25007 24089
rect 25314 24080 25320 24092
rect 25372 24080 25378 24132
rect 26602 24120 26608 24132
rect 26252 24092 26608 24120
rect 4157 24055 4215 24061
rect 4157 24021 4169 24055
rect 4203 24052 4215 24055
rect 5534 24052 5540 24064
rect 4203 24024 5540 24052
rect 4203 24021 4215 24024
rect 4157 24015 4215 24021
rect 5534 24012 5540 24024
rect 5592 24012 5598 24064
rect 6733 24055 6791 24061
rect 6733 24021 6745 24055
rect 6779 24052 6791 24055
rect 7466 24052 7472 24064
rect 6779 24024 7472 24052
rect 6779 24021 6791 24024
rect 6733 24015 6791 24021
rect 7466 24012 7472 24024
rect 7524 24012 7530 24064
rect 9122 24012 9128 24064
rect 9180 24012 9186 24064
rect 11146 24012 11152 24064
rect 11204 24052 11210 24064
rect 11701 24055 11759 24061
rect 11701 24052 11713 24055
rect 11204 24024 11713 24052
rect 11204 24012 11210 24024
rect 11701 24021 11713 24024
rect 11747 24021 11759 24055
rect 11701 24015 11759 24021
rect 11790 24012 11796 24064
rect 11848 24052 11854 24064
rect 14277 24055 14335 24061
rect 14277 24052 14289 24055
rect 11848 24024 14289 24052
rect 11848 24012 11854 24024
rect 14277 24021 14289 24024
rect 14323 24021 14335 24055
rect 14277 24015 14335 24021
rect 17037 24055 17095 24061
rect 17037 24021 17049 24055
rect 17083 24052 17095 24055
rect 18414 24052 18420 24064
rect 17083 24024 18420 24052
rect 17083 24021 17095 24024
rect 17037 24015 17095 24021
rect 18414 24012 18420 24024
rect 18472 24012 18478 24064
rect 19426 24012 19432 24064
rect 19484 24012 19490 24064
rect 20254 24012 20260 24064
rect 20312 24052 20318 24064
rect 23842 24052 23848 24064
rect 20312 24024 23848 24052
rect 20312 24012 20318 24024
rect 23842 24012 23848 24024
rect 23900 24012 23906 24064
rect 24029 24055 24087 24061
rect 24029 24021 24041 24055
rect 24075 24052 24087 24055
rect 24670 24052 24676 24064
rect 24075 24024 24676 24052
rect 24075 24021 24087 24024
rect 24029 24015 24087 24021
rect 24670 24012 24676 24024
rect 24728 24012 24734 24064
rect 25041 24055 25099 24061
rect 25041 24021 25053 24055
rect 25087 24052 25099 24055
rect 26252 24052 26280 24092
rect 26602 24080 26608 24092
rect 26660 24080 26666 24132
rect 26789 24123 26847 24129
rect 26789 24089 26801 24123
rect 26835 24120 26847 24123
rect 27246 24120 27252 24132
rect 26835 24092 27252 24120
rect 26835 24089 26847 24092
rect 26789 24083 26847 24089
rect 27246 24080 27252 24092
rect 27304 24080 27310 24132
rect 27338 24080 27344 24132
rect 27396 24080 27402 24132
rect 27908 24120 27936 24151
rect 28997 24123 29055 24129
rect 28997 24120 29009 24123
rect 27908 24092 29009 24120
rect 28997 24089 29009 24092
rect 29043 24089 29055 24123
rect 29932 24120 29960 24151
rect 30374 24148 30380 24200
rect 30432 24148 30438 24200
rect 30944 24188 30972 24296
rect 31665 24293 31677 24296
rect 31711 24293 31723 24327
rect 31665 24287 31723 24293
rect 32953 24327 33011 24333
rect 32953 24293 32965 24327
rect 32999 24293 33011 24327
rect 32953 24287 33011 24293
rect 31110 24216 31116 24268
rect 31168 24256 31174 24268
rect 32968 24256 32996 24287
rect 33502 24284 33508 24336
rect 33560 24324 33566 24336
rect 37292 24324 37320 24364
rect 33560 24296 37320 24324
rect 33560 24284 33566 24296
rect 35084 24265 35112 24296
rect 31168 24228 32996 24256
rect 34241 24259 34299 24265
rect 31168 24216 31174 24228
rect 34241 24225 34253 24259
rect 34287 24225 34299 24259
rect 34241 24219 34299 24225
rect 35069 24259 35127 24265
rect 35069 24225 35081 24259
rect 35115 24225 35127 24259
rect 35069 24219 35127 24225
rect 31021 24191 31079 24197
rect 31021 24188 31033 24191
rect 30944 24160 31033 24188
rect 31021 24157 31033 24160
rect 31067 24157 31079 24191
rect 31021 24151 31079 24157
rect 31570 24148 31576 24200
rect 31628 24188 31634 24200
rect 32493 24191 32551 24197
rect 32493 24188 32505 24191
rect 31628 24160 32505 24188
rect 31628 24148 31634 24160
rect 32493 24157 32505 24160
rect 32539 24157 32551 24191
rect 32493 24151 32551 24157
rect 33137 24191 33195 24197
rect 33137 24157 33149 24191
rect 33183 24188 33195 24191
rect 33318 24188 33324 24200
rect 33183 24160 33324 24188
rect 33183 24157 33195 24160
rect 33137 24151 33195 24157
rect 33318 24148 33324 24160
rect 33376 24148 33382 24200
rect 34256 24188 34284 24219
rect 36722 24216 36728 24268
rect 36780 24216 36786 24268
rect 37274 24216 37280 24268
rect 37332 24256 37338 24268
rect 37553 24259 37611 24265
rect 37553 24256 37565 24259
rect 37332 24228 37565 24256
rect 37332 24216 37338 24228
rect 37553 24225 37565 24228
rect 37599 24225 37611 24259
rect 37826 24256 37832 24268
rect 37553 24219 37611 24225
rect 37660 24228 37832 24256
rect 36354 24188 36360 24200
rect 34256 24160 36360 24188
rect 36354 24148 36360 24160
rect 36412 24148 36418 24200
rect 36541 24191 36599 24197
rect 36541 24157 36553 24191
rect 36587 24188 36599 24191
rect 37660 24188 37688 24228
rect 37826 24216 37832 24228
rect 37884 24216 37890 24268
rect 37936 24256 37964 24364
rect 38654 24352 38660 24404
rect 38712 24352 38718 24404
rect 39298 24352 39304 24404
rect 39356 24352 39362 24404
rect 39850 24352 39856 24404
rect 39908 24392 39914 24404
rect 41049 24395 41107 24401
rect 41049 24392 41061 24395
rect 39908 24364 41061 24392
rect 39908 24352 39914 24364
rect 41049 24361 41061 24364
rect 41095 24392 41107 24395
rect 42242 24392 42248 24404
rect 41095 24364 42248 24392
rect 41095 24361 41107 24364
rect 41049 24355 41107 24361
rect 42242 24352 42248 24364
rect 42300 24352 42306 24404
rect 42610 24352 42616 24404
rect 42668 24392 42674 24404
rect 43717 24395 43775 24401
rect 43717 24392 43729 24395
rect 42668 24364 43729 24392
rect 42668 24352 42674 24364
rect 43717 24361 43729 24364
rect 43763 24361 43775 24395
rect 43717 24355 43775 24361
rect 43898 24352 43904 24404
rect 43956 24392 43962 24404
rect 44361 24395 44419 24401
rect 44361 24392 44373 24395
rect 43956 24364 44373 24392
rect 43956 24352 43962 24364
rect 44361 24361 44373 24364
rect 44407 24361 44419 24395
rect 44361 24355 44419 24361
rect 38197 24327 38255 24333
rect 38197 24293 38209 24327
rect 38243 24324 38255 24327
rect 39758 24324 39764 24336
rect 38243 24296 39764 24324
rect 38243 24293 38255 24296
rect 38197 24287 38255 24293
rect 39758 24284 39764 24296
rect 39816 24284 39822 24336
rect 42518 24284 42524 24336
rect 42576 24324 42582 24336
rect 46661 24327 46719 24333
rect 46661 24324 46673 24327
rect 42576 24296 46673 24324
rect 42576 24284 42582 24296
rect 46661 24293 46673 24296
rect 46707 24293 46719 24327
rect 46661 24287 46719 24293
rect 40589 24259 40647 24265
rect 40589 24256 40601 24259
rect 37936 24228 40601 24256
rect 40589 24225 40601 24228
rect 40635 24225 40647 24259
rect 40589 24219 40647 24225
rect 41417 24259 41475 24265
rect 41417 24225 41429 24259
rect 41463 24256 41475 24259
rect 45370 24256 45376 24268
rect 41463 24228 45376 24256
rect 41463 24225 41475 24228
rect 41417 24219 41475 24225
rect 45370 24216 45376 24228
rect 45428 24216 45434 24268
rect 47486 24216 47492 24268
rect 47544 24256 47550 24268
rect 48222 24256 48228 24268
rect 47544 24228 48228 24256
rect 47544 24216 47550 24228
rect 48222 24216 48228 24228
rect 48280 24256 48286 24268
rect 48501 24259 48559 24265
rect 48501 24256 48513 24259
rect 48280 24228 48513 24256
rect 48280 24216 48286 24228
rect 48501 24225 48513 24228
rect 48547 24225 48559 24259
rect 48501 24219 48559 24225
rect 36587 24160 37688 24188
rect 36587 24157 36599 24160
rect 36541 24151 36599 24157
rect 37734 24148 37740 24200
rect 37792 24148 37798 24200
rect 37918 24148 37924 24200
rect 37976 24188 37982 24200
rect 38841 24191 38899 24197
rect 38841 24188 38853 24191
rect 37976 24160 38853 24188
rect 37976 24148 37982 24160
rect 38841 24157 38853 24160
rect 38887 24157 38899 24191
rect 38841 24151 38899 24157
rect 33965 24123 34023 24129
rect 29932 24092 33640 24120
rect 28997 24083 29055 24089
rect 25087 24024 26280 24052
rect 25087 24021 25099 24024
rect 25041 24015 25099 24021
rect 26970 24012 26976 24064
rect 27028 24052 27034 24064
rect 27798 24052 27804 24064
rect 27028 24024 27804 24052
rect 27028 24012 27034 24024
rect 27798 24012 27804 24024
rect 27856 24012 27862 24064
rect 28077 24055 28135 24061
rect 28077 24021 28089 24055
rect 28123 24052 28135 24055
rect 28534 24052 28540 24064
rect 28123 24024 28540 24052
rect 28123 24021 28135 24024
rect 28077 24015 28135 24021
rect 28534 24012 28540 24024
rect 28592 24012 28598 24064
rect 28718 24012 28724 24064
rect 28776 24012 28782 24064
rect 30558 24012 30564 24064
rect 30616 24012 30622 24064
rect 30926 24012 30932 24064
rect 30984 24052 30990 24064
rect 31205 24055 31263 24061
rect 31205 24052 31217 24055
rect 30984 24024 31217 24052
rect 30984 24012 30990 24024
rect 31205 24021 31217 24024
rect 31251 24021 31263 24055
rect 31205 24015 31263 24021
rect 31941 24055 31999 24061
rect 31941 24021 31953 24055
rect 31987 24052 31999 24055
rect 32122 24052 32128 24064
rect 31987 24024 32128 24052
rect 31987 24021 31999 24024
rect 31941 24015 31999 24021
rect 32122 24012 32128 24024
rect 32180 24012 32186 24064
rect 32306 24012 32312 24064
rect 32364 24012 32370 24064
rect 33612 24061 33640 24092
rect 33965 24089 33977 24123
rect 34011 24120 34023 24123
rect 34146 24120 34152 24132
rect 34011 24092 34152 24120
rect 34011 24089 34023 24092
rect 33965 24083 34023 24089
rect 34146 24080 34152 24092
rect 34204 24080 34210 24132
rect 34606 24080 34612 24132
rect 34664 24120 34670 24132
rect 35158 24120 35164 24132
rect 34664 24092 35164 24120
rect 34664 24080 34670 24092
rect 35158 24080 35164 24092
rect 35216 24080 35222 24132
rect 36449 24123 36507 24129
rect 36449 24089 36461 24123
rect 36495 24120 36507 24123
rect 36814 24120 36820 24132
rect 36495 24092 36820 24120
rect 36495 24089 36507 24092
rect 36449 24083 36507 24089
rect 36814 24080 36820 24092
rect 36872 24080 36878 24132
rect 37752 24120 37780 24148
rect 37829 24123 37887 24129
rect 37829 24120 37841 24123
rect 37752 24092 37841 24120
rect 37829 24089 37841 24092
rect 37875 24089 37887 24123
rect 37829 24083 37887 24089
rect 38102 24080 38108 24132
rect 38160 24120 38166 24132
rect 38856 24120 38884 24151
rect 39482 24148 39488 24200
rect 39540 24188 39546 24200
rect 40126 24188 40132 24200
rect 39540 24160 40132 24188
rect 39540 24148 39546 24160
rect 40126 24148 40132 24160
rect 40184 24148 40190 24200
rect 40405 24191 40463 24197
rect 40405 24157 40417 24191
rect 40451 24188 40463 24191
rect 42061 24191 42119 24197
rect 40451 24160 42012 24188
rect 40451 24157 40463 24160
rect 40405 24151 40463 24157
rect 39666 24120 39672 24132
rect 38160 24092 38792 24120
rect 38856 24092 39672 24120
rect 38160 24080 38166 24092
rect 33597 24055 33655 24061
rect 33597 24021 33609 24055
rect 33643 24021 33655 24055
rect 33597 24015 33655 24021
rect 34054 24012 34060 24064
rect 34112 24012 34118 24064
rect 34790 24012 34796 24064
rect 34848 24052 34854 24064
rect 35250 24052 35256 24064
rect 34848 24024 35256 24052
rect 34848 24012 34854 24024
rect 35250 24012 35256 24024
rect 35308 24012 35314 24064
rect 35618 24012 35624 24064
rect 35676 24012 35682 24064
rect 36078 24012 36084 24064
rect 36136 24012 36142 24064
rect 37734 24012 37740 24064
rect 37792 24052 37798 24064
rect 38654 24052 38660 24064
rect 37792 24024 38660 24052
rect 37792 24012 37798 24024
rect 38654 24012 38660 24024
rect 38712 24012 38718 24064
rect 38764 24052 38792 24092
rect 39666 24080 39672 24092
rect 39724 24080 39730 24132
rect 40497 24123 40555 24129
rect 40497 24089 40509 24123
rect 40543 24120 40555 24123
rect 41138 24120 41144 24132
rect 40543 24092 41144 24120
rect 40543 24089 40555 24092
rect 40497 24083 40555 24089
rect 41138 24080 41144 24092
rect 41196 24080 41202 24132
rect 41984 24120 42012 24160
rect 42061 24157 42073 24191
rect 42107 24188 42119 24191
rect 42613 24191 42671 24197
rect 42613 24188 42625 24191
rect 42107 24160 42625 24188
rect 42107 24157 42119 24160
rect 42061 24151 42119 24157
rect 42613 24157 42625 24160
rect 42659 24157 42671 24191
rect 42613 24151 42671 24157
rect 42794 24148 42800 24200
rect 42852 24188 42858 24200
rect 43257 24191 43315 24197
rect 43257 24188 43269 24191
rect 42852 24160 43269 24188
rect 42852 24148 42858 24160
rect 43257 24157 43269 24160
rect 43303 24188 43315 24191
rect 43806 24188 43812 24200
rect 43303 24160 43812 24188
rect 43303 24157 43315 24160
rect 43257 24151 43315 24157
rect 43806 24148 43812 24160
rect 43864 24148 43870 24200
rect 43898 24148 43904 24200
rect 43956 24148 43962 24200
rect 44450 24148 44456 24200
rect 44508 24188 44514 24200
rect 44545 24191 44603 24197
rect 44545 24188 44557 24191
rect 44508 24160 44557 24188
rect 44508 24148 44514 24160
rect 44545 24157 44557 24160
rect 44591 24157 44603 24191
rect 44545 24151 44603 24157
rect 45554 24148 45560 24200
rect 45612 24188 45618 24200
rect 46198 24188 46204 24200
rect 45612 24160 46204 24188
rect 45612 24148 45618 24160
rect 46198 24148 46204 24160
rect 46256 24148 46262 24200
rect 46290 24148 46296 24200
rect 46348 24188 46354 24200
rect 46845 24191 46903 24197
rect 46845 24188 46857 24191
rect 46348 24160 46857 24188
rect 46348 24148 46354 24160
rect 46845 24157 46857 24160
rect 46891 24188 46903 24191
rect 47213 24191 47271 24197
rect 47213 24188 47225 24191
rect 46891 24160 47225 24188
rect 46891 24157 46903 24160
rect 46845 24151 46903 24157
rect 47213 24157 47225 24160
rect 47259 24157 47271 24191
rect 47213 24151 47271 24157
rect 48038 24148 48044 24200
rect 48096 24148 48102 24200
rect 48774 24148 48780 24200
rect 48832 24148 48838 24200
rect 44266 24120 44272 24132
rect 41984 24092 44272 24120
rect 44266 24080 44272 24092
rect 44324 24080 44330 24132
rect 44726 24080 44732 24132
rect 44784 24120 44790 24132
rect 45373 24123 45431 24129
rect 45373 24120 45385 24123
rect 44784 24092 45385 24120
rect 44784 24080 44790 24092
rect 45373 24089 45385 24092
rect 45419 24120 45431 24123
rect 47394 24120 47400 24132
rect 45419 24092 47400 24120
rect 45419 24089 45431 24092
rect 45373 24083 45431 24089
rect 47394 24080 47400 24092
rect 47452 24080 47458 24132
rect 39850 24052 39856 24064
rect 38764 24024 39856 24052
rect 39850 24012 39856 24024
rect 39908 24012 39914 24064
rect 40034 24012 40040 24064
rect 40092 24012 40098 24064
rect 40310 24012 40316 24064
rect 40368 24052 40374 24064
rect 42610 24052 42616 24064
rect 40368 24024 42616 24052
rect 40368 24012 40374 24024
rect 42610 24012 42616 24024
rect 42668 24012 42674 24064
rect 42702 24012 42708 24064
rect 42760 24052 42766 24064
rect 45281 24055 45339 24061
rect 45281 24052 45293 24055
rect 42760 24024 45293 24052
rect 42760 24012 42766 24024
rect 45281 24021 45293 24024
rect 45327 24021 45339 24055
rect 45281 24015 45339 24021
rect 46014 24012 46020 24064
rect 46072 24012 46078 24064
rect 46106 24012 46112 24064
rect 46164 24052 46170 24064
rect 47857 24055 47915 24061
rect 47857 24052 47869 24055
rect 46164 24024 47869 24052
rect 46164 24012 46170 24024
rect 47857 24021 47869 24024
rect 47903 24021 47915 24055
rect 47857 24015 47915 24021
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 2317 23851 2375 23857
rect 2317 23817 2329 23851
rect 2363 23848 2375 23851
rect 4614 23848 4620 23860
rect 2363 23820 4620 23848
rect 2363 23817 2375 23820
rect 2317 23811 2375 23817
rect 4614 23808 4620 23820
rect 4672 23808 4678 23860
rect 10318 23848 10324 23860
rect 6886 23820 10324 23848
rect 6886 23780 6914 23820
rect 10318 23808 10324 23820
rect 10376 23808 10382 23860
rect 19610 23848 19616 23860
rect 16316 23820 19616 23848
rect 11790 23780 11796 23792
rect 2148 23752 6914 23780
rect 9324 23752 11796 23780
rect 2148 23721 2176 23752
rect 2133 23715 2191 23721
rect 2133 23681 2145 23715
rect 2179 23681 2191 23715
rect 2133 23675 2191 23681
rect 4062 23672 4068 23724
rect 4120 23672 4126 23724
rect 4706 23672 4712 23724
rect 4764 23672 4770 23724
rect 6825 23715 6883 23721
rect 6825 23681 6837 23715
rect 6871 23681 6883 23715
rect 6825 23675 6883 23681
rect 7285 23715 7343 23721
rect 7285 23681 7297 23715
rect 7331 23712 7343 23715
rect 8478 23712 8484 23724
rect 7331 23684 8484 23712
rect 7331 23681 7343 23684
rect 7285 23675 7343 23681
rect 3697 23647 3755 23653
rect 3697 23613 3709 23647
rect 3743 23644 3755 23647
rect 4154 23644 4160 23656
rect 3743 23616 4160 23644
rect 3743 23613 3755 23616
rect 3697 23607 3755 23613
rect 4154 23604 4160 23616
rect 4212 23604 4218 23656
rect 5442 23604 5448 23656
rect 5500 23604 5506 23656
rect 6840 23644 6868 23675
rect 8478 23672 8484 23684
rect 8536 23672 8542 23724
rect 9324 23721 9352 23752
rect 11790 23740 11796 23752
rect 11848 23740 11854 23792
rect 14182 23780 14188 23792
rect 13004 23752 14188 23780
rect 9309 23715 9367 23721
rect 9309 23681 9321 23715
rect 9355 23681 9367 23715
rect 9309 23675 9367 23681
rect 11149 23715 11207 23721
rect 11149 23681 11161 23715
rect 11195 23681 11207 23715
rect 11149 23675 11207 23681
rect 8386 23644 8392 23656
rect 6840 23616 8392 23644
rect 8386 23604 8392 23616
rect 8444 23604 8450 23656
rect 8849 23647 8907 23653
rect 8849 23613 8861 23647
rect 8895 23644 8907 23647
rect 9214 23644 9220 23656
rect 8895 23616 9220 23644
rect 8895 23613 8907 23616
rect 8849 23607 8907 23613
rect 9214 23604 9220 23616
rect 9272 23604 9278 23656
rect 10594 23604 10600 23656
rect 10652 23604 10658 23656
rect 11164 23644 11192 23675
rect 12342 23672 12348 23724
rect 12400 23672 12406 23724
rect 12710 23712 12716 23724
rect 12544 23684 12716 23712
rect 12544 23644 12572 23684
rect 12710 23672 12716 23684
rect 12768 23672 12774 23724
rect 11164 23616 12572 23644
rect 12621 23647 12679 23653
rect 12621 23613 12633 23647
rect 12667 23644 12679 23647
rect 13004 23644 13032 23752
rect 14182 23740 14188 23752
rect 14240 23740 14246 23792
rect 14277 23783 14335 23789
rect 14277 23749 14289 23783
rect 14323 23780 14335 23783
rect 14366 23780 14372 23792
rect 14323 23752 14372 23780
rect 14323 23749 14335 23752
rect 14277 23743 14335 23749
rect 14366 23740 14372 23752
rect 14424 23740 14430 23792
rect 16316 23721 16344 23820
rect 19610 23808 19616 23820
rect 19668 23808 19674 23860
rect 20180 23820 21036 23848
rect 20180 23780 20208 23820
rect 19826 23752 20208 23780
rect 20254 23740 20260 23792
rect 20312 23740 20318 23792
rect 21008 23789 21036 23820
rect 21450 23808 21456 23860
rect 21508 23808 21514 23860
rect 23753 23851 23811 23857
rect 23753 23817 23765 23851
rect 23799 23848 23811 23851
rect 27890 23848 27896 23860
rect 23799 23820 27896 23848
rect 23799 23817 23811 23820
rect 23753 23811 23811 23817
rect 27890 23808 27896 23820
rect 27948 23808 27954 23860
rect 28442 23808 28448 23860
rect 28500 23808 28506 23860
rect 32309 23851 32367 23857
rect 32309 23848 32321 23851
rect 28644 23820 32321 23848
rect 20993 23783 21051 23789
rect 20993 23749 21005 23783
rect 21039 23780 21051 23783
rect 21634 23780 21640 23792
rect 21039 23752 21640 23780
rect 21039 23749 21051 23752
rect 20993 23743 21051 23749
rect 21634 23740 21640 23752
rect 21692 23740 21698 23792
rect 24489 23783 24547 23789
rect 24489 23780 24501 23783
rect 23492 23752 24501 23780
rect 23492 23724 23520 23752
rect 24489 23749 24501 23752
rect 24535 23749 24547 23783
rect 24489 23743 24547 23749
rect 25866 23740 25872 23792
rect 25924 23740 25930 23792
rect 26329 23783 26387 23789
rect 26329 23749 26341 23783
rect 26375 23780 26387 23783
rect 27706 23780 27712 23792
rect 26375 23752 27712 23780
rect 26375 23749 26387 23752
rect 26329 23743 26387 23749
rect 27706 23740 27712 23752
rect 27764 23740 27770 23792
rect 28258 23780 28264 23792
rect 27816 23752 28264 23780
rect 27816 23724 27844 23752
rect 28258 23740 28264 23752
rect 28316 23740 28322 23792
rect 13081 23715 13139 23721
rect 13081 23681 13093 23715
rect 13127 23681 13139 23715
rect 13081 23675 13139 23681
rect 16301 23715 16359 23721
rect 16301 23681 16313 23715
rect 16347 23681 16359 23715
rect 16301 23675 16359 23681
rect 18233 23715 18291 23721
rect 18233 23681 18245 23715
rect 18279 23712 18291 23715
rect 18279 23684 19104 23712
rect 18279 23681 18291 23684
rect 18233 23675 18291 23681
rect 12667 23616 13032 23644
rect 12667 23613 12679 23616
rect 12621 23607 12679 23613
rect 3418 23536 3424 23588
rect 3476 23576 3482 23588
rect 5810 23576 5816 23588
rect 3476 23548 5816 23576
rect 3476 23536 3482 23548
rect 5810 23536 5816 23548
rect 5868 23536 5874 23588
rect 7469 23579 7527 23585
rect 7469 23545 7481 23579
rect 7515 23576 7527 23579
rect 13096 23576 13124 23675
rect 15841 23647 15899 23653
rect 15841 23613 15853 23647
rect 15887 23644 15899 23647
rect 16390 23644 16396 23656
rect 15887 23616 16396 23644
rect 15887 23613 15899 23616
rect 15841 23607 15899 23613
rect 16390 23604 16396 23616
rect 16448 23604 16454 23656
rect 17865 23647 17923 23653
rect 17865 23613 17877 23647
rect 17911 23644 17923 23647
rect 18322 23644 18328 23656
rect 17911 23616 18328 23644
rect 17911 23613 17923 23616
rect 17865 23607 17923 23613
rect 18322 23604 18328 23616
rect 18380 23604 18386 23656
rect 7515 23548 13124 23576
rect 7515 23545 7527 23548
rect 7469 23539 7527 23545
rect 2774 23468 2780 23520
rect 2832 23508 2838 23520
rect 5718 23508 5724 23520
rect 2832 23480 5724 23508
rect 2832 23468 2838 23480
rect 5718 23468 5724 23480
rect 5776 23468 5782 23520
rect 5994 23468 6000 23520
rect 6052 23508 6058 23520
rect 6641 23511 6699 23517
rect 6641 23508 6653 23511
rect 6052 23480 6653 23508
rect 6052 23468 6058 23480
rect 6641 23477 6653 23480
rect 6687 23477 6699 23511
rect 6641 23471 6699 23477
rect 18782 23468 18788 23520
rect 18840 23468 18846 23520
rect 19076 23508 19104 23684
rect 21266 23672 21272 23724
rect 21324 23672 21330 23724
rect 22833 23715 22891 23721
rect 22833 23681 22845 23715
rect 22879 23712 22891 23715
rect 23474 23712 23480 23724
rect 22879 23684 23480 23712
rect 22879 23681 22891 23684
rect 22833 23675 22891 23681
rect 23474 23672 23480 23684
rect 23532 23672 23538 23724
rect 23658 23672 23664 23724
rect 23716 23672 23722 23724
rect 27341 23715 27399 23721
rect 27341 23681 27353 23715
rect 27387 23712 27399 23715
rect 27387 23684 27614 23712
rect 27387 23681 27399 23684
rect 27341 23675 27399 23681
rect 20533 23647 20591 23653
rect 20533 23613 20545 23647
rect 20579 23644 20591 23647
rect 21726 23644 21732 23656
rect 20579 23616 21732 23644
rect 20579 23613 20591 23616
rect 20533 23607 20591 23613
rect 21726 23604 21732 23616
rect 21784 23604 21790 23656
rect 22554 23604 22560 23656
rect 22612 23604 22618 23656
rect 23842 23604 23848 23656
rect 23900 23604 23906 23656
rect 26602 23604 26608 23656
rect 26660 23604 26666 23656
rect 23382 23576 23388 23588
rect 20456 23548 23388 23576
rect 20456 23508 20484 23548
rect 23382 23536 23388 23548
rect 23440 23536 23446 23588
rect 27586 23576 27614 23684
rect 27798 23672 27804 23724
rect 27856 23672 27862 23724
rect 28644 23721 28672 23820
rect 32309 23817 32321 23820
rect 32355 23817 32367 23851
rect 32309 23811 32367 23817
rect 32769 23851 32827 23857
rect 32769 23817 32781 23851
rect 32815 23848 32827 23851
rect 37461 23851 37519 23857
rect 37461 23848 37473 23851
rect 32815 23820 37473 23848
rect 32815 23817 32827 23820
rect 32769 23811 32827 23817
rect 37461 23817 37473 23820
rect 37507 23817 37519 23851
rect 37461 23811 37519 23817
rect 37829 23851 37887 23857
rect 37829 23817 37841 23851
rect 37875 23848 37887 23851
rect 40034 23848 40040 23860
rect 37875 23820 40040 23848
rect 37875 23817 37887 23820
rect 37829 23811 37887 23817
rect 40034 23808 40040 23820
rect 40092 23808 40098 23860
rect 40126 23808 40132 23860
rect 40184 23848 40190 23860
rect 41969 23851 42027 23857
rect 41969 23848 41981 23851
rect 40184 23820 41981 23848
rect 40184 23808 40190 23820
rect 41969 23817 41981 23820
rect 42015 23817 42027 23851
rect 41969 23811 42027 23817
rect 42242 23808 42248 23860
rect 42300 23848 42306 23860
rect 42300 23820 46060 23848
rect 42300 23808 42306 23820
rect 31481 23783 31539 23789
rect 31481 23749 31493 23783
rect 31527 23780 31539 23783
rect 32398 23780 32404 23792
rect 31527 23752 32404 23780
rect 31527 23749 31539 23752
rect 31481 23743 31539 23749
rect 32398 23740 32404 23752
rect 32456 23780 32462 23792
rect 32456 23752 33732 23780
rect 32456 23740 32462 23752
rect 28629 23715 28687 23721
rect 28629 23681 28641 23715
rect 28675 23681 28687 23715
rect 28629 23675 28687 23681
rect 29089 23715 29147 23721
rect 29089 23681 29101 23715
rect 29135 23712 29147 23715
rect 29549 23715 29607 23721
rect 29549 23712 29561 23715
rect 29135 23684 29561 23712
rect 29135 23681 29147 23684
rect 29089 23675 29147 23681
rect 29549 23681 29561 23684
rect 29595 23681 29607 23715
rect 29549 23675 29607 23681
rect 28350 23604 28356 23656
rect 28408 23644 28414 23656
rect 29104 23644 29132 23675
rect 30374 23672 30380 23724
rect 30432 23672 30438 23724
rect 32674 23672 32680 23724
rect 32732 23672 32738 23724
rect 28408 23616 29132 23644
rect 28408 23604 28414 23616
rect 29362 23604 29368 23656
rect 29420 23644 29426 23656
rect 29420 23616 31708 23644
rect 29420 23604 29426 23616
rect 29638 23576 29644 23588
rect 24044 23548 25360 23576
rect 27586 23548 29644 23576
rect 19076 23480 20484 23508
rect 20990 23468 20996 23520
rect 21048 23508 21054 23520
rect 23293 23511 23351 23517
rect 23293 23508 23305 23511
rect 21048 23480 23305 23508
rect 21048 23468 21054 23480
rect 23293 23477 23305 23480
rect 23339 23477 23351 23511
rect 23293 23471 23351 23477
rect 23474 23468 23480 23520
rect 23532 23508 23538 23520
rect 24044 23508 24072 23548
rect 23532 23480 24072 23508
rect 23532 23468 23538 23480
rect 24394 23468 24400 23520
rect 24452 23468 24458 23520
rect 24854 23468 24860 23520
rect 24912 23468 24918 23520
rect 25332 23508 25360 23548
rect 29638 23536 29644 23548
rect 29696 23536 29702 23588
rect 31680 23576 31708 23616
rect 31754 23604 31760 23656
rect 31812 23604 31818 23656
rect 32953 23647 33011 23653
rect 32953 23613 32965 23647
rect 32999 23644 33011 23647
rect 33704 23644 33732 23752
rect 33778 23740 33784 23792
rect 33836 23780 33842 23792
rect 33836 23752 33902 23780
rect 33836 23740 33842 23752
rect 34974 23740 34980 23792
rect 35032 23780 35038 23792
rect 35032 23752 35480 23780
rect 35032 23740 35038 23752
rect 34974 23644 34980 23656
rect 32999 23616 33640 23644
rect 33704 23616 34980 23644
rect 32999 23613 33011 23616
rect 32953 23607 33011 23613
rect 32306 23576 32312 23588
rect 31680 23548 32312 23576
rect 32306 23536 32312 23548
rect 32364 23536 32370 23588
rect 27157 23511 27215 23517
rect 27157 23508 27169 23511
rect 25332 23480 27169 23508
rect 27157 23477 27169 23480
rect 27203 23477 27215 23511
rect 27157 23471 27215 23477
rect 27798 23468 27804 23520
rect 27856 23508 27862 23520
rect 27985 23511 28043 23517
rect 27985 23508 27997 23511
rect 27856 23480 27997 23508
rect 27856 23468 27862 23480
rect 27985 23477 27997 23480
rect 28031 23477 28043 23511
rect 27985 23471 28043 23477
rect 29086 23468 29092 23520
rect 29144 23508 29150 23520
rect 29273 23511 29331 23517
rect 29273 23508 29285 23511
rect 29144 23480 29285 23508
rect 29144 23468 29150 23480
rect 29273 23477 29285 23480
rect 29319 23477 29331 23511
rect 29273 23471 29331 23477
rect 30009 23511 30067 23517
rect 30009 23477 30021 23511
rect 30055 23508 30067 23511
rect 30282 23508 30288 23520
rect 30055 23480 30288 23508
rect 30055 23477 30067 23480
rect 30009 23471 30067 23477
rect 30282 23468 30288 23480
rect 30340 23468 30346 23520
rect 33612 23517 33640 23616
rect 34974 23604 34980 23616
rect 35032 23604 35038 23656
rect 35069 23647 35127 23653
rect 35069 23613 35081 23647
rect 35115 23644 35127 23647
rect 35115 23616 35296 23644
rect 35115 23613 35127 23616
rect 35069 23607 35127 23613
rect 33597 23511 33655 23517
rect 33597 23477 33609 23511
rect 33643 23508 33655 23511
rect 34514 23508 34520 23520
rect 33643 23480 34520 23508
rect 33643 23477 33655 23480
rect 33597 23471 33655 23477
rect 34514 23468 34520 23480
rect 34572 23468 34578 23520
rect 35268 23508 35296 23616
rect 35342 23604 35348 23656
rect 35400 23604 35406 23656
rect 35452 23644 35480 23752
rect 35618 23740 35624 23792
rect 35676 23780 35682 23792
rect 37921 23783 37979 23789
rect 37921 23780 37933 23783
rect 35676 23752 37933 23780
rect 35676 23740 35682 23752
rect 37921 23749 37933 23752
rect 37967 23749 37979 23783
rect 37921 23743 37979 23749
rect 39666 23740 39672 23792
rect 39724 23780 39730 23792
rect 41785 23783 41843 23789
rect 41785 23780 41797 23783
rect 39724 23752 41797 23780
rect 39724 23740 39730 23752
rect 41785 23749 41797 23752
rect 41831 23749 41843 23783
rect 41785 23743 41843 23749
rect 42521 23783 42579 23789
rect 42521 23749 42533 23783
rect 42567 23780 42579 23783
rect 42702 23780 42708 23792
rect 42567 23752 42708 23780
rect 42567 23749 42579 23752
rect 42521 23743 42579 23749
rect 42702 23740 42708 23752
rect 42760 23740 42766 23792
rect 35986 23672 35992 23724
rect 36044 23712 36050 23724
rect 36265 23715 36323 23721
rect 36044 23684 36124 23712
rect 36044 23672 36050 23684
rect 36096 23644 36124 23684
rect 36265 23681 36277 23715
rect 36311 23712 36323 23715
rect 36311 23684 38148 23712
rect 36311 23681 36323 23684
rect 36265 23675 36323 23681
rect 36357 23647 36415 23653
rect 36357 23644 36369 23647
rect 35452 23616 36032 23644
rect 36096 23616 36369 23644
rect 35434 23536 35440 23588
rect 35492 23576 35498 23588
rect 35897 23579 35955 23585
rect 35897 23576 35909 23579
rect 35492 23548 35909 23576
rect 35492 23536 35498 23548
rect 35897 23545 35909 23548
rect 35943 23545 35955 23579
rect 36004 23576 36032 23616
rect 36357 23613 36369 23616
rect 36403 23613 36415 23647
rect 36357 23607 36415 23613
rect 36449 23647 36507 23653
rect 36449 23613 36461 23647
rect 36495 23613 36507 23647
rect 38013 23647 38071 23653
rect 38013 23644 38025 23647
rect 36449 23607 36507 23613
rect 36556 23616 38025 23644
rect 36464 23576 36492 23607
rect 36004 23548 36492 23576
rect 35897 23539 35955 23545
rect 35526 23508 35532 23520
rect 35268 23480 35532 23508
rect 35526 23468 35532 23480
rect 35584 23508 35590 23520
rect 36556 23508 36584 23616
rect 38013 23613 38025 23616
rect 38059 23613 38071 23647
rect 38013 23607 38071 23613
rect 38120 23576 38148 23684
rect 39206 23672 39212 23724
rect 39264 23672 39270 23724
rect 39942 23672 39948 23724
rect 40000 23712 40006 23724
rect 40221 23715 40279 23721
rect 40221 23712 40233 23715
rect 40000 23684 40233 23712
rect 40000 23672 40006 23684
rect 40221 23681 40233 23684
rect 40267 23681 40279 23715
rect 40221 23675 40279 23681
rect 38562 23604 38568 23656
rect 38620 23604 38626 23656
rect 39301 23647 39359 23653
rect 39301 23613 39313 23647
rect 39347 23644 39359 23647
rect 39390 23644 39396 23656
rect 39347 23616 39396 23644
rect 39347 23613 39359 23616
rect 39301 23607 39359 23613
rect 39390 23604 39396 23616
rect 39448 23604 39454 23656
rect 39482 23604 39488 23656
rect 39540 23604 39546 23656
rect 40236 23644 40264 23675
rect 40310 23672 40316 23724
rect 40368 23712 40374 23724
rect 40957 23715 41015 23721
rect 40957 23712 40969 23715
rect 40368 23684 40969 23712
rect 40368 23672 40374 23684
rect 40957 23681 40969 23684
rect 41003 23681 41015 23715
rect 42613 23715 42671 23721
rect 42613 23712 42625 23715
rect 40957 23675 41015 23681
rect 41064 23684 42625 23712
rect 40586 23644 40592 23656
rect 40236 23616 40592 23644
rect 40586 23604 40592 23616
rect 40644 23604 40650 23656
rect 40681 23647 40739 23653
rect 40681 23613 40693 23647
rect 40727 23613 40739 23647
rect 40681 23607 40739 23613
rect 38841 23579 38899 23585
rect 38841 23576 38853 23579
rect 38120 23548 38853 23576
rect 38841 23545 38853 23548
rect 38887 23545 38899 23579
rect 38841 23539 38899 23545
rect 40037 23579 40095 23585
rect 40037 23545 40049 23579
rect 40083 23576 40095 23579
rect 40218 23576 40224 23588
rect 40083 23548 40224 23576
rect 40083 23545 40095 23548
rect 40037 23539 40095 23545
rect 40218 23536 40224 23548
rect 40276 23536 40282 23588
rect 40696 23576 40724 23607
rect 40770 23604 40776 23656
rect 40828 23644 40834 23656
rect 41064 23644 41092 23684
rect 42613 23681 42625 23684
rect 42659 23681 42671 23715
rect 42613 23675 42671 23681
rect 42794 23672 42800 23724
rect 42852 23712 42858 23724
rect 43073 23715 43131 23721
rect 43073 23712 43085 23715
rect 42852 23684 43085 23712
rect 42852 23672 42858 23684
rect 43073 23681 43085 23684
rect 43119 23681 43131 23715
rect 43073 23675 43131 23681
rect 44818 23672 44824 23724
rect 44876 23672 44882 23724
rect 45922 23672 45928 23724
rect 45980 23672 45986 23724
rect 46032 23712 46060 23820
rect 46198 23808 46204 23860
rect 46256 23848 46262 23860
rect 47581 23851 47639 23857
rect 47581 23848 47593 23851
rect 46256 23820 47593 23848
rect 46256 23808 46262 23820
rect 47581 23817 47593 23820
rect 47627 23817 47639 23851
rect 47581 23811 47639 23817
rect 47854 23808 47860 23860
rect 47912 23848 47918 23860
rect 49329 23851 49387 23857
rect 49329 23848 49341 23851
rect 47912 23820 49341 23848
rect 47912 23808 47918 23820
rect 49329 23817 49341 23820
rect 49375 23817 49387 23851
rect 49329 23811 49387 23817
rect 46934 23740 46940 23792
rect 46992 23780 46998 23792
rect 47765 23783 47823 23789
rect 47765 23780 47777 23783
rect 46992 23752 47777 23780
rect 46992 23740 46998 23752
rect 47765 23749 47777 23752
rect 47811 23749 47823 23783
rect 47765 23743 47823 23749
rect 46753 23715 46811 23721
rect 46753 23712 46765 23715
rect 46032 23684 46765 23712
rect 46753 23681 46765 23684
rect 46799 23681 46811 23715
rect 46753 23675 46811 23681
rect 47394 23672 47400 23724
rect 47452 23672 47458 23724
rect 48869 23715 48927 23721
rect 48869 23681 48881 23715
rect 48915 23712 48927 23715
rect 49234 23712 49240 23724
rect 48915 23684 49240 23712
rect 48915 23681 48927 23684
rect 48869 23675 48927 23681
rect 49234 23672 49240 23684
rect 49292 23672 49298 23724
rect 46385 23647 46443 23653
rect 46385 23644 46397 23647
rect 40828 23616 41092 23644
rect 41156 23616 46397 23644
rect 40828 23604 40834 23616
rect 41156 23576 41184 23616
rect 46385 23613 46397 23616
rect 46431 23613 46443 23647
rect 46385 23607 46443 23613
rect 47302 23604 47308 23656
rect 47360 23644 47366 23656
rect 49145 23647 49203 23653
rect 49145 23644 49157 23647
rect 47360 23616 49157 23644
rect 47360 23604 47366 23616
rect 49145 23613 49157 23616
rect 49191 23613 49203 23647
rect 49145 23607 49203 23613
rect 40604 23548 41184 23576
rect 35584 23480 36584 23508
rect 35584 23468 35590 23480
rect 36906 23468 36912 23520
rect 36964 23468 36970 23520
rect 37366 23468 37372 23520
rect 37424 23508 37430 23520
rect 40604 23508 40632 23548
rect 42702 23536 42708 23588
rect 42760 23536 42766 23588
rect 45922 23536 45928 23588
rect 45980 23576 45986 23588
rect 46934 23576 46940 23588
rect 45980 23548 46940 23576
rect 45980 23536 45986 23548
rect 46934 23536 46940 23548
rect 46992 23536 46998 23588
rect 47118 23536 47124 23588
rect 47176 23576 47182 23588
rect 48225 23579 48283 23585
rect 48225 23576 48237 23579
rect 47176 23548 48237 23576
rect 47176 23536 47182 23548
rect 48225 23545 48237 23548
rect 48271 23545 48283 23579
rect 48225 23539 48283 23545
rect 37424 23480 40632 23508
rect 37424 23468 37430 23480
rect 40678 23468 40684 23520
rect 40736 23508 40742 23520
rect 42720 23508 42748 23536
rect 40736 23480 42748 23508
rect 40736 23468 40742 23480
rect 43530 23468 43536 23520
rect 43588 23508 43594 23520
rect 45281 23511 45339 23517
rect 45281 23508 45293 23511
rect 43588 23480 45293 23508
rect 43588 23468 43594 23480
rect 45281 23477 45293 23480
rect 45327 23477 45339 23511
rect 45281 23471 45339 23477
rect 46198 23468 46204 23520
rect 46256 23468 46262 23520
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 4706 23264 4712 23316
rect 4764 23264 4770 23316
rect 15838 23304 15844 23316
rect 10060 23276 15844 23304
rect 5258 23196 5264 23248
rect 5316 23236 5322 23248
rect 9125 23239 9183 23245
rect 9125 23236 9137 23239
rect 5316 23208 9137 23236
rect 5316 23196 5322 23208
rect 9125 23205 9137 23208
rect 9171 23205 9183 23239
rect 9125 23199 9183 23205
rect 5626 23168 5632 23180
rect 2976 23140 5632 23168
rect 2976 23109 3004 23140
rect 5626 23128 5632 23140
rect 5684 23128 5690 23180
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 10060 23177 10088 23276
rect 15838 23264 15844 23276
rect 15896 23264 15902 23316
rect 16224 23276 19748 23304
rect 14182 23196 14188 23248
rect 14240 23236 14246 23248
rect 16224 23236 16252 23276
rect 14240 23208 16252 23236
rect 14240 23196 14246 23208
rect 19610 23196 19616 23248
rect 19668 23196 19674 23248
rect 19720 23236 19748 23276
rect 19886 23264 19892 23316
rect 19944 23304 19950 23316
rect 20254 23304 20260 23316
rect 19944 23276 20260 23304
rect 19944 23264 19950 23276
rect 20254 23264 20260 23276
rect 20312 23304 20318 23316
rect 20349 23307 20407 23313
rect 20349 23304 20361 23307
rect 20312 23276 20361 23304
rect 20312 23264 20318 23276
rect 20349 23273 20361 23276
rect 20395 23273 20407 23307
rect 22830 23304 22836 23316
rect 20349 23267 20407 23273
rect 20456 23276 22836 23304
rect 20456 23236 20484 23276
rect 22830 23264 22836 23276
rect 22888 23264 22894 23316
rect 25130 23304 25136 23316
rect 23308 23276 25136 23304
rect 23308 23236 23336 23276
rect 25130 23264 25136 23276
rect 25188 23264 25194 23316
rect 25225 23307 25283 23313
rect 25225 23273 25237 23307
rect 25271 23304 25283 23307
rect 25406 23304 25412 23316
rect 25271 23276 25412 23304
rect 25271 23273 25283 23276
rect 25225 23267 25283 23273
rect 25406 23264 25412 23276
rect 25464 23264 25470 23316
rect 27890 23264 27896 23316
rect 27948 23264 27954 23316
rect 28350 23264 28356 23316
rect 28408 23304 28414 23316
rect 29089 23307 29147 23313
rect 29089 23304 29101 23307
rect 28408 23276 29101 23304
rect 28408 23264 28414 23276
rect 29089 23273 29101 23276
rect 29135 23304 29147 23307
rect 30374 23304 30380 23316
rect 29135 23276 30380 23304
rect 29135 23273 29147 23276
rect 29089 23267 29147 23273
rect 30374 23264 30380 23276
rect 30432 23304 30438 23316
rect 30745 23307 30803 23313
rect 30745 23304 30757 23307
rect 30432 23276 30757 23304
rect 30432 23264 30438 23276
rect 30745 23273 30757 23276
rect 30791 23273 30803 23307
rect 30745 23267 30803 23273
rect 31113 23307 31171 23313
rect 31113 23273 31125 23307
rect 31159 23304 31171 23307
rect 31478 23304 31484 23316
rect 31159 23276 31484 23304
rect 31159 23273 31171 23276
rect 31113 23267 31171 23273
rect 31478 23264 31484 23276
rect 31536 23264 31542 23316
rect 33318 23264 33324 23316
rect 33376 23304 33382 23316
rect 34149 23307 34207 23313
rect 34149 23304 34161 23307
rect 33376 23276 34161 23304
rect 33376 23264 33382 23276
rect 34149 23273 34161 23276
rect 34195 23273 34207 23307
rect 34149 23267 34207 23273
rect 35066 23264 35072 23316
rect 35124 23304 35130 23316
rect 37366 23304 37372 23316
rect 35124 23276 37372 23304
rect 35124 23264 35130 23276
rect 37366 23264 37372 23276
rect 37424 23264 37430 23316
rect 37458 23264 37464 23316
rect 37516 23304 37522 23316
rect 38767 23307 38825 23313
rect 38767 23304 38779 23307
rect 37516 23276 38779 23304
rect 37516 23264 37522 23276
rect 38767 23273 38779 23276
rect 38813 23304 38825 23307
rect 38813 23276 40632 23304
rect 38813 23273 38825 23276
rect 38767 23267 38825 23273
rect 19720 23208 20484 23236
rect 22756 23208 23336 23236
rect 10045 23171 10103 23177
rect 10045 23137 10057 23171
rect 10091 23137 10103 23171
rect 10045 23131 10103 23137
rect 11238 23128 11244 23180
rect 11296 23128 11302 23180
rect 13265 23171 13323 23177
rect 13265 23137 13277 23171
rect 13311 23168 13323 23171
rect 13354 23168 13360 23180
rect 13311 23140 13360 23168
rect 13311 23137 13323 23140
rect 13265 23131 13323 23137
rect 13354 23128 13360 23140
rect 13412 23128 13418 23180
rect 15746 23128 15752 23180
rect 15804 23128 15810 23180
rect 19518 23168 19524 23180
rect 16684 23140 19524 23168
rect 2961 23103 3019 23109
rect 2961 23069 2973 23103
rect 3007 23069 3019 23103
rect 2961 23063 3019 23069
rect 4249 23103 4307 23109
rect 4249 23069 4261 23103
rect 4295 23100 4307 23103
rect 4430 23100 4436 23112
rect 4295 23072 4436 23100
rect 4295 23069 4307 23072
rect 4249 23063 4307 23069
rect 4430 23060 4436 23072
rect 4488 23060 4494 23112
rect 4893 23103 4951 23109
rect 4893 23069 4905 23103
rect 4939 23069 4951 23103
rect 4893 23063 4951 23069
rect 1762 22992 1768 23044
rect 1820 22992 1826 23044
rect 4065 22967 4123 22973
rect 4065 22933 4077 22967
rect 4111 22964 4123 22967
rect 4614 22964 4620 22976
rect 4111 22936 4620 22964
rect 4111 22933 4123 22936
rect 4065 22927 4123 22933
rect 4614 22924 4620 22936
rect 4672 22924 4678 22976
rect 4908 22964 4936 23063
rect 5350 23060 5356 23112
rect 5408 23060 5414 23112
rect 5534 23060 5540 23112
rect 5592 23100 5598 23112
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 5592 23072 7205 23100
rect 5592 23060 5598 23072
rect 7193 23069 7205 23072
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 9122 23060 9128 23112
rect 9180 23100 9186 23112
rect 9309 23103 9367 23109
rect 9309 23100 9321 23103
rect 9180 23072 9321 23100
rect 9180 23060 9186 23072
rect 9309 23069 9321 23072
rect 9355 23069 9367 23103
rect 9309 23063 9367 23069
rect 11882 23060 11888 23112
rect 11940 23060 11946 23112
rect 13725 23103 13783 23109
rect 13725 23069 13737 23103
rect 13771 23100 13783 23103
rect 13814 23100 13820 23112
rect 13771 23072 13820 23100
rect 13771 23069 13783 23072
rect 13725 23063 13783 23069
rect 13814 23060 13820 23072
rect 13872 23060 13878 23112
rect 16684 23109 16712 23140
rect 19518 23128 19524 23140
rect 19576 23128 19582 23180
rect 21726 23128 21732 23180
rect 21784 23168 21790 23180
rect 22097 23171 22155 23177
rect 22097 23168 22109 23171
rect 21784 23140 22109 23168
rect 21784 23128 21790 23140
rect 22097 23137 22109 23140
rect 22143 23137 22155 23171
rect 22097 23131 22155 23137
rect 14829 23103 14887 23109
rect 14829 23069 14841 23103
rect 14875 23069 14887 23103
rect 14829 23063 14887 23069
rect 16669 23103 16727 23109
rect 16669 23069 16681 23103
rect 16715 23069 16727 23103
rect 16669 23063 16727 23069
rect 18877 23103 18935 23109
rect 18877 23069 18889 23103
rect 18923 23100 18935 23103
rect 19334 23100 19340 23112
rect 18923 23072 19340 23100
rect 18923 23069 18935 23072
rect 18877 23063 18935 23069
rect 14844 23032 14872 23063
rect 19334 23060 19340 23072
rect 19392 23060 19398 23112
rect 22756 23109 22784 23208
rect 23382 23196 23388 23248
rect 23440 23236 23446 23248
rect 24581 23239 24639 23245
rect 24581 23236 24593 23239
rect 23440 23208 24593 23236
rect 23440 23196 23446 23208
rect 24581 23205 24593 23208
rect 24627 23205 24639 23239
rect 24581 23199 24639 23205
rect 28258 23196 28264 23248
rect 28316 23236 28322 23248
rect 28997 23239 29055 23245
rect 28997 23236 29009 23239
rect 28316 23208 29009 23236
rect 28316 23196 28322 23208
rect 28997 23205 29009 23208
rect 29043 23205 29055 23239
rect 29733 23239 29791 23245
rect 29733 23236 29745 23239
rect 28997 23199 29055 23205
rect 29656 23208 29745 23236
rect 29656 23180 29684 23208
rect 29733 23205 29745 23208
rect 29779 23205 29791 23239
rect 29733 23199 29791 23205
rect 33778 23196 33784 23248
rect 33836 23236 33842 23248
rect 34425 23239 34483 23245
rect 34425 23236 34437 23239
rect 33836 23208 34437 23236
rect 33836 23196 33842 23208
rect 34425 23205 34437 23208
rect 34471 23236 34483 23239
rect 34606 23236 34612 23248
rect 34471 23208 34612 23236
rect 34471 23205 34483 23208
rect 34425 23199 34483 23205
rect 34606 23196 34612 23208
rect 34664 23196 34670 23248
rect 36354 23196 36360 23248
rect 36412 23236 36418 23248
rect 37182 23236 37188 23248
rect 36412 23208 37188 23236
rect 36412 23196 36418 23208
rect 37182 23196 37188 23208
rect 37240 23236 37246 23248
rect 37277 23239 37335 23245
rect 37277 23236 37289 23239
rect 37240 23208 37289 23236
rect 37240 23196 37246 23208
rect 37277 23205 37289 23208
rect 37323 23205 37335 23239
rect 37277 23199 37335 23205
rect 40034 23196 40040 23248
rect 40092 23196 40098 23248
rect 23937 23171 23995 23177
rect 23937 23137 23949 23171
rect 23983 23168 23995 23171
rect 24854 23168 24860 23180
rect 23983 23140 24860 23168
rect 23983 23137 23995 23140
rect 23937 23131 23995 23137
rect 24854 23128 24860 23140
rect 24912 23168 24918 23180
rect 25961 23171 26019 23177
rect 25961 23168 25973 23171
rect 24912 23140 25973 23168
rect 24912 23128 24918 23140
rect 25961 23137 25973 23140
rect 26007 23137 26019 23171
rect 25961 23131 26019 23137
rect 26050 23128 26056 23180
rect 26108 23168 26114 23180
rect 28445 23171 28503 23177
rect 28445 23168 28457 23171
rect 26108 23140 28457 23168
rect 26108 23128 26114 23140
rect 28445 23137 28457 23140
rect 28491 23137 28503 23171
rect 28445 23131 28503 23137
rect 29638 23128 29644 23180
rect 29696 23128 29702 23180
rect 30190 23128 30196 23180
rect 30248 23128 30254 23180
rect 30282 23128 30288 23180
rect 30340 23128 30346 23180
rect 31754 23168 31760 23180
rect 31404 23140 31760 23168
rect 22741 23103 22799 23109
rect 22741 23069 22753 23103
rect 22787 23069 22799 23103
rect 22741 23063 22799 23069
rect 23661 23103 23719 23109
rect 23661 23069 23673 23103
rect 23707 23100 23719 23103
rect 23707 23072 25636 23100
rect 23707 23069 23719 23072
rect 23661 23063 23719 23069
rect 16574 23032 16580 23044
rect 14844 23004 16580 23032
rect 16574 22992 16580 23004
rect 16632 22992 16638 23044
rect 17862 22992 17868 23044
rect 17920 22992 17926 23044
rect 18598 22992 18604 23044
rect 18656 22992 18662 23044
rect 19794 22992 19800 23044
rect 19852 22992 19858 23044
rect 21726 23032 21732 23044
rect 21390 23004 21732 23032
rect 21726 22992 21732 23004
rect 21784 22992 21790 23044
rect 21818 22992 21824 23044
rect 21876 22992 21882 23044
rect 22554 22992 22560 23044
rect 22612 22992 22618 23044
rect 24762 22992 24768 23044
rect 24820 22992 24826 23044
rect 25608 23032 25636 23072
rect 25682 23060 25688 23112
rect 25740 23060 25746 23112
rect 28353 23103 28411 23109
rect 28353 23069 28365 23103
rect 28399 23100 28411 23103
rect 29365 23103 29423 23109
rect 29365 23100 29377 23103
rect 28399 23072 29377 23100
rect 28399 23069 28411 23072
rect 28353 23063 28411 23069
rect 29365 23069 29377 23072
rect 29411 23100 29423 23103
rect 30098 23100 30104 23112
rect 29411 23072 30104 23100
rect 29411 23069 29423 23072
rect 29365 23063 29423 23069
rect 30098 23060 30104 23072
rect 30156 23060 30162 23112
rect 26234 23032 26240 23044
rect 25608 23004 26240 23032
rect 26234 22992 26240 23004
rect 26292 22992 26298 23044
rect 27246 23032 27252 23044
rect 27186 23004 27252 23032
rect 27246 22992 27252 23004
rect 27304 22992 27310 23044
rect 29914 23032 29920 23044
rect 27448 23004 29920 23032
rect 9214 22964 9220 22976
rect 4908 22936 9220 22964
rect 9214 22924 9220 22936
rect 9272 22924 9278 22976
rect 14366 22924 14372 22976
rect 14424 22924 14430 22976
rect 14642 22924 14648 22976
rect 14700 22924 14706 22976
rect 17126 22924 17132 22976
rect 17184 22924 17190 22976
rect 18874 22924 18880 22976
rect 18932 22964 18938 22976
rect 19337 22967 19395 22973
rect 19337 22964 19349 22967
rect 18932 22936 19349 22964
rect 18932 22924 18938 22936
rect 19337 22933 19349 22936
rect 19383 22964 19395 22967
rect 20806 22964 20812 22976
rect 19383 22936 20812 22964
rect 19383 22933 19395 22936
rect 19337 22927 19395 22933
rect 20806 22924 20812 22936
rect 20864 22924 20870 22976
rect 21542 22924 21548 22976
rect 21600 22964 21606 22976
rect 23198 22964 23204 22976
rect 21600 22936 23204 22964
rect 21600 22924 21606 22936
rect 23198 22924 23204 22936
rect 23256 22924 23262 22976
rect 23290 22924 23296 22976
rect 23348 22924 23354 22976
rect 23750 22924 23756 22976
rect 23808 22924 23814 22976
rect 25314 22924 25320 22976
rect 25372 22924 25378 22976
rect 25406 22924 25412 22976
rect 25464 22964 25470 22976
rect 26050 22964 26056 22976
rect 25464 22936 26056 22964
rect 25464 22924 25470 22936
rect 26050 22924 26056 22936
rect 26108 22924 26114 22976
rect 26326 22924 26332 22976
rect 26384 22964 26390 22976
rect 27448 22973 27476 23004
rect 29914 22992 29920 23004
rect 29972 22992 29978 23044
rect 30300 23032 30328 23128
rect 31404 23112 31432 23140
rect 31754 23128 31760 23140
rect 31812 23128 31818 23180
rect 33137 23171 33195 23177
rect 33137 23137 33149 23171
rect 33183 23168 33195 23171
rect 33502 23168 33508 23180
rect 33183 23140 33508 23168
rect 33183 23137 33195 23140
rect 33137 23131 33195 23137
rect 33502 23128 33508 23140
rect 33560 23128 33566 23180
rect 34330 23128 34336 23180
rect 34388 23168 34394 23180
rect 35069 23171 35127 23177
rect 35069 23168 35081 23171
rect 34388 23140 35081 23168
rect 34388 23128 34394 23140
rect 35069 23137 35081 23140
rect 35115 23168 35127 23171
rect 35342 23168 35348 23180
rect 35115 23140 35348 23168
rect 35115 23137 35127 23140
rect 35069 23131 35127 23137
rect 35342 23128 35348 23140
rect 35400 23128 35406 23180
rect 35710 23128 35716 23180
rect 35768 23168 35774 23180
rect 38378 23168 38384 23180
rect 35768 23140 38384 23168
rect 35768 23128 35774 23140
rect 38378 23128 38384 23140
rect 38436 23128 38442 23180
rect 38654 23128 38660 23180
rect 38712 23168 38718 23180
rect 39025 23171 39083 23177
rect 39025 23168 39037 23171
rect 38712 23140 39037 23168
rect 38712 23128 38718 23140
rect 39025 23137 39037 23140
rect 39071 23168 39083 23171
rect 39482 23168 39488 23180
rect 39071 23140 39488 23168
rect 39071 23137 39083 23140
rect 39025 23131 39083 23137
rect 39482 23128 39488 23140
rect 39540 23128 39546 23180
rect 40604 23177 40632 23276
rect 42794 23264 42800 23316
rect 42852 23304 42858 23316
rect 44269 23307 44327 23313
rect 44269 23304 44281 23307
rect 42852 23276 44281 23304
rect 42852 23264 42858 23276
rect 44269 23273 44281 23276
rect 44315 23273 44327 23307
rect 44269 23267 44327 23273
rect 44818 23264 44824 23316
rect 44876 23304 44882 23316
rect 45189 23307 45247 23313
rect 45189 23304 45201 23307
rect 44876 23276 45201 23304
rect 44876 23264 44882 23276
rect 45189 23273 45201 23276
rect 45235 23273 45247 23307
rect 45189 23267 45247 23273
rect 46658 23264 46664 23316
rect 46716 23264 46722 23316
rect 46934 23264 46940 23316
rect 46992 23264 46998 23316
rect 43714 23196 43720 23248
rect 43772 23236 43778 23248
rect 44729 23239 44787 23245
rect 44729 23236 44741 23239
rect 43772 23208 44741 23236
rect 43772 23196 43778 23208
rect 44729 23205 44741 23208
rect 44775 23236 44787 23239
rect 46106 23236 46112 23248
rect 44775 23208 46112 23236
rect 44775 23205 44787 23208
rect 44729 23199 44787 23205
rect 46106 23196 46112 23208
rect 46164 23196 46170 23248
rect 40589 23171 40647 23177
rect 40589 23137 40601 23171
rect 40635 23137 40647 23171
rect 43533 23171 43591 23177
rect 43533 23168 43545 23171
rect 40589 23131 40647 23137
rect 41064 23140 43545 23168
rect 31386 23060 31392 23112
rect 31444 23060 31450 23112
rect 33873 23103 33931 23109
rect 33873 23100 33885 23103
rect 33060 23072 33885 23100
rect 31665 23035 31723 23041
rect 31665 23032 31677 23035
rect 30024 23004 30236 23032
rect 30300 23004 31677 23032
rect 27433 22967 27491 22973
rect 27433 22964 27445 22967
rect 26384 22936 27445 22964
rect 26384 22924 26390 22936
rect 27433 22933 27445 22936
rect 27479 22933 27491 22967
rect 27433 22927 27491 22933
rect 28261 22967 28319 22973
rect 28261 22933 28273 22967
rect 28307 22964 28319 22967
rect 30024 22964 30052 23004
rect 28307 22936 30052 22964
rect 28307 22933 28319 22936
rect 28261 22927 28319 22933
rect 30098 22924 30104 22976
rect 30156 22924 30162 22976
rect 30208 22964 30236 23004
rect 31665 23001 31677 23004
rect 31711 23001 31723 23035
rect 31665 22995 31723 23001
rect 32122 22992 32128 23044
rect 32180 22992 32186 23044
rect 30374 22964 30380 22976
rect 30208 22936 30380 22964
rect 30374 22924 30380 22936
rect 30432 22924 30438 22976
rect 31202 22924 31208 22976
rect 31260 22964 31266 22976
rect 33060 22964 33088 23072
rect 33873 23069 33885 23072
rect 33919 23100 33931 23103
rect 34701 23103 34759 23109
rect 34701 23100 34713 23103
rect 33919 23072 34713 23100
rect 33919 23069 33931 23072
rect 33873 23063 33931 23069
rect 34701 23069 34713 23072
rect 34747 23069 34759 23103
rect 39500 23100 39528 23128
rect 41064 23109 41092 23140
rect 43533 23137 43545 23140
rect 43579 23168 43591 23171
rect 45649 23171 45707 23177
rect 45649 23168 45661 23171
rect 43579 23140 45661 23168
rect 43579 23137 43591 23140
rect 43533 23131 43591 23137
rect 45649 23137 45661 23140
rect 45695 23137 45707 23171
rect 45649 23131 45707 23137
rect 41049 23103 41107 23109
rect 41049 23100 41061 23103
rect 39500 23072 41061 23100
rect 34701 23063 34759 23069
rect 41049 23069 41061 23072
rect 41095 23069 41107 23103
rect 41049 23063 41107 23069
rect 44082 23060 44088 23112
rect 44140 23100 44146 23112
rect 44361 23103 44419 23109
rect 44361 23100 44373 23103
rect 44140 23072 44373 23100
rect 44140 23060 44146 23072
rect 44361 23069 44373 23072
rect 44407 23069 44419 23103
rect 44361 23063 44419 23069
rect 45370 23060 45376 23112
rect 45428 23060 45434 23112
rect 46293 23103 46351 23109
rect 46293 23069 46305 23103
rect 46339 23100 46351 23103
rect 46658 23100 46664 23112
rect 46339 23072 46664 23100
rect 46339 23069 46351 23072
rect 46293 23063 46351 23069
rect 46658 23060 46664 23072
rect 46716 23060 46722 23112
rect 47118 23060 47124 23112
rect 47176 23060 47182 23112
rect 47302 23060 47308 23112
rect 47360 23100 47366 23112
rect 47857 23103 47915 23109
rect 47857 23100 47869 23103
rect 47360 23072 47869 23100
rect 47360 23060 47366 23072
rect 47857 23069 47869 23072
rect 47903 23069 47915 23103
rect 47857 23063 47915 23069
rect 48593 23103 48651 23109
rect 48593 23069 48605 23103
rect 48639 23100 48651 23103
rect 48682 23100 48688 23112
rect 48639 23072 48688 23100
rect 48639 23069 48651 23072
rect 48593 23063 48651 23069
rect 48682 23060 48688 23072
rect 48740 23060 48746 23112
rect 49329 23103 49387 23109
rect 49329 23069 49341 23103
rect 49375 23100 49387 23103
rect 49418 23100 49424 23112
rect 49375 23072 49424 23100
rect 49375 23069 49387 23072
rect 49329 23063 49387 23069
rect 49418 23060 49424 23072
rect 49476 23060 49482 23112
rect 33410 22992 33416 23044
rect 33468 23032 33474 23044
rect 33468 23004 33916 23032
rect 33468 22992 33474 23004
rect 31260 22936 33088 22964
rect 33689 22967 33747 22973
rect 31260 22924 31266 22936
rect 33689 22933 33701 22967
rect 33735 22964 33747 22967
rect 33778 22964 33784 22976
rect 33735 22936 33784 22964
rect 33735 22933 33747 22936
rect 33689 22927 33747 22933
rect 33778 22924 33784 22936
rect 33836 22924 33842 22976
rect 33888 22964 33916 23004
rect 34514 22992 34520 23044
rect 34572 23032 34578 23044
rect 35345 23035 35403 23041
rect 35345 23032 35357 23035
rect 34572 23004 35357 23032
rect 34572 22992 34578 23004
rect 35345 23001 35357 23004
rect 35391 23001 35403 23035
rect 36906 23032 36912 23044
rect 36570 23004 36912 23032
rect 35345 22995 35403 23001
rect 36906 22992 36912 23004
rect 36964 23032 36970 23044
rect 36964 23004 37504 23032
rect 38318 23004 38654 23032
rect 36964 22992 36970 23004
rect 35158 22964 35164 22976
rect 33888 22936 35164 22964
rect 35158 22924 35164 22936
rect 35216 22924 35222 22976
rect 36817 22967 36875 22973
rect 36817 22933 36829 22967
rect 36863 22964 36875 22967
rect 37090 22964 37096 22976
rect 36863 22936 37096 22964
rect 36863 22933 36875 22936
rect 36817 22927 36875 22933
rect 37090 22924 37096 22936
rect 37148 22924 37154 22976
rect 37476 22964 37504 23004
rect 38396 22964 38424 23004
rect 37476 22936 38424 22964
rect 38626 22976 38654 23004
rect 40218 22992 40224 23044
rect 40276 23032 40282 23044
rect 40497 23035 40555 23041
rect 40497 23032 40509 23035
rect 40276 23004 40509 23032
rect 40276 22992 40282 23004
rect 40497 23001 40509 23004
rect 40543 23001 40555 23035
rect 40497 22995 40555 23001
rect 41506 22992 41512 23044
rect 41564 22992 41570 23044
rect 42702 22992 42708 23044
rect 42760 22992 42766 23044
rect 43257 23035 43315 23041
rect 43257 23001 43269 23035
rect 43303 23032 43315 23035
rect 43530 23032 43536 23044
rect 43303 23004 43536 23032
rect 43303 23001 43315 23004
rect 43257 22995 43315 23001
rect 43530 22992 43536 23004
rect 43588 22992 43594 23044
rect 43622 22992 43628 23044
rect 43680 23032 43686 23044
rect 43680 23004 49188 23032
rect 43680 22992 43686 23004
rect 38626 22936 38660 22976
rect 38654 22924 38660 22936
rect 38712 22964 38718 22976
rect 39393 22967 39451 22973
rect 39393 22964 39405 22967
rect 38712 22936 39405 22964
rect 38712 22924 38718 22936
rect 39393 22933 39405 22936
rect 39439 22964 39451 22967
rect 39666 22964 39672 22976
rect 39439 22936 39672 22964
rect 39439 22933 39451 22936
rect 39393 22927 39451 22933
rect 39666 22924 39672 22936
rect 39724 22924 39730 22976
rect 40405 22967 40463 22973
rect 40405 22933 40417 22967
rect 40451 22964 40463 22967
rect 41230 22964 41236 22976
rect 40451 22936 41236 22964
rect 40451 22933 40463 22936
rect 40405 22927 40463 22933
rect 41230 22924 41236 22936
rect 41288 22924 41294 22976
rect 41524 22964 41552 22992
rect 43809 22967 43867 22973
rect 43809 22964 43821 22967
rect 41524 22936 43821 22964
rect 43809 22933 43821 22936
rect 43855 22933 43867 22967
rect 43809 22927 43867 22933
rect 46106 22924 46112 22976
rect 46164 22924 46170 22976
rect 47026 22924 47032 22976
rect 47084 22964 47090 22976
rect 47486 22964 47492 22976
rect 47084 22936 47492 22964
rect 47084 22924 47090 22936
rect 47486 22924 47492 22936
rect 47544 22924 47550 22976
rect 47670 22924 47676 22976
rect 47728 22924 47734 22976
rect 48406 22924 48412 22976
rect 48464 22924 48470 22976
rect 49160 22973 49188 23004
rect 49145 22967 49203 22973
rect 49145 22933 49157 22967
rect 49191 22933 49203 22967
rect 49145 22927 49203 22933
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 1578 22720 1584 22772
rect 1636 22760 1642 22772
rect 3418 22760 3424 22772
rect 1636 22732 3424 22760
rect 1636 22720 1642 22732
rect 3418 22720 3424 22732
rect 3476 22720 3482 22772
rect 3602 22720 3608 22772
rect 3660 22760 3666 22772
rect 5350 22760 5356 22772
rect 3660 22732 5356 22760
rect 3660 22720 3666 22732
rect 5350 22720 5356 22732
rect 5408 22720 5414 22772
rect 7190 22720 7196 22772
rect 7248 22720 7254 22772
rect 15746 22760 15752 22772
rect 7300 22732 15752 22760
rect 4798 22652 4804 22704
rect 4856 22652 4862 22704
rect 7098 22692 7104 22704
rect 5644 22664 7104 22692
rect 2961 22627 3019 22633
rect 2961 22593 2973 22627
rect 3007 22593 3019 22627
rect 2961 22587 3019 22593
rect 3973 22627 4031 22633
rect 3973 22593 3985 22627
rect 4019 22624 4031 22627
rect 5644 22624 5672 22664
rect 7098 22652 7104 22664
rect 7156 22652 7162 22704
rect 4019 22596 5672 22624
rect 4019 22593 4031 22596
rect 3973 22587 4031 22593
rect 2501 22559 2559 22565
rect 2501 22525 2513 22559
rect 2547 22556 2559 22559
rect 2774 22556 2780 22568
rect 2547 22528 2780 22556
rect 2547 22525 2559 22528
rect 2501 22519 2559 22525
rect 2774 22516 2780 22528
rect 2832 22516 2838 22568
rect 2976 22556 3004 22587
rect 5994 22584 6000 22636
rect 6052 22584 6058 22636
rect 6641 22627 6699 22633
rect 6641 22593 6653 22627
rect 6687 22624 6699 22627
rect 7190 22624 7196 22636
rect 6687 22596 7196 22624
rect 6687 22593 6699 22596
rect 6641 22587 6699 22593
rect 7190 22584 7196 22596
rect 7248 22584 7254 22636
rect 7300 22556 7328 22732
rect 15746 22720 15752 22732
rect 15804 22720 15810 22772
rect 18598 22720 18604 22772
rect 18656 22720 18662 22772
rect 19153 22763 19211 22769
rect 19153 22729 19165 22763
rect 19199 22760 19211 22763
rect 19334 22760 19340 22772
rect 19199 22732 19340 22760
rect 19199 22729 19211 22732
rect 19153 22723 19211 22729
rect 19334 22720 19340 22732
rect 19392 22720 19398 22772
rect 21177 22763 21235 22769
rect 19904 22732 21036 22760
rect 9950 22652 9956 22704
rect 10008 22652 10014 22704
rect 11885 22695 11943 22701
rect 11885 22692 11897 22695
rect 11072 22664 11897 22692
rect 7466 22584 7472 22636
rect 7524 22584 7530 22636
rect 9309 22627 9367 22633
rect 9309 22593 9321 22627
rect 9355 22624 9367 22627
rect 11072 22624 11100 22664
rect 11885 22661 11897 22664
rect 11931 22661 11943 22695
rect 11885 22655 11943 22661
rect 9355 22596 11100 22624
rect 9355 22593 9367 22596
rect 9309 22587 9367 22593
rect 11146 22584 11152 22636
rect 11204 22584 11210 22636
rect 11900 22624 11928 22655
rect 12802 22652 12808 22704
rect 12860 22652 12866 22704
rect 15102 22652 15108 22704
rect 15160 22652 15166 22704
rect 15194 22652 15200 22704
rect 15252 22692 15258 22704
rect 17129 22695 17187 22701
rect 17129 22692 17141 22695
rect 15252 22664 17141 22692
rect 15252 22652 15258 22664
rect 17129 22661 17141 22664
rect 17175 22661 17187 22695
rect 17129 22655 17187 22661
rect 17862 22652 17868 22704
rect 17920 22652 17926 22704
rect 19904 22692 19932 22732
rect 19352 22664 19932 22692
rect 13446 22624 13452 22636
rect 11900 22596 13452 22624
rect 13446 22584 13452 22596
rect 13504 22584 13510 22636
rect 14001 22627 14059 22633
rect 14001 22593 14013 22627
rect 14047 22624 14059 22627
rect 14642 22624 14648 22636
rect 14047 22596 14648 22624
rect 14047 22593 14059 22596
rect 14001 22587 14059 22593
rect 14642 22584 14648 22596
rect 14700 22584 14706 22636
rect 16301 22627 16359 22633
rect 16301 22593 16313 22627
rect 16347 22624 16359 22627
rect 16347 22596 16712 22624
rect 16347 22593 16359 22596
rect 16301 22587 16359 22593
rect 2976 22528 7328 22556
rect 7374 22516 7380 22568
rect 7432 22556 7438 22568
rect 7929 22559 7987 22565
rect 7929 22556 7941 22559
rect 7432 22528 7941 22556
rect 7432 22516 7438 22528
rect 7929 22525 7941 22528
rect 7975 22525 7987 22559
rect 7929 22519 7987 22525
rect 9493 22559 9551 22565
rect 9493 22525 9505 22559
rect 9539 22556 9551 22559
rect 11790 22556 11796 22568
rect 9539 22528 11796 22556
rect 9539 22525 9551 22528
rect 9493 22519 9551 22525
rect 11790 22516 11796 22528
rect 11848 22516 11854 22568
rect 4157 22491 4215 22497
rect 4157 22457 4169 22491
rect 4203 22488 4215 22491
rect 5442 22488 5448 22500
rect 4203 22460 5448 22488
rect 4203 22457 4215 22460
rect 4157 22451 4215 22457
rect 5442 22448 5448 22460
rect 5500 22448 5506 22500
rect 6825 22491 6883 22497
rect 6825 22457 6837 22491
rect 6871 22488 6883 22491
rect 9122 22488 9128 22500
rect 6871 22460 9128 22488
rect 6871 22457 6883 22460
rect 6825 22451 6883 22457
rect 9122 22448 9128 22460
rect 9180 22448 9186 22500
rect 11054 22448 11060 22500
rect 11112 22488 11118 22500
rect 11701 22491 11759 22497
rect 11701 22488 11713 22491
rect 11112 22460 11713 22488
rect 11112 22448 11118 22460
rect 11701 22457 11713 22460
rect 11747 22457 11759 22491
rect 11701 22451 11759 22457
rect 13906 22448 13912 22500
rect 13964 22488 13970 22500
rect 14553 22491 14611 22497
rect 14553 22488 14565 22491
rect 13964 22460 14565 22488
rect 13964 22448 13970 22460
rect 14553 22457 14565 22460
rect 14599 22457 14611 22491
rect 14553 22451 14611 22457
rect 3050 22380 3056 22432
rect 3108 22420 3114 22432
rect 5994 22420 6000 22432
rect 3108 22392 6000 22420
rect 3108 22380 3114 22392
rect 5994 22380 6000 22392
rect 6052 22380 6058 22432
rect 12066 22380 12072 22432
rect 12124 22420 12130 22432
rect 12253 22423 12311 22429
rect 12253 22420 12265 22423
rect 12124 22392 12265 22420
rect 12124 22380 12130 22392
rect 12253 22389 12265 22392
rect 12299 22389 12311 22423
rect 12253 22383 12311 22389
rect 14366 22380 14372 22432
rect 14424 22380 14430 22432
rect 16684 22420 16712 22596
rect 18782 22584 18788 22636
rect 18840 22624 18846 22636
rect 19352 22624 19380 22664
rect 18840 22596 19380 22624
rect 18840 22584 18846 22596
rect 20806 22584 20812 22636
rect 20864 22584 20870 22636
rect 21008 22624 21036 22732
rect 21177 22729 21189 22763
rect 21223 22760 21235 22763
rect 21358 22760 21364 22772
rect 21223 22732 21364 22760
rect 21223 22729 21235 22732
rect 21177 22723 21235 22729
rect 21358 22720 21364 22732
rect 21416 22760 21422 22772
rect 21818 22760 21824 22772
rect 21416 22732 21824 22760
rect 21416 22720 21422 22732
rect 21818 22720 21824 22732
rect 21876 22720 21882 22772
rect 23198 22720 23204 22772
rect 23256 22760 23262 22772
rect 25498 22760 25504 22772
rect 23256 22732 25504 22760
rect 23256 22720 23262 22732
rect 25498 22720 25504 22732
rect 25556 22720 25562 22772
rect 25976 22732 26464 22760
rect 22281 22695 22339 22701
rect 22281 22692 22293 22695
rect 21744 22664 22293 22692
rect 21744 22624 21772 22664
rect 22281 22661 22293 22664
rect 22327 22661 22339 22695
rect 22281 22655 22339 22661
rect 24026 22652 24032 22704
rect 24084 22692 24090 22704
rect 24121 22695 24179 22701
rect 24121 22692 24133 22695
rect 24084 22664 24133 22692
rect 24084 22652 24090 22664
rect 24121 22661 24133 22664
rect 24167 22692 24179 22695
rect 24854 22692 24860 22704
rect 24167 22664 24860 22692
rect 24167 22661 24179 22664
rect 24121 22655 24179 22661
rect 24854 22652 24860 22664
rect 24912 22652 24918 22704
rect 25866 22652 25872 22704
rect 25924 22692 25930 22704
rect 25976 22692 26004 22732
rect 25924 22664 26004 22692
rect 25924 22652 25930 22664
rect 26326 22652 26332 22704
rect 26384 22652 26390 22704
rect 26436 22692 26464 22732
rect 26602 22720 26608 22772
rect 26660 22760 26666 22772
rect 31386 22760 31392 22772
rect 26660 22732 31392 22760
rect 26660 22720 26666 22732
rect 27246 22692 27252 22704
rect 26436 22664 27252 22692
rect 27246 22652 27252 22664
rect 27304 22652 27310 22704
rect 27614 22652 27620 22704
rect 27672 22692 27678 22704
rect 27709 22695 27767 22701
rect 27709 22692 27721 22695
rect 27672 22664 27721 22692
rect 27672 22652 27678 22664
rect 27709 22661 27721 22664
rect 27755 22692 27767 22695
rect 27890 22692 27896 22704
rect 27755 22664 27896 22692
rect 27755 22661 27767 22664
rect 27709 22655 27767 22661
rect 27890 22652 27896 22664
rect 27948 22692 27954 22704
rect 28258 22692 28264 22704
rect 27948 22664 28264 22692
rect 27948 22652 27954 22664
rect 28258 22652 28264 22664
rect 28316 22692 28322 22704
rect 28316 22664 28382 22692
rect 28316 22652 28322 22664
rect 21008 22596 21772 22624
rect 21910 22584 21916 22636
rect 21968 22624 21974 22636
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 21968 22596 22017 22624
rect 21968 22584 21974 22596
rect 22005 22593 22017 22596
rect 22051 22593 22063 22627
rect 24394 22624 24400 22636
rect 23414 22596 24400 22624
rect 22005 22587 22063 22593
rect 24394 22584 24400 22596
rect 24452 22624 24458 22636
rect 24452 22610 25254 22624
rect 24452 22596 25268 22610
rect 24452 22584 24458 22596
rect 16758 22516 16764 22568
rect 16816 22556 16822 22568
rect 16853 22559 16911 22565
rect 16853 22556 16865 22559
rect 16816 22528 16865 22556
rect 16816 22516 16822 22528
rect 16853 22525 16865 22528
rect 16899 22525 16911 22559
rect 16853 22519 16911 22525
rect 17862 22516 17868 22568
rect 17920 22556 17926 22568
rect 18874 22556 18880 22568
rect 17920 22528 18880 22556
rect 17920 22516 17926 22528
rect 18874 22516 18880 22528
rect 18932 22516 18938 22568
rect 19436 22559 19494 22565
rect 19436 22525 19448 22559
rect 19482 22556 19494 22559
rect 19482 22528 19564 22556
rect 19482 22525 19494 22528
rect 19436 22519 19494 22525
rect 18156 22460 19012 22488
rect 18156 22420 18184 22460
rect 16684 22392 18184 22420
rect 18984 22420 19012 22460
rect 19334 22448 19340 22500
rect 19392 22488 19398 22500
rect 19536 22488 19564 22528
rect 19702 22516 19708 22568
rect 19760 22516 19766 22568
rect 23290 22556 23296 22568
rect 20732 22528 23296 22556
rect 19392 22460 19564 22488
rect 19392 22448 19398 22460
rect 20732 22420 20760 22528
rect 23290 22516 23296 22528
rect 23348 22516 23354 22568
rect 23566 22516 23572 22568
rect 23624 22556 23630 22568
rect 24857 22559 24915 22565
rect 24857 22556 24869 22559
rect 23624 22528 24869 22556
rect 23624 22516 23630 22528
rect 24857 22525 24869 22528
rect 24903 22556 24915 22559
rect 25240 22556 25268 22596
rect 26602 22584 26608 22636
rect 26660 22584 26666 22636
rect 29840 22633 29868 22732
rect 31386 22720 31392 22732
rect 31444 22720 31450 22772
rect 32309 22763 32367 22769
rect 32309 22760 32321 22763
rect 31496 22732 32321 22760
rect 30650 22652 30656 22704
rect 30708 22652 30714 22704
rect 30742 22652 30748 22704
rect 30800 22652 30806 22704
rect 27157 22627 27215 22633
rect 27157 22593 27169 22627
rect 27203 22624 27215 22627
rect 29825 22627 29883 22633
rect 27203 22596 28396 22624
rect 27203 22593 27215 22596
rect 27157 22587 27215 22593
rect 28368 22568 28396 22596
rect 29825 22593 29837 22627
rect 29871 22593 29883 22627
rect 29825 22587 29883 22593
rect 30466 22584 30472 22636
rect 30524 22624 30530 22636
rect 31496 22624 31524 22732
rect 32309 22729 32321 22732
rect 32355 22729 32367 22763
rect 32309 22723 32367 22729
rect 32769 22763 32827 22769
rect 32769 22729 32781 22763
rect 32815 22760 32827 22763
rect 34238 22760 34244 22772
rect 32815 22732 34244 22760
rect 32815 22729 32827 22732
rect 32769 22723 32827 22729
rect 34238 22720 34244 22732
rect 34296 22720 34302 22772
rect 34330 22720 34336 22772
rect 34388 22720 34394 22772
rect 35437 22763 35495 22769
rect 35437 22729 35449 22763
rect 35483 22760 35495 22763
rect 35526 22760 35532 22772
rect 35483 22732 35532 22760
rect 35483 22729 35495 22732
rect 35437 22723 35495 22729
rect 35526 22720 35532 22732
rect 35584 22720 35590 22772
rect 37458 22720 37464 22772
rect 37516 22720 37522 22772
rect 37642 22720 37648 22772
rect 37700 22760 37706 22772
rect 38562 22760 38568 22772
rect 37700 22732 38568 22760
rect 37700 22720 37706 22732
rect 38562 22720 38568 22732
rect 38620 22720 38626 22772
rect 38746 22720 38752 22772
rect 38804 22760 38810 22772
rect 40497 22763 40555 22769
rect 38804 22732 39804 22760
rect 38804 22720 38810 22732
rect 33594 22692 33600 22704
rect 31680 22664 33600 22692
rect 31680 22633 31708 22664
rect 33594 22652 33600 22664
rect 33652 22652 33658 22704
rect 34348 22692 34376 22720
rect 33704 22664 34376 22692
rect 30524 22596 31524 22624
rect 31665 22627 31723 22633
rect 30524 22584 30530 22596
rect 31665 22593 31677 22627
rect 31711 22593 31723 22627
rect 31665 22587 31723 22593
rect 32677 22627 32735 22633
rect 32677 22593 32689 22627
rect 32723 22624 32735 22627
rect 32766 22624 32772 22636
rect 32723 22596 32772 22624
rect 32723 22593 32735 22596
rect 32677 22587 32735 22593
rect 32766 22584 32772 22596
rect 32824 22584 32830 22636
rect 33410 22584 33416 22636
rect 33468 22584 33474 22636
rect 33704 22633 33732 22664
rect 34606 22652 34612 22704
rect 34664 22652 34670 22704
rect 33689 22627 33747 22633
rect 33689 22593 33701 22627
rect 33735 22593 33747 22627
rect 33689 22587 33747 22593
rect 35250 22584 35256 22636
rect 35308 22624 35314 22636
rect 36449 22627 36507 22633
rect 36449 22624 36461 22627
rect 35308 22596 36461 22624
rect 35308 22584 35314 22596
rect 36449 22593 36461 22596
rect 36495 22593 36507 22627
rect 36449 22587 36507 22593
rect 25774 22556 25780 22568
rect 24903 22528 25176 22556
rect 25240 22528 25780 22556
rect 24903 22525 24915 22528
rect 24857 22519 24915 22525
rect 21818 22448 21824 22500
rect 21876 22488 21882 22500
rect 23753 22491 23811 22497
rect 21876 22460 22094 22488
rect 21876 22448 21882 22460
rect 18984 22392 20760 22420
rect 20806 22380 20812 22432
rect 20864 22420 20870 22432
rect 21634 22420 21640 22432
rect 20864 22392 21640 22420
rect 20864 22380 20870 22392
rect 21634 22380 21640 22392
rect 21692 22380 21698 22432
rect 22066 22420 22094 22460
rect 23753 22457 23765 22491
rect 23799 22488 23811 22491
rect 24210 22488 24216 22500
rect 23799 22460 24216 22488
rect 23799 22457 23811 22460
rect 23753 22451 23811 22457
rect 24210 22448 24216 22460
rect 24268 22448 24274 22500
rect 24946 22488 24952 22500
rect 24320 22460 24952 22488
rect 24320 22420 24348 22460
rect 24946 22448 24952 22460
rect 25004 22448 25010 22500
rect 22066 22392 24348 22420
rect 24486 22380 24492 22432
rect 24544 22380 24550 22432
rect 25148 22420 25176 22528
rect 25774 22516 25780 22528
rect 25832 22516 25838 22568
rect 27246 22516 27252 22568
rect 27304 22556 27310 22568
rect 27614 22556 27620 22568
rect 27304 22528 27620 22556
rect 27304 22516 27310 22528
rect 27614 22516 27620 22528
rect 27672 22516 27678 22568
rect 27706 22516 27712 22568
rect 27764 22556 27770 22568
rect 28074 22556 28080 22568
rect 27764 22528 28080 22556
rect 27764 22516 27770 22528
rect 28074 22516 28080 22528
rect 28132 22516 28138 22568
rect 28350 22516 28356 22568
rect 28408 22516 28414 22568
rect 29178 22516 29184 22568
rect 29236 22556 29242 22568
rect 29549 22559 29607 22565
rect 29549 22556 29561 22559
rect 29236 22528 29561 22556
rect 29236 22516 29242 22528
rect 29549 22525 29561 22528
rect 29595 22556 29607 22559
rect 29595 22528 29868 22556
rect 29595 22525 29607 22528
rect 29549 22519 29607 22525
rect 27338 22448 27344 22500
rect 27396 22448 27402 22500
rect 29840 22488 29868 22528
rect 29914 22516 29920 22568
rect 29972 22556 29978 22568
rect 30837 22559 30895 22565
rect 30837 22556 30849 22559
rect 29972 22528 30849 22556
rect 29972 22516 29978 22528
rect 30837 22525 30849 22528
rect 30883 22525 30895 22559
rect 32861 22559 32919 22565
rect 30837 22519 30895 22525
rect 30944 22528 31754 22556
rect 30944 22488 30972 22528
rect 29840 22460 30972 22488
rect 31018 22448 31024 22500
rect 31076 22488 31082 22500
rect 31726 22488 31754 22528
rect 32861 22525 32873 22559
rect 32907 22525 32919 22559
rect 32861 22519 32919 22525
rect 32876 22488 32904 22519
rect 31076 22460 31616 22488
rect 31726 22460 32904 22488
rect 31076 22448 31082 22460
rect 26326 22420 26332 22432
rect 25148 22392 26332 22420
rect 26326 22380 26332 22392
rect 26384 22380 26390 22432
rect 26602 22380 26608 22432
rect 26660 22420 26666 22432
rect 30285 22423 30343 22429
rect 30285 22420 30297 22423
rect 26660 22392 30297 22420
rect 26660 22380 26666 22392
rect 30285 22389 30297 22392
rect 30331 22389 30343 22423
rect 30285 22383 30343 22389
rect 30374 22380 30380 22432
rect 30432 22420 30438 22432
rect 31110 22420 31116 22432
rect 30432 22392 31116 22420
rect 30432 22380 30438 22392
rect 31110 22380 31116 22392
rect 31168 22380 31174 22432
rect 31478 22380 31484 22432
rect 31536 22380 31542 22432
rect 31588 22420 31616 22460
rect 33428 22420 33456 22584
rect 33502 22516 33508 22568
rect 33560 22556 33566 22568
rect 33965 22559 34023 22565
rect 33965 22556 33977 22559
rect 33560 22528 33977 22556
rect 33560 22516 33566 22528
rect 33965 22525 33977 22528
rect 34011 22525 34023 22559
rect 33965 22519 34023 22525
rect 34054 22516 34060 22568
rect 34112 22556 34118 22568
rect 36541 22559 36599 22565
rect 36541 22556 36553 22559
rect 34112 22528 36553 22556
rect 34112 22516 34118 22528
rect 36541 22525 36553 22528
rect 36587 22525 36599 22559
rect 36541 22519 36599 22525
rect 36725 22559 36783 22565
rect 36725 22525 36737 22559
rect 36771 22556 36783 22559
rect 37476 22556 37504 22720
rect 38654 22692 38660 22704
rect 38502 22664 38660 22692
rect 38654 22652 38660 22664
rect 38712 22652 38718 22704
rect 38838 22652 38844 22704
rect 38896 22692 38902 22704
rect 38933 22695 38991 22701
rect 38933 22692 38945 22695
rect 38896 22664 38945 22692
rect 38896 22652 38902 22664
rect 38933 22661 38945 22664
rect 38979 22661 38991 22695
rect 38933 22655 38991 22661
rect 39209 22627 39267 22633
rect 39209 22593 39221 22627
rect 39255 22624 39267 22627
rect 39482 22624 39488 22636
rect 39255 22596 39488 22624
rect 39255 22593 39267 22596
rect 39209 22587 39267 22593
rect 39482 22584 39488 22596
rect 39540 22584 39546 22636
rect 39776 22633 39804 22732
rect 40497 22729 40509 22763
rect 40543 22760 40555 22763
rect 46385 22763 46443 22769
rect 40543 22732 41828 22760
rect 40543 22729 40555 22732
rect 40497 22723 40555 22729
rect 40405 22695 40463 22701
rect 40405 22661 40417 22695
rect 40451 22692 40463 22695
rect 40586 22692 40592 22704
rect 40451 22664 40592 22692
rect 40451 22661 40463 22664
rect 40405 22655 40463 22661
rect 40586 22652 40592 22664
rect 40644 22652 40650 22704
rect 41800 22692 41828 22732
rect 46385 22729 46397 22763
rect 46431 22760 46443 22763
rect 48682 22760 48688 22772
rect 46431 22732 48688 22760
rect 46431 22729 46443 22732
rect 46385 22723 46443 22729
rect 48682 22720 48688 22732
rect 48740 22720 48746 22772
rect 46106 22692 46112 22704
rect 41800 22664 46112 22692
rect 46106 22652 46112 22664
rect 46164 22652 46170 22704
rect 46750 22652 46756 22704
rect 46808 22692 46814 22704
rect 47581 22695 47639 22701
rect 47581 22692 47593 22695
rect 46808 22664 47593 22692
rect 46808 22652 46814 22664
rect 39761 22627 39819 22633
rect 39761 22593 39773 22627
rect 39807 22624 39819 22627
rect 40678 22624 40684 22636
rect 39807 22596 40684 22624
rect 39807 22593 39819 22596
rect 39761 22587 39819 22593
rect 40678 22584 40684 22596
rect 40736 22584 40742 22636
rect 41414 22584 41420 22636
rect 41472 22584 41478 22636
rect 42058 22584 42064 22636
rect 42116 22584 42122 22636
rect 43990 22584 43996 22636
rect 44048 22624 44054 22636
rect 44085 22627 44143 22633
rect 44085 22624 44097 22627
rect 44048 22596 44097 22624
rect 44048 22584 44054 22596
rect 44085 22593 44097 22596
rect 44131 22593 44143 22627
rect 44085 22587 44143 22593
rect 44726 22584 44732 22636
rect 44784 22584 44790 22636
rect 45278 22584 45284 22636
rect 45336 22624 45342 22636
rect 47228 22633 47256 22664
rect 47581 22661 47593 22664
rect 47627 22661 47639 22695
rect 47581 22655 47639 22661
rect 45373 22627 45431 22633
rect 45373 22624 45385 22627
rect 45336 22596 45385 22624
rect 45336 22584 45342 22596
rect 45373 22593 45385 22596
rect 45419 22624 45431 22627
rect 45649 22627 45707 22633
rect 45649 22624 45661 22627
rect 45419 22596 45661 22624
rect 45419 22593 45431 22596
rect 45373 22587 45431 22593
rect 45649 22593 45661 22596
rect 45695 22593 45707 22627
rect 45649 22587 45707 22593
rect 47213 22627 47271 22633
rect 47213 22593 47225 22627
rect 47259 22624 47271 22627
rect 47259 22596 47293 22624
rect 47259 22593 47271 22596
rect 47213 22587 47271 22593
rect 47762 22584 47768 22636
rect 47820 22624 47826 22636
rect 48593 22627 48651 22633
rect 48593 22624 48605 22627
rect 47820 22596 48605 22624
rect 47820 22584 47826 22596
rect 48593 22593 48605 22596
rect 48639 22593 48651 22627
rect 48593 22587 48651 22593
rect 49326 22584 49332 22636
rect 49384 22584 49390 22636
rect 40589 22559 40647 22565
rect 40589 22556 40601 22559
rect 36771 22528 37504 22556
rect 37568 22528 40601 22556
rect 36771 22525 36783 22528
rect 36725 22519 36783 22525
rect 36081 22491 36139 22497
rect 36081 22488 36093 22491
rect 35084 22460 36093 22488
rect 31588 22392 33456 22420
rect 34146 22380 34152 22432
rect 34204 22420 34210 22432
rect 35084 22420 35112 22460
rect 36081 22457 36093 22460
rect 36127 22457 36139 22491
rect 36081 22451 36139 22457
rect 36354 22448 36360 22500
rect 36412 22488 36418 22500
rect 37090 22488 37096 22500
rect 36412 22460 37096 22488
rect 36412 22448 36418 22460
rect 37090 22448 37096 22460
rect 37148 22488 37154 22500
rect 37568 22488 37596 22528
rect 40589 22525 40601 22528
rect 40635 22525 40647 22559
rect 40589 22519 40647 22525
rect 42610 22516 42616 22568
rect 42668 22516 42674 22568
rect 42889 22559 42947 22565
rect 42889 22525 42901 22559
rect 42935 22556 42947 22559
rect 43438 22556 43444 22568
rect 42935 22528 43444 22556
rect 42935 22525 42947 22528
rect 42889 22519 42947 22525
rect 43438 22516 43444 22528
rect 43496 22516 43502 22568
rect 46753 22559 46811 22565
rect 46753 22525 46765 22559
rect 46799 22556 46811 22559
rect 49344 22556 49372 22584
rect 46799 22528 49372 22556
rect 46799 22525 46811 22528
rect 46753 22519 46811 22525
rect 37148 22460 37596 22488
rect 37148 22448 37154 22460
rect 41874 22448 41880 22500
rect 41932 22448 41938 22500
rect 45186 22448 45192 22500
rect 45244 22448 45250 22500
rect 46569 22491 46627 22497
rect 46569 22457 46581 22491
rect 46615 22488 46627 22491
rect 46615 22460 47532 22488
rect 46615 22457 46627 22460
rect 46569 22451 46627 22457
rect 34204 22392 35112 22420
rect 34204 22380 34210 22392
rect 35158 22380 35164 22432
rect 35216 22420 35222 22432
rect 35805 22423 35863 22429
rect 35805 22420 35817 22423
rect 35216 22392 35817 22420
rect 35216 22380 35222 22392
rect 35805 22389 35817 22392
rect 35851 22420 35863 22423
rect 37550 22420 37556 22432
rect 35851 22392 37556 22420
rect 35851 22389 35863 22392
rect 35805 22383 35863 22389
rect 37550 22380 37556 22392
rect 37608 22380 37614 22432
rect 38746 22380 38752 22432
rect 38804 22420 38810 22432
rect 39114 22420 39120 22432
rect 38804 22392 39120 22420
rect 38804 22380 38810 22392
rect 39114 22380 39120 22392
rect 39172 22380 39178 22432
rect 40034 22380 40040 22432
rect 40092 22380 40098 22432
rect 41230 22380 41236 22432
rect 41288 22380 41294 22432
rect 43898 22380 43904 22432
rect 43956 22380 43962 22432
rect 44542 22380 44548 22432
rect 44600 22380 44606 22432
rect 45370 22380 45376 22432
rect 45428 22420 45434 22432
rect 45833 22423 45891 22429
rect 45833 22420 45845 22423
rect 45428 22392 45845 22420
rect 45428 22380 45434 22392
rect 45833 22389 45845 22392
rect 45879 22389 45891 22423
rect 45833 22383 45891 22389
rect 46934 22380 46940 22432
rect 46992 22420 46998 22432
rect 47029 22423 47087 22429
rect 47029 22420 47041 22423
rect 46992 22392 47041 22420
rect 46992 22380 46998 22392
rect 47029 22389 47041 22392
rect 47075 22389 47087 22423
rect 47504 22420 47532 22460
rect 47578 22448 47584 22500
rect 47636 22488 47642 22500
rect 47949 22491 48007 22497
rect 47949 22488 47961 22491
rect 47636 22460 47961 22488
rect 47636 22448 47642 22460
rect 47949 22457 47961 22460
rect 47995 22457 48007 22491
rect 49234 22488 49240 22500
rect 47949 22451 48007 22457
rect 48240 22460 49240 22488
rect 48240 22420 48268 22460
rect 49234 22448 49240 22460
rect 49292 22448 49298 22500
rect 47504 22392 48268 22420
rect 47029 22383 47087 22389
rect 48314 22380 48320 22432
rect 48372 22420 48378 22432
rect 48409 22423 48467 22429
rect 48409 22420 48421 22423
rect 48372 22392 48421 22420
rect 48372 22380 48378 22392
rect 48409 22389 48421 22392
rect 48455 22389 48467 22423
rect 48409 22383 48467 22389
rect 48682 22380 48688 22432
rect 48740 22420 48746 22432
rect 49145 22423 49203 22429
rect 49145 22420 49157 22423
rect 48740 22392 49157 22420
rect 48740 22380 48746 22392
rect 49145 22389 49157 22392
rect 49191 22389 49203 22423
rect 49145 22383 49203 22389
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 2222 22176 2228 22228
rect 2280 22216 2286 22228
rect 4246 22216 4252 22228
rect 2280 22188 4252 22216
rect 2280 22176 2286 22188
rect 4246 22176 4252 22188
rect 4304 22176 4310 22228
rect 11882 22176 11888 22228
rect 11940 22216 11946 22228
rect 12345 22219 12403 22225
rect 12345 22216 12357 22219
rect 11940 22188 12357 22216
rect 11940 22176 11946 22188
rect 12345 22185 12357 22188
rect 12391 22185 12403 22219
rect 12345 22179 12403 22185
rect 13648 22188 15240 22216
rect 2866 22108 2872 22160
rect 2924 22148 2930 22160
rect 2924 22120 6040 22148
rect 2924 22108 2930 22120
rect 6012 22094 6040 22120
rect 7098 22108 7104 22160
rect 7156 22148 7162 22160
rect 7834 22148 7840 22160
rect 7156 22120 7840 22148
rect 7156 22108 7162 22120
rect 7834 22108 7840 22120
rect 7892 22108 7898 22160
rect 10226 22108 10232 22160
rect 10284 22148 10290 22160
rect 10284 22120 13400 22148
rect 10284 22108 10290 22120
rect 6012 22089 6077 22094
rect 5997 22083 6077 22089
rect 2976 22052 5488 22080
rect 2976 22021 3004 22052
rect 2961 22015 3019 22021
rect 2961 21981 2973 22015
rect 3007 21981 3019 22015
rect 2961 21975 3019 21981
rect 5353 22015 5411 22021
rect 5353 21981 5365 22015
rect 5399 21981 5411 22015
rect 5460 22012 5488 22052
rect 5997 22049 6009 22083
rect 6043 22066 6077 22083
rect 9674 22080 9680 22092
rect 6043 22049 6055 22066
rect 5997 22043 6055 22049
rect 7852 22052 9680 22080
rect 6730 22012 6736 22024
rect 5460 21984 6736 22012
rect 5353 21975 5411 21981
rect 1026 21904 1032 21956
rect 1084 21944 1090 21956
rect 1765 21947 1823 21953
rect 1765 21944 1777 21947
rect 1084 21916 1777 21944
rect 1084 21904 1090 21916
rect 1765 21913 1777 21916
rect 1811 21913 1823 21947
rect 1765 21907 1823 21913
rect 3234 21904 3240 21956
rect 3292 21944 3298 21956
rect 4157 21947 4215 21953
rect 4157 21944 4169 21947
rect 3292 21916 4169 21944
rect 3292 21904 3298 21916
rect 4157 21913 4169 21916
rect 4203 21913 4215 21947
rect 4157 21907 4215 21913
rect 5368 21876 5396 21975
rect 6730 21972 6736 21984
rect 6788 21972 6794 22024
rect 7193 22015 7251 22021
rect 7193 21981 7205 22015
rect 7239 22012 7251 22015
rect 7742 22012 7748 22024
rect 7239 21984 7748 22012
rect 7239 21981 7251 21984
rect 7193 21975 7251 21981
rect 7742 21972 7748 21984
rect 7800 21972 7806 22024
rect 7852 22021 7880 22052
rect 9674 22040 9680 22052
rect 9732 22040 9738 22092
rect 9766 22040 9772 22092
rect 9824 22040 9830 22092
rect 11882 22040 11888 22092
rect 11940 22040 11946 22092
rect 7837 22015 7895 22021
rect 7837 21981 7849 22015
rect 7883 21981 7895 22015
rect 7837 21975 7895 21981
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 22012 8631 22015
rect 8619 21984 9076 22012
rect 8619 21981 8631 21984
rect 8573 21975 8631 21981
rect 5626 21904 5632 21956
rect 5684 21944 5690 21956
rect 7653 21947 7711 21953
rect 7653 21944 7665 21947
rect 5684 21916 7665 21944
rect 5684 21904 5690 21916
rect 7653 21913 7665 21916
rect 7699 21913 7711 21947
rect 7653 21907 7711 21913
rect 8312 21916 8524 21944
rect 8312 21876 8340 21916
rect 5368 21848 8340 21876
rect 8386 21836 8392 21888
rect 8444 21836 8450 21888
rect 8496 21876 8524 21916
rect 8938 21876 8944 21888
rect 8496 21848 8944 21876
rect 8938 21836 8944 21848
rect 8996 21836 9002 21888
rect 9048 21876 9076 21984
rect 9122 21972 9128 22024
rect 9180 21972 9186 22024
rect 11609 22015 11667 22021
rect 11609 21981 11621 22015
rect 11655 22012 11667 22015
rect 11655 21984 12434 22012
rect 11655 21981 11667 21984
rect 11609 21975 11667 21981
rect 12406 21944 12434 21984
rect 12526 21972 12532 22024
rect 12584 21972 12590 22024
rect 13372 22021 13400 22120
rect 13648 22089 13676 22188
rect 14182 22108 14188 22160
rect 14240 22148 14246 22160
rect 14366 22148 14372 22160
rect 14240 22120 14372 22148
rect 14240 22108 14246 22120
rect 14366 22108 14372 22120
rect 14424 22148 14430 22160
rect 15102 22148 15108 22160
rect 14424 22120 15108 22148
rect 14424 22108 14430 22120
rect 15102 22108 15108 22120
rect 15160 22108 15166 22160
rect 15212 22092 15240 22188
rect 19610 22176 19616 22228
rect 19668 22216 19674 22228
rect 22186 22216 22192 22228
rect 19668 22188 22192 22216
rect 19668 22176 19674 22188
rect 22186 22176 22192 22188
rect 22244 22176 22250 22228
rect 24670 22176 24676 22228
rect 24728 22216 24734 22228
rect 25593 22219 25651 22225
rect 25593 22216 25605 22219
rect 24728 22188 25605 22216
rect 24728 22176 24734 22188
rect 25593 22185 25605 22188
rect 25639 22185 25651 22219
rect 25593 22179 25651 22185
rect 15654 22148 15660 22160
rect 15304 22120 15660 22148
rect 13633 22083 13691 22089
rect 13633 22049 13645 22083
rect 13679 22080 13691 22083
rect 13679 22052 13713 22080
rect 13679 22049 13691 22052
rect 13633 22043 13691 22049
rect 14274 22040 14280 22092
rect 14332 22080 14338 22092
rect 14461 22083 14519 22089
rect 14461 22080 14473 22083
rect 14332 22052 14473 22080
rect 14332 22040 14338 22052
rect 14461 22049 14473 22052
rect 14507 22049 14519 22083
rect 14461 22043 14519 22049
rect 15194 22040 15200 22092
rect 15252 22040 15258 22092
rect 13357 22015 13415 22021
rect 13357 21981 13369 22015
rect 13403 21981 13415 22015
rect 13357 21975 13415 21981
rect 13449 22015 13507 22021
rect 13449 21981 13461 22015
rect 13495 22012 13507 22015
rect 15304 22012 15332 22120
rect 15654 22108 15660 22120
rect 15712 22108 15718 22160
rect 17034 22108 17040 22160
rect 17092 22148 17098 22160
rect 17092 22120 17632 22148
rect 17092 22108 17098 22120
rect 15378 22040 15384 22092
rect 15436 22080 15442 22092
rect 17604 22089 17632 22120
rect 20162 22108 20168 22160
rect 20220 22148 20226 22160
rect 24581 22151 24639 22157
rect 20220 22120 22048 22148
rect 20220 22108 20226 22120
rect 16945 22083 17003 22089
rect 16945 22080 16957 22083
rect 15436 22052 16957 22080
rect 15436 22040 15442 22052
rect 16945 22049 16957 22052
rect 16991 22049 17003 22083
rect 16945 22043 17003 22049
rect 17589 22083 17647 22089
rect 17589 22049 17601 22083
rect 17635 22049 17647 22083
rect 17589 22043 17647 22049
rect 17788 22052 18920 22080
rect 13495 21984 15332 22012
rect 13495 21981 13507 21984
rect 13449 21975 13507 21981
rect 17126 21972 17132 22024
rect 17184 22012 17190 22024
rect 17788 22012 17816 22052
rect 17184 21984 17816 22012
rect 18785 22015 18843 22021
rect 17184 21972 17190 21984
rect 18785 21981 18797 22015
rect 18831 21981 18843 22015
rect 18892 22012 18920 22052
rect 18966 22040 18972 22092
rect 19024 22080 19030 22092
rect 22020 22089 22048 22120
rect 24581 22117 24593 22151
rect 24627 22148 24639 22151
rect 24854 22148 24860 22160
rect 24627 22120 24661 22148
rect 24780 22120 24860 22148
rect 24627 22117 24639 22120
rect 24581 22111 24639 22117
rect 19889 22083 19947 22089
rect 19889 22080 19901 22083
rect 19024 22052 19901 22080
rect 19024 22040 19030 22052
rect 19889 22049 19901 22052
rect 19935 22049 19947 22083
rect 19889 22043 19947 22049
rect 22005 22083 22063 22089
rect 22005 22049 22017 22083
rect 22051 22049 22063 22083
rect 22005 22043 22063 22049
rect 22738 22040 22744 22092
rect 22796 22080 22802 22092
rect 23201 22083 23259 22089
rect 23201 22080 23213 22083
rect 22796 22052 23213 22080
rect 22796 22040 22802 22052
rect 23201 22049 23213 22052
rect 23247 22080 23259 22083
rect 23566 22080 23572 22092
rect 23247 22052 23572 22080
rect 23247 22049 23259 22052
rect 23201 22043 23259 22049
rect 23566 22040 23572 22052
rect 23624 22040 23630 22092
rect 23658 22040 23664 22092
rect 23716 22080 23722 22092
rect 24596 22080 24624 22111
rect 23716 22052 24624 22080
rect 24780 22080 24808 22120
rect 24854 22108 24860 22120
rect 24912 22108 24918 22160
rect 24946 22108 24952 22160
rect 25004 22108 25010 22160
rect 24964 22080 24992 22108
rect 25133 22083 25191 22089
rect 25133 22080 25145 22083
rect 24780 22052 24900 22080
rect 24964 22052 25145 22080
rect 23716 22040 23722 22052
rect 19242 22012 19248 22024
rect 18892 21984 19248 22012
rect 18785 21975 18843 21981
rect 12406 21916 14596 21944
rect 12989 21879 13047 21885
rect 12989 21876 13001 21879
rect 9048 21848 13001 21876
rect 12989 21845 13001 21848
rect 13035 21845 13047 21879
rect 14568 21876 14596 21916
rect 14642 21904 14648 21956
rect 14700 21904 14706 21956
rect 16114 21904 16120 21956
rect 16172 21904 16178 21956
rect 16666 21904 16672 21956
rect 16724 21904 16730 21956
rect 18800 21944 18828 21975
rect 19242 21972 19248 21984
rect 19300 21972 19306 22024
rect 19426 21972 19432 22024
rect 19484 21972 19490 22024
rect 22554 22012 22560 22024
rect 19904 21984 22560 22012
rect 19904 21944 19932 21984
rect 22554 21972 22560 21984
rect 22612 21972 22618 22024
rect 24026 21972 24032 22024
rect 24084 21972 24090 22024
rect 24872 22012 24900 22052
rect 25133 22049 25145 22052
rect 25179 22080 25191 22083
rect 25406 22080 25412 22092
rect 25179 22052 25412 22080
rect 25179 22049 25191 22052
rect 25133 22043 25191 22049
rect 25406 22040 25412 22052
rect 25464 22040 25470 22092
rect 25041 22015 25099 22021
rect 25041 22012 25053 22015
rect 24872 21984 25053 22012
rect 25041 21981 25053 21984
rect 25087 22012 25099 22015
rect 25314 22012 25320 22024
rect 25087 21984 25320 22012
rect 25087 21981 25099 21984
rect 25041 21975 25099 21981
rect 25314 21972 25320 21984
rect 25372 21972 25378 22024
rect 25608 22012 25636 22179
rect 28258 22176 28264 22228
rect 28316 22216 28322 22228
rect 28353 22219 28411 22225
rect 28353 22216 28365 22219
rect 28316 22188 28365 22216
rect 28316 22176 28322 22188
rect 28353 22185 28365 22188
rect 28399 22185 28411 22219
rect 28718 22216 28724 22228
rect 28353 22179 28411 22185
rect 28460 22188 28724 22216
rect 26694 22108 26700 22160
rect 26752 22148 26758 22160
rect 28460 22148 28488 22188
rect 28718 22176 28724 22188
rect 28776 22176 28782 22228
rect 30190 22176 30196 22228
rect 30248 22216 30254 22228
rect 30285 22219 30343 22225
rect 30285 22216 30297 22219
rect 30248 22188 30297 22216
rect 30248 22176 30254 22188
rect 30285 22185 30297 22188
rect 30331 22216 30343 22219
rect 31846 22216 31852 22228
rect 30331 22188 31852 22216
rect 30331 22185 30343 22188
rect 30285 22179 30343 22185
rect 31846 22176 31852 22188
rect 31904 22176 31910 22228
rect 32766 22176 32772 22228
rect 32824 22216 32830 22228
rect 35434 22216 35440 22228
rect 32824 22188 35440 22216
rect 32824 22176 32830 22188
rect 35434 22176 35440 22188
rect 35492 22176 35498 22228
rect 35526 22176 35532 22228
rect 35584 22176 35590 22228
rect 38654 22216 38660 22228
rect 36280 22188 38660 22216
rect 35544 22148 35572 22176
rect 26752 22120 28488 22148
rect 33704 22120 35572 22148
rect 26752 22108 26758 22120
rect 26326 22040 26332 22092
rect 26384 22080 26390 22092
rect 26513 22083 26571 22089
rect 26513 22080 26525 22083
rect 26384 22052 26525 22080
rect 26384 22040 26390 22052
rect 26513 22049 26525 22052
rect 26559 22049 26571 22083
rect 26513 22043 26571 22049
rect 27614 22040 27620 22092
rect 27672 22040 27678 22092
rect 27706 22040 27712 22092
rect 27764 22040 27770 22092
rect 28074 22040 28080 22092
rect 28132 22080 28138 22092
rect 28902 22080 28908 22092
rect 28132 22052 28908 22080
rect 28132 22040 28138 22052
rect 28902 22040 28908 22052
rect 28960 22040 28966 22092
rect 29546 22040 29552 22092
rect 29604 22080 29610 22092
rect 30558 22080 30564 22092
rect 29604 22052 30564 22080
rect 29604 22040 29610 22052
rect 30558 22040 30564 22052
rect 30616 22040 30622 22092
rect 31478 22080 31484 22092
rect 30852 22052 31484 22080
rect 30852 22024 30880 22052
rect 31478 22040 31484 22052
rect 31536 22040 31542 22092
rect 32306 22040 32312 22092
rect 32364 22080 32370 22092
rect 33704 22089 33732 22120
rect 33505 22083 33563 22089
rect 33505 22080 33517 22083
rect 32364 22052 33517 22080
rect 32364 22040 32370 22052
rect 33505 22049 33517 22052
rect 33551 22049 33563 22083
rect 33505 22043 33563 22049
rect 33689 22083 33747 22089
rect 33689 22049 33701 22083
rect 33735 22080 33747 22083
rect 33735 22052 33769 22080
rect 33735 22049 33747 22052
rect 33689 22043 33747 22049
rect 33870 22040 33876 22092
rect 33928 22080 33934 22092
rect 34790 22080 34796 22092
rect 33928 22052 34796 22080
rect 33928 22040 33934 22052
rect 34790 22040 34796 22052
rect 34848 22040 34854 22092
rect 34974 22040 34980 22092
rect 35032 22040 35038 22092
rect 36280 22089 36308 22188
rect 38654 22176 38660 22188
rect 38712 22176 38718 22228
rect 38838 22176 38844 22228
rect 38896 22216 38902 22228
rect 38896 22188 39068 22216
rect 38896 22176 38902 22188
rect 39040 22148 39068 22188
rect 39482 22176 39488 22228
rect 39540 22176 39546 22228
rect 40218 22176 40224 22228
rect 40276 22176 40282 22228
rect 41046 22176 41052 22228
rect 41104 22216 41110 22228
rect 42702 22216 42708 22228
rect 41104 22188 42708 22216
rect 41104 22176 41110 22188
rect 42702 22176 42708 22188
rect 42760 22216 42766 22228
rect 43530 22216 43536 22228
rect 42760 22188 43536 22216
rect 42760 22176 42766 22188
rect 43530 22176 43536 22188
rect 43588 22176 43594 22228
rect 44082 22176 44088 22228
rect 44140 22216 44146 22228
rect 44729 22219 44787 22225
rect 44729 22216 44741 22219
rect 44140 22188 44741 22216
rect 44140 22176 44146 22188
rect 44729 22185 44741 22188
rect 44775 22185 44787 22219
rect 44729 22179 44787 22185
rect 47026 22176 47032 22228
rect 47084 22176 47090 22228
rect 47213 22219 47271 22225
rect 47213 22185 47225 22219
rect 47259 22216 47271 22219
rect 49418 22216 49424 22228
rect 47259 22188 49424 22216
rect 47259 22185 47271 22188
rect 47213 22179 47271 22185
rect 49418 22176 49424 22188
rect 49476 22176 49482 22228
rect 43714 22148 43720 22160
rect 39040 22120 42012 22148
rect 36265 22083 36323 22089
rect 36265 22049 36277 22083
rect 36311 22049 36323 22083
rect 36265 22043 36323 22049
rect 38838 22040 38844 22092
rect 38896 22040 38902 22092
rect 39117 22083 39175 22089
rect 39117 22049 39129 22083
rect 39163 22080 39175 22083
rect 39163 22052 39252 22080
rect 39163 22049 39175 22052
rect 39117 22043 39175 22049
rect 26421 22015 26479 22021
rect 25608 21984 26372 22012
rect 26344 21956 26372 21984
rect 26421 21981 26433 22015
rect 26467 22012 26479 22015
rect 26602 22012 26608 22024
rect 26467 21984 26608 22012
rect 26467 21981 26479 21984
rect 26421 21975 26479 21981
rect 26602 21972 26608 21984
rect 26660 21972 26666 22024
rect 27525 22015 27583 22021
rect 27525 21981 27537 22015
rect 27571 22012 27583 22015
rect 27798 22012 27804 22024
rect 27571 21984 27804 22012
rect 27571 21981 27583 21984
rect 27525 21975 27583 21981
rect 27798 21972 27804 21984
rect 27856 22012 27862 22024
rect 29822 22012 29828 22024
rect 27856 21984 29828 22012
rect 27856 21972 27862 21984
rect 29822 21972 29828 21984
rect 29880 21972 29886 22024
rect 29917 22015 29975 22021
rect 29917 21981 29929 22015
rect 29963 22012 29975 22015
rect 30650 22012 30656 22024
rect 29963 21984 30656 22012
rect 29963 21981 29975 21984
rect 29917 21975 29975 21981
rect 30650 21972 30656 21984
rect 30708 21972 30714 22024
rect 30834 21972 30840 22024
rect 30892 21972 30898 22024
rect 32122 21972 32128 22024
rect 32180 22012 32186 22024
rect 34057 22015 34115 22021
rect 34057 22012 34069 22015
rect 32180 21984 34069 22012
rect 32180 21972 32186 21984
rect 34057 21981 34069 21984
rect 34103 22012 34115 22015
rect 34425 22015 34483 22021
rect 34425 22012 34437 22015
rect 34103 21984 34437 22012
rect 34103 21981 34115 21984
rect 34057 21975 34115 21981
rect 34425 21981 34437 21984
rect 34471 21981 34483 22015
rect 39224 22012 39252 22052
rect 39390 22040 39396 22092
rect 39448 22080 39454 22092
rect 40880 22089 40908 22120
rect 41984 22089 42012 22120
rect 42536 22120 43720 22148
rect 40865 22083 40923 22089
rect 39448 22052 39712 22080
rect 39448 22040 39454 22052
rect 39574 22012 39580 22024
rect 34425 21975 34483 21981
rect 35176 21984 36400 22012
rect 39224 21984 39580 22012
rect 18800 21916 19932 21944
rect 21177 21947 21235 21953
rect 21177 21913 21189 21947
rect 21223 21944 21235 21947
rect 21542 21944 21548 21956
rect 21223 21916 21548 21944
rect 21223 21913 21235 21916
rect 21177 21907 21235 21913
rect 21542 21904 21548 21916
rect 21600 21904 21606 21956
rect 21821 21947 21879 21953
rect 21821 21913 21833 21947
rect 21867 21944 21879 21947
rect 22922 21944 22928 21956
rect 21867 21916 22928 21944
rect 21867 21913 21879 21916
rect 21821 21907 21879 21913
rect 22922 21904 22928 21916
rect 22980 21904 22986 21956
rect 23017 21947 23075 21953
rect 23017 21913 23029 21947
rect 23063 21944 23075 21947
rect 24578 21944 24584 21956
rect 23063 21916 24584 21944
rect 23063 21913 23075 21916
rect 23017 21907 23075 21913
rect 24578 21904 24584 21916
rect 24636 21904 24642 21956
rect 24946 21904 24952 21956
rect 25004 21944 25010 21956
rect 26050 21944 26056 21956
rect 25004 21916 26056 21944
rect 25004 21904 25010 21916
rect 26050 21904 26056 21916
rect 26108 21904 26114 21956
rect 26326 21904 26332 21956
rect 26384 21904 26390 21956
rect 28813 21947 28871 21953
rect 28813 21913 28825 21947
rect 28859 21944 28871 21947
rect 30466 21944 30472 21956
rect 28859 21916 30472 21944
rect 28859 21913 28871 21916
rect 28813 21907 28871 21913
rect 30466 21904 30472 21916
rect 30524 21904 30530 21956
rect 31018 21904 31024 21956
rect 31076 21944 31082 21956
rect 31113 21947 31171 21953
rect 31113 21944 31125 21947
rect 31076 21916 31125 21944
rect 31076 21904 31082 21916
rect 31113 21913 31125 21916
rect 31159 21913 31171 21947
rect 31113 21907 31171 21913
rect 31386 21904 31392 21956
rect 31444 21944 31450 21956
rect 31444 21916 31602 21944
rect 31444 21904 31450 21916
rect 21266 21876 21272 21888
rect 14568 21848 21272 21876
rect 12989 21839 13047 21845
rect 21266 21836 21272 21848
rect 21324 21836 21330 21888
rect 21450 21836 21456 21888
rect 21508 21836 21514 21888
rect 21910 21836 21916 21888
rect 21968 21836 21974 21888
rect 22646 21836 22652 21888
rect 22704 21836 22710 21888
rect 23106 21836 23112 21888
rect 23164 21836 23170 21888
rect 23750 21836 23756 21888
rect 23808 21876 23814 21888
rect 23845 21879 23903 21885
rect 23845 21876 23857 21879
rect 23808 21848 23857 21876
rect 23808 21836 23814 21848
rect 23845 21845 23857 21848
rect 23891 21845 23903 21879
rect 23845 21839 23903 21845
rect 25958 21836 25964 21888
rect 26016 21836 26022 21888
rect 26142 21836 26148 21888
rect 26200 21876 26206 21888
rect 27157 21879 27215 21885
rect 27157 21876 27169 21879
rect 26200 21848 27169 21876
rect 26200 21836 26206 21848
rect 27157 21845 27169 21848
rect 27203 21845 27215 21879
rect 27157 21839 27215 21845
rect 28721 21879 28779 21885
rect 28721 21845 28733 21879
rect 28767 21876 28779 21879
rect 29546 21876 29552 21888
rect 28767 21848 29552 21876
rect 28767 21845 28779 21848
rect 28721 21839 28779 21845
rect 29546 21836 29552 21848
rect 29604 21836 29610 21888
rect 29730 21836 29736 21888
rect 29788 21836 29794 21888
rect 30374 21836 30380 21888
rect 30432 21836 30438 21888
rect 31496 21876 31524 21916
rect 32122 21876 32128 21888
rect 31496 21848 32128 21876
rect 32122 21836 32128 21848
rect 32180 21836 32186 21888
rect 32398 21836 32404 21888
rect 32456 21876 32462 21888
rect 32585 21879 32643 21885
rect 32585 21876 32597 21879
rect 32456 21848 32597 21876
rect 32456 21836 32462 21848
rect 32585 21845 32597 21848
rect 32631 21845 32643 21879
rect 32585 21839 32643 21845
rect 32674 21836 32680 21888
rect 32732 21876 32738 21888
rect 33045 21879 33103 21885
rect 33045 21876 33057 21879
rect 32732 21848 33057 21876
rect 32732 21836 32738 21848
rect 33045 21845 33057 21848
rect 33091 21845 33103 21879
rect 33045 21839 33103 21845
rect 33410 21836 33416 21888
rect 33468 21836 33474 21888
rect 34330 21836 34336 21888
rect 34388 21836 34394 21888
rect 34606 21836 34612 21888
rect 34664 21876 34670 21888
rect 35176 21885 35204 21984
rect 35253 21947 35311 21953
rect 35253 21913 35265 21947
rect 35299 21944 35311 21947
rect 35802 21944 35808 21956
rect 35299 21916 35808 21944
rect 35299 21913 35311 21916
rect 35253 21907 35311 21913
rect 35802 21904 35808 21916
rect 35860 21904 35866 21956
rect 36372 21944 36400 21984
rect 39574 21972 39580 21984
rect 39632 21972 39638 22024
rect 39684 22012 39712 22052
rect 40865 22049 40877 22083
rect 40911 22049 40923 22083
rect 40865 22043 40923 22049
rect 41969 22083 42027 22089
rect 41969 22049 41981 22083
rect 42015 22049 42027 22083
rect 41969 22043 42027 22049
rect 41877 22015 41935 22021
rect 41877 22012 41889 22015
rect 39684 21984 41889 22012
rect 41877 21981 41889 21984
rect 41923 22012 41935 22015
rect 42426 22012 42432 22024
rect 41923 21984 42432 22012
rect 41923 21981 41935 21984
rect 41877 21975 41935 21981
rect 42426 21972 42432 21984
rect 42484 22012 42490 22024
rect 42536 22012 42564 22120
rect 43714 22108 43720 22120
rect 43772 22108 43778 22160
rect 44266 22108 44272 22160
rect 44324 22148 44330 22160
rect 47673 22151 47731 22157
rect 47673 22148 47685 22151
rect 44324 22120 47685 22148
rect 44324 22108 44330 22120
rect 47673 22117 47685 22120
rect 47719 22117 47731 22151
rect 47673 22111 47731 22117
rect 42886 22040 42892 22092
rect 42944 22080 42950 22092
rect 43533 22083 43591 22089
rect 43533 22080 43545 22083
rect 42944 22052 43545 22080
rect 42944 22040 42950 22052
rect 43533 22049 43545 22052
rect 43579 22049 43591 22083
rect 43533 22043 43591 22049
rect 43806 22040 43812 22092
rect 43864 22080 43870 22092
rect 44361 22083 44419 22089
rect 44361 22080 44373 22083
rect 43864 22052 44373 22080
rect 43864 22040 43870 22052
rect 44361 22049 44373 22052
rect 44407 22049 44419 22083
rect 44361 22043 44419 22049
rect 44637 22083 44695 22089
rect 44637 22049 44649 22083
rect 44683 22080 44695 22083
rect 44726 22080 44732 22092
rect 44683 22052 44732 22080
rect 44683 22049 44695 22052
rect 44637 22043 44695 22049
rect 44726 22040 44732 22052
rect 44784 22040 44790 22092
rect 46845 22083 46903 22089
rect 46845 22049 46857 22083
rect 46891 22080 46903 22083
rect 46891 22052 49280 22080
rect 46891 22049 46903 22052
rect 46845 22043 46903 22049
rect 42484 21984 42564 22012
rect 42484 21972 42490 21984
rect 42794 21972 42800 22024
rect 42852 21972 42858 22024
rect 43254 21972 43260 22024
rect 43312 21972 43318 22024
rect 47578 21972 47584 22024
rect 47636 22012 47642 22024
rect 47857 22015 47915 22021
rect 47857 22012 47869 22015
rect 47636 21984 47869 22012
rect 47636 21972 47642 21984
rect 47857 21981 47869 21984
rect 47903 21981 47915 22015
rect 47857 21975 47915 21981
rect 48498 21972 48504 22024
rect 48556 21972 48562 22024
rect 37182 21944 37188 21956
rect 36372 21916 37188 21944
rect 37182 21904 37188 21916
rect 37240 21944 37246 21956
rect 37550 21944 37556 21956
rect 37240 21916 37556 21944
rect 37240 21904 37246 21916
rect 37550 21904 37556 21916
rect 37608 21904 37614 21956
rect 38378 21904 38384 21956
rect 38436 21904 38442 21956
rect 40034 21944 40040 21956
rect 39224 21916 40040 21944
rect 35161 21879 35219 21885
rect 35161 21876 35173 21879
rect 34664 21848 35173 21876
rect 34664 21836 34670 21848
rect 35161 21845 35173 21848
rect 35207 21845 35219 21879
rect 35161 21839 35219 21845
rect 35621 21879 35679 21885
rect 35621 21845 35633 21879
rect 35667 21876 35679 21879
rect 35986 21876 35992 21888
rect 35667 21848 35992 21876
rect 35667 21845 35679 21848
rect 35621 21839 35679 21845
rect 35986 21836 35992 21848
rect 36044 21836 36050 21888
rect 36262 21836 36268 21888
rect 36320 21876 36326 21888
rect 36357 21879 36415 21885
rect 36357 21876 36369 21879
rect 36320 21848 36369 21876
rect 36320 21836 36326 21848
rect 36357 21845 36369 21848
rect 36403 21845 36415 21879
rect 36357 21839 36415 21845
rect 36449 21879 36507 21885
rect 36449 21845 36461 21879
rect 36495 21876 36507 21879
rect 36538 21876 36544 21888
rect 36495 21848 36544 21876
rect 36495 21845 36507 21848
rect 36449 21839 36507 21845
rect 36538 21836 36544 21848
rect 36596 21836 36602 21888
rect 36814 21836 36820 21888
rect 36872 21836 36878 21888
rect 37274 21836 37280 21888
rect 37332 21876 37338 21888
rect 37369 21879 37427 21885
rect 37369 21876 37381 21879
rect 37332 21848 37381 21876
rect 37332 21836 37338 21848
rect 37369 21845 37381 21848
rect 37415 21845 37427 21879
rect 37369 21839 37427 21845
rect 37458 21836 37464 21888
rect 37516 21876 37522 21888
rect 39224 21876 39252 21916
rect 40034 21904 40040 21916
rect 40092 21904 40098 21956
rect 40681 21947 40739 21953
rect 40681 21913 40693 21947
rect 40727 21944 40739 21947
rect 42702 21944 42708 21956
rect 40727 21916 41092 21944
rect 40727 21913 40739 21916
rect 40681 21907 40739 21913
rect 37516 21848 39252 21876
rect 37516 21836 37522 21848
rect 39666 21836 39672 21888
rect 39724 21876 39730 21888
rect 39853 21879 39911 21885
rect 39853 21876 39865 21879
rect 39724 21848 39865 21876
rect 39724 21836 39730 21848
rect 39853 21845 39865 21848
rect 39899 21845 39911 21879
rect 39853 21839 39911 21845
rect 39942 21836 39948 21888
rect 40000 21876 40006 21888
rect 40589 21879 40647 21885
rect 40589 21876 40601 21879
rect 40000 21848 40601 21876
rect 40000 21836 40006 21848
rect 40589 21845 40601 21848
rect 40635 21876 40647 21879
rect 40862 21876 40868 21888
rect 40635 21848 40868 21876
rect 40635 21845 40647 21848
rect 40589 21839 40647 21845
rect 40862 21836 40868 21848
rect 40920 21836 40926 21888
rect 40954 21836 40960 21888
rect 41012 21876 41018 21888
rect 41064 21876 41092 21916
rect 41248 21916 42708 21944
rect 41248 21876 41276 21916
rect 42702 21904 42708 21916
rect 42760 21904 42766 21956
rect 47397 21947 47455 21953
rect 47397 21913 47409 21947
rect 47443 21944 47455 21947
rect 48516 21944 48544 21972
rect 49252 21956 49280 22052
rect 47443 21916 48544 21944
rect 47443 21913 47455 21916
rect 47397 21907 47455 21913
rect 49050 21904 49056 21956
rect 49108 21904 49114 21956
rect 49234 21904 49240 21956
rect 49292 21904 49298 21956
rect 41012 21848 41276 21876
rect 41012 21836 41018 21848
rect 41322 21836 41328 21888
rect 41380 21876 41386 21888
rect 41417 21879 41475 21885
rect 41417 21876 41429 21879
rect 41380 21848 41429 21876
rect 41380 21836 41386 21848
rect 41417 21845 41429 21848
rect 41463 21845 41475 21879
rect 41417 21839 41475 21845
rect 41782 21836 41788 21888
rect 41840 21836 41846 21888
rect 41874 21836 41880 21888
rect 41932 21876 41938 21888
rect 42613 21879 42671 21885
rect 42613 21876 42625 21879
rect 41932 21848 42625 21876
rect 41932 21836 41938 21848
rect 42613 21845 42625 21848
rect 42659 21845 42671 21879
rect 42613 21839 42671 21845
rect 47854 21836 47860 21888
rect 47912 21876 47918 21888
rect 48409 21879 48467 21885
rect 48409 21876 48421 21879
rect 47912 21848 48421 21876
rect 47912 21836 47918 21848
rect 48409 21845 48421 21848
rect 48455 21845 48467 21879
rect 48409 21839 48467 21845
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 9582 21632 9588 21684
rect 9640 21672 9646 21684
rect 10505 21675 10563 21681
rect 10505 21672 10517 21675
rect 9640 21644 10517 21672
rect 9640 21632 9646 21644
rect 10505 21641 10517 21644
rect 10551 21641 10563 21675
rect 12434 21672 12440 21684
rect 10505 21635 10563 21641
rect 10612 21644 12440 21672
rect 3326 21564 3332 21616
rect 3384 21604 3390 21616
rect 3605 21607 3663 21613
rect 3605 21604 3617 21607
rect 3384 21576 3617 21604
rect 3384 21564 3390 21576
rect 3605 21573 3617 21576
rect 3651 21573 3663 21607
rect 3605 21567 3663 21573
rect 6730 21564 6736 21616
rect 6788 21604 6794 21616
rect 6788 21576 8984 21604
rect 6788 21564 6794 21576
rect 2961 21539 3019 21545
rect 2961 21505 2973 21539
rect 3007 21505 3019 21539
rect 2961 21499 3019 21505
rect 1762 21428 1768 21480
rect 1820 21428 1826 21480
rect 2976 21468 3004 21499
rect 4614 21496 4620 21548
rect 4672 21496 4678 21548
rect 5721 21539 5779 21545
rect 5721 21505 5733 21539
rect 5767 21536 5779 21539
rect 6546 21536 6552 21548
rect 5767 21508 6552 21536
rect 5767 21505 5779 21508
rect 5721 21499 5779 21505
rect 6546 21496 6552 21508
rect 6604 21496 6610 21548
rect 6638 21496 6644 21548
rect 6696 21496 6702 21548
rect 8481 21539 8539 21545
rect 8481 21505 8493 21539
rect 8527 21505 8539 21539
rect 8481 21499 8539 21505
rect 5626 21468 5632 21480
rect 2976 21440 5632 21468
rect 5626 21428 5632 21440
rect 5684 21428 5690 21480
rect 5810 21428 5816 21480
rect 5868 21468 5874 21480
rect 7009 21471 7067 21477
rect 7009 21468 7021 21471
rect 5868 21440 7021 21468
rect 5868 21428 5874 21440
rect 7009 21437 7021 21440
rect 7055 21437 7067 21471
rect 7009 21431 7067 21437
rect 5905 21403 5963 21409
rect 5905 21369 5917 21403
rect 5951 21400 5963 21403
rect 8496 21400 8524 21499
rect 8849 21471 8907 21477
rect 8849 21437 8861 21471
rect 8895 21437 8907 21471
rect 8956 21468 8984 21576
rect 9030 21496 9036 21548
rect 9088 21536 9094 21548
rect 9950 21536 9956 21548
rect 9088 21508 9956 21536
rect 9088 21496 9094 21508
rect 9950 21496 9956 21508
rect 10008 21496 10014 21548
rect 10612 21468 10640 21644
rect 12434 21632 12440 21644
rect 12492 21632 12498 21684
rect 12544 21644 13216 21672
rect 10962 21564 10968 21616
rect 11020 21604 11026 21616
rect 12544 21604 12572 21644
rect 11020 21576 12572 21604
rect 11020 21564 11026 21576
rect 12618 21564 12624 21616
rect 12676 21604 12682 21616
rect 13081 21607 13139 21613
rect 13081 21604 13093 21607
rect 12676 21576 13093 21604
rect 12676 21564 12682 21576
rect 13081 21573 13093 21576
rect 13127 21573 13139 21607
rect 13188 21604 13216 21644
rect 13814 21632 13820 21684
rect 13872 21672 13878 21684
rect 13909 21675 13967 21681
rect 13909 21672 13921 21675
rect 13872 21644 13921 21672
rect 13872 21632 13878 21644
rect 13909 21641 13921 21644
rect 13955 21641 13967 21675
rect 17405 21675 17463 21681
rect 17405 21672 17417 21675
rect 13909 21635 13967 21641
rect 14200 21644 17417 21672
rect 14200 21604 14228 21644
rect 17405 21641 17417 21644
rect 17451 21641 17463 21675
rect 17405 21635 17463 21641
rect 17865 21675 17923 21681
rect 17865 21641 17877 21675
rect 17911 21672 17923 21675
rect 20990 21672 20996 21684
rect 17911 21644 20996 21672
rect 17911 21641 17923 21644
rect 17865 21635 17923 21641
rect 20990 21632 20996 21644
rect 21048 21632 21054 21684
rect 21910 21632 21916 21684
rect 21968 21672 21974 21684
rect 22554 21672 22560 21684
rect 21968 21644 22560 21672
rect 21968 21632 21974 21644
rect 22554 21632 22560 21644
rect 22612 21632 22618 21684
rect 22922 21632 22928 21684
rect 22980 21672 22986 21684
rect 24765 21675 24823 21681
rect 24765 21672 24777 21675
rect 22980 21644 24777 21672
rect 22980 21632 22986 21644
rect 24765 21641 24777 21644
rect 24811 21641 24823 21675
rect 27062 21672 27068 21684
rect 24765 21635 24823 21641
rect 24872 21644 27068 21672
rect 13188 21576 14228 21604
rect 13081 21567 13139 21573
rect 14274 21564 14280 21616
rect 14332 21604 14338 21616
rect 14829 21607 14887 21613
rect 14829 21604 14841 21607
rect 14332 21576 14841 21604
rect 14332 21564 14338 21576
rect 14829 21573 14841 21576
rect 14875 21573 14887 21607
rect 16114 21604 16120 21616
rect 16054 21590 16120 21604
rect 14829 21567 14887 21573
rect 16040 21576 16120 21590
rect 10689 21539 10747 21545
rect 10689 21505 10701 21539
rect 10735 21505 10747 21539
rect 10689 21499 10747 21505
rect 11149 21539 11207 21545
rect 11149 21505 11161 21539
rect 11195 21536 11207 21539
rect 12066 21536 12072 21548
rect 11195 21508 12072 21536
rect 11195 21505 11207 21508
rect 11149 21499 11207 21505
rect 8956 21440 10640 21468
rect 8849 21431 8907 21437
rect 5951 21372 8524 21400
rect 5951 21369 5963 21372
rect 5905 21363 5963 21369
rect 3786 21292 3792 21344
rect 3844 21332 3850 21344
rect 8864 21332 8892 21431
rect 10704 21400 10732 21499
rect 12066 21496 12072 21508
rect 12124 21496 12130 21548
rect 12158 21496 12164 21548
rect 12216 21536 12222 21548
rect 12345 21539 12403 21545
rect 12345 21536 12357 21539
rect 12216 21508 12357 21536
rect 12216 21496 12222 21508
rect 12345 21505 12357 21508
rect 12391 21505 12403 21539
rect 12345 21499 12403 21505
rect 13265 21539 13323 21545
rect 13265 21505 13277 21539
rect 13311 21536 13323 21539
rect 13998 21536 14004 21548
rect 13311 21508 14004 21536
rect 13311 21505 13323 21508
rect 13265 21499 13323 21505
rect 13998 21496 14004 21508
rect 14056 21496 14062 21548
rect 14093 21539 14151 21545
rect 14093 21505 14105 21539
rect 14139 21536 14151 21539
rect 14366 21536 14372 21548
rect 14139 21508 14372 21536
rect 14139 21505 14151 21508
rect 14093 21499 14151 21505
rect 14366 21496 14372 21508
rect 14424 21496 14430 21548
rect 11422 21428 11428 21480
rect 11480 21468 11486 21480
rect 11698 21468 11704 21480
rect 11480 21440 11704 21468
rect 11480 21428 11486 21440
rect 11698 21428 11704 21440
rect 11756 21428 11762 21480
rect 11885 21471 11943 21477
rect 11885 21437 11897 21471
rect 11931 21468 11943 21471
rect 12618 21468 12624 21480
rect 11931 21440 12624 21468
rect 11931 21437 11943 21440
rect 11885 21431 11943 21437
rect 12618 21428 12624 21440
rect 12676 21428 12682 21480
rect 12802 21428 12808 21480
rect 12860 21468 12866 21480
rect 13906 21468 13912 21480
rect 12860 21440 13912 21468
rect 12860 21428 12866 21440
rect 13906 21428 13912 21440
rect 13964 21468 13970 21480
rect 14553 21471 14611 21477
rect 14553 21468 14565 21471
rect 13964 21440 14565 21468
rect 13964 21428 13970 21440
rect 14553 21437 14565 21440
rect 14599 21468 14611 21471
rect 14599 21440 14688 21468
rect 14599 21437 14611 21440
rect 14553 21431 14611 21437
rect 13722 21400 13728 21412
rect 10704 21372 13728 21400
rect 13722 21360 13728 21372
rect 13780 21360 13786 21412
rect 3844 21304 8892 21332
rect 3844 21292 3850 21304
rect 8938 21292 8944 21344
rect 8996 21332 9002 21344
rect 10870 21332 10876 21344
rect 8996 21304 10876 21332
rect 8996 21292 9002 21304
rect 10870 21292 10876 21304
rect 10928 21292 10934 21344
rect 11333 21335 11391 21341
rect 11333 21301 11345 21335
rect 11379 21332 11391 21335
rect 11790 21332 11796 21344
rect 11379 21304 11796 21332
rect 11379 21301 11391 21304
rect 11333 21295 11391 21301
rect 11790 21292 11796 21304
rect 11848 21292 11854 21344
rect 12250 21292 12256 21344
rect 12308 21292 12314 21344
rect 14660 21332 14688 21440
rect 15194 21428 15200 21480
rect 15252 21468 15258 21480
rect 16040 21468 16068 21576
rect 16114 21564 16120 21576
rect 16172 21604 16178 21616
rect 16942 21604 16948 21616
rect 16172 21576 16948 21604
rect 16172 21564 16178 21576
rect 16942 21564 16948 21576
rect 17000 21564 17006 21616
rect 18782 21604 18788 21616
rect 18432 21576 18788 21604
rect 17773 21539 17831 21545
rect 17773 21505 17785 21539
rect 17819 21536 17831 21539
rect 18322 21536 18328 21548
rect 17819 21508 18328 21536
rect 17819 21505 17831 21508
rect 17773 21499 17831 21505
rect 18322 21496 18328 21508
rect 18380 21496 18386 21548
rect 15252 21440 16068 21468
rect 16301 21471 16359 21477
rect 15252 21428 15258 21440
rect 16301 21437 16313 21471
rect 16347 21468 16359 21471
rect 16666 21468 16672 21480
rect 16347 21440 16672 21468
rect 16347 21437 16359 21440
rect 16301 21431 16359 21437
rect 16666 21428 16672 21440
rect 16724 21468 16730 21480
rect 17494 21468 17500 21480
rect 16724 21440 17500 21468
rect 16724 21428 16730 21440
rect 17494 21428 17500 21440
rect 17552 21428 17558 21480
rect 18049 21471 18107 21477
rect 18049 21437 18061 21471
rect 18095 21468 18107 21471
rect 18432 21468 18460 21576
rect 18782 21564 18788 21576
rect 18840 21564 18846 21616
rect 19150 21564 19156 21616
rect 19208 21604 19214 21616
rect 19208 21576 19366 21604
rect 19208 21564 19214 21576
rect 20622 21564 20628 21616
rect 20680 21604 20686 21616
rect 21177 21607 21235 21613
rect 21177 21604 21189 21607
rect 20680 21576 21189 21604
rect 20680 21564 20686 21576
rect 21177 21573 21189 21576
rect 21223 21573 21235 21607
rect 22741 21607 22799 21613
rect 22741 21604 22753 21607
rect 21177 21567 21235 21573
rect 21284 21576 22753 21604
rect 18095 21440 18460 21468
rect 18601 21471 18659 21477
rect 18095 21437 18107 21440
rect 18049 21431 18107 21437
rect 18601 21437 18613 21471
rect 18647 21437 18659 21471
rect 18601 21431 18659 21437
rect 16758 21360 16764 21412
rect 16816 21400 16822 21412
rect 17129 21403 17187 21409
rect 17129 21400 17141 21403
rect 16816 21372 17141 21400
rect 16816 21360 16822 21372
rect 17129 21369 17141 21372
rect 17175 21400 17187 21403
rect 18616 21400 18644 21431
rect 18874 21428 18880 21480
rect 18932 21428 18938 21480
rect 19242 21428 19248 21480
rect 19300 21468 19306 21480
rect 21284 21468 21312 21576
rect 22741 21573 22753 21576
rect 22787 21573 22799 21607
rect 24872 21604 24900 21644
rect 27062 21632 27068 21644
rect 27120 21632 27126 21684
rect 27157 21675 27215 21681
rect 27157 21641 27169 21675
rect 27203 21641 27215 21675
rect 27157 21635 27215 21641
rect 22741 21567 22799 21573
rect 24228 21576 24900 21604
rect 21361 21539 21419 21545
rect 21361 21505 21373 21539
rect 21407 21505 21419 21539
rect 22278 21536 22284 21548
rect 21361 21499 21419 21505
rect 22066 21508 22284 21536
rect 19300 21440 21312 21468
rect 19300 21428 19306 21440
rect 17175 21372 18644 21400
rect 17175 21369 17187 21372
rect 17129 21363 17187 21369
rect 16776 21332 16804 21360
rect 14660 21304 16804 21332
rect 16942 21292 16948 21344
rect 17000 21332 17006 21344
rect 17862 21332 17868 21344
rect 17000 21304 17868 21332
rect 17000 21292 17006 21304
rect 17862 21292 17868 21304
rect 17920 21292 17926 21344
rect 18616 21332 18644 21372
rect 20349 21403 20407 21409
rect 20349 21369 20361 21403
rect 20395 21400 20407 21403
rect 21082 21400 21088 21412
rect 20395 21372 21088 21400
rect 20395 21369 20407 21372
rect 20349 21363 20407 21369
rect 21082 21360 21088 21372
rect 21140 21360 21146 21412
rect 21376 21400 21404 21499
rect 21542 21428 21548 21480
rect 21600 21468 21606 21480
rect 22066 21468 22094 21508
rect 22278 21496 22284 21508
rect 22336 21496 22342 21548
rect 23842 21496 23848 21548
rect 23900 21496 23906 21548
rect 21600 21440 22094 21468
rect 21600 21428 21606 21440
rect 22186 21428 22192 21480
rect 22244 21468 22250 21480
rect 24228 21477 24256 21576
rect 25038 21564 25044 21616
rect 25096 21604 25102 21616
rect 27172 21604 27200 21635
rect 27430 21632 27436 21684
rect 27488 21672 27494 21684
rect 27617 21675 27675 21681
rect 27617 21672 27629 21675
rect 27488 21644 27629 21672
rect 27488 21632 27494 21644
rect 27617 21641 27629 21644
rect 27663 21641 27675 21675
rect 27617 21635 27675 21641
rect 30009 21675 30067 21681
rect 30009 21641 30021 21675
rect 30055 21672 30067 21675
rect 31754 21672 31760 21684
rect 30055 21644 31760 21672
rect 30055 21641 30067 21644
rect 30009 21635 30067 21641
rect 31754 21632 31760 21644
rect 31812 21632 31818 21684
rect 32769 21675 32827 21681
rect 32769 21641 32781 21675
rect 32815 21672 32827 21675
rect 33410 21672 33416 21684
rect 32815 21644 33416 21672
rect 32815 21641 32827 21644
rect 32769 21635 32827 21641
rect 33410 21632 33416 21644
rect 33468 21632 33474 21684
rect 33965 21675 34023 21681
rect 33965 21641 33977 21675
rect 34011 21672 34023 21675
rect 35894 21672 35900 21684
rect 34011 21644 35900 21672
rect 34011 21641 34023 21644
rect 33965 21635 34023 21641
rect 35894 21632 35900 21644
rect 35952 21632 35958 21684
rect 36081 21675 36139 21681
rect 36081 21641 36093 21675
rect 36127 21672 36139 21675
rect 37458 21672 37464 21684
rect 36127 21644 37464 21672
rect 36127 21641 36139 21644
rect 36081 21635 36139 21641
rect 37458 21632 37464 21644
rect 37516 21632 37522 21684
rect 37550 21632 37556 21684
rect 37608 21672 37614 21684
rect 39114 21672 39120 21684
rect 37608 21644 39120 21672
rect 37608 21632 37614 21644
rect 39114 21632 39120 21644
rect 39172 21632 39178 21684
rect 39206 21632 39212 21684
rect 39264 21672 39270 21684
rect 39942 21672 39948 21684
rect 39264 21644 39948 21672
rect 39264 21632 39270 21644
rect 39942 21632 39948 21644
rect 40000 21632 40006 21684
rect 40129 21675 40187 21681
rect 40129 21641 40141 21675
rect 40175 21672 40187 21675
rect 40313 21675 40371 21681
rect 40313 21672 40325 21675
rect 40175 21644 40325 21672
rect 40175 21641 40187 21644
rect 40129 21635 40187 21641
rect 40313 21641 40325 21644
rect 40359 21672 40371 21675
rect 40497 21675 40555 21681
rect 40497 21672 40509 21675
rect 40359 21644 40509 21672
rect 40359 21641 40371 21644
rect 40313 21635 40371 21641
rect 40497 21641 40509 21644
rect 40543 21672 40555 21675
rect 40681 21675 40739 21681
rect 40681 21672 40693 21675
rect 40543 21644 40693 21672
rect 40543 21641 40555 21644
rect 40497 21635 40555 21641
rect 40681 21641 40693 21644
rect 40727 21672 40739 21675
rect 41046 21672 41052 21684
rect 40727 21644 41052 21672
rect 40727 21641 40739 21644
rect 40681 21635 40739 21641
rect 25096 21576 27200 21604
rect 27525 21607 27583 21613
rect 25096 21564 25102 21576
rect 27525 21573 27537 21607
rect 27571 21604 27583 21607
rect 29362 21604 29368 21616
rect 27571 21576 29368 21604
rect 27571 21573 27583 21576
rect 27525 21567 27583 21573
rect 29362 21564 29368 21576
rect 29420 21564 29426 21616
rect 31113 21607 31171 21613
rect 31113 21573 31125 21607
rect 31159 21604 31171 21607
rect 33597 21607 33655 21613
rect 33597 21604 33609 21607
rect 31159 21576 33609 21604
rect 31159 21573 31171 21576
rect 31113 21567 31171 21573
rect 33597 21573 33609 21576
rect 33643 21604 33655 21607
rect 33686 21604 33692 21616
rect 33643 21576 33692 21604
rect 33643 21573 33655 21576
rect 33597 21567 33655 21573
rect 33686 21564 33692 21576
rect 33744 21564 33750 21616
rect 34793 21607 34851 21613
rect 34793 21573 34805 21607
rect 34839 21604 34851 21607
rect 34882 21604 34888 21616
rect 34839 21576 34888 21604
rect 34839 21573 34851 21576
rect 34793 21567 34851 21573
rect 34882 21564 34888 21576
rect 34940 21564 34946 21616
rect 37274 21564 37280 21616
rect 37332 21604 37338 21616
rect 38286 21604 38292 21616
rect 37332 21576 38292 21604
rect 37332 21564 37338 21576
rect 38286 21564 38292 21576
rect 38344 21564 38350 21616
rect 39666 21604 39672 21616
rect 39514 21576 39672 21604
rect 39666 21564 39672 21576
rect 39724 21604 39730 21616
rect 40144 21604 40172 21635
rect 41046 21632 41052 21644
rect 41104 21632 41110 21684
rect 42058 21632 42064 21684
rect 42116 21672 42122 21684
rect 43349 21675 43407 21681
rect 43349 21672 43361 21675
rect 42116 21644 43361 21672
rect 42116 21632 42122 21644
rect 43349 21641 43361 21644
rect 43395 21641 43407 21675
rect 43349 21635 43407 21641
rect 43530 21632 43536 21684
rect 43588 21672 43594 21684
rect 43625 21675 43683 21681
rect 43625 21672 43637 21675
rect 43588 21644 43637 21672
rect 43588 21632 43594 21644
rect 43625 21641 43637 21644
rect 43671 21641 43683 21675
rect 43625 21635 43683 21641
rect 43901 21675 43959 21681
rect 43901 21641 43913 21675
rect 43947 21672 43959 21675
rect 43990 21672 43996 21684
rect 43947 21644 43996 21672
rect 43947 21641 43959 21644
rect 43901 21635 43959 21641
rect 43990 21632 43996 21644
rect 44048 21632 44054 21684
rect 46198 21632 46204 21684
rect 46256 21672 46262 21684
rect 47854 21672 47860 21684
rect 46256 21644 47860 21672
rect 46256 21632 46262 21644
rect 47854 21632 47860 21644
rect 47912 21632 47918 21684
rect 39724 21576 40172 21604
rect 39724 21564 39730 21576
rect 40862 21564 40868 21616
rect 40920 21604 40926 21616
rect 42518 21604 42524 21616
rect 40920 21576 42524 21604
rect 40920 21564 40926 21576
rect 42518 21564 42524 21576
rect 42576 21564 42582 21616
rect 42702 21564 42708 21616
rect 42760 21564 42766 21616
rect 42794 21564 42800 21616
rect 42852 21604 42858 21616
rect 42981 21607 43039 21613
rect 42981 21604 42993 21607
rect 42852 21576 42993 21604
rect 42852 21564 42858 21576
rect 42981 21573 42993 21576
rect 43027 21573 43039 21607
rect 42981 21567 43039 21573
rect 25133 21539 25191 21545
rect 25133 21505 25145 21539
rect 25179 21536 25191 21539
rect 25866 21536 25872 21548
rect 25179 21508 25872 21536
rect 25179 21505 25191 21508
rect 25133 21499 25191 21505
rect 25866 21496 25872 21508
rect 25924 21496 25930 21548
rect 26050 21496 26056 21548
rect 26108 21496 26114 21548
rect 26605 21539 26663 21545
rect 26605 21505 26617 21539
rect 26651 21536 26663 21539
rect 26651 21508 27844 21536
rect 26651 21505 26663 21508
rect 26605 21499 26663 21505
rect 22465 21471 22523 21477
rect 22465 21468 22477 21471
rect 22244 21440 22477 21468
rect 22244 21428 22250 21440
rect 22465 21437 22477 21440
rect 22511 21437 22523 21471
rect 24213 21471 24271 21477
rect 22465 21431 22523 21437
rect 22572 21440 23796 21468
rect 22572 21400 22600 21440
rect 21376 21372 22600 21400
rect 23768 21400 23796 21440
rect 24213 21437 24225 21471
rect 24259 21437 24271 21471
rect 24213 21431 24271 21437
rect 24486 21428 24492 21480
rect 24544 21468 24550 21480
rect 25225 21471 25283 21477
rect 25225 21468 25237 21471
rect 24544 21440 25237 21468
rect 24544 21428 24550 21440
rect 25148 21412 25176 21440
rect 25225 21437 25237 21440
rect 25271 21437 25283 21471
rect 25225 21431 25283 21437
rect 25406 21428 25412 21480
rect 25464 21468 25470 21480
rect 27709 21471 27767 21477
rect 27709 21468 27721 21471
rect 25464 21440 27721 21468
rect 25464 21428 25470 21440
rect 27709 21437 27721 21440
rect 27755 21437 27767 21471
rect 27709 21431 27767 21437
rect 23768 21372 24808 21400
rect 19334 21332 19340 21344
rect 18616 21304 19340 21332
rect 19334 21292 19340 21304
rect 19392 21292 19398 21344
rect 19610 21292 19616 21344
rect 19668 21332 19674 21344
rect 20717 21335 20775 21341
rect 20717 21332 20729 21335
rect 19668 21304 20729 21332
rect 19668 21292 19674 21304
rect 20717 21301 20729 21304
rect 20763 21332 20775 21335
rect 20901 21335 20959 21341
rect 20901 21332 20913 21335
rect 20763 21304 20913 21332
rect 20763 21301 20775 21304
rect 20717 21295 20775 21301
rect 20901 21301 20913 21304
rect 20947 21332 20959 21335
rect 21634 21332 21640 21344
rect 20947 21304 21640 21332
rect 20947 21301 20959 21304
rect 20901 21295 20959 21301
rect 21634 21292 21640 21304
rect 21692 21332 21698 21344
rect 22005 21335 22063 21341
rect 22005 21332 22017 21335
rect 21692 21304 22017 21332
rect 21692 21292 21698 21304
rect 22005 21301 22017 21304
rect 22051 21332 22063 21335
rect 22189 21335 22247 21341
rect 22189 21332 22201 21335
rect 22051 21304 22201 21332
rect 22051 21301 22063 21304
rect 22005 21295 22063 21301
rect 22189 21301 22201 21304
rect 22235 21332 22247 21335
rect 22370 21332 22376 21344
rect 22235 21304 22376 21332
rect 22235 21301 22247 21304
rect 22189 21295 22247 21301
rect 22370 21292 22376 21304
rect 22428 21292 22434 21344
rect 22554 21292 22560 21344
rect 22612 21332 22618 21344
rect 24670 21332 24676 21344
rect 22612 21304 24676 21332
rect 22612 21292 22618 21304
rect 24670 21292 24676 21304
rect 24728 21292 24734 21344
rect 24780 21332 24808 21372
rect 25130 21360 25136 21412
rect 25188 21360 25194 21412
rect 26421 21403 26479 21409
rect 26421 21400 26433 21403
rect 25516 21372 26433 21400
rect 25516 21332 25544 21372
rect 26421 21369 26433 21372
rect 26467 21369 26479 21403
rect 27816 21400 27844 21508
rect 27890 21496 27896 21548
rect 27948 21536 27954 21548
rect 28721 21539 28779 21545
rect 28721 21536 28733 21539
rect 27948 21508 28733 21536
rect 27948 21496 27954 21508
rect 28721 21505 28733 21508
rect 28767 21505 28779 21539
rect 28721 21499 28779 21505
rect 29917 21539 29975 21545
rect 29917 21505 29929 21539
rect 29963 21536 29975 21539
rect 30742 21536 30748 21548
rect 29963 21508 30748 21536
rect 29963 21505 29975 21508
rect 29917 21499 29975 21505
rect 30742 21496 30748 21508
rect 30800 21496 30806 21548
rect 31202 21496 31208 21548
rect 31260 21496 31266 21548
rect 33502 21496 33508 21548
rect 33560 21496 33566 21548
rect 34701 21539 34759 21545
rect 34701 21505 34713 21539
rect 34747 21505 34759 21539
rect 37734 21536 37740 21548
rect 34701 21499 34759 21505
rect 34808 21508 37740 21536
rect 28810 21428 28816 21480
rect 28868 21428 28874 21480
rect 28902 21428 28908 21480
rect 28960 21428 28966 21480
rect 29730 21428 29736 21480
rect 29788 21468 29794 21480
rect 30101 21471 30159 21477
rect 30101 21468 30113 21471
rect 29788 21440 30113 21468
rect 29788 21428 29794 21440
rect 30101 21437 30113 21440
rect 30147 21437 30159 21471
rect 30101 21431 30159 21437
rect 31389 21471 31447 21477
rect 31389 21437 31401 21471
rect 31435 21468 31447 21471
rect 31570 21468 31576 21480
rect 31435 21440 31576 21468
rect 31435 21437 31447 21440
rect 31389 21431 31447 21437
rect 31570 21428 31576 21440
rect 31628 21468 31634 21480
rect 31757 21471 31815 21477
rect 31757 21468 31769 21471
rect 31628 21440 31769 21468
rect 31628 21428 31634 21440
rect 31757 21437 31769 21440
rect 31803 21437 31815 21471
rect 31757 21431 31815 21437
rect 33410 21428 33416 21480
rect 33468 21428 33474 21480
rect 34238 21428 34244 21480
rect 34296 21468 34302 21480
rect 34517 21471 34575 21477
rect 34517 21468 34529 21471
rect 34296 21440 34529 21468
rect 34296 21428 34302 21440
rect 34517 21437 34529 21440
rect 34563 21437 34575 21471
rect 34517 21431 34575 21437
rect 34716 21412 34744 21499
rect 30466 21400 30472 21412
rect 27816 21372 30472 21400
rect 26421 21363 26479 21369
rect 30466 21360 30472 21372
rect 30524 21360 30530 21412
rect 30558 21360 30564 21412
rect 30616 21400 30622 21412
rect 31478 21400 31484 21412
rect 30616 21372 31484 21400
rect 30616 21360 30622 21372
rect 31478 21360 31484 21372
rect 31536 21360 31542 21412
rect 34698 21360 34704 21412
rect 34756 21360 34762 21412
rect 24780 21304 25544 21332
rect 25866 21292 25872 21344
rect 25924 21292 25930 21344
rect 26234 21292 26240 21344
rect 26292 21332 26298 21344
rect 28353 21335 28411 21341
rect 28353 21332 28365 21335
rect 26292 21304 28365 21332
rect 26292 21292 26298 21304
rect 28353 21301 28365 21304
rect 28399 21301 28411 21335
rect 28353 21295 28411 21301
rect 29546 21292 29552 21344
rect 29604 21292 29610 21344
rect 29638 21292 29644 21344
rect 29696 21332 29702 21344
rect 29914 21332 29920 21344
rect 29696 21304 29920 21332
rect 29696 21292 29702 21304
rect 29914 21292 29920 21304
rect 29972 21292 29978 21344
rect 30742 21292 30748 21344
rect 30800 21292 30806 21344
rect 31938 21292 31944 21344
rect 31996 21332 32002 21344
rect 34808 21332 34836 21508
rect 37734 21496 37740 21508
rect 37792 21496 37798 21548
rect 40678 21496 40684 21548
rect 40736 21536 40742 21548
rect 43254 21536 43260 21548
rect 40736 21508 43260 21536
rect 40736 21496 40742 21508
rect 43254 21496 43260 21508
rect 43312 21496 43318 21548
rect 46842 21496 46848 21548
rect 46900 21536 46906 21548
rect 47949 21539 48007 21545
rect 47949 21536 47961 21539
rect 46900 21508 47961 21536
rect 46900 21496 46906 21508
rect 47949 21505 47961 21508
rect 47995 21505 48007 21539
rect 47949 21499 48007 21505
rect 48590 21496 48596 21548
rect 48648 21496 48654 21548
rect 49326 21496 49332 21548
rect 49384 21496 49390 21548
rect 34882 21428 34888 21480
rect 34940 21468 34946 21480
rect 34940 21440 36124 21468
rect 34940 21428 34946 21440
rect 36096 21400 36124 21440
rect 36170 21428 36176 21480
rect 36228 21428 36234 21480
rect 36265 21471 36323 21477
rect 36265 21437 36277 21471
rect 36311 21437 36323 21471
rect 36265 21431 36323 21437
rect 36817 21471 36875 21477
rect 36817 21437 36829 21471
rect 36863 21468 36875 21471
rect 36906 21468 36912 21480
rect 36863 21440 36912 21468
rect 36863 21437 36875 21440
rect 36817 21431 36875 21437
rect 36280 21400 36308 21431
rect 36906 21428 36912 21440
rect 36964 21428 36970 21480
rect 37182 21428 37188 21480
rect 37240 21468 37246 21480
rect 37277 21471 37335 21477
rect 37277 21468 37289 21471
rect 37240 21440 37289 21468
rect 37240 21428 37246 21440
rect 37277 21437 37289 21440
rect 37323 21437 37335 21471
rect 37277 21431 37335 21437
rect 37550 21428 37556 21480
rect 37608 21468 37614 21480
rect 37645 21471 37703 21477
rect 37645 21468 37657 21471
rect 37608 21440 37657 21468
rect 37608 21428 37614 21440
rect 37645 21437 37657 21440
rect 37691 21468 37703 21471
rect 38002 21471 38060 21477
rect 38002 21468 38014 21471
rect 37691 21440 38014 21468
rect 37691 21437 37703 21440
rect 37645 21431 37703 21437
rect 38002 21437 38014 21440
rect 38048 21437 38060 21471
rect 40310 21468 40316 21480
rect 38002 21431 38060 21437
rect 38120 21440 40316 21468
rect 38120 21400 38148 21440
rect 40310 21428 40316 21440
rect 40368 21428 40374 21480
rect 41233 21471 41291 21477
rect 41233 21437 41245 21471
rect 41279 21437 41291 21471
rect 41233 21431 41291 21437
rect 36096 21372 36308 21400
rect 38028 21372 38148 21400
rect 31996 21304 34836 21332
rect 31996 21292 32002 21304
rect 35158 21292 35164 21344
rect 35216 21292 35222 21344
rect 35710 21292 35716 21344
rect 35768 21292 35774 21344
rect 35802 21292 35808 21344
rect 35860 21332 35866 21344
rect 36909 21335 36967 21341
rect 36909 21332 36921 21335
rect 35860 21304 36921 21332
rect 35860 21292 35866 21304
rect 36909 21301 36921 21304
rect 36955 21301 36967 21335
rect 36909 21295 36967 21301
rect 37550 21292 37556 21344
rect 37608 21292 37614 21344
rect 37734 21292 37740 21344
rect 37792 21332 37798 21344
rect 38028 21332 38056 21372
rect 37792 21304 38056 21332
rect 37792 21292 37798 21304
rect 38102 21292 38108 21344
rect 38160 21332 38166 21344
rect 38838 21332 38844 21344
rect 38160 21304 38844 21332
rect 38160 21292 38166 21304
rect 38838 21292 38844 21304
rect 38896 21292 38902 21344
rect 39022 21292 39028 21344
rect 39080 21332 39086 21344
rect 39761 21335 39819 21341
rect 39761 21332 39773 21335
rect 39080 21304 39773 21332
rect 39080 21292 39086 21304
rect 39761 21301 39773 21304
rect 39807 21301 39819 21335
rect 39761 21295 39819 21301
rect 40862 21292 40868 21344
rect 40920 21332 40926 21344
rect 41248 21332 41276 21431
rect 41506 21428 41512 21480
rect 41564 21428 41570 21480
rect 41598 21428 41604 21480
rect 41656 21468 41662 21480
rect 41656 21440 48452 21468
rect 41656 21428 41662 21440
rect 41782 21360 41788 21412
rect 41840 21400 41846 21412
rect 48424 21409 48452 21440
rect 47765 21403 47823 21409
rect 47765 21400 47777 21403
rect 41840 21372 47777 21400
rect 41840 21360 41846 21372
rect 47765 21369 47777 21372
rect 47811 21369 47823 21403
rect 47765 21363 47823 21369
rect 48409 21403 48467 21409
rect 48409 21369 48421 21403
rect 48455 21369 48467 21403
rect 48409 21363 48467 21369
rect 40920 21304 41276 21332
rect 40920 21292 40926 21304
rect 41322 21292 41328 21344
rect 41380 21332 41386 21344
rect 42797 21335 42855 21341
rect 42797 21332 42809 21335
rect 41380 21304 42809 21332
rect 41380 21292 41386 21304
rect 42797 21301 42809 21304
rect 42843 21332 42855 21335
rect 43530 21332 43536 21344
rect 42843 21304 43536 21332
rect 42843 21301 42855 21304
rect 42797 21295 42855 21301
rect 43530 21292 43536 21304
rect 43588 21292 43594 21344
rect 49142 21292 49148 21344
rect 49200 21292 49206 21344
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 9122 21128 9128 21140
rect 2976 21100 9128 21128
rect 2501 20995 2559 21001
rect 2501 20961 2513 20995
rect 2547 20992 2559 20995
rect 2866 20992 2872 21004
rect 2547 20964 2872 20992
rect 2547 20961 2559 20964
rect 2501 20955 2559 20961
rect 2866 20952 2872 20964
rect 2924 20952 2930 21004
rect 2976 20933 3004 21100
rect 9122 21088 9128 21100
rect 9180 21088 9186 21140
rect 9214 21088 9220 21140
rect 9272 21088 9278 21140
rect 12250 21128 12256 21140
rect 9324 21100 12256 21128
rect 9324 21060 9352 21100
rect 12250 21088 12256 21100
rect 12308 21088 12314 21140
rect 12437 21131 12495 21137
rect 12437 21097 12449 21131
rect 12483 21128 12495 21131
rect 12802 21128 12808 21140
rect 12483 21100 12808 21128
rect 12483 21097 12495 21100
rect 12437 21091 12495 21097
rect 12802 21088 12808 21100
rect 12860 21088 12866 21140
rect 14274 21088 14280 21140
rect 14332 21088 14338 21140
rect 14366 21088 14372 21140
rect 14424 21128 14430 21140
rect 15286 21128 15292 21140
rect 14424 21100 15292 21128
rect 14424 21088 14430 21100
rect 15286 21088 15292 21100
rect 15344 21088 15350 21140
rect 16298 21088 16304 21140
rect 16356 21128 16362 21140
rect 17129 21131 17187 21137
rect 17129 21128 17141 21131
rect 16356 21100 17141 21128
rect 16356 21088 16362 21100
rect 17129 21097 17141 21100
rect 17175 21128 17187 21131
rect 19702 21128 19708 21140
rect 17175 21100 19708 21128
rect 17175 21097 17187 21100
rect 17129 21091 17187 21097
rect 19702 21088 19708 21100
rect 19760 21088 19766 21140
rect 22554 21088 22560 21140
rect 22612 21128 22618 21140
rect 24029 21131 24087 21137
rect 22612 21100 23888 21128
rect 22612 21088 22618 21100
rect 23860 21072 23888 21100
rect 24029 21097 24041 21131
rect 24075 21128 24087 21131
rect 24118 21128 24124 21140
rect 24075 21100 24124 21128
rect 24075 21097 24087 21100
rect 24029 21091 24087 21097
rect 24118 21088 24124 21100
rect 24176 21088 24182 21140
rect 24213 21131 24271 21137
rect 24213 21097 24225 21131
rect 24259 21128 24271 21131
rect 24259 21100 25268 21128
rect 24259 21097 24271 21100
rect 24213 21091 24271 21097
rect 11793 21063 11851 21069
rect 11793 21060 11805 21063
rect 5368 21032 9352 21060
rect 9646 21032 11805 21060
rect 4154 20952 4160 21004
rect 4212 20952 4218 21004
rect 5368 20933 5396 21032
rect 5994 20952 6000 21004
rect 6052 20952 6058 21004
rect 7742 20952 7748 21004
rect 7800 20992 7806 21004
rect 7800 20964 9536 20992
rect 7800 20952 7806 20964
rect 2961 20927 3019 20933
rect 2961 20893 2973 20927
rect 3007 20893 3019 20927
rect 2961 20887 3019 20893
rect 5353 20927 5411 20933
rect 5353 20893 5365 20927
rect 5399 20893 5411 20927
rect 5353 20887 5411 20893
rect 7193 20927 7251 20933
rect 7193 20893 7205 20927
rect 7239 20924 7251 20927
rect 8021 20927 8079 20933
rect 7239 20896 7880 20924
rect 7239 20893 7251 20896
rect 7193 20887 7251 20893
rect 7282 20748 7288 20800
rect 7340 20788 7346 20800
rect 7558 20788 7564 20800
rect 7340 20760 7564 20788
rect 7340 20748 7346 20760
rect 7558 20748 7564 20760
rect 7616 20748 7622 20800
rect 7852 20797 7880 20896
rect 8021 20893 8033 20927
rect 8067 20893 8079 20927
rect 8021 20887 8079 20893
rect 8036 20856 8064 20887
rect 8386 20884 8392 20936
rect 8444 20884 8450 20936
rect 9401 20927 9459 20933
rect 9401 20893 9413 20927
rect 9447 20893 9459 20927
rect 9508 20924 9536 20964
rect 9646 20924 9674 21032
rect 11793 21029 11805 21032
rect 11839 21029 11851 21063
rect 11793 21023 11851 21029
rect 19242 21020 19248 21072
rect 19300 21060 19306 21072
rect 19610 21060 19616 21072
rect 19300 21032 19616 21060
rect 19300 21020 19306 21032
rect 19610 21020 19616 21032
rect 19668 21020 19674 21072
rect 19981 21063 20039 21069
rect 19981 21029 19993 21063
rect 20027 21029 20039 21063
rect 21177 21063 21235 21069
rect 21177 21060 21189 21063
rect 19981 21023 20039 21029
rect 20548 21032 21189 21060
rect 10045 20995 10103 21001
rect 10045 20961 10057 20995
rect 10091 20992 10103 20995
rect 10226 20992 10232 21004
rect 10091 20964 10232 20992
rect 10091 20961 10103 20964
rect 10045 20955 10103 20961
rect 10226 20952 10232 20964
rect 10284 20952 10290 21004
rect 12710 20952 12716 21004
rect 12768 20952 12774 21004
rect 19996 20992 20024 21023
rect 20548 21001 20576 21032
rect 21177 21029 21189 21032
rect 21223 21029 21235 21063
rect 21177 21023 21235 21029
rect 23290 21020 23296 21072
rect 23348 21060 23354 21072
rect 23385 21063 23443 21069
rect 23385 21060 23397 21063
rect 23348 21032 23397 21060
rect 23348 21020 23354 21032
rect 23385 21029 23397 21032
rect 23431 21029 23443 21063
rect 23385 21023 23443 21029
rect 23842 21020 23848 21072
rect 23900 21060 23906 21072
rect 24228 21060 24256 21091
rect 25240 21072 25268 21100
rect 25498 21088 25504 21140
rect 25556 21128 25562 21140
rect 26881 21131 26939 21137
rect 26881 21128 26893 21131
rect 25556 21100 26893 21128
rect 25556 21088 25562 21100
rect 26881 21097 26893 21100
rect 26927 21097 26939 21131
rect 26881 21091 26939 21097
rect 27062 21088 27068 21140
rect 27120 21128 27126 21140
rect 29454 21128 29460 21140
rect 27120 21100 29460 21128
rect 27120 21088 27126 21100
rect 29454 21088 29460 21100
rect 29512 21128 29518 21140
rect 29733 21131 29791 21137
rect 29512 21100 29684 21128
rect 29512 21088 29518 21100
rect 23900 21032 24256 21060
rect 24765 21063 24823 21069
rect 23900 21020 23906 21032
rect 24765 21029 24777 21063
rect 24811 21029 24823 21063
rect 24765 21023 24823 21029
rect 20533 20995 20591 21001
rect 20533 20992 20545 20995
rect 13740 20964 20024 20992
rect 20272 20964 20545 20992
rect 9508 20896 9674 20924
rect 9401 20887 9459 20893
rect 9416 20856 9444 20887
rect 11330 20884 11336 20936
rect 11388 20884 11394 20936
rect 12618 20924 12624 20936
rect 11900 20896 12624 20924
rect 11333 20883 11391 20884
rect 8036 20828 9352 20856
rect 9416 20828 11284 20856
rect 7837 20791 7895 20797
rect 7837 20757 7849 20791
rect 7883 20757 7895 20791
rect 9324 20788 9352 20828
rect 10594 20788 10600 20800
rect 9324 20760 10600 20788
rect 7837 20751 7895 20757
rect 10594 20748 10600 20760
rect 10652 20748 10658 20800
rect 10686 20748 10692 20800
rect 10744 20748 10750 20800
rect 11054 20748 11060 20800
rect 11112 20788 11118 20800
rect 11149 20791 11207 20797
rect 11149 20788 11161 20791
rect 11112 20760 11161 20788
rect 11112 20748 11118 20760
rect 11149 20757 11161 20760
rect 11195 20757 11207 20791
rect 11256 20788 11284 20828
rect 11900 20788 11928 20896
rect 12618 20884 12624 20896
rect 12676 20884 12682 20936
rect 13740 20933 13768 20964
rect 13725 20927 13783 20933
rect 13725 20893 13737 20927
rect 13771 20893 13783 20927
rect 13725 20887 13783 20893
rect 16025 20927 16083 20933
rect 16025 20893 16037 20927
rect 16071 20924 16083 20927
rect 16758 20924 16764 20936
rect 16071 20896 16764 20924
rect 16071 20893 16083 20896
rect 16025 20887 16083 20893
rect 16758 20884 16764 20896
rect 16816 20884 16822 20936
rect 18877 20927 18935 20933
rect 18877 20893 18889 20927
rect 18923 20924 18935 20927
rect 19334 20924 19340 20936
rect 18923 20896 19340 20924
rect 18923 20893 18935 20896
rect 18877 20887 18935 20893
rect 19334 20884 19340 20896
rect 19392 20924 19398 20936
rect 19392 20896 19564 20924
rect 19392 20884 19398 20896
rect 11977 20859 12035 20865
rect 11977 20825 11989 20859
rect 12023 20856 12035 20859
rect 12066 20856 12072 20868
rect 12023 20828 12072 20856
rect 12023 20825 12035 20828
rect 11977 20819 12035 20825
rect 12066 20816 12072 20828
rect 12124 20816 12130 20868
rect 12897 20859 12955 20865
rect 12897 20825 12909 20859
rect 12943 20825 12955 20859
rect 12897 20819 12955 20825
rect 11256 20760 11928 20788
rect 11149 20751 11207 20757
rect 12618 20748 12624 20800
rect 12676 20788 12682 20800
rect 12912 20788 12940 20819
rect 15194 20816 15200 20868
rect 15252 20816 15258 20868
rect 15749 20859 15807 20865
rect 15749 20825 15761 20859
rect 15795 20856 15807 20859
rect 16114 20856 16120 20868
rect 15795 20828 16120 20856
rect 15795 20825 15807 20828
rect 15749 20819 15807 20825
rect 16114 20816 16120 20828
rect 16172 20816 16178 20868
rect 16669 20859 16727 20865
rect 16669 20825 16681 20859
rect 16715 20856 16727 20859
rect 16715 20828 17356 20856
rect 16715 20825 16727 20828
rect 16669 20819 16727 20825
rect 12676 20760 12940 20788
rect 12676 20748 12682 20760
rect 13538 20748 13544 20800
rect 13596 20748 13602 20800
rect 17328 20788 17356 20828
rect 17862 20816 17868 20868
rect 17920 20816 17926 20868
rect 18601 20859 18659 20865
rect 18601 20825 18613 20859
rect 18647 20856 18659 20859
rect 19426 20856 19432 20868
rect 18647 20828 19432 20856
rect 18647 20825 18659 20828
rect 18601 20819 18659 20825
rect 19426 20816 19432 20828
rect 19484 20816 19490 20868
rect 18506 20788 18512 20800
rect 17328 20760 18512 20788
rect 18506 20748 18512 20760
rect 18564 20748 18570 20800
rect 19334 20748 19340 20800
rect 19392 20748 19398 20800
rect 19536 20797 19564 20896
rect 19794 20884 19800 20936
rect 19852 20924 19858 20936
rect 20272 20924 20300 20964
rect 20533 20961 20545 20964
rect 20579 20961 20591 20995
rect 22646 20992 22652 21004
rect 20533 20955 20591 20961
rect 21192 20964 22652 20992
rect 19852 20896 20300 20924
rect 20349 20927 20407 20933
rect 19852 20884 19858 20896
rect 20349 20893 20361 20927
rect 20395 20924 20407 20927
rect 21192 20924 21220 20964
rect 22646 20952 22652 20964
rect 22704 20952 22710 21004
rect 24780 20992 24808 21023
rect 25222 21020 25228 21072
rect 25280 21060 25286 21072
rect 25409 21063 25467 21069
rect 25409 21060 25421 21063
rect 25280 21032 25421 21060
rect 25280 21020 25286 21032
rect 25409 21029 25421 21032
rect 25455 21060 25467 21063
rect 25774 21060 25780 21072
rect 25455 21032 25780 21060
rect 25455 21029 25467 21032
rect 25409 21023 25467 21029
rect 25774 21020 25780 21032
rect 25832 21020 25838 21072
rect 26142 21020 26148 21072
rect 26200 21060 26206 21072
rect 29546 21060 29552 21072
rect 26200 21032 29552 21060
rect 26200 21020 26206 21032
rect 29546 21020 29552 21032
rect 29604 21020 29610 21072
rect 29656 21060 29684 21100
rect 29733 21097 29745 21131
rect 29779 21128 29791 21131
rect 29914 21128 29920 21140
rect 29779 21100 29920 21128
rect 29779 21097 29791 21100
rect 29733 21091 29791 21097
rect 29914 21088 29920 21100
rect 29972 21088 29978 21140
rect 30006 21088 30012 21140
rect 30064 21128 30070 21140
rect 30193 21131 30251 21137
rect 30193 21128 30205 21131
rect 30064 21100 30205 21128
rect 30064 21088 30070 21100
rect 30193 21097 30205 21100
rect 30239 21097 30251 21131
rect 35710 21128 35716 21140
rect 30193 21091 30251 21097
rect 31312 21100 35716 21128
rect 30377 21063 30435 21069
rect 30377 21060 30389 21063
rect 29656 21032 30389 21060
rect 30377 21029 30389 21032
rect 30423 21029 30435 21063
rect 30377 21023 30435 21029
rect 26234 20992 26240 21004
rect 24780 20964 26240 20992
rect 26234 20952 26240 20964
rect 26292 20952 26298 21004
rect 26326 20952 26332 21004
rect 26384 20952 26390 21004
rect 27890 20952 27896 21004
rect 27948 20952 27954 21004
rect 31312 21001 31340 21100
rect 35710 21088 35716 21100
rect 35768 21088 35774 21140
rect 36722 21088 36728 21140
rect 36780 21128 36786 21140
rect 37642 21128 37648 21140
rect 36780 21100 37648 21128
rect 36780 21088 36786 21100
rect 37642 21088 37648 21100
rect 37700 21088 37706 21140
rect 38378 21128 38384 21140
rect 37752 21100 38384 21128
rect 31938 21020 31944 21072
rect 31996 21020 32002 21072
rect 34882 21020 34888 21072
rect 34940 21020 34946 21072
rect 37369 21063 37427 21069
rect 37369 21029 37381 21063
rect 37415 21060 37427 21063
rect 37752 21060 37780 21100
rect 38378 21088 38384 21100
rect 38436 21088 38442 21140
rect 40037 21131 40095 21137
rect 40037 21097 40049 21131
rect 40083 21128 40095 21131
rect 40126 21128 40132 21140
rect 40083 21100 40132 21128
rect 40083 21097 40095 21100
rect 40037 21091 40095 21097
rect 40126 21088 40132 21100
rect 40184 21088 40190 21140
rect 40494 21088 40500 21140
rect 40552 21128 40558 21140
rect 41322 21128 41328 21140
rect 40552 21100 41328 21128
rect 40552 21088 40558 21100
rect 41322 21088 41328 21100
rect 41380 21088 41386 21140
rect 41414 21088 41420 21140
rect 41472 21128 41478 21140
rect 42429 21131 42487 21137
rect 42429 21128 42441 21131
rect 41472 21100 42441 21128
rect 41472 21088 41478 21100
rect 42429 21097 42441 21100
rect 42475 21097 42487 21131
rect 42429 21091 42487 21097
rect 42610 21088 42616 21140
rect 42668 21128 42674 21140
rect 42981 21131 43039 21137
rect 42981 21128 42993 21131
rect 42668 21100 42993 21128
rect 42668 21088 42674 21100
rect 42981 21097 42993 21100
rect 43027 21097 43039 21131
rect 42981 21091 43039 21097
rect 46842 21088 46848 21140
rect 46900 21128 46906 21140
rect 48041 21131 48099 21137
rect 48041 21128 48053 21131
rect 46900 21100 48053 21128
rect 46900 21088 46906 21100
rect 48041 21097 48053 21100
rect 48087 21097 48099 21131
rect 48041 21091 48099 21097
rect 48590 21088 48596 21140
rect 48648 21088 48654 21140
rect 37415 21032 37780 21060
rect 37415 21029 37427 21032
rect 37369 21023 37427 21029
rect 40218 21020 40224 21072
rect 40276 21060 40282 21072
rect 41046 21060 41052 21072
rect 40276 21032 41052 21060
rect 40276 21020 40282 21032
rect 41046 21020 41052 21032
rect 41104 21060 41110 21072
rect 49145 21063 49203 21069
rect 49145 21060 49157 21063
rect 41104 21032 49157 21060
rect 41104 21020 41110 21032
rect 49145 21029 49157 21032
rect 49191 21029 49203 21063
rect 49145 21023 49203 21029
rect 49326 21020 49332 21072
rect 49384 21020 49390 21072
rect 28537 20995 28595 21001
rect 28537 20961 28549 20995
rect 28583 20992 28595 20995
rect 31297 20995 31355 21001
rect 28583 20964 30144 20992
rect 28583 20961 28595 20964
rect 28537 20955 28595 20961
rect 20395 20896 21220 20924
rect 20395 20893 20407 20896
rect 20349 20887 20407 20893
rect 22922 20884 22928 20936
rect 22980 20884 22986 20936
rect 24118 20884 24124 20936
rect 24176 20924 24182 20936
rect 24581 20927 24639 20933
rect 24581 20924 24593 20927
rect 24176 20896 24593 20924
rect 24176 20884 24182 20896
rect 24581 20893 24593 20896
rect 24627 20893 24639 20927
rect 24581 20887 24639 20893
rect 26970 20884 26976 20936
rect 27028 20924 27034 20936
rect 29730 20924 29736 20936
rect 27028 20896 29736 20924
rect 27028 20884 27034 20896
rect 29730 20884 29736 20896
rect 29788 20884 29794 20936
rect 29914 20884 29920 20936
rect 29972 20884 29978 20936
rect 30116 20924 30144 20964
rect 31297 20961 31309 20995
rect 31343 20961 31355 20995
rect 31297 20955 31355 20961
rect 31481 20995 31539 21001
rect 31481 20961 31493 20995
rect 31527 20992 31539 20995
rect 32306 20992 32312 21004
rect 31527 20964 32312 20992
rect 31527 20961 31539 20964
rect 31481 20955 31539 20961
rect 32306 20952 32312 20964
rect 32364 20992 32370 21004
rect 32769 20995 32827 21001
rect 32769 20992 32781 20995
rect 32364 20964 32781 20992
rect 32364 20952 32370 20964
rect 32769 20961 32781 20964
rect 32815 20961 32827 20995
rect 32769 20955 32827 20961
rect 33134 20952 33140 21004
rect 33192 20992 33198 21004
rect 33502 20992 33508 21004
rect 33192 20964 33508 20992
rect 33192 20952 33198 20964
rect 33502 20952 33508 20964
rect 33560 20952 33566 21004
rect 34330 20952 34336 21004
rect 34388 20992 34394 21004
rect 38654 20992 38660 21004
rect 34388 20964 36676 20992
rect 34388 20952 34394 20964
rect 32398 20924 32404 20936
rect 30116 20896 32404 20924
rect 32398 20884 32404 20896
rect 32456 20884 32462 20936
rect 32490 20884 32496 20936
rect 32548 20884 32554 20936
rect 36648 20933 36676 20964
rect 37660 20964 38660 20992
rect 36633 20927 36691 20933
rect 36633 20893 36645 20927
rect 36679 20924 36691 20927
rect 36679 20896 37228 20924
rect 36679 20893 36691 20896
rect 36633 20887 36691 20893
rect 20441 20859 20499 20865
rect 20441 20825 20453 20859
rect 20487 20856 20499 20859
rect 22370 20856 22376 20868
rect 20487 20828 21312 20856
rect 22218 20828 22376 20856
rect 20487 20825 20499 20828
rect 20441 20819 20499 20825
rect 19521 20791 19579 20797
rect 19521 20757 19533 20791
rect 19567 20788 19579 20791
rect 19610 20788 19616 20800
rect 19567 20760 19616 20788
rect 19567 20757 19579 20760
rect 19521 20751 19579 20757
rect 19610 20748 19616 20760
rect 19668 20748 19674 20800
rect 21284 20788 21312 20828
rect 22370 20816 22376 20828
rect 22428 20856 22434 20868
rect 22554 20856 22560 20868
rect 22428 20828 22560 20856
rect 22428 20816 22434 20828
rect 22554 20816 22560 20828
rect 22612 20816 22618 20868
rect 22649 20859 22707 20865
rect 22649 20825 22661 20859
rect 22695 20856 22707 20859
rect 22738 20856 22744 20868
rect 22695 20828 22744 20856
rect 22695 20825 22707 20828
rect 22649 20819 22707 20825
rect 22738 20816 22744 20828
rect 22796 20816 22802 20868
rect 23566 20816 23572 20868
rect 23624 20816 23630 20868
rect 25958 20856 25964 20868
rect 24044 20828 25964 20856
rect 24044 20788 24072 20828
rect 25958 20816 25964 20828
rect 26016 20816 26022 20868
rect 26053 20859 26111 20865
rect 26053 20825 26065 20859
rect 26099 20856 26111 20859
rect 26786 20856 26792 20868
rect 26099 20828 26792 20856
rect 26099 20825 26111 20828
rect 26053 20819 26111 20825
rect 26786 20816 26792 20828
rect 26844 20816 26850 20868
rect 27430 20816 27436 20868
rect 27488 20816 27494 20868
rect 28350 20816 28356 20868
rect 28408 20856 28414 20868
rect 28408 20828 30880 20856
rect 28408 20816 28414 20828
rect 21284 20760 24072 20788
rect 24118 20748 24124 20800
rect 24176 20788 24182 20800
rect 25685 20791 25743 20797
rect 25685 20788 25697 20791
rect 24176 20760 25697 20788
rect 24176 20748 24182 20760
rect 25685 20757 25697 20760
rect 25731 20757 25743 20791
rect 25685 20751 25743 20757
rect 26142 20748 26148 20800
rect 26200 20748 26206 20800
rect 26697 20791 26755 20797
rect 26697 20757 26709 20791
rect 26743 20788 26755 20791
rect 26878 20788 26884 20800
rect 26743 20760 26884 20788
rect 26743 20757 26755 20760
rect 26697 20751 26755 20757
rect 26878 20748 26884 20760
rect 26936 20788 26942 20800
rect 27154 20788 27160 20800
rect 26936 20760 27160 20788
rect 26936 20748 26942 20760
rect 27154 20748 27160 20760
rect 27212 20748 27218 20800
rect 27614 20748 27620 20800
rect 27672 20788 27678 20800
rect 28629 20791 28687 20797
rect 28629 20788 28641 20791
rect 27672 20760 28641 20788
rect 27672 20748 27678 20760
rect 28629 20757 28641 20760
rect 28675 20757 28687 20791
rect 28629 20751 28687 20757
rect 28718 20748 28724 20800
rect 28776 20748 28782 20800
rect 29089 20791 29147 20797
rect 29089 20757 29101 20791
rect 29135 20788 29147 20791
rect 30098 20788 30104 20800
rect 29135 20760 30104 20788
rect 29135 20757 29147 20760
rect 29089 20751 29147 20757
rect 30098 20748 30104 20760
rect 30156 20748 30162 20800
rect 30852 20797 30880 20828
rect 32122 20816 32128 20868
rect 32180 20856 32186 20868
rect 35066 20856 35072 20868
rect 32180 20828 33258 20856
rect 34072 20828 35072 20856
rect 32180 20816 32186 20828
rect 30837 20791 30895 20797
rect 30837 20757 30849 20791
rect 30883 20757 30895 20791
rect 30837 20751 30895 20757
rect 31202 20748 31208 20800
rect 31260 20748 31266 20800
rect 31478 20748 31484 20800
rect 31536 20788 31542 20800
rect 32950 20788 32956 20800
rect 31536 20760 32956 20788
rect 31536 20748 31542 20760
rect 32950 20748 32956 20760
rect 33008 20748 33014 20800
rect 33152 20788 33180 20828
rect 34072 20788 34100 20828
rect 35066 20816 35072 20828
rect 35124 20856 35130 20868
rect 35124 20828 35190 20856
rect 35124 20816 35130 20828
rect 36354 20816 36360 20868
rect 36412 20816 36418 20868
rect 37200 20865 37228 20896
rect 37185 20859 37243 20865
rect 36464 20828 37136 20856
rect 33152 20760 34100 20788
rect 34241 20791 34299 20797
rect 34241 20757 34253 20791
rect 34287 20788 34299 20791
rect 34330 20788 34336 20800
rect 34287 20760 34336 20788
rect 34287 20757 34299 20760
rect 34241 20751 34299 20757
rect 34330 20748 34336 20760
rect 34388 20788 34394 20800
rect 36464 20788 36492 20828
rect 34388 20760 36492 20788
rect 34388 20748 34394 20760
rect 36998 20748 37004 20800
rect 37056 20748 37062 20800
rect 37108 20788 37136 20828
rect 37185 20825 37197 20859
rect 37231 20856 37243 20859
rect 37550 20856 37556 20868
rect 37231 20828 37556 20856
rect 37231 20825 37243 20828
rect 37185 20819 37243 20825
rect 37550 20816 37556 20828
rect 37608 20816 37614 20868
rect 37660 20788 37688 20964
rect 38654 20952 38660 20964
rect 38712 20952 38718 21004
rect 39114 20952 39120 21004
rect 39172 20992 39178 21004
rect 39393 20995 39451 21001
rect 39393 20992 39405 20995
rect 39172 20964 39405 20992
rect 39172 20952 39178 20964
rect 39393 20961 39405 20964
rect 39439 20992 39451 20995
rect 39574 20992 39580 21004
rect 39439 20964 39580 20992
rect 39439 20961 39451 20964
rect 39393 20955 39451 20961
rect 39574 20952 39580 20964
rect 39632 20952 39638 21004
rect 39758 20952 39764 21004
rect 39816 20992 39822 21004
rect 40497 20995 40555 21001
rect 40497 20992 40509 20995
rect 39816 20964 40509 20992
rect 39816 20952 39822 20964
rect 40497 20961 40509 20964
rect 40543 20961 40555 20995
rect 40497 20955 40555 20961
rect 40589 20995 40647 21001
rect 40589 20961 40601 20995
rect 40635 20961 40647 20995
rect 40589 20955 40647 20961
rect 40604 20924 40632 20955
rect 40678 20952 40684 21004
rect 40736 20992 40742 21004
rect 41785 20995 41843 21001
rect 41785 20992 41797 20995
rect 40736 20964 41797 20992
rect 40736 20952 40742 20964
rect 41785 20961 41797 20964
rect 41831 20961 41843 20995
rect 41785 20955 41843 20961
rect 42426 20952 42432 21004
rect 42484 20992 42490 21004
rect 42613 20995 42671 21001
rect 42613 20992 42625 20995
rect 42484 20964 42625 20992
rect 42484 20952 42490 20964
rect 42613 20961 42625 20964
rect 42659 20961 42671 20995
rect 42613 20955 42671 20961
rect 42889 20995 42947 21001
rect 42889 20961 42901 20995
rect 42935 20992 42947 20995
rect 43346 20992 43352 21004
rect 42935 20964 43352 20992
rect 42935 20961 42947 20964
rect 42889 20955 42947 20961
rect 43346 20952 43352 20964
rect 43404 20952 43410 21004
rect 47949 20995 48007 21001
rect 47949 20961 47961 20995
rect 47995 20992 48007 20995
rect 49344 20992 49372 21020
rect 47995 20964 49372 20992
rect 47995 20961 48007 20964
rect 47949 20955 48007 20961
rect 40328 20896 40632 20924
rect 38378 20816 38384 20868
rect 38436 20816 38442 20868
rect 39022 20816 39028 20868
rect 39080 20856 39086 20868
rect 39117 20859 39175 20865
rect 39117 20856 39129 20859
rect 39080 20828 39129 20856
rect 39080 20816 39086 20828
rect 39117 20825 39129 20828
rect 39163 20856 39175 20859
rect 40328 20856 40356 20896
rect 41598 20884 41604 20936
rect 41656 20884 41662 20936
rect 48409 20927 48467 20933
rect 48409 20893 48421 20927
rect 48455 20924 48467 20927
rect 49326 20924 49332 20936
rect 48455 20896 49332 20924
rect 48455 20893 48467 20896
rect 48409 20887 48467 20893
rect 49326 20884 49332 20896
rect 49384 20884 49390 20936
rect 39163 20828 40356 20856
rect 40405 20859 40463 20865
rect 39163 20825 39175 20828
rect 39117 20819 39175 20825
rect 40405 20825 40417 20859
rect 40451 20856 40463 20859
rect 48777 20859 48835 20865
rect 40451 20828 41276 20856
rect 40451 20825 40463 20828
rect 40405 20819 40463 20825
rect 37108 20760 37688 20788
rect 38286 20748 38292 20800
rect 38344 20788 38350 20800
rect 40678 20788 40684 20800
rect 38344 20760 40684 20788
rect 38344 20748 38350 20760
rect 40678 20748 40684 20760
rect 40736 20748 40742 20800
rect 41248 20797 41276 20828
rect 48777 20825 48789 20859
rect 48823 20856 48835 20859
rect 49418 20856 49424 20868
rect 48823 20828 49424 20856
rect 48823 20825 48835 20828
rect 48777 20819 48835 20825
rect 49418 20816 49424 20828
rect 49476 20816 49482 20868
rect 41233 20791 41291 20797
rect 41233 20757 41245 20791
rect 41279 20757 41291 20791
rect 41233 20751 41291 20757
rect 41322 20748 41328 20800
rect 41380 20788 41386 20800
rect 41693 20791 41751 20797
rect 41693 20788 41705 20791
rect 41380 20760 41705 20788
rect 41380 20748 41386 20760
rect 41693 20757 41705 20760
rect 41739 20788 41751 20791
rect 42245 20791 42303 20797
rect 42245 20788 42257 20791
rect 41739 20760 42257 20788
rect 41739 20757 41751 20760
rect 41693 20751 41751 20757
rect 42245 20757 42257 20760
rect 42291 20788 42303 20791
rect 46198 20788 46204 20800
rect 42291 20760 46204 20788
rect 42291 20757 42303 20760
rect 42245 20751 42303 20757
rect 46198 20748 46204 20760
rect 46256 20748 46262 20800
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 5445 20587 5503 20593
rect 5445 20553 5457 20587
rect 5491 20584 5503 20587
rect 6638 20584 6644 20596
rect 5491 20556 6644 20584
rect 5491 20553 5503 20556
rect 5445 20547 5503 20553
rect 6638 20544 6644 20556
rect 6696 20544 6702 20596
rect 9674 20544 9680 20596
rect 9732 20544 9738 20596
rect 10318 20544 10324 20596
rect 10376 20544 10382 20596
rect 11149 20587 11207 20593
rect 11149 20553 11161 20587
rect 11195 20584 11207 20587
rect 11195 20556 12664 20584
rect 11195 20553 11207 20556
rect 11149 20547 11207 20553
rect 1302 20476 1308 20528
rect 1360 20516 1366 20528
rect 3605 20519 3663 20525
rect 3605 20516 3617 20519
rect 1360 20488 3617 20516
rect 1360 20476 1366 20488
rect 3605 20485 3617 20488
rect 3651 20485 3663 20519
rect 8294 20516 8300 20528
rect 3605 20479 3663 20485
rect 5276 20488 8300 20516
rect 2961 20451 3019 20457
rect 2961 20417 2973 20451
rect 3007 20448 3019 20451
rect 3970 20448 3976 20460
rect 3007 20420 3976 20448
rect 3007 20417 3019 20420
rect 2961 20411 3019 20417
rect 3970 20408 3976 20420
rect 4028 20408 4034 20460
rect 4798 20408 4804 20460
rect 4856 20408 4862 20460
rect 5276 20457 5304 20488
rect 8294 20476 8300 20488
rect 8352 20476 8358 20528
rect 10962 20516 10968 20528
rect 9876 20488 10968 20516
rect 5261 20451 5319 20457
rect 5261 20417 5273 20451
rect 5307 20417 5319 20451
rect 5261 20411 5319 20417
rect 5442 20408 5448 20460
rect 5500 20448 5506 20460
rect 6549 20451 6607 20457
rect 6549 20448 6561 20451
rect 5500 20420 6561 20448
rect 5500 20408 5506 20420
rect 6549 20417 6561 20420
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 9217 20451 9275 20457
rect 9217 20417 9229 20451
rect 9263 20448 9275 20451
rect 9674 20448 9680 20460
rect 9263 20420 9680 20448
rect 9263 20417 9275 20420
rect 9217 20411 9275 20417
rect 9674 20408 9680 20420
rect 9732 20408 9738 20460
rect 9876 20457 9904 20488
rect 10962 20476 10968 20488
rect 11020 20476 11026 20528
rect 12342 20476 12348 20528
rect 12400 20516 12406 20528
rect 12437 20519 12495 20525
rect 12437 20516 12449 20519
rect 12400 20488 12449 20516
rect 12400 20476 12406 20488
rect 12437 20485 12449 20488
rect 12483 20485 12495 20519
rect 12636 20516 12664 20556
rect 12710 20544 12716 20596
rect 12768 20584 12774 20596
rect 13725 20587 13783 20593
rect 13725 20584 13737 20587
rect 12768 20556 13737 20584
rect 12768 20544 12774 20556
rect 13725 20553 13737 20556
rect 13771 20553 13783 20587
rect 13725 20547 13783 20553
rect 14090 20544 14096 20596
rect 14148 20544 14154 20596
rect 14918 20544 14924 20596
rect 14976 20544 14982 20596
rect 15470 20544 15476 20596
rect 15528 20584 15534 20596
rect 15565 20587 15623 20593
rect 15565 20584 15577 20587
rect 15528 20556 15577 20584
rect 15528 20544 15534 20556
rect 15565 20553 15577 20556
rect 15611 20553 15623 20587
rect 15565 20547 15623 20553
rect 15838 20544 15844 20596
rect 15896 20584 15902 20596
rect 15933 20587 15991 20593
rect 15933 20584 15945 20587
rect 15896 20556 15945 20584
rect 15896 20544 15902 20556
rect 15933 20553 15945 20556
rect 15979 20553 15991 20587
rect 15933 20547 15991 20553
rect 16022 20544 16028 20596
rect 16080 20544 16086 20596
rect 16390 20584 16396 20596
rect 16132 20556 16396 20584
rect 13906 20516 13912 20528
rect 12636 20488 13912 20516
rect 12437 20479 12495 20485
rect 13906 20476 13912 20488
rect 13964 20476 13970 20528
rect 16132 20516 16160 20556
rect 16390 20544 16396 20556
rect 16448 20544 16454 20596
rect 17126 20544 17132 20596
rect 17184 20544 17190 20596
rect 17954 20544 17960 20596
rect 18012 20584 18018 20596
rect 18785 20587 18843 20593
rect 18012 20556 18644 20584
rect 18012 20544 18018 20556
rect 17144 20516 17172 20544
rect 18616 20516 18644 20556
rect 18785 20553 18797 20587
rect 18831 20584 18843 20587
rect 18874 20584 18880 20596
rect 18831 20556 18880 20584
rect 18831 20553 18843 20556
rect 18785 20547 18843 20553
rect 18874 20544 18880 20556
rect 18932 20544 18938 20596
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 19702 20584 19708 20596
rect 19484 20556 19708 20584
rect 19484 20544 19490 20556
rect 19702 20544 19708 20556
rect 19760 20584 19766 20596
rect 20162 20584 20168 20596
rect 19760 20556 20168 20584
rect 19760 20544 19766 20556
rect 20162 20544 20168 20556
rect 20220 20544 20226 20596
rect 21082 20544 21088 20596
rect 21140 20584 21146 20596
rect 21726 20584 21732 20596
rect 21140 20556 21732 20584
rect 21140 20544 21146 20556
rect 21726 20544 21732 20556
rect 21784 20584 21790 20596
rect 22738 20584 22744 20596
rect 21784 20556 22744 20584
rect 21784 20544 21790 20556
rect 22738 20544 22744 20556
rect 22796 20544 22802 20596
rect 22922 20544 22928 20596
rect 22980 20584 22986 20596
rect 25682 20584 25688 20596
rect 22980 20556 25688 20584
rect 22980 20544 22986 20556
rect 19058 20516 19064 20528
rect 14016 20488 16160 20516
rect 16224 20488 17172 20516
rect 18538 20488 19064 20516
rect 9861 20451 9919 20457
rect 9861 20417 9873 20451
rect 9907 20417 9919 20451
rect 9861 20411 9919 20417
rect 10505 20451 10563 20457
rect 10505 20417 10517 20451
rect 10551 20417 10563 20451
rect 10505 20411 10563 20417
rect 2501 20383 2559 20389
rect 2501 20349 2513 20383
rect 2547 20380 2559 20383
rect 2547 20352 2774 20380
rect 2547 20349 2559 20352
rect 2501 20343 2559 20349
rect 2746 20324 2774 20352
rect 5902 20340 5908 20392
rect 5960 20380 5966 20392
rect 7009 20383 7067 20389
rect 7009 20380 7021 20383
rect 5960 20352 7021 20380
rect 5960 20340 5966 20352
rect 7009 20349 7021 20352
rect 7055 20349 7067 20383
rect 10520 20380 10548 20411
rect 10870 20408 10876 20460
rect 10928 20448 10934 20460
rect 11701 20451 11759 20457
rect 11701 20448 11713 20451
rect 10928 20420 11713 20448
rect 10928 20408 10934 20420
rect 11701 20417 11713 20420
rect 11747 20417 11759 20451
rect 11701 20411 11759 20417
rect 11790 20408 11796 20460
rect 11848 20448 11854 20460
rect 11885 20451 11943 20457
rect 11885 20448 11897 20451
rect 11848 20420 11897 20448
rect 11848 20408 11854 20420
rect 11885 20417 11897 20420
rect 11931 20448 11943 20451
rect 12621 20451 12679 20457
rect 11931 20420 12572 20448
rect 11931 20417 11943 20420
rect 11885 20411 11943 20417
rect 12342 20380 12348 20392
rect 10520 20352 12348 20380
rect 7009 20343 7067 20349
rect 12342 20340 12348 20352
rect 12400 20340 12406 20392
rect 12544 20380 12572 20420
rect 12621 20417 12633 20451
rect 12667 20448 12679 20451
rect 12894 20448 12900 20460
rect 12667 20420 12900 20448
rect 12667 20417 12679 20420
rect 12621 20411 12679 20417
rect 12894 20408 12900 20420
rect 12952 20408 12958 20460
rect 14016 20380 14044 20488
rect 14185 20451 14243 20457
rect 14185 20417 14197 20451
rect 14231 20448 14243 20451
rect 15010 20448 15016 20460
rect 14231 20420 15016 20448
rect 14231 20417 14243 20420
rect 14185 20411 14243 20417
rect 15010 20408 15016 20420
rect 15068 20408 15074 20460
rect 15105 20451 15163 20457
rect 15105 20417 15117 20451
rect 15151 20417 15163 20451
rect 15105 20411 15163 20417
rect 12544 20352 14044 20380
rect 14274 20340 14280 20392
rect 14332 20340 14338 20392
rect 2746 20284 2780 20324
rect 2774 20272 2780 20284
rect 2832 20272 2838 20324
rect 3326 20272 3332 20324
rect 3384 20312 3390 20324
rect 14918 20312 14924 20324
rect 3384 20284 9674 20312
rect 3384 20272 3390 20284
rect 4154 20204 4160 20256
rect 4212 20244 4218 20256
rect 9033 20247 9091 20253
rect 9033 20244 9045 20247
rect 4212 20216 9045 20244
rect 4212 20204 4218 20216
rect 9033 20213 9045 20216
rect 9079 20213 9091 20247
rect 9646 20244 9674 20284
rect 12636 20284 14924 20312
rect 12636 20244 12664 20284
rect 14918 20272 14924 20284
rect 14976 20272 14982 20324
rect 15120 20312 15148 20411
rect 16224 20389 16252 20488
rect 19058 20476 19064 20488
rect 19116 20516 19122 20528
rect 19334 20516 19340 20528
rect 19116 20488 19340 20516
rect 19116 20476 19122 20488
rect 19334 20476 19340 20488
rect 19392 20516 19398 20528
rect 22373 20519 22431 20525
rect 19392 20488 20010 20516
rect 19392 20476 19398 20488
rect 22373 20485 22385 20519
rect 22419 20516 22431 20519
rect 23750 20516 23756 20528
rect 22419 20488 23756 20516
rect 22419 20485 22431 20488
rect 22373 20479 22431 20485
rect 23750 20476 23756 20488
rect 23808 20476 23814 20528
rect 16758 20408 16764 20460
rect 16816 20448 16822 20460
rect 17037 20451 17095 20457
rect 17037 20448 17049 20451
rect 16816 20420 17049 20448
rect 16816 20408 16822 20420
rect 17037 20417 17049 20420
rect 17083 20417 17095 20451
rect 17037 20411 17095 20417
rect 21453 20451 21511 20457
rect 21453 20417 21465 20451
rect 21499 20448 21511 20451
rect 22186 20448 22192 20460
rect 21499 20420 22192 20448
rect 21499 20417 21511 20420
rect 21453 20411 21511 20417
rect 22186 20408 22192 20420
rect 22244 20408 22250 20460
rect 23382 20408 23388 20460
rect 23440 20408 23446 20460
rect 23860 20457 23888 20556
rect 25682 20544 25688 20556
rect 25740 20544 25746 20596
rect 25774 20544 25780 20596
rect 25832 20584 25838 20596
rect 26326 20584 26332 20596
rect 25832 20556 26332 20584
rect 25832 20544 25838 20556
rect 26326 20544 26332 20556
rect 26384 20544 26390 20596
rect 30834 20584 30840 20596
rect 27264 20556 30840 20584
rect 26970 20516 26976 20528
rect 25424 20488 26976 20516
rect 23845 20451 23903 20457
rect 23845 20417 23857 20451
rect 23891 20417 23903 20451
rect 23845 20411 23903 20417
rect 25222 20408 25228 20460
rect 25280 20408 25286 20460
rect 16209 20383 16267 20389
rect 16209 20349 16221 20383
rect 16255 20349 16267 20383
rect 16209 20343 16267 20349
rect 16850 20340 16856 20392
rect 16908 20380 16914 20392
rect 17313 20383 17371 20389
rect 17313 20380 17325 20383
rect 16908 20352 17325 20380
rect 16908 20340 16914 20352
rect 17313 20349 17325 20352
rect 17359 20380 17371 20383
rect 20438 20380 20444 20392
rect 17359 20352 20444 20380
rect 17359 20349 17371 20352
rect 17313 20343 17371 20349
rect 20438 20340 20444 20352
rect 20496 20340 20502 20392
rect 21174 20340 21180 20392
rect 21232 20380 21238 20392
rect 21232 20352 22416 20380
rect 21232 20340 21238 20352
rect 16482 20312 16488 20324
rect 15120 20284 16488 20312
rect 16482 20272 16488 20284
rect 16540 20272 16546 20324
rect 19058 20272 19064 20324
rect 19116 20272 19122 20324
rect 22388 20312 22416 20352
rect 22462 20340 22468 20392
rect 22520 20340 22526 20392
rect 22554 20340 22560 20392
rect 22612 20340 22618 20392
rect 24121 20383 24179 20389
rect 24121 20349 24133 20383
rect 24167 20380 24179 20383
rect 24210 20380 24216 20392
rect 24167 20352 24216 20380
rect 24167 20349 24179 20352
rect 24121 20343 24179 20349
rect 24210 20340 24216 20352
rect 24268 20380 24274 20392
rect 25424 20380 25452 20488
rect 26970 20476 26976 20488
rect 27028 20476 27034 20528
rect 25498 20408 25504 20460
rect 25556 20448 25562 20460
rect 27264 20457 27292 20556
rect 30834 20544 30840 20556
rect 30892 20584 30898 20596
rect 31478 20584 31484 20596
rect 30892 20556 31484 20584
rect 30892 20544 30898 20556
rect 31478 20544 31484 20556
rect 31536 20584 31542 20596
rect 32490 20584 32496 20596
rect 31536 20556 32496 20584
rect 31536 20544 31542 20556
rect 32490 20544 32496 20556
rect 32548 20584 32554 20596
rect 35253 20587 35311 20593
rect 32548 20556 34100 20584
rect 32548 20544 32554 20556
rect 27798 20476 27804 20528
rect 27856 20516 27862 20528
rect 27856 20488 28014 20516
rect 27856 20476 27862 20488
rect 29822 20476 29828 20528
rect 29880 20476 29886 20528
rect 31021 20519 31079 20525
rect 31021 20485 31033 20519
rect 31067 20516 31079 20519
rect 31110 20516 31116 20528
rect 31067 20488 31116 20516
rect 31067 20485 31079 20488
rect 31021 20479 31079 20485
rect 31110 20476 31116 20488
rect 31168 20476 31174 20528
rect 31757 20519 31815 20525
rect 31757 20485 31769 20519
rect 31803 20516 31815 20519
rect 31846 20516 31852 20528
rect 31803 20488 31852 20516
rect 31803 20485 31815 20488
rect 31757 20479 31815 20485
rect 31846 20476 31852 20488
rect 31904 20476 31910 20528
rect 32122 20476 32128 20528
rect 32180 20516 32186 20528
rect 32180 20488 32614 20516
rect 32180 20476 32186 20488
rect 26053 20451 26111 20457
rect 26053 20448 26065 20451
rect 25556 20420 26065 20448
rect 25556 20408 25562 20420
rect 26053 20417 26065 20420
rect 26099 20417 26111 20451
rect 26053 20411 26111 20417
rect 27249 20451 27307 20457
rect 27249 20417 27261 20451
rect 27295 20417 27307 20451
rect 27249 20411 27307 20417
rect 28902 20408 28908 20460
rect 28960 20448 28966 20460
rect 29733 20451 29791 20457
rect 28960 20420 29684 20448
rect 28960 20408 28966 20420
rect 24268 20352 25452 20380
rect 24268 20340 24274 20352
rect 25590 20340 25596 20392
rect 25648 20380 25654 20392
rect 25774 20380 25780 20392
rect 25648 20352 25780 20380
rect 25648 20340 25654 20352
rect 25774 20340 25780 20352
rect 25832 20340 25838 20392
rect 25866 20340 25872 20392
rect 25924 20380 25930 20392
rect 27525 20383 27583 20389
rect 27525 20380 27537 20383
rect 25924 20352 27537 20380
rect 25924 20340 25930 20352
rect 27525 20349 27537 20352
rect 27571 20349 27583 20383
rect 27525 20343 27583 20349
rect 28997 20383 29055 20389
rect 28997 20349 29009 20383
rect 29043 20380 29055 20383
rect 29270 20380 29276 20392
rect 29043 20352 29276 20380
rect 29043 20349 29055 20352
rect 28997 20343 29055 20349
rect 29270 20340 29276 20352
rect 29328 20340 29334 20392
rect 29454 20340 29460 20392
rect 29512 20380 29518 20392
rect 29549 20383 29607 20389
rect 29549 20380 29561 20383
rect 29512 20352 29561 20380
rect 29512 20340 29518 20352
rect 29549 20349 29561 20352
rect 29595 20349 29607 20383
rect 29656 20380 29684 20420
rect 29733 20417 29745 20451
rect 29779 20448 29791 20451
rect 30190 20448 30196 20460
rect 29779 20420 30196 20448
rect 29779 20417 29791 20420
rect 29733 20411 29791 20417
rect 30190 20408 30196 20420
rect 30248 20408 30254 20460
rect 30282 20408 30288 20460
rect 30340 20448 30346 20460
rect 31938 20448 31944 20460
rect 30340 20420 31944 20448
rect 30340 20408 30346 20420
rect 31018 20380 31024 20392
rect 29656 20352 31024 20380
rect 29549 20343 29607 20349
rect 31018 20340 31024 20352
rect 31076 20340 31082 20392
rect 31128 20389 31156 20420
rect 31938 20408 31944 20420
rect 31996 20408 32002 20460
rect 31113 20383 31171 20389
rect 31113 20349 31125 20383
rect 31159 20349 31171 20383
rect 31113 20343 31171 20349
rect 31294 20340 31300 20392
rect 31352 20340 31358 20392
rect 32306 20340 32312 20392
rect 32364 20340 32370 20392
rect 32582 20340 32588 20392
rect 32640 20380 32646 20392
rect 34072 20389 34100 20556
rect 35253 20553 35265 20587
rect 35299 20584 35311 20587
rect 36170 20584 36176 20596
rect 35299 20556 36176 20584
rect 35299 20553 35311 20556
rect 35253 20547 35311 20553
rect 36170 20544 36176 20556
rect 36228 20544 36234 20596
rect 36630 20544 36636 20596
rect 36688 20584 36694 20596
rect 40313 20587 40371 20593
rect 40313 20584 40325 20587
rect 36688 20556 40325 20584
rect 36688 20544 36694 20556
rect 36354 20516 36360 20528
rect 34716 20488 36360 20516
rect 33781 20383 33839 20389
rect 33781 20380 33793 20383
rect 32640 20352 33793 20380
rect 32640 20340 32646 20352
rect 33781 20349 33793 20352
rect 33827 20380 33839 20383
rect 34057 20383 34115 20389
rect 33827 20352 34008 20380
rect 33827 20349 33839 20352
rect 33781 20343 33839 20349
rect 19260 20284 20208 20312
rect 22388 20284 22600 20312
rect 9646 20216 12664 20244
rect 13081 20247 13139 20253
rect 9033 20207 9091 20213
rect 13081 20213 13093 20247
rect 13127 20244 13139 20247
rect 13265 20247 13323 20253
rect 13265 20244 13277 20247
rect 13127 20216 13277 20244
rect 13127 20213 13139 20216
rect 13081 20207 13139 20213
rect 13265 20213 13277 20216
rect 13311 20244 13323 20247
rect 13354 20244 13360 20256
rect 13311 20216 13360 20244
rect 13311 20213 13323 20216
rect 13265 20207 13323 20213
rect 13354 20204 13360 20216
rect 13412 20204 13418 20256
rect 13449 20247 13507 20253
rect 13449 20213 13461 20247
rect 13495 20244 13507 20247
rect 15562 20244 15568 20256
rect 13495 20216 15568 20244
rect 13495 20213 13507 20216
rect 13449 20207 13507 20213
rect 15562 20204 15568 20216
rect 15620 20204 15626 20256
rect 16761 20247 16819 20253
rect 16761 20213 16773 20247
rect 16807 20244 16819 20247
rect 17034 20244 17040 20256
rect 16807 20216 17040 20244
rect 16807 20213 16819 20216
rect 16761 20207 16819 20213
rect 17034 20204 17040 20216
rect 17092 20204 17098 20256
rect 17126 20204 17132 20256
rect 17184 20244 17190 20256
rect 19260 20244 19288 20284
rect 17184 20216 19288 20244
rect 19337 20247 19395 20253
rect 17184 20204 17190 20216
rect 19337 20213 19349 20247
rect 19383 20244 19395 20247
rect 19610 20244 19616 20256
rect 19383 20216 19616 20244
rect 19383 20213 19395 20216
rect 19337 20207 19395 20213
rect 19610 20204 19616 20216
rect 19668 20204 19674 20256
rect 20180 20244 20208 20284
rect 21450 20244 21456 20256
rect 20180 20216 21456 20244
rect 21450 20204 21456 20216
rect 21508 20204 21514 20256
rect 22002 20204 22008 20256
rect 22060 20204 22066 20256
rect 22572 20244 22600 20284
rect 22646 20272 22652 20324
rect 22704 20312 22710 20324
rect 23201 20315 23259 20321
rect 23201 20312 23213 20315
rect 22704 20284 23213 20312
rect 22704 20272 22710 20284
rect 23201 20281 23213 20284
rect 23247 20281 23259 20315
rect 23201 20275 23259 20281
rect 26142 20272 26148 20324
rect 26200 20312 26206 20324
rect 26605 20315 26663 20321
rect 26605 20312 26617 20315
rect 26200 20284 26617 20312
rect 26200 20272 26206 20284
rect 26605 20281 26617 20284
rect 26651 20281 26663 20315
rect 26605 20275 26663 20281
rect 28626 20272 28632 20324
rect 28684 20312 28690 20324
rect 30926 20312 30932 20324
rect 28684 20284 30932 20312
rect 28684 20272 28690 20284
rect 30926 20272 30932 20284
rect 30984 20312 30990 20324
rect 31386 20312 31392 20324
rect 30984 20284 31392 20312
rect 30984 20272 30990 20284
rect 31386 20272 31392 20284
rect 31444 20272 31450 20324
rect 31941 20315 31999 20321
rect 31941 20312 31953 20315
rect 31726 20284 31953 20312
rect 25406 20244 25412 20256
rect 22572 20216 25412 20244
rect 25406 20204 25412 20216
rect 25464 20204 25470 20256
rect 26234 20204 26240 20256
rect 26292 20204 26298 20256
rect 26326 20204 26332 20256
rect 26384 20244 26390 20256
rect 27246 20244 27252 20256
rect 26384 20216 27252 20244
rect 26384 20204 26390 20216
rect 27246 20204 27252 20216
rect 27304 20204 27310 20256
rect 30193 20247 30251 20253
rect 30193 20213 30205 20247
rect 30239 20244 30251 20247
rect 30282 20244 30288 20256
rect 30239 20216 30288 20244
rect 30239 20213 30251 20216
rect 30193 20207 30251 20213
rect 30282 20204 30288 20216
rect 30340 20204 30346 20256
rect 30653 20247 30711 20253
rect 30653 20213 30665 20247
rect 30699 20244 30711 20247
rect 30834 20244 30840 20256
rect 30699 20216 30840 20244
rect 30699 20213 30711 20216
rect 30653 20207 30711 20213
rect 30834 20204 30840 20216
rect 30892 20204 30898 20256
rect 31110 20204 31116 20256
rect 31168 20244 31174 20256
rect 31726 20244 31754 20284
rect 31941 20281 31953 20284
rect 31987 20312 31999 20315
rect 32766 20312 32772 20324
rect 31987 20284 32772 20312
rect 31987 20281 31999 20284
rect 31941 20275 31999 20281
rect 32766 20272 32772 20284
rect 32824 20272 32830 20324
rect 33980 20312 34008 20352
rect 34057 20349 34069 20383
rect 34103 20380 34115 20383
rect 34514 20380 34520 20392
rect 34103 20352 34520 20380
rect 34103 20349 34115 20352
rect 34057 20343 34115 20349
rect 34514 20340 34520 20352
rect 34572 20340 34578 20392
rect 34716 20389 34744 20488
rect 36354 20476 36360 20488
rect 36412 20476 36418 20528
rect 36541 20519 36599 20525
rect 36541 20485 36553 20519
rect 36587 20516 36599 20519
rect 37090 20516 37096 20528
rect 36587 20488 37096 20516
rect 36587 20485 36599 20488
rect 36541 20479 36599 20485
rect 37090 20476 37096 20488
rect 37148 20476 37154 20528
rect 38470 20476 38476 20528
rect 38528 20476 38534 20528
rect 34885 20451 34943 20457
rect 34885 20417 34897 20451
rect 34931 20417 34943 20451
rect 34885 20411 34943 20417
rect 34701 20383 34759 20389
rect 34701 20349 34713 20383
rect 34747 20349 34759 20383
rect 34701 20343 34759 20349
rect 34790 20340 34796 20392
rect 34848 20340 34854 20392
rect 34900 20380 34928 20411
rect 35066 20408 35072 20460
rect 35124 20448 35130 20460
rect 35529 20451 35587 20457
rect 35529 20448 35541 20451
rect 35124 20420 35541 20448
rect 35124 20408 35130 20420
rect 35529 20417 35541 20420
rect 35575 20417 35587 20451
rect 35529 20411 35587 20417
rect 36449 20451 36507 20457
rect 36449 20417 36461 20451
rect 36495 20448 36507 20451
rect 37182 20448 37188 20460
rect 36495 20420 37188 20448
rect 36495 20417 36507 20420
rect 36449 20411 36507 20417
rect 37182 20408 37188 20420
rect 37240 20408 37246 20460
rect 39485 20451 39543 20457
rect 39485 20417 39497 20451
rect 39531 20448 39543 20451
rect 39574 20448 39580 20460
rect 39531 20420 39580 20448
rect 39531 20417 39543 20420
rect 39485 20411 39543 20417
rect 39574 20408 39580 20420
rect 39632 20408 39638 20460
rect 40144 20448 40172 20556
rect 40313 20553 40325 20556
rect 40359 20553 40371 20587
rect 40313 20547 40371 20553
rect 40402 20544 40408 20596
rect 40460 20584 40466 20596
rect 49142 20584 49148 20596
rect 40460 20556 49148 20584
rect 40460 20544 40466 20556
rect 49142 20544 49148 20556
rect 49200 20544 49206 20596
rect 40221 20519 40279 20525
rect 40221 20485 40233 20519
rect 40267 20516 40279 20519
rect 40586 20516 40592 20528
rect 40267 20488 40592 20516
rect 40267 20485 40279 20488
rect 40221 20479 40279 20485
rect 40586 20476 40592 20488
rect 40644 20516 40650 20528
rect 41785 20519 41843 20525
rect 41785 20516 41797 20519
rect 40644 20488 41797 20516
rect 40644 20476 40650 20488
rect 41785 20485 41797 20488
rect 41831 20485 41843 20519
rect 41785 20479 41843 20485
rect 41601 20451 41659 20457
rect 41601 20448 41613 20451
rect 40144 20420 41613 20448
rect 41601 20417 41613 20420
rect 41647 20417 41659 20451
rect 41601 20411 41659 20417
rect 48593 20451 48651 20457
rect 48593 20417 48605 20451
rect 48639 20448 48651 20451
rect 48774 20448 48780 20460
rect 48639 20420 48780 20448
rect 48639 20417 48651 20420
rect 48593 20411 48651 20417
rect 35342 20380 35348 20392
rect 34900 20352 35348 20380
rect 35342 20340 35348 20352
rect 35400 20340 35406 20392
rect 36630 20380 36636 20392
rect 35452 20352 36636 20380
rect 34882 20312 34888 20324
rect 33980 20284 34888 20312
rect 34882 20272 34888 20284
rect 34940 20272 34946 20324
rect 34974 20272 34980 20324
rect 35032 20312 35038 20324
rect 35452 20312 35480 20352
rect 36630 20340 36636 20352
rect 36688 20340 36694 20392
rect 36725 20383 36783 20389
rect 36725 20349 36737 20383
rect 36771 20380 36783 20383
rect 37458 20380 37464 20392
rect 36771 20352 37464 20380
rect 36771 20349 36783 20352
rect 36725 20343 36783 20349
rect 37458 20340 37464 20352
rect 37516 20340 37522 20392
rect 37642 20340 37648 20392
rect 37700 20380 37706 20392
rect 39209 20383 39267 20389
rect 39209 20380 39221 20383
rect 37700 20352 39221 20380
rect 37700 20340 37706 20352
rect 39209 20349 39221 20352
rect 39255 20349 39267 20383
rect 39209 20343 39267 20349
rect 40126 20340 40132 20392
rect 40184 20340 40190 20392
rect 41141 20383 41199 20389
rect 41141 20380 41153 20383
rect 40236 20352 41153 20380
rect 35032 20284 35480 20312
rect 35032 20272 35038 20284
rect 36078 20272 36084 20324
rect 36136 20272 36142 20324
rect 36538 20272 36544 20324
rect 36596 20312 36602 20324
rect 36596 20284 37872 20312
rect 36596 20272 36602 20284
rect 31168 20216 31754 20244
rect 31168 20204 31174 20216
rect 35710 20204 35716 20256
rect 35768 20204 35774 20256
rect 36814 20204 36820 20256
rect 36872 20244 36878 20256
rect 37277 20247 37335 20253
rect 37277 20244 37289 20247
rect 36872 20216 37289 20244
rect 36872 20204 36878 20216
rect 37277 20213 37289 20216
rect 37323 20213 37335 20247
rect 37277 20207 37335 20213
rect 37734 20204 37740 20256
rect 37792 20204 37798 20256
rect 37844 20244 37872 20284
rect 40236 20244 40264 20352
rect 41141 20349 41153 20352
rect 41187 20349 41199 20383
rect 41141 20343 41199 20349
rect 41616 20312 41644 20411
rect 48774 20408 48780 20420
rect 48832 20408 48838 20460
rect 49329 20451 49387 20457
rect 49329 20417 49341 20451
rect 49375 20448 49387 20451
rect 49418 20448 49424 20460
rect 49375 20420 49424 20448
rect 49375 20417 49387 20420
rect 49329 20411 49387 20417
rect 49418 20408 49424 20420
rect 49476 20408 49482 20460
rect 49145 20315 49203 20321
rect 49145 20312 49157 20315
rect 41616 20284 49157 20312
rect 49145 20281 49157 20284
rect 49191 20281 49203 20315
rect 49145 20275 49203 20281
rect 37844 20216 40264 20244
rect 40678 20204 40684 20256
rect 40736 20204 40742 20256
rect 48406 20204 48412 20256
rect 48464 20204 48470 20256
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 4798 20000 4804 20052
rect 4856 20040 4862 20052
rect 11333 20043 11391 20049
rect 11333 20040 11345 20043
rect 4856 20012 11345 20040
rect 4856 20000 4862 20012
rect 11333 20009 11345 20012
rect 11379 20009 11391 20043
rect 11333 20003 11391 20009
rect 11624 20012 11928 20040
rect 9950 19932 9956 19984
rect 10008 19932 10014 19984
rect 10594 19932 10600 19984
rect 10652 19932 10658 19984
rect 4246 19864 4252 19916
rect 4304 19864 4310 19916
rect 5718 19864 5724 19916
rect 5776 19904 5782 19916
rect 5997 19907 6055 19913
rect 5997 19904 6009 19907
rect 5776 19876 6009 19904
rect 5776 19864 5782 19876
rect 5997 19873 6009 19876
rect 6043 19873 6055 19907
rect 11624 19904 11652 20012
rect 11900 19972 11928 20012
rect 11974 20000 11980 20052
rect 12032 20040 12038 20052
rect 12802 20040 12808 20052
rect 12032 20012 12808 20040
rect 12032 20000 12038 20012
rect 12802 20000 12808 20012
rect 12860 20000 12866 20052
rect 14458 20000 14464 20052
rect 14516 20000 14522 20052
rect 16853 20043 16911 20049
rect 16853 20040 16865 20043
rect 14568 20012 16865 20040
rect 14568 19972 14596 20012
rect 16853 20009 16865 20012
rect 16899 20009 16911 20043
rect 16853 20003 16911 20009
rect 16960 20012 19932 20040
rect 11900 19944 12112 19972
rect 5997 19867 6055 19873
rect 10152 19876 11652 19904
rect 2961 19839 3019 19845
rect 2961 19805 2973 19839
rect 3007 19836 3019 19839
rect 3326 19836 3332 19848
rect 3007 19808 3332 19836
rect 3007 19805 3019 19808
rect 2961 19799 3019 19805
rect 3326 19796 3332 19808
rect 3384 19796 3390 19848
rect 5258 19796 5264 19848
rect 5316 19796 5322 19848
rect 7193 19839 7251 19845
rect 7193 19805 7205 19839
rect 7239 19805 7251 19839
rect 7193 19799 7251 19805
rect 7929 19839 7987 19845
rect 7929 19805 7941 19839
rect 7975 19836 7987 19839
rect 9582 19836 9588 19848
rect 7975 19808 9588 19836
rect 7975 19805 7987 19808
rect 7929 19799 7987 19805
rect 1486 19728 1492 19780
rect 1544 19768 1550 19780
rect 1765 19771 1823 19777
rect 1765 19768 1777 19771
rect 1544 19740 1777 19768
rect 1544 19728 1550 19740
rect 1765 19737 1777 19740
rect 1811 19737 1823 19771
rect 1765 19731 1823 19737
rect 7208 19700 7236 19799
rect 9582 19796 9588 19808
rect 9640 19796 9646 19848
rect 10152 19845 10180 19876
rect 11974 19864 11980 19916
rect 12032 19864 12038 19916
rect 12084 19904 12112 19944
rect 13556 19944 14596 19972
rect 13556 19904 13584 19944
rect 14918 19932 14924 19984
rect 14976 19932 14982 19984
rect 15657 19975 15715 19981
rect 15657 19941 15669 19975
rect 15703 19941 15715 19975
rect 15657 19935 15715 19941
rect 12084 19876 13584 19904
rect 13630 19864 13636 19916
rect 13688 19904 13694 19916
rect 15672 19904 15700 19935
rect 13688 19876 15700 19904
rect 13688 19864 13694 19876
rect 16298 19864 16304 19916
rect 16356 19864 16362 19916
rect 10137 19839 10195 19845
rect 10137 19805 10149 19839
rect 10183 19805 10195 19839
rect 10137 19799 10195 19805
rect 10781 19839 10839 19845
rect 10781 19805 10793 19839
rect 10827 19805 10839 19839
rect 10781 19799 10839 19805
rect 7745 19703 7803 19709
rect 7745 19700 7757 19703
rect 7208 19672 7757 19700
rect 7745 19669 7757 19672
rect 7791 19669 7803 19703
rect 10796 19700 10824 19799
rect 10962 19796 10968 19848
rect 11020 19836 11026 19848
rect 11020 19808 11560 19836
rect 11020 19796 11026 19808
rect 11422 19728 11428 19780
rect 11480 19728 11486 19780
rect 11532 19768 11560 19808
rect 13354 19796 13360 19848
rect 13412 19836 13418 19848
rect 14182 19836 14188 19848
rect 13412 19808 14188 19836
rect 13412 19796 13418 19808
rect 14182 19796 14188 19808
rect 14240 19796 14246 19848
rect 14274 19796 14280 19848
rect 14332 19796 14338 19848
rect 15105 19839 15163 19845
rect 15105 19805 15117 19839
rect 15151 19836 15163 19839
rect 15562 19836 15568 19848
rect 15151 19808 15568 19836
rect 15151 19805 15163 19808
rect 15105 19799 15163 19805
rect 15562 19796 15568 19808
rect 15620 19796 15626 19848
rect 16960 19836 16988 20012
rect 18874 19972 18880 19984
rect 17420 19944 18880 19972
rect 17420 19913 17448 19944
rect 18874 19932 18880 19944
rect 18932 19932 18938 19984
rect 19518 19932 19524 19984
rect 19576 19972 19582 19984
rect 19613 19975 19671 19981
rect 19613 19972 19625 19975
rect 19576 19944 19625 19972
rect 19576 19932 19582 19944
rect 19613 19941 19625 19944
rect 19659 19941 19671 19975
rect 19904 19972 19932 20012
rect 19978 20000 19984 20052
rect 20036 20040 20042 20052
rect 22002 20040 22008 20052
rect 20036 20012 22008 20040
rect 20036 20000 20042 20012
rect 22002 20000 22008 20012
rect 22060 20000 22066 20052
rect 22462 20000 22468 20052
rect 22520 20040 22526 20052
rect 25593 20043 25651 20049
rect 25593 20040 25605 20043
rect 22520 20012 25605 20040
rect 22520 20000 22526 20012
rect 25593 20009 25605 20012
rect 25639 20009 25651 20043
rect 25593 20003 25651 20009
rect 26786 20000 26792 20052
rect 26844 20000 26850 20052
rect 27062 20000 27068 20052
rect 27120 20040 27126 20052
rect 29089 20043 29147 20049
rect 29089 20040 29101 20043
rect 27120 20012 29101 20040
rect 27120 20000 27126 20012
rect 29089 20009 29101 20012
rect 29135 20040 29147 20043
rect 34974 20040 34980 20052
rect 29135 20012 34980 20040
rect 29135 20009 29147 20012
rect 29089 20003 29147 20009
rect 34974 20000 34980 20012
rect 35032 20000 35038 20052
rect 35434 20000 35440 20052
rect 35492 20040 35498 20052
rect 36998 20040 37004 20052
rect 35492 20012 37004 20040
rect 35492 20000 35498 20012
rect 36998 20000 37004 20012
rect 37056 20040 37062 20052
rect 38378 20040 38384 20052
rect 37056 20012 38384 20040
rect 37056 20000 37062 20012
rect 38378 20000 38384 20012
rect 38436 20000 38442 20052
rect 38838 20000 38844 20052
rect 38896 20040 38902 20052
rect 38896 20012 40356 20040
rect 38896 20000 38902 20012
rect 22925 19975 22983 19981
rect 22925 19972 22937 19975
rect 19904 19944 21036 19972
rect 19613 19935 19671 19941
rect 17405 19907 17463 19913
rect 17405 19873 17417 19907
rect 17451 19873 17463 19907
rect 18785 19907 18843 19913
rect 17405 19867 17463 19873
rect 18524 19876 18736 19904
rect 15672 19808 16988 19836
rect 17313 19839 17371 19845
rect 12253 19771 12311 19777
rect 12253 19768 12265 19771
rect 11532 19740 12265 19768
rect 12253 19737 12265 19740
rect 12299 19737 12311 19771
rect 12253 19731 12311 19737
rect 13814 19728 13820 19780
rect 13872 19768 13878 19780
rect 15672 19768 15700 19808
rect 17313 19805 17325 19839
rect 17359 19836 17371 19839
rect 18524 19836 18552 19876
rect 17359 19808 18552 19836
rect 18708 19836 18736 19876
rect 18785 19873 18797 19907
rect 18831 19904 18843 19907
rect 19886 19904 19892 19916
rect 18831 19876 19892 19904
rect 18831 19873 18843 19876
rect 18785 19867 18843 19873
rect 19886 19864 19892 19876
rect 19944 19864 19950 19916
rect 21008 19904 21036 19944
rect 22204 19944 22937 19972
rect 22204 19904 22232 19944
rect 22925 19941 22937 19944
rect 22971 19972 22983 19975
rect 23934 19972 23940 19984
rect 22971 19944 23940 19972
rect 22971 19941 22983 19944
rect 22925 19935 22983 19941
rect 21008 19876 22232 19904
rect 22281 19907 22339 19913
rect 22281 19873 22293 19907
rect 22327 19873 22339 19907
rect 22830 19904 22836 19916
rect 22281 19867 22339 19873
rect 22664 19876 22836 19904
rect 19518 19836 19524 19848
rect 18708 19808 19524 19836
rect 17359 19805 17371 19808
rect 17313 19799 17371 19805
rect 19518 19796 19524 19808
rect 19576 19796 19582 19848
rect 20530 19836 20536 19848
rect 19720 19808 20536 19836
rect 13872 19740 15700 19768
rect 16025 19771 16083 19777
rect 13872 19728 13878 19740
rect 16025 19737 16037 19771
rect 16071 19768 16083 19771
rect 17862 19768 17868 19780
rect 16071 19740 17868 19768
rect 16071 19737 16083 19740
rect 16025 19731 16083 19737
rect 17862 19728 17868 19740
rect 17920 19728 17926 19780
rect 19720 19768 19748 19808
rect 20530 19796 20536 19808
rect 20588 19796 20594 19848
rect 22296 19836 22324 19867
rect 22664 19836 22692 19876
rect 22830 19864 22836 19876
rect 22888 19864 22894 19916
rect 23382 19864 23388 19916
rect 23440 19864 23446 19916
rect 23584 19913 23612 19944
rect 23934 19932 23940 19944
rect 23992 19932 23998 19984
rect 24029 19975 24087 19981
rect 24029 19941 24041 19975
rect 24075 19972 24087 19975
rect 27614 19972 27620 19984
rect 24075 19944 27620 19972
rect 24075 19941 24087 19944
rect 24029 19935 24087 19941
rect 27614 19932 27620 19944
rect 27672 19932 27678 19984
rect 27982 19932 27988 19984
rect 28040 19972 28046 19984
rect 29822 19972 29828 19984
rect 28040 19944 29828 19972
rect 28040 19932 28046 19944
rect 29822 19932 29828 19944
rect 29880 19932 29886 19984
rect 29932 19944 32720 19972
rect 23569 19907 23627 19913
rect 23569 19873 23581 19907
rect 23615 19873 23627 19907
rect 23569 19867 23627 19873
rect 24578 19864 24584 19916
rect 24636 19864 24642 19916
rect 25038 19864 25044 19916
rect 25096 19904 25102 19916
rect 25317 19907 25375 19913
rect 25317 19904 25329 19907
rect 25096 19876 25329 19904
rect 25096 19864 25102 19876
rect 25317 19873 25329 19876
rect 25363 19873 25375 19907
rect 25317 19867 25375 19873
rect 26145 19907 26203 19913
rect 26145 19873 26157 19907
rect 26191 19873 26203 19907
rect 26145 19867 26203 19873
rect 22296 19808 22692 19836
rect 22738 19796 22744 19848
rect 22796 19836 22802 19848
rect 25222 19836 25228 19848
rect 22796 19808 25228 19836
rect 22796 19796 22802 19808
rect 25222 19796 25228 19808
rect 25280 19836 25286 19848
rect 26160 19836 26188 19867
rect 26970 19864 26976 19916
rect 27028 19904 27034 19916
rect 27341 19907 27399 19913
rect 27341 19904 27353 19907
rect 27028 19876 27353 19904
rect 27028 19864 27034 19876
rect 27341 19873 27353 19876
rect 27387 19873 27399 19907
rect 27341 19867 27399 19873
rect 28350 19864 28356 19916
rect 28408 19904 28414 19916
rect 28537 19907 28595 19913
rect 28537 19904 28549 19907
rect 28408 19876 28549 19904
rect 28408 19864 28414 19876
rect 28537 19873 28549 19876
rect 28583 19873 28595 19907
rect 28537 19867 28595 19873
rect 28994 19864 29000 19916
rect 29052 19904 29058 19916
rect 29932 19904 29960 19944
rect 29052 19876 29960 19904
rect 30377 19907 30435 19913
rect 29052 19864 29058 19876
rect 30377 19873 30389 19907
rect 30423 19904 30435 19907
rect 30576 19904 30604 19944
rect 32692 19913 32720 19944
rect 33318 19932 33324 19984
rect 33376 19972 33382 19984
rect 36081 19975 36139 19981
rect 36081 19972 36093 19975
rect 33376 19944 36093 19972
rect 33376 19932 33382 19944
rect 36081 19941 36093 19944
rect 36127 19941 36139 19975
rect 36081 19935 36139 19941
rect 36372 19944 38148 19972
rect 30423 19876 30604 19904
rect 31113 19907 31171 19913
rect 30423 19873 30435 19876
rect 30377 19867 30435 19873
rect 31113 19873 31125 19907
rect 31159 19904 31171 19907
rect 32677 19907 32735 19913
rect 31159 19876 32451 19904
rect 31159 19873 31171 19876
rect 31113 19867 31171 19873
rect 25280 19808 26188 19836
rect 25280 19796 25286 19808
rect 27246 19796 27252 19848
rect 27304 19836 27310 19848
rect 30190 19836 30196 19848
rect 27304 19808 30196 19836
rect 27304 19796 27310 19808
rect 30190 19796 30196 19808
rect 30248 19796 30254 19848
rect 30558 19796 30564 19848
rect 30616 19836 30622 19848
rect 31294 19836 31300 19848
rect 30616 19808 31300 19836
rect 30616 19796 30622 19808
rect 31294 19796 31300 19808
rect 31352 19796 31358 19848
rect 18616 19740 19748 19768
rect 19797 19771 19855 19777
rect 13630 19700 13636 19712
rect 10796 19672 13636 19700
rect 7745 19663 7803 19669
rect 13630 19660 13636 19672
rect 13688 19660 13694 19712
rect 13725 19703 13783 19709
rect 13725 19669 13737 19703
rect 13771 19700 13783 19703
rect 15930 19700 15936 19712
rect 13771 19672 15936 19700
rect 13771 19669 13783 19672
rect 13725 19663 13783 19669
rect 15930 19660 15936 19672
rect 15988 19660 15994 19712
rect 16117 19703 16175 19709
rect 16117 19669 16129 19703
rect 16163 19700 16175 19703
rect 17126 19700 17132 19712
rect 16163 19672 17132 19700
rect 16163 19669 16175 19672
rect 16117 19663 16175 19669
rect 17126 19660 17132 19672
rect 17184 19660 17190 19712
rect 17218 19660 17224 19712
rect 17276 19660 17282 19712
rect 18141 19703 18199 19709
rect 18141 19669 18153 19703
rect 18187 19700 18199 19703
rect 18322 19700 18328 19712
rect 18187 19672 18328 19700
rect 18187 19669 18199 19672
rect 18141 19663 18199 19669
rect 18322 19660 18328 19672
rect 18380 19660 18386 19712
rect 18414 19660 18420 19712
rect 18472 19700 18478 19712
rect 18616 19709 18644 19740
rect 19797 19737 19809 19771
rect 19843 19768 19855 19771
rect 20346 19768 20352 19780
rect 19843 19740 20352 19768
rect 19843 19737 19855 19740
rect 19797 19731 19855 19737
rect 20346 19728 20352 19740
rect 20404 19728 20410 19780
rect 21542 19728 21548 19780
rect 21600 19728 21606 19780
rect 22005 19771 22063 19777
rect 22005 19737 22017 19771
rect 22051 19768 22063 19771
rect 22094 19768 22100 19780
rect 22051 19740 22100 19768
rect 22051 19737 22063 19740
rect 22005 19731 22063 19737
rect 22094 19728 22100 19740
rect 22152 19728 22158 19780
rect 25961 19771 26019 19777
rect 25961 19737 25973 19771
rect 26007 19768 26019 19771
rect 26694 19768 26700 19780
rect 26007 19740 26700 19768
rect 26007 19737 26019 19740
rect 25961 19731 26019 19737
rect 26694 19728 26700 19740
rect 26752 19728 26758 19780
rect 28445 19771 28503 19777
rect 28445 19737 28457 19771
rect 28491 19768 28503 19771
rect 30006 19768 30012 19780
rect 28491 19740 30012 19768
rect 28491 19737 28503 19740
rect 28445 19731 28503 19737
rect 30006 19728 30012 19740
rect 30064 19728 30070 19780
rect 30098 19728 30104 19780
rect 30156 19728 30162 19780
rect 32214 19768 32220 19780
rect 31680 19740 32220 19768
rect 18509 19703 18567 19709
rect 18509 19700 18521 19703
rect 18472 19672 18521 19700
rect 18472 19660 18478 19672
rect 18509 19669 18521 19672
rect 18555 19669 18567 19703
rect 18509 19663 18567 19669
rect 18601 19703 18659 19709
rect 18601 19669 18613 19703
rect 18647 19669 18659 19703
rect 18601 19663 18659 19669
rect 19334 19660 19340 19712
rect 19392 19660 19398 19712
rect 20254 19660 20260 19712
rect 20312 19660 20318 19712
rect 20438 19660 20444 19712
rect 20496 19700 20502 19712
rect 20533 19703 20591 19709
rect 20533 19700 20545 19703
rect 20496 19672 20545 19700
rect 20496 19660 20502 19672
rect 20533 19669 20545 19672
rect 20579 19669 20591 19703
rect 20533 19663 20591 19669
rect 22646 19660 22652 19712
rect 22704 19660 22710 19712
rect 22833 19703 22891 19709
rect 22833 19669 22845 19703
rect 22879 19700 22891 19703
rect 23382 19700 23388 19712
rect 22879 19672 23388 19700
rect 22879 19669 22891 19672
rect 22833 19663 22891 19669
rect 23382 19660 23388 19672
rect 23440 19660 23446 19712
rect 23474 19660 23480 19712
rect 23532 19700 23538 19712
rect 23661 19703 23719 19709
rect 23661 19700 23673 19703
rect 23532 19672 23673 19700
rect 23532 19660 23538 19672
rect 23661 19669 23673 19672
rect 23707 19669 23719 19703
rect 23661 19663 23719 19669
rect 25133 19703 25191 19709
rect 25133 19669 25145 19703
rect 25179 19700 25191 19703
rect 26053 19703 26111 19709
rect 26053 19700 26065 19703
rect 25179 19672 26065 19700
rect 25179 19669 25191 19672
rect 25133 19663 25191 19669
rect 26053 19669 26065 19672
rect 26099 19700 26111 19703
rect 26326 19700 26332 19712
rect 26099 19672 26332 19700
rect 26099 19669 26111 19672
rect 26053 19663 26111 19669
rect 26326 19660 26332 19672
rect 26384 19660 26390 19712
rect 27062 19660 27068 19712
rect 27120 19700 27126 19712
rect 27157 19703 27215 19709
rect 27157 19700 27169 19703
rect 27120 19672 27169 19700
rect 27120 19660 27126 19672
rect 27157 19669 27169 19672
rect 27203 19669 27215 19703
rect 27157 19663 27215 19669
rect 27246 19660 27252 19712
rect 27304 19660 27310 19712
rect 27614 19660 27620 19712
rect 27672 19700 27678 19712
rect 27985 19703 28043 19709
rect 27985 19700 27997 19703
rect 27672 19672 27997 19700
rect 27672 19660 27678 19672
rect 27985 19669 27997 19672
rect 28031 19669 28043 19703
rect 27985 19663 28043 19669
rect 28353 19703 28411 19709
rect 28353 19669 28365 19703
rect 28399 19700 28411 19703
rect 28626 19700 28632 19712
rect 28399 19672 28632 19700
rect 28399 19669 28411 19672
rect 28353 19663 28411 19669
rect 28626 19660 28632 19672
rect 28684 19660 28690 19712
rect 28902 19660 28908 19712
rect 28960 19700 28966 19712
rect 29273 19703 29331 19709
rect 29273 19700 29285 19703
rect 28960 19672 29285 19700
rect 28960 19660 28966 19672
rect 29273 19669 29285 19672
rect 29319 19669 29331 19703
rect 29273 19663 29331 19669
rect 29730 19660 29736 19712
rect 29788 19660 29794 19712
rect 30116 19700 30144 19728
rect 30926 19700 30932 19712
rect 30116 19672 30932 19700
rect 30926 19660 30932 19672
rect 30984 19660 30990 19712
rect 31110 19660 31116 19712
rect 31168 19700 31174 19712
rect 31205 19703 31263 19709
rect 31205 19700 31217 19703
rect 31168 19672 31217 19700
rect 31168 19660 31174 19672
rect 31205 19669 31217 19672
rect 31251 19669 31263 19703
rect 31205 19663 31263 19669
rect 31297 19703 31355 19709
rect 31297 19669 31309 19703
rect 31343 19700 31355 19703
rect 31570 19700 31576 19712
rect 31343 19672 31576 19700
rect 31343 19669 31355 19672
rect 31297 19663 31355 19669
rect 31570 19660 31576 19672
rect 31628 19660 31634 19712
rect 31680 19709 31708 19740
rect 32214 19728 32220 19740
rect 32272 19728 32278 19780
rect 31665 19703 31723 19709
rect 31665 19669 31677 19703
rect 31711 19669 31723 19703
rect 31665 19663 31723 19669
rect 32122 19660 32128 19712
rect 32180 19660 32186 19712
rect 32423 19700 32451 19876
rect 32677 19873 32689 19907
rect 32723 19873 32735 19907
rect 32677 19867 32735 19873
rect 33597 19907 33655 19913
rect 33597 19873 33609 19907
rect 33643 19904 33655 19907
rect 34054 19904 34060 19916
rect 33643 19876 34060 19904
rect 33643 19873 33655 19876
rect 33597 19867 33655 19873
rect 34054 19864 34060 19876
rect 34112 19904 34118 19916
rect 34425 19907 34483 19913
rect 34425 19904 34437 19907
rect 34112 19876 34437 19904
rect 34112 19864 34118 19876
rect 34425 19873 34437 19876
rect 34471 19873 34483 19907
rect 34425 19867 34483 19873
rect 35066 19864 35072 19916
rect 35124 19904 35130 19916
rect 35710 19904 35716 19916
rect 35124 19876 35716 19904
rect 35124 19864 35130 19876
rect 35710 19864 35716 19876
rect 35768 19864 35774 19916
rect 35802 19864 35808 19916
rect 35860 19904 35866 19916
rect 36372 19904 36400 19944
rect 35860 19876 36400 19904
rect 35860 19864 35866 19876
rect 36446 19864 36452 19916
rect 36504 19904 36510 19916
rect 36633 19907 36691 19913
rect 36633 19904 36645 19907
rect 36504 19876 36645 19904
rect 36504 19864 36510 19876
rect 36633 19873 36645 19876
rect 36679 19873 36691 19907
rect 36633 19867 36691 19873
rect 37642 19864 37648 19916
rect 37700 19904 37706 19916
rect 38120 19913 38148 19944
rect 38470 19932 38476 19984
rect 38528 19972 38534 19984
rect 39577 19975 39635 19981
rect 39577 19972 39589 19975
rect 38528 19944 39589 19972
rect 38528 19932 38534 19944
rect 39577 19941 39589 19944
rect 39623 19941 39635 19975
rect 39577 19935 39635 19941
rect 37921 19907 37979 19913
rect 37921 19904 37933 19907
rect 37700 19876 37933 19904
rect 37700 19864 37706 19876
rect 37921 19873 37933 19876
rect 37967 19873 37979 19907
rect 37921 19867 37979 19873
rect 38105 19907 38163 19913
rect 38105 19873 38117 19907
rect 38151 19904 38163 19907
rect 39025 19907 39083 19913
rect 39025 19904 39037 19907
rect 38151 19876 39037 19904
rect 38151 19873 38163 19876
rect 38105 19867 38163 19873
rect 39025 19873 39037 19876
rect 39071 19904 39083 19907
rect 39206 19904 39212 19916
rect 39071 19876 39212 19904
rect 39071 19873 39083 19876
rect 39025 19867 39083 19873
rect 39206 19864 39212 19876
rect 39264 19864 39270 19916
rect 39390 19864 39396 19916
rect 39448 19904 39454 19916
rect 40328 19913 40356 20012
rect 41046 20000 41052 20052
rect 41104 20000 41110 20052
rect 48774 20000 48780 20052
rect 48832 20000 48838 20052
rect 40954 19932 40960 19984
rect 41012 19972 41018 19984
rect 41233 19975 41291 19981
rect 41233 19972 41245 19975
rect 41012 19944 41245 19972
rect 41012 19932 41018 19944
rect 41233 19941 41245 19944
rect 41279 19941 41291 19975
rect 41233 19935 41291 19941
rect 40129 19907 40187 19913
rect 40129 19904 40141 19907
rect 39448 19876 40141 19904
rect 39448 19864 39454 19876
rect 40129 19873 40141 19876
rect 40175 19873 40187 19907
rect 40129 19867 40187 19873
rect 40313 19907 40371 19913
rect 40313 19873 40325 19907
rect 40359 19904 40371 19907
rect 40972 19904 41000 19932
rect 40359 19876 41000 19904
rect 40359 19873 40371 19876
rect 40313 19867 40371 19873
rect 32493 19839 32551 19845
rect 32493 19805 32505 19839
rect 32539 19836 32551 19839
rect 33778 19836 33784 19848
rect 32539 19808 33784 19836
rect 32539 19805 32551 19808
rect 32493 19799 32551 19805
rect 33778 19796 33784 19808
rect 33836 19796 33842 19848
rect 34146 19796 34152 19848
rect 34204 19836 34210 19848
rect 35161 19839 35219 19845
rect 35161 19836 35173 19839
rect 34204 19808 35173 19836
rect 34204 19796 34210 19808
rect 35161 19805 35173 19808
rect 35207 19805 35219 19839
rect 35161 19799 35219 19805
rect 35253 19839 35311 19845
rect 35253 19805 35265 19839
rect 35299 19836 35311 19839
rect 35526 19836 35532 19848
rect 35299 19808 35532 19836
rect 35299 19805 35311 19808
rect 35253 19799 35311 19805
rect 35526 19796 35532 19808
rect 35584 19796 35590 19848
rect 37366 19796 37372 19848
rect 37424 19836 37430 19848
rect 38197 19839 38255 19845
rect 38197 19836 38209 19839
rect 37424 19808 38209 19836
rect 37424 19796 37430 19808
rect 38197 19805 38209 19808
rect 38243 19836 38255 19839
rect 38841 19839 38899 19845
rect 38841 19836 38853 19839
rect 38243 19808 38853 19836
rect 38243 19805 38255 19808
rect 38197 19799 38255 19805
rect 38841 19805 38853 19808
rect 38887 19836 38899 19839
rect 40862 19836 40868 19848
rect 38887 19808 40868 19836
rect 38887 19805 38899 19808
rect 38841 19799 38899 19805
rect 40862 19796 40868 19808
rect 40920 19796 40926 19848
rect 32585 19771 32643 19777
rect 32585 19737 32597 19771
rect 32631 19768 32643 19771
rect 33689 19771 33747 19777
rect 33689 19768 33701 19771
rect 32631 19740 33701 19768
rect 32631 19737 32643 19740
rect 32585 19731 32643 19737
rect 33689 19737 33701 19740
rect 33735 19768 33747 19771
rect 34882 19768 34888 19780
rect 33735 19740 34888 19768
rect 33735 19737 33747 19740
rect 33689 19731 33747 19737
rect 34882 19728 34888 19740
rect 34940 19728 34946 19780
rect 34974 19728 34980 19780
rect 35032 19768 35038 19780
rect 36262 19768 36268 19780
rect 35032 19740 36268 19768
rect 35032 19728 35038 19740
rect 36262 19728 36268 19740
rect 36320 19728 36326 19780
rect 36449 19771 36507 19777
rect 36449 19737 36461 19771
rect 36495 19768 36507 19771
rect 40034 19768 40040 19780
rect 36495 19740 40040 19768
rect 36495 19737 36507 19740
rect 36449 19731 36507 19737
rect 40034 19728 40040 19740
rect 40092 19728 40098 19780
rect 40405 19771 40463 19777
rect 40405 19737 40417 19771
rect 40451 19768 40463 19771
rect 41046 19768 41052 19780
rect 40451 19740 41052 19768
rect 40451 19737 40463 19740
rect 40405 19731 40463 19737
rect 41046 19728 41052 19740
rect 41104 19728 41110 19780
rect 48593 19771 48651 19777
rect 48593 19737 48605 19771
rect 48639 19768 48651 19771
rect 49237 19771 49295 19777
rect 49237 19768 49249 19771
rect 48639 19740 49249 19768
rect 48639 19737 48651 19740
rect 48593 19731 48651 19737
rect 49237 19737 49249 19740
rect 49283 19768 49295 19771
rect 49326 19768 49332 19780
rect 49283 19740 49332 19768
rect 49283 19737 49295 19740
rect 49237 19731 49295 19737
rect 49326 19728 49332 19740
rect 49384 19728 49390 19780
rect 33410 19700 33416 19712
rect 32423 19672 33416 19700
rect 33410 19660 33416 19672
rect 33468 19660 33474 19712
rect 34146 19660 34152 19712
rect 34204 19660 34210 19712
rect 35621 19703 35679 19709
rect 35621 19669 35633 19703
rect 35667 19700 35679 19703
rect 35986 19700 35992 19712
rect 35667 19672 35992 19700
rect 35667 19669 35679 19672
rect 35621 19663 35679 19669
rect 35986 19660 35992 19672
rect 36044 19660 36050 19712
rect 36538 19660 36544 19712
rect 36596 19660 36602 19712
rect 37369 19703 37427 19709
rect 37369 19669 37381 19703
rect 37415 19700 37427 19703
rect 37550 19700 37556 19712
rect 37415 19672 37556 19700
rect 37415 19669 37427 19672
rect 37369 19663 37427 19669
rect 37550 19660 37556 19672
rect 37608 19660 37614 19712
rect 38378 19660 38384 19712
rect 38436 19700 38442 19712
rect 38565 19703 38623 19709
rect 38565 19700 38577 19703
rect 38436 19672 38577 19700
rect 38436 19660 38442 19672
rect 38565 19669 38577 19672
rect 38611 19669 38623 19703
rect 38565 19663 38623 19669
rect 40770 19660 40776 19712
rect 40828 19660 40834 19712
rect 49142 19660 49148 19712
rect 49200 19660 49206 19712
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 7834 19456 7840 19508
rect 7892 19496 7898 19508
rect 10965 19499 11023 19505
rect 10965 19496 10977 19499
rect 7892 19468 10977 19496
rect 7892 19456 7898 19468
rect 10965 19465 10977 19468
rect 11011 19465 11023 19499
rect 10965 19459 11023 19465
rect 13446 19456 13452 19508
rect 13504 19496 13510 19508
rect 13504 19468 14504 19496
rect 13504 19456 13510 19468
rect 3418 19388 3424 19440
rect 3476 19428 3482 19440
rect 3605 19431 3663 19437
rect 3605 19428 3617 19431
rect 3476 19400 3617 19428
rect 3476 19388 3482 19400
rect 3605 19397 3617 19400
rect 3651 19397 3663 19431
rect 9214 19428 9220 19440
rect 3605 19391 3663 19397
rect 4540 19400 9220 19428
rect 1762 19320 1768 19372
rect 1820 19320 1826 19372
rect 2961 19363 3019 19369
rect 2961 19329 2973 19363
rect 3007 19360 3019 19363
rect 4540 19360 4568 19400
rect 9214 19388 9220 19400
rect 9272 19388 9278 19440
rect 10505 19431 10563 19437
rect 10505 19397 10517 19431
rect 10551 19428 10563 19431
rect 12802 19428 12808 19440
rect 10551 19400 12808 19428
rect 10551 19397 10563 19400
rect 10505 19391 10563 19397
rect 12802 19388 12808 19400
rect 12860 19388 12866 19440
rect 14182 19428 14188 19440
rect 13754 19400 14188 19428
rect 14182 19388 14188 19400
rect 14240 19388 14246 19440
rect 3007 19332 4568 19360
rect 4801 19363 4859 19369
rect 3007 19329 3019 19332
rect 2961 19323 3019 19329
rect 4801 19329 4813 19363
rect 4847 19360 4859 19363
rect 5445 19363 5503 19369
rect 4847 19332 5396 19360
rect 4847 19329 4859 19332
rect 4801 19323 4859 19329
rect 3878 19252 3884 19304
rect 3936 19292 3942 19304
rect 5261 19295 5319 19301
rect 5261 19292 5273 19295
rect 3936 19264 5273 19292
rect 3936 19252 3942 19264
rect 5261 19261 5273 19264
rect 5307 19261 5319 19295
rect 5368 19292 5396 19332
rect 5445 19329 5457 19363
rect 5491 19360 5503 19363
rect 5902 19360 5908 19372
rect 5491 19332 5908 19360
rect 5491 19329 5503 19332
rect 5445 19323 5503 19329
rect 5902 19320 5908 19332
rect 5960 19320 5966 19372
rect 9122 19320 9128 19372
rect 9180 19360 9186 19372
rect 9180 19332 11100 19360
rect 9180 19320 9186 19332
rect 6822 19292 6828 19304
rect 5368 19264 6828 19292
rect 5261 19255 5319 19261
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 9858 19252 9864 19304
rect 9916 19252 9922 19304
rect 11072 19292 11100 19332
rect 11146 19320 11152 19372
rect 11204 19320 11210 19372
rect 11701 19363 11759 19369
rect 11701 19329 11713 19363
rect 11747 19360 11759 19363
rect 12158 19360 12164 19372
rect 11747 19332 12164 19360
rect 11747 19329 11759 19332
rect 11701 19323 11759 19329
rect 12158 19320 12164 19332
rect 12216 19320 12222 19372
rect 14476 19369 14504 19468
rect 15010 19456 15016 19508
rect 15068 19496 15074 19508
rect 16853 19499 16911 19505
rect 16853 19496 16865 19499
rect 15068 19468 16865 19496
rect 15068 19456 15074 19468
rect 16853 19465 16865 19468
rect 16899 19465 16911 19499
rect 16853 19459 16911 19465
rect 17313 19499 17371 19505
rect 17313 19465 17325 19499
rect 17359 19496 17371 19499
rect 19426 19496 19432 19508
rect 17359 19468 19432 19496
rect 17359 19465 17371 19468
rect 17313 19459 17371 19465
rect 19426 19456 19432 19468
rect 19484 19456 19490 19508
rect 20717 19499 20775 19505
rect 20717 19465 20729 19499
rect 20763 19496 20775 19499
rect 20806 19496 20812 19508
rect 20763 19468 20812 19496
rect 20763 19465 20775 19468
rect 20717 19459 20775 19465
rect 20806 19456 20812 19468
rect 20864 19456 20870 19508
rect 21177 19499 21235 19505
rect 21177 19465 21189 19499
rect 21223 19496 21235 19499
rect 21266 19496 21272 19508
rect 21223 19468 21272 19496
rect 21223 19465 21235 19468
rect 21177 19459 21235 19465
rect 21266 19456 21272 19468
rect 21324 19456 21330 19508
rect 23474 19496 23480 19508
rect 22572 19468 23480 19496
rect 14921 19431 14979 19437
rect 14921 19397 14933 19431
rect 14967 19428 14979 19431
rect 16206 19428 16212 19440
rect 14967 19400 16212 19428
rect 14967 19397 14979 19400
rect 14921 19391 14979 19397
rect 16206 19388 16212 19400
rect 16264 19388 16270 19440
rect 19058 19388 19064 19440
rect 19116 19388 19122 19440
rect 20254 19388 20260 19440
rect 20312 19428 20318 19440
rect 22572 19428 22600 19468
rect 23474 19456 23480 19468
rect 23532 19456 23538 19508
rect 23676 19468 26096 19496
rect 20312 19400 22600 19428
rect 20312 19388 20318 19400
rect 22646 19388 22652 19440
rect 22704 19428 22710 19440
rect 22925 19431 22983 19437
rect 22925 19428 22937 19431
rect 22704 19400 22937 19428
rect 22704 19388 22710 19400
rect 22925 19397 22937 19400
rect 22971 19397 22983 19431
rect 22925 19391 22983 19397
rect 23382 19388 23388 19440
rect 23440 19428 23446 19440
rect 23676 19428 23704 19468
rect 23440 19400 23704 19428
rect 23440 19388 23446 19400
rect 24486 19388 24492 19440
rect 24544 19388 24550 19440
rect 24854 19388 24860 19440
rect 24912 19428 24918 19440
rect 24912 19400 25820 19428
rect 24912 19388 24918 19400
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19360 14519 19363
rect 15378 19360 15384 19372
rect 14507 19332 15384 19360
rect 14507 19329 14519 19332
rect 14461 19323 14519 19329
rect 15378 19320 15384 19332
rect 15436 19320 15442 19372
rect 15470 19320 15476 19372
rect 15528 19320 15534 19372
rect 17034 19320 17040 19372
rect 17092 19360 17098 19372
rect 17221 19363 17279 19369
rect 17221 19360 17233 19363
rect 17092 19332 17233 19360
rect 17092 19320 17098 19332
rect 17221 19329 17233 19332
rect 17267 19329 17279 19363
rect 17221 19323 17279 19329
rect 18049 19363 18107 19369
rect 18049 19329 18061 19363
rect 18095 19360 18107 19363
rect 18414 19360 18420 19372
rect 18095 19332 18420 19360
rect 18095 19329 18107 19332
rect 18049 19323 18107 19329
rect 18414 19320 18420 19332
rect 18472 19320 18478 19372
rect 21085 19363 21143 19369
rect 21085 19329 21097 19363
rect 21131 19360 21143 19363
rect 21131 19332 22140 19360
rect 21131 19329 21143 19332
rect 21085 19323 21143 19329
rect 11977 19295 12035 19301
rect 11977 19292 11989 19295
rect 11072 19264 11989 19292
rect 11977 19261 11989 19264
rect 12023 19261 12035 19295
rect 12710 19292 12716 19304
rect 11977 19255 12035 19261
rect 12452 19264 12716 19292
rect 7558 19184 7564 19236
rect 7616 19224 7622 19236
rect 12066 19224 12072 19236
rect 7616 19196 12072 19224
rect 7616 19184 7622 19196
rect 12066 19184 12072 19196
rect 12124 19184 12130 19236
rect 12452 19168 12480 19264
rect 12710 19252 12716 19264
rect 12768 19252 12774 19304
rect 14185 19295 14243 19301
rect 14185 19261 14197 19295
rect 14231 19292 14243 19295
rect 15194 19292 15200 19304
rect 14231 19264 15200 19292
rect 14231 19261 14243 19264
rect 14185 19255 14243 19261
rect 15194 19252 15200 19264
rect 15252 19252 15258 19304
rect 15289 19295 15347 19301
rect 15289 19261 15301 19295
rect 15335 19292 15347 19295
rect 15746 19292 15752 19304
rect 15335 19264 15752 19292
rect 15335 19261 15347 19264
rect 15289 19255 15347 19261
rect 15746 19252 15752 19264
rect 15804 19252 15810 19304
rect 16022 19252 16028 19304
rect 16080 19252 16086 19304
rect 16114 19252 16120 19304
rect 16172 19292 16178 19304
rect 17405 19295 17463 19301
rect 17405 19292 17417 19295
rect 16172 19264 17417 19292
rect 16172 19252 16178 19264
rect 17405 19261 17417 19264
rect 17451 19261 17463 19295
rect 19426 19292 19432 19304
rect 17405 19255 17463 19261
rect 18800 19264 19432 19292
rect 14829 19227 14887 19233
rect 14829 19193 14841 19227
rect 14875 19224 14887 19227
rect 15470 19224 15476 19236
rect 14875 19196 15476 19224
rect 14875 19193 14887 19196
rect 14829 19187 14887 19193
rect 15470 19184 15476 19196
rect 15528 19184 15534 19236
rect 18800 19224 18828 19264
rect 19426 19252 19432 19264
rect 19484 19252 19490 19304
rect 19794 19252 19800 19304
rect 19852 19252 19858 19304
rect 20073 19295 20131 19301
rect 20073 19292 20085 19295
rect 19996 19264 20085 19292
rect 16408 19196 18828 19224
rect 5902 19116 5908 19168
rect 5960 19116 5966 19168
rect 8294 19116 8300 19168
rect 8352 19156 8358 19168
rect 11882 19156 11888 19168
rect 8352 19128 11888 19156
rect 8352 19116 8358 19128
rect 11882 19116 11888 19128
rect 11940 19116 11946 19168
rect 12434 19116 12440 19168
rect 12492 19116 12498 19168
rect 12710 19116 12716 19168
rect 12768 19116 12774 19168
rect 15102 19116 15108 19168
rect 15160 19156 15166 19168
rect 16408 19156 16436 19196
rect 15160 19128 16436 19156
rect 15160 19116 15166 19128
rect 16482 19116 16488 19168
rect 16540 19156 16546 19168
rect 19058 19156 19064 19168
rect 16540 19128 19064 19156
rect 16540 19116 16546 19128
rect 19058 19116 19064 19128
rect 19116 19116 19122 19168
rect 19610 19116 19616 19168
rect 19668 19156 19674 19168
rect 19996 19156 20024 19264
rect 20073 19261 20085 19264
rect 20119 19261 20131 19295
rect 20073 19255 20131 19261
rect 21361 19295 21419 19301
rect 21361 19261 21373 19295
rect 21407 19261 21419 19295
rect 22112 19292 22140 19332
rect 22186 19320 22192 19372
rect 22244 19320 22250 19372
rect 25225 19363 25283 19369
rect 25225 19329 25237 19363
rect 25271 19360 25283 19363
rect 25682 19360 25688 19372
rect 25271 19332 25688 19360
rect 25271 19329 25283 19332
rect 25225 19323 25283 19329
rect 25682 19320 25688 19332
rect 25740 19320 25746 19372
rect 22278 19292 22284 19304
rect 22112 19264 22284 19292
rect 21361 19255 21419 19261
rect 21376 19224 21404 19255
rect 22278 19252 22284 19264
rect 22336 19252 22342 19304
rect 22830 19252 22836 19304
rect 22888 19292 22894 19304
rect 24854 19292 24860 19304
rect 22888 19264 24860 19292
rect 22888 19252 22894 19264
rect 24854 19252 24860 19264
rect 24912 19252 24918 19304
rect 24946 19252 24952 19304
rect 25004 19292 25010 19304
rect 25590 19292 25596 19304
rect 25004 19264 25596 19292
rect 25004 19252 25010 19264
rect 25590 19252 25596 19264
rect 25648 19252 25654 19304
rect 25792 19292 25820 19400
rect 26068 19360 26096 19468
rect 26142 19456 26148 19508
rect 26200 19456 26206 19508
rect 26234 19456 26240 19508
rect 26292 19496 26298 19508
rect 27338 19496 27344 19508
rect 26292 19468 27344 19496
rect 26292 19456 26298 19468
rect 27338 19456 27344 19468
rect 27396 19456 27402 19508
rect 27430 19456 27436 19508
rect 27488 19496 27494 19508
rect 28350 19496 28356 19508
rect 27488 19468 28356 19496
rect 27488 19456 27494 19468
rect 28350 19456 28356 19468
rect 28408 19456 28414 19508
rect 28445 19499 28503 19505
rect 28445 19465 28457 19499
rect 28491 19496 28503 19499
rect 28718 19496 28724 19508
rect 28491 19468 28724 19496
rect 28491 19465 28503 19468
rect 28445 19459 28503 19465
rect 28718 19456 28724 19468
rect 28776 19456 28782 19508
rect 30190 19456 30196 19508
rect 30248 19496 30254 19508
rect 31846 19496 31852 19508
rect 30248 19468 31852 19496
rect 30248 19456 30254 19468
rect 31846 19456 31852 19468
rect 31904 19456 31910 19508
rect 32490 19456 32496 19508
rect 32548 19496 32554 19508
rect 33045 19499 33103 19505
rect 33045 19496 33057 19499
rect 32548 19468 33057 19496
rect 32548 19456 32554 19468
rect 33045 19465 33057 19468
rect 33091 19465 33103 19499
rect 33045 19459 33103 19465
rect 34241 19499 34299 19505
rect 34241 19465 34253 19499
rect 34287 19496 34299 19499
rect 34974 19496 34980 19508
rect 34287 19468 34980 19496
rect 34287 19465 34299 19468
rect 34241 19459 34299 19465
rect 34974 19456 34980 19468
rect 35032 19456 35038 19508
rect 35437 19499 35495 19505
rect 35437 19465 35449 19499
rect 35483 19496 35495 19499
rect 36538 19496 36544 19508
rect 35483 19468 36544 19496
rect 35483 19465 35495 19468
rect 35437 19459 35495 19465
rect 36538 19456 36544 19468
rect 36596 19456 36602 19508
rect 36998 19456 37004 19508
rect 37056 19496 37062 19508
rect 37277 19499 37335 19505
rect 37277 19496 37289 19499
rect 37056 19468 37289 19496
rect 37056 19456 37062 19468
rect 37277 19465 37289 19468
rect 37323 19465 37335 19499
rect 38470 19496 38476 19508
rect 37277 19459 37335 19465
rect 38304 19468 38476 19496
rect 26160 19428 26188 19456
rect 26160 19400 30880 19428
rect 27617 19363 27675 19369
rect 26068 19332 27568 19360
rect 26421 19295 26479 19301
rect 26421 19292 26433 19295
rect 25792 19264 26433 19292
rect 26421 19261 26433 19264
rect 26467 19292 26479 19295
rect 27430 19292 27436 19304
rect 26467 19264 27436 19292
rect 26467 19261 26479 19264
rect 26421 19255 26479 19261
rect 27430 19252 27436 19264
rect 27488 19252 27494 19304
rect 27540 19292 27568 19332
rect 27617 19329 27629 19363
rect 27663 19360 27675 19363
rect 28442 19360 28448 19372
rect 27663 19332 28448 19360
rect 27663 19329 27675 19332
rect 27617 19323 27675 19329
rect 28442 19320 28448 19332
rect 28500 19320 28506 19372
rect 28813 19363 28871 19369
rect 28813 19329 28825 19363
rect 28859 19360 28871 19363
rect 29733 19363 29791 19369
rect 29733 19360 29745 19363
rect 28859 19332 29745 19360
rect 28859 19329 28871 19332
rect 28813 19323 28871 19329
rect 29733 19329 29745 19332
rect 29779 19329 29791 19363
rect 29733 19323 29791 19329
rect 29932 19332 30328 19360
rect 27709 19295 27767 19301
rect 27540 19264 27660 19292
rect 21376 19196 22094 19224
rect 19668 19128 20024 19156
rect 20441 19159 20499 19165
rect 19668 19116 19674 19128
rect 20441 19125 20453 19159
rect 20487 19156 20499 19159
rect 21174 19156 21180 19168
rect 20487 19128 21180 19156
rect 20487 19125 20499 19128
rect 20441 19119 20499 19125
rect 21174 19116 21180 19128
rect 21232 19116 21238 19168
rect 22066 19156 22094 19196
rect 23477 19159 23535 19165
rect 23477 19156 23489 19159
rect 22066 19128 23489 19156
rect 23477 19125 23489 19128
rect 23523 19156 23535 19159
rect 23842 19156 23848 19168
rect 23523 19128 23848 19156
rect 23523 19125 23535 19128
rect 23477 19119 23535 19125
rect 23842 19116 23848 19128
rect 23900 19116 23906 19168
rect 25774 19116 25780 19168
rect 25832 19116 25838 19168
rect 27246 19116 27252 19168
rect 27304 19116 27310 19168
rect 27632 19156 27660 19264
rect 27709 19261 27721 19295
rect 27755 19261 27767 19295
rect 27709 19255 27767 19261
rect 27893 19295 27951 19301
rect 27893 19261 27905 19295
rect 27939 19292 27951 19295
rect 28074 19292 28080 19304
rect 27939 19264 28080 19292
rect 27939 19261 27951 19264
rect 27893 19255 27951 19261
rect 27724 19224 27752 19255
rect 28074 19252 28080 19264
rect 28132 19252 28138 19304
rect 28626 19252 28632 19304
rect 28684 19292 28690 19304
rect 28905 19295 28963 19301
rect 28905 19292 28917 19295
rect 28684 19264 28917 19292
rect 28684 19252 28690 19264
rect 28905 19261 28917 19264
rect 28951 19261 28963 19295
rect 28905 19255 28963 19261
rect 28997 19295 29055 19301
rect 28997 19261 29009 19295
rect 29043 19261 29055 19295
rect 28997 19255 29055 19261
rect 28534 19224 28540 19236
rect 27724 19196 28540 19224
rect 28534 19184 28540 19196
rect 28592 19184 28598 19236
rect 29012 19224 29040 19255
rect 29270 19252 29276 19304
rect 29328 19292 29334 19304
rect 29932 19292 29960 19332
rect 29328 19264 29960 19292
rect 30300 19292 30328 19332
rect 30374 19320 30380 19372
rect 30432 19360 30438 19372
rect 30745 19363 30803 19369
rect 30745 19360 30757 19363
rect 30432 19332 30757 19360
rect 30432 19320 30438 19332
rect 30745 19329 30757 19332
rect 30791 19329 30803 19363
rect 30852 19360 30880 19400
rect 31478 19388 31484 19440
rect 31536 19388 31542 19440
rect 31754 19388 31760 19440
rect 31812 19428 31818 19440
rect 32585 19431 32643 19437
rect 32585 19428 32597 19431
rect 31812 19400 32597 19428
rect 31812 19388 31818 19400
rect 32585 19397 32597 19400
rect 32631 19397 32643 19431
rect 32585 19391 32643 19397
rect 32677 19431 32735 19437
rect 32677 19397 32689 19431
rect 32723 19428 32735 19431
rect 32858 19428 32864 19440
rect 32723 19400 32864 19428
rect 32723 19397 32735 19400
rect 32677 19391 32735 19397
rect 32858 19388 32864 19400
rect 32916 19388 32922 19440
rect 33781 19431 33839 19437
rect 33781 19397 33793 19431
rect 33827 19428 33839 19431
rect 34698 19428 34704 19440
rect 33827 19400 34704 19428
rect 33827 19397 33839 19400
rect 33781 19391 33839 19397
rect 33796 19360 33824 19391
rect 34698 19388 34704 19400
rect 34756 19388 34762 19440
rect 34790 19388 34796 19440
rect 34848 19428 34854 19440
rect 35069 19431 35127 19437
rect 34848 19400 35020 19428
rect 34848 19388 34854 19400
rect 34992 19372 35020 19400
rect 35069 19397 35081 19431
rect 35115 19428 35127 19431
rect 35342 19428 35348 19440
rect 35115 19400 35348 19428
rect 35115 19397 35127 19400
rect 35069 19391 35127 19397
rect 35342 19388 35348 19400
rect 35400 19388 35406 19440
rect 35894 19388 35900 19440
rect 35952 19428 35958 19440
rect 36173 19431 36231 19437
rect 36173 19428 36185 19431
rect 35952 19400 36185 19428
rect 35952 19388 35958 19400
rect 36173 19397 36185 19400
rect 36219 19397 36231 19431
rect 36173 19391 36231 19397
rect 30852 19332 33824 19360
rect 33873 19363 33931 19369
rect 30745 19323 30803 19329
rect 33873 19329 33885 19363
rect 33919 19360 33931 19363
rect 34238 19360 34244 19372
rect 33919 19332 34244 19360
rect 33919 19329 33931 19332
rect 33873 19323 33931 19329
rect 34238 19320 34244 19332
rect 34296 19320 34302 19372
rect 34882 19360 34888 19372
rect 34440 19332 34888 19360
rect 31662 19292 31668 19304
rect 30300 19264 31668 19292
rect 29328 19252 29334 19264
rect 31662 19252 31668 19264
rect 31720 19252 31726 19304
rect 32398 19252 32404 19304
rect 32456 19252 32462 19304
rect 33689 19295 33747 19301
rect 33689 19261 33701 19295
rect 33735 19292 33747 19295
rect 34440 19292 34468 19332
rect 34882 19320 34888 19332
rect 34940 19320 34946 19372
rect 34974 19320 34980 19372
rect 35032 19320 35038 19372
rect 35526 19320 35532 19372
rect 35584 19360 35590 19372
rect 36265 19363 36323 19369
rect 36265 19360 36277 19363
rect 35584 19332 36277 19360
rect 35584 19320 35590 19332
rect 36265 19329 36277 19332
rect 36311 19329 36323 19363
rect 36265 19323 36323 19329
rect 36722 19320 36728 19372
rect 36780 19360 36786 19372
rect 37366 19360 37372 19372
rect 36780 19332 37372 19360
rect 36780 19320 36786 19332
rect 37366 19320 37372 19332
rect 37424 19360 37430 19372
rect 37553 19363 37611 19369
rect 37553 19360 37565 19363
rect 37424 19332 37565 19360
rect 37424 19320 37430 19332
rect 37553 19329 37565 19332
rect 37599 19360 37611 19363
rect 38304 19360 38332 19468
rect 38470 19456 38476 19468
rect 38528 19456 38534 19508
rect 40034 19456 40040 19508
rect 40092 19496 40098 19508
rect 40129 19499 40187 19505
rect 40129 19496 40141 19499
rect 40092 19468 40141 19496
rect 40092 19456 40098 19468
rect 40129 19465 40141 19468
rect 40175 19465 40187 19499
rect 40129 19459 40187 19465
rect 40402 19456 40408 19508
rect 40460 19496 40466 19508
rect 40589 19499 40647 19505
rect 40589 19496 40601 19499
rect 40460 19468 40601 19496
rect 40460 19456 40466 19468
rect 40589 19465 40601 19468
rect 40635 19496 40647 19499
rect 41325 19499 41383 19505
rect 41325 19496 41337 19499
rect 40635 19468 41337 19496
rect 40635 19465 40647 19468
rect 40589 19459 40647 19465
rect 41325 19465 41337 19468
rect 41371 19465 41383 19499
rect 41325 19459 41383 19465
rect 39390 19388 39396 19440
rect 39448 19388 39454 19440
rect 40497 19431 40555 19437
rect 40497 19397 40509 19431
rect 40543 19428 40555 19431
rect 48406 19428 48412 19440
rect 40543 19400 48412 19428
rect 40543 19397 40555 19400
rect 40497 19391 40555 19397
rect 48406 19388 48412 19400
rect 48464 19388 48470 19440
rect 37599 19346 38332 19360
rect 37599 19332 38318 19346
rect 37599 19329 37611 19332
rect 37553 19323 37611 19329
rect 39666 19320 39672 19372
rect 39724 19320 39730 19372
rect 48593 19363 48651 19369
rect 48593 19329 48605 19363
rect 48639 19360 48651 19363
rect 49234 19360 49240 19372
rect 48639 19332 49240 19360
rect 48639 19329 48651 19332
rect 48593 19323 48651 19329
rect 49234 19320 49240 19332
rect 49292 19320 49298 19372
rect 34793 19295 34851 19301
rect 34793 19292 34805 19295
rect 33735 19264 34468 19292
rect 34532 19264 34805 19292
rect 33735 19261 33747 19264
rect 33689 19255 33747 19261
rect 28920 19196 29040 19224
rect 28920 19168 28948 19196
rect 29914 19184 29920 19236
rect 29972 19224 29978 19236
rect 34422 19224 34428 19236
rect 29972 19196 34428 19224
rect 29972 19184 29978 19196
rect 34422 19184 34428 19196
rect 34480 19184 34486 19236
rect 28902 19156 28908 19168
rect 27632 19128 28908 19156
rect 28902 19116 28908 19128
rect 28960 19116 28966 19168
rect 30006 19116 30012 19168
rect 30064 19156 30070 19168
rect 30193 19159 30251 19165
rect 30193 19156 30205 19159
rect 30064 19128 30205 19156
rect 30064 19116 30070 19128
rect 30193 19125 30205 19128
rect 30239 19125 30251 19159
rect 30193 19119 30251 19125
rect 30374 19116 30380 19168
rect 30432 19116 30438 19168
rect 34532 19156 34560 19264
rect 34793 19261 34805 19264
rect 34839 19261 34851 19295
rect 34793 19255 34851 19261
rect 35894 19252 35900 19304
rect 35952 19292 35958 19304
rect 35989 19295 36047 19301
rect 35989 19292 36001 19295
rect 35952 19264 36001 19292
rect 35952 19252 35958 19264
rect 35989 19261 36001 19264
rect 36035 19261 36047 19295
rect 35989 19255 36047 19261
rect 36078 19252 36084 19304
rect 36136 19292 36142 19304
rect 40310 19292 40316 19304
rect 36136 19264 40316 19292
rect 36136 19252 36142 19264
rect 40310 19252 40316 19264
rect 40368 19252 40374 19304
rect 40681 19295 40739 19301
rect 40681 19261 40693 19295
rect 40727 19261 40739 19295
rect 40681 19255 40739 19261
rect 37734 19224 37740 19236
rect 35268 19196 37740 19224
rect 35268 19156 35296 19196
rect 37734 19184 37740 19196
rect 37792 19224 37798 19236
rect 37792 19196 38056 19224
rect 37792 19184 37798 19196
rect 34532 19128 35296 19156
rect 36630 19116 36636 19168
rect 36688 19116 36694 19168
rect 36814 19116 36820 19168
rect 36872 19156 36878 19168
rect 36909 19159 36967 19165
rect 36909 19156 36921 19159
rect 36872 19128 36921 19156
rect 36872 19116 36878 19128
rect 36909 19125 36921 19128
rect 36955 19125 36967 19159
rect 36909 19119 36967 19125
rect 37826 19116 37832 19168
rect 37884 19156 37890 19168
rect 37921 19159 37979 19165
rect 37921 19156 37933 19159
rect 37884 19128 37933 19156
rect 37884 19116 37890 19128
rect 37921 19125 37933 19128
rect 37967 19125 37979 19159
rect 38028 19156 38056 19196
rect 40696 19156 40724 19255
rect 40862 19184 40868 19236
rect 40920 19224 40926 19236
rect 49053 19227 49111 19233
rect 49053 19224 49065 19227
rect 40920 19196 49065 19224
rect 40920 19184 40926 19196
rect 49053 19193 49065 19196
rect 49099 19193 49111 19227
rect 49053 19187 49111 19193
rect 38028 19128 40724 19156
rect 37921 19119 37979 19125
rect 41046 19116 41052 19168
rect 41104 19156 41110 19168
rect 41233 19159 41291 19165
rect 41233 19156 41245 19159
rect 41104 19128 41245 19156
rect 41104 19116 41110 19128
rect 41233 19125 41245 19128
rect 41279 19156 41291 19159
rect 42058 19156 42064 19168
rect 41279 19128 42064 19156
rect 41279 19125 41291 19128
rect 41233 19119 41291 19125
rect 42058 19116 42064 19128
rect 42116 19116 42122 19168
rect 48777 19159 48835 19165
rect 48777 19125 48789 19159
rect 48823 19156 48835 19159
rect 49418 19156 49424 19168
rect 48823 19128 49424 19156
rect 48823 19125 48835 19128
rect 48777 19119 48835 19125
rect 49418 19116 49424 19128
rect 49476 19116 49482 19168
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 6822 18912 6828 18964
rect 6880 18952 6886 18964
rect 9217 18955 9275 18961
rect 9217 18952 9229 18955
rect 6880 18924 9229 18952
rect 6880 18912 6886 18924
rect 9217 18921 9229 18924
rect 9263 18952 9275 18955
rect 10870 18952 10876 18964
rect 9263 18924 10876 18952
rect 9263 18921 9275 18924
rect 9217 18915 9275 18921
rect 10870 18912 10876 18924
rect 10928 18912 10934 18964
rect 11882 18912 11888 18964
rect 11940 18912 11946 18964
rect 12342 18912 12348 18964
rect 12400 18952 12406 18964
rect 12529 18955 12587 18961
rect 12529 18952 12541 18955
rect 12400 18924 12541 18952
rect 12400 18912 12406 18924
rect 12529 18921 12541 18924
rect 12575 18921 12587 18955
rect 15102 18952 15108 18964
rect 12529 18915 12587 18921
rect 12636 18924 15108 18952
rect 11054 18884 11060 18896
rect 10888 18856 11060 18884
rect 3510 18776 3516 18828
rect 3568 18816 3574 18828
rect 4157 18819 4215 18825
rect 4157 18816 4169 18819
rect 3568 18788 4169 18816
rect 3568 18776 3574 18788
rect 4157 18785 4169 18788
rect 4203 18785 4215 18819
rect 10888 18816 10916 18856
rect 11054 18844 11060 18856
rect 11112 18844 11118 18896
rect 4157 18779 4215 18785
rect 8312 18788 10916 18816
rect 10965 18819 11023 18825
rect 2961 18751 3019 18757
rect 2961 18717 2973 18751
rect 3007 18717 3019 18751
rect 2961 18711 3019 18717
rect 1394 18640 1400 18692
rect 1452 18680 1458 18692
rect 1765 18683 1823 18689
rect 1765 18680 1777 18683
rect 1452 18652 1777 18680
rect 1452 18640 1458 18652
rect 1765 18649 1777 18652
rect 1811 18649 1823 18683
rect 1765 18643 1823 18649
rect 2976 18612 3004 18711
rect 5350 18708 5356 18760
rect 5408 18708 5414 18760
rect 8312 18757 8340 18788
rect 10965 18785 10977 18819
rect 11011 18816 11023 18819
rect 12526 18816 12532 18828
rect 11011 18788 12532 18816
rect 11011 18785 11023 18788
rect 10965 18779 11023 18785
rect 12526 18776 12532 18788
rect 12584 18776 12590 18828
rect 8297 18751 8355 18757
rect 8297 18717 8309 18751
rect 8343 18717 8355 18751
rect 8297 18711 8355 18717
rect 12069 18751 12127 18757
rect 12069 18717 12081 18751
rect 12115 18748 12127 18751
rect 12434 18748 12440 18760
rect 12115 18720 12440 18748
rect 12115 18717 12127 18720
rect 12069 18711 12127 18717
rect 12434 18708 12440 18720
rect 12492 18708 12498 18760
rect 4338 18640 4344 18692
rect 4396 18680 4402 18692
rect 8113 18683 8171 18689
rect 8113 18680 8125 18683
rect 4396 18652 8125 18680
rect 4396 18640 4402 18652
rect 8113 18649 8125 18652
rect 8159 18649 8171 18683
rect 8113 18643 8171 18649
rect 10134 18640 10140 18692
rect 10192 18640 10198 18692
rect 10226 18640 10232 18692
rect 10284 18680 10290 18692
rect 10284 18652 10640 18680
rect 10284 18640 10290 18652
rect 10410 18612 10416 18624
rect 2976 18584 10416 18612
rect 10410 18572 10416 18584
rect 10468 18572 10474 18624
rect 10612 18612 10640 18652
rect 10686 18640 10692 18692
rect 10744 18640 10750 18692
rect 12158 18640 12164 18692
rect 12216 18680 12222 18692
rect 12636 18680 12664 18924
rect 15102 18912 15108 18924
rect 15160 18912 15166 18964
rect 15194 18912 15200 18964
rect 15252 18952 15258 18964
rect 16025 18955 16083 18961
rect 16025 18952 16037 18955
rect 15252 18924 16037 18952
rect 15252 18912 15258 18924
rect 16025 18921 16037 18924
rect 16071 18952 16083 18955
rect 16114 18952 16120 18964
rect 16071 18924 16120 18952
rect 16071 18921 16083 18924
rect 16025 18915 16083 18921
rect 16114 18912 16120 18924
rect 16172 18912 16178 18964
rect 16945 18955 17003 18961
rect 16945 18921 16957 18955
rect 16991 18921 17003 18955
rect 16945 18915 17003 18921
rect 13354 18844 13360 18896
rect 13412 18884 13418 18896
rect 13725 18887 13783 18893
rect 13725 18884 13737 18887
rect 13412 18856 13737 18884
rect 13412 18844 13418 18856
rect 13725 18853 13737 18856
rect 13771 18884 13783 18887
rect 13814 18884 13820 18896
rect 13771 18856 13820 18884
rect 13771 18853 13783 18856
rect 13725 18847 13783 18853
rect 13814 18844 13820 18856
rect 13872 18844 13878 18896
rect 15654 18844 15660 18896
rect 15712 18884 15718 18896
rect 16960 18884 16988 18915
rect 17862 18912 17868 18964
rect 17920 18952 17926 18964
rect 18141 18955 18199 18961
rect 18141 18952 18153 18955
rect 17920 18924 18153 18952
rect 17920 18912 17926 18924
rect 18141 18921 18153 18924
rect 18187 18921 18199 18955
rect 18141 18915 18199 18921
rect 19518 18912 19524 18964
rect 19576 18952 19582 18964
rect 19889 18955 19947 18961
rect 19889 18952 19901 18955
rect 19576 18924 19901 18952
rect 19576 18912 19582 18924
rect 19889 18921 19901 18924
rect 19935 18921 19947 18955
rect 19889 18915 19947 18921
rect 20714 18912 20720 18964
rect 20772 18952 20778 18964
rect 21085 18955 21143 18961
rect 21085 18952 21097 18955
rect 20772 18924 21097 18952
rect 20772 18912 20778 18924
rect 21085 18921 21097 18924
rect 21131 18921 21143 18955
rect 21085 18915 21143 18921
rect 23106 18912 23112 18964
rect 23164 18952 23170 18964
rect 27614 18952 27620 18964
rect 23164 18924 27620 18952
rect 23164 18912 23170 18924
rect 27614 18912 27620 18924
rect 27672 18912 27678 18964
rect 27706 18912 27712 18964
rect 27764 18952 27770 18964
rect 28077 18955 28135 18961
rect 28077 18952 28089 18955
rect 27764 18924 28089 18952
rect 27764 18912 27770 18924
rect 28077 18921 28089 18924
rect 28123 18952 28135 18955
rect 30190 18952 30196 18964
rect 28123 18924 30196 18952
rect 28123 18921 28135 18924
rect 28077 18915 28135 18921
rect 30190 18912 30196 18924
rect 30248 18912 30254 18964
rect 30466 18912 30472 18964
rect 30524 18952 30530 18964
rect 31481 18955 31539 18961
rect 31481 18952 31493 18955
rect 30524 18924 31493 18952
rect 30524 18912 30530 18924
rect 31481 18921 31493 18924
rect 31527 18921 31539 18955
rect 33318 18952 33324 18964
rect 31481 18915 31539 18921
rect 31956 18924 33324 18952
rect 20622 18884 20628 18896
rect 15712 18856 16988 18884
rect 20364 18856 20628 18884
rect 15712 18844 15718 18856
rect 12710 18776 12716 18828
rect 12768 18816 12774 18828
rect 13081 18819 13139 18825
rect 13081 18816 13093 18819
rect 12768 18788 13093 18816
rect 12768 18776 12774 18788
rect 13081 18785 13093 18788
rect 13127 18816 13139 18819
rect 13170 18816 13176 18828
rect 13127 18788 13176 18816
rect 13127 18785 13139 18788
rect 13081 18779 13139 18785
rect 13170 18776 13176 18788
rect 13228 18776 13234 18828
rect 14277 18819 14335 18825
rect 14277 18785 14289 18819
rect 14323 18816 14335 18819
rect 16942 18816 16948 18828
rect 14323 18788 16948 18816
rect 14323 18785 14335 18788
rect 14277 18779 14335 18785
rect 16942 18776 16948 18788
rect 17000 18776 17006 18828
rect 17494 18776 17500 18828
rect 17552 18776 17558 18828
rect 18785 18819 18843 18825
rect 18785 18785 18797 18819
rect 18831 18816 18843 18819
rect 19702 18816 19708 18828
rect 18831 18788 19708 18816
rect 18831 18785 18843 18788
rect 18785 18779 18843 18785
rect 19702 18776 19708 18788
rect 19760 18776 19766 18828
rect 20364 18825 20392 18856
rect 20622 18844 20628 18856
rect 20680 18844 20686 18896
rect 27525 18887 27583 18893
rect 25148 18856 25912 18884
rect 20349 18819 20407 18825
rect 20349 18785 20361 18819
rect 20395 18785 20407 18819
rect 20349 18779 20407 18785
rect 20438 18776 20444 18828
rect 20496 18776 20502 18828
rect 21358 18776 21364 18828
rect 21416 18816 21422 18828
rect 21637 18819 21695 18825
rect 21637 18816 21649 18819
rect 21416 18788 21649 18816
rect 21416 18776 21422 18788
rect 21637 18785 21649 18788
rect 21683 18785 21695 18819
rect 21637 18779 21695 18785
rect 23014 18776 23020 18828
rect 23072 18816 23078 18828
rect 25148 18816 25176 18856
rect 23072 18788 25176 18816
rect 25225 18819 25283 18825
rect 23072 18776 23078 18788
rect 25225 18785 25237 18819
rect 25271 18816 25283 18819
rect 25590 18816 25596 18828
rect 25271 18788 25596 18816
rect 25271 18785 25283 18788
rect 25225 18779 25283 18785
rect 25590 18776 25596 18788
rect 25648 18776 25654 18828
rect 25682 18776 25688 18828
rect 25740 18816 25746 18828
rect 25777 18819 25835 18825
rect 25777 18816 25789 18819
rect 25740 18788 25789 18816
rect 25740 18776 25746 18788
rect 25777 18785 25789 18788
rect 25823 18785 25835 18819
rect 25884 18816 25912 18856
rect 27525 18853 27537 18887
rect 27571 18884 27583 18887
rect 28902 18884 28908 18896
rect 27571 18856 28908 18884
rect 27571 18853 27583 18856
rect 27525 18847 27583 18853
rect 28902 18844 28908 18856
rect 28960 18844 28966 18896
rect 28994 18844 29000 18896
rect 29052 18844 29058 18896
rect 29178 18844 29184 18896
rect 29236 18884 29242 18896
rect 30742 18884 30748 18896
rect 29236 18856 30748 18884
rect 29236 18844 29242 18856
rect 30742 18844 30748 18856
rect 30800 18844 30806 18896
rect 30926 18844 30932 18896
rect 30984 18844 30990 18896
rect 27062 18816 27068 18828
rect 25884 18788 27068 18816
rect 25777 18779 25835 18785
rect 27062 18776 27068 18788
rect 27120 18776 27126 18828
rect 27430 18816 27436 18828
rect 27172 18788 27436 18816
rect 12802 18708 12808 18760
rect 12860 18748 12866 18760
rect 12897 18751 12955 18757
rect 12897 18748 12909 18751
rect 12860 18720 12909 18748
rect 12860 18708 12866 18720
rect 12897 18717 12909 18720
rect 12943 18717 12955 18751
rect 12897 18711 12955 18717
rect 18506 18708 18512 18760
rect 18564 18708 18570 18760
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18748 18659 18751
rect 21082 18748 21088 18760
rect 18647 18720 21088 18748
rect 18647 18717 18659 18720
rect 18601 18711 18659 18717
rect 21082 18708 21088 18720
rect 21140 18708 21146 18760
rect 21453 18751 21511 18757
rect 21453 18717 21465 18751
rect 21499 18748 21511 18751
rect 21818 18748 21824 18760
rect 21499 18720 21824 18748
rect 21499 18717 21511 18720
rect 21453 18711 21511 18717
rect 21818 18708 21824 18720
rect 21876 18708 21882 18760
rect 24029 18751 24087 18757
rect 24029 18717 24041 18751
rect 24075 18748 24087 18751
rect 24118 18748 24124 18760
rect 24075 18720 24124 18748
rect 24075 18717 24087 18720
rect 24029 18711 24087 18717
rect 24118 18708 24124 18720
rect 24176 18748 24182 18760
rect 25700 18748 25728 18776
rect 24176 18720 25728 18748
rect 27172 18734 27200 18788
rect 27430 18776 27436 18788
rect 27488 18816 27494 18828
rect 27801 18819 27859 18825
rect 27801 18816 27813 18819
rect 27488 18788 27813 18816
rect 27488 18776 27494 18788
rect 27801 18785 27813 18788
rect 27847 18816 27859 18819
rect 27982 18816 27988 18828
rect 27847 18788 27988 18816
rect 27847 18785 27859 18788
rect 27801 18779 27859 18785
rect 27982 18776 27988 18788
rect 28040 18776 28046 18828
rect 28442 18776 28448 18828
rect 28500 18776 28506 18828
rect 29270 18816 29276 18828
rect 28966 18788 29276 18816
rect 24176 18708 24182 18720
rect 28074 18708 28080 18760
rect 28132 18748 28138 18760
rect 28966 18748 28994 18788
rect 29270 18776 29276 18788
rect 29328 18776 29334 18828
rect 29546 18776 29552 18828
rect 29604 18816 29610 18828
rect 31956 18825 31984 18924
rect 33318 18912 33324 18924
rect 33376 18912 33382 18964
rect 33413 18955 33471 18961
rect 33413 18921 33425 18955
rect 33459 18952 33471 18955
rect 33962 18952 33968 18964
rect 33459 18924 33968 18952
rect 33459 18921 33471 18924
rect 33413 18915 33471 18921
rect 33962 18912 33968 18924
rect 34020 18912 34026 18964
rect 34330 18912 34336 18964
rect 34388 18912 34394 18964
rect 34422 18912 34428 18964
rect 34480 18952 34486 18964
rect 37369 18955 37427 18961
rect 34480 18924 36952 18952
rect 34480 18912 34486 18924
rect 32048 18856 32996 18884
rect 29825 18819 29883 18825
rect 29825 18816 29837 18819
rect 29604 18788 29837 18816
rect 29604 18776 29610 18788
rect 29825 18785 29837 18788
rect 29871 18785 29883 18819
rect 29825 18779 29883 18785
rect 31941 18819 31999 18825
rect 31941 18785 31953 18819
rect 31987 18785 31999 18819
rect 31941 18779 31999 18785
rect 28132 18720 28994 18748
rect 29181 18751 29239 18757
rect 28132 18708 28138 18720
rect 29181 18717 29193 18751
rect 29227 18748 29239 18751
rect 31018 18748 31024 18760
rect 29227 18720 31024 18748
rect 29227 18717 29239 18720
rect 29181 18711 29239 18717
rect 31018 18708 31024 18720
rect 31076 18708 31082 18760
rect 31110 18708 31116 18760
rect 31168 18748 31174 18760
rect 31168 18720 31432 18748
rect 31168 18708 31174 18720
rect 12216 18652 12664 18680
rect 12989 18683 13047 18689
rect 12216 18640 12222 18652
rect 12989 18649 13001 18683
rect 13035 18680 13047 18683
rect 13035 18652 14504 18680
rect 13035 18649 13047 18652
rect 12989 18643 13047 18649
rect 11241 18615 11299 18621
rect 11241 18612 11253 18615
rect 10612 18584 11253 18612
rect 11241 18581 11253 18584
rect 11287 18612 11299 18615
rect 11514 18612 11520 18624
rect 11287 18584 11520 18612
rect 11287 18581 11299 18584
rect 11241 18575 11299 18581
rect 11514 18572 11520 18584
rect 11572 18572 11578 18624
rect 13909 18615 13967 18621
rect 13909 18581 13921 18615
rect 13955 18612 13967 18615
rect 14090 18612 14096 18624
rect 13955 18584 14096 18612
rect 13955 18581 13967 18584
rect 13909 18575 13967 18581
rect 14090 18572 14096 18584
rect 14148 18572 14154 18624
rect 14476 18612 14504 18652
rect 14550 18640 14556 18692
rect 14608 18640 14614 18692
rect 14826 18640 14832 18692
rect 14884 18680 14890 18692
rect 14884 18652 15042 18680
rect 14884 18640 14890 18652
rect 16298 18640 16304 18692
rect 16356 18640 16362 18692
rect 17402 18640 17408 18692
rect 17460 18640 17466 18692
rect 19334 18640 19340 18692
rect 19392 18640 19398 18692
rect 19426 18640 19432 18692
rect 19484 18680 19490 18692
rect 20257 18683 20315 18689
rect 19484 18652 20208 18680
rect 19484 18640 19490 18652
rect 15562 18612 15568 18624
rect 14476 18584 15568 18612
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 16666 18572 16672 18624
rect 16724 18612 16730 18624
rect 17313 18615 17371 18621
rect 17313 18612 17325 18615
rect 16724 18584 17325 18612
rect 16724 18572 16730 18584
rect 17313 18581 17325 18584
rect 17359 18581 17371 18615
rect 17313 18575 17371 18581
rect 19610 18572 19616 18624
rect 19668 18572 19674 18624
rect 20180 18612 20208 18652
rect 20257 18649 20269 18683
rect 20303 18680 20315 18683
rect 20303 18652 22508 18680
rect 20303 18649 20315 18652
rect 20257 18643 20315 18649
rect 21450 18612 21456 18624
rect 20180 18584 21456 18612
rect 21450 18572 21456 18584
rect 21508 18572 21514 18624
rect 21545 18615 21603 18621
rect 21545 18581 21557 18615
rect 21591 18612 21603 18615
rect 22002 18612 22008 18624
rect 21591 18584 22008 18612
rect 21591 18581 21603 18584
rect 21545 18575 21603 18581
rect 22002 18572 22008 18584
rect 22060 18572 22066 18624
rect 22094 18572 22100 18624
rect 22152 18612 22158 18624
rect 22281 18615 22339 18621
rect 22281 18612 22293 18615
rect 22152 18584 22293 18612
rect 22152 18572 22158 18584
rect 22281 18581 22293 18584
rect 22327 18612 22339 18615
rect 22370 18612 22376 18624
rect 22327 18584 22376 18612
rect 22327 18581 22339 18584
rect 22281 18575 22339 18581
rect 22370 18572 22376 18584
rect 22428 18572 22434 18624
rect 22480 18612 22508 18652
rect 23290 18640 23296 18692
rect 23348 18640 23354 18692
rect 23474 18640 23480 18692
rect 23532 18680 23538 18692
rect 23753 18683 23811 18689
rect 23753 18680 23765 18683
rect 23532 18652 23765 18680
rect 23532 18640 23538 18652
rect 23753 18649 23765 18652
rect 23799 18649 23811 18683
rect 23753 18643 23811 18649
rect 23842 18640 23848 18692
rect 23900 18680 23906 18692
rect 26053 18683 26111 18689
rect 26053 18680 26065 18683
rect 23900 18652 26065 18680
rect 23900 18640 23906 18652
rect 26053 18649 26065 18652
rect 26099 18649 26111 18683
rect 26053 18643 26111 18649
rect 27356 18652 29224 18680
rect 24581 18615 24639 18621
rect 24581 18612 24593 18615
rect 22480 18584 24593 18612
rect 24581 18581 24593 18584
rect 24627 18581 24639 18615
rect 24581 18575 24639 18581
rect 24854 18572 24860 18624
rect 24912 18612 24918 18624
rect 24949 18615 25007 18621
rect 24949 18612 24961 18615
rect 24912 18584 24961 18612
rect 24912 18572 24918 18584
rect 24949 18581 24961 18584
rect 24995 18581 25007 18615
rect 24949 18575 25007 18581
rect 25038 18572 25044 18624
rect 25096 18572 25102 18624
rect 26326 18572 26332 18624
rect 26384 18612 26390 18624
rect 27356 18612 27384 18652
rect 29196 18624 29224 18652
rect 29362 18640 29368 18692
rect 29420 18680 29426 18692
rect 30101 18683 30159 18689
rect 30101 18680 30113 18683
rect 29420 18652 30113 18680
rect 29420 18640 29426 18652
rect 30101 18649 30113 18652
rect 30147 18649 30159 18683
rect 30745 18683 30803 18689
rect 30745 18680 30757 18683
rect 30101 18643 30159 18649
rect 30208 18652 30757 18680
rect 26384 18584 27384 18612
rect 26384 18572 26390 18584
rect 27614 18572 27620 18624
rect 27672 18612 27678 18624
rect 28074 18612 28080 18624
rect 27672 18584 28080 18612
rect 27672 18572 27678 18584
rect 28074 18572 28080 18584
rect 28132 18612 28138 18624
rect 28169 18615 28227 18621
rect 28169 18612 28181 18615
rect 28132 18584 28181 18612
rect 28132 18572 28138 18584
rect 28169 18581 28181 18584
rect 28215 18581 28227 18615
rect 28169 18575 28227 18581
rect 28626 18572 28632 18624
rect 28684 18572 28690 18624
rect 29178 18572 29184 18624
rect 29236 18572 29242 18624
rect 29638 18572 29644 18624
rect 29696 18612 29702 18624
rect 30009 18615 30067 18621
rect 30009 18612 30021 18615
rect 29696 18584 30021 18612
rect 29696 18572 29702 18584
rect 30009 18581 30021 18584
rect 30055 18612 30067 18615
rect 30208 18612 30236 18652
rect 30745 18649 30757 18652
rect 30791 18680 30803 18683
rect 31294 18680 31300 18692
rect 30791 18652 31300 18680
rect 30791 18649 30803 18652
rect 30745 18643 30803 18649
rect 31294 18640 31300 18652
rect 31352 18640 31358 18692
rect 31404 18680 31432 18720
rect 31662 18708 31668 18760
rect 31720 18748 31726 18760
rect 31849 18751 31907 18757
rect 31849 18748 31861 18751
rect 31720 18720 31861 18748
rect 31720 18708 31726 18720
rect 31849 18717 31861 18720
rect 31895 18717 31907 18751
rect 31849 18711 31907 18717
rect 32048 18680 32076 18856
rect 32968 18825 32996 18856
rect 33042 18844 33048 18896
rect 33100 18884 33106 18896
rect 33873 18887 33931 18893
rect 33873 18884 33885 18887
rect 33100 18856 33885 18884
rect 33100 18844 33106 18856
rect 33873 18853 33885 18856
rect 33919 18853 33931 18887
rect 34348 18884 34376 18912
rect 36924 18884 36952 18924
rect 37369 18921 37381 18955
rect 37415 18952 37427 18955
rect 39390 18952 39396 18964
rect 37415 18924 39396 18952
rect 37415 18921 37427 18924
rect 37369 18915 37427 18921
rect 39390 18912 39396 18924
rect 39448 18912 39454 18964
rect 42058 18912 42064 18964
rect 42116 18912 42122 18964
rect 38013 18887 38071 18893
rect 38013 18884 38025 18887
rect 34348 18856 34468 18884
rect 36924 18856 38025 18884
rect 33873 18847 33931 18853
rect 32125 18819 32183 18825
rect 32125 18785 32137 18819
rect 32171 18785 32183 18819
rect 32125 18779 32183 18785
rect 32861 18819 32919 18825
rect 32861 18785 32873 18819
rect 32907 18785 32919 18819
rect 32861 18779 32919 18785
rect 32953 18819 33011 18825
rect 32953 18785 32965 18819
rect 32999 18816 33011 18819
rect 34149 18819 34207 18825
rect 34149 18816 34161 18819
rect 32999 18788 34161 18816
rect 32999 18785 33011 18788
rect 32953 18779 33011 18785
rect 34149 18785 34161 18788
rect 34195 18816 34207 18819
rect 34330 18816 34336 18828
rect 34195 18788 34336 18816
rect 34195 18785 34207 18788
rect 34149 18779 34207 18785
rect 31404 18652 32076 18680
rect 32140 18680 32168 18779
rect 32876 18748 32904 18779
rect 34330 18776 34336 18788
rect 34388 18776 34394 18828
rect 34440 18748 34468 18856
rect 38013 18853 38025 18856
rect 38059 18853 38071 18887
rect 38013 18847 38071 18853
rect 34514 18776 34520 18828
rect 34572 18816 34578 18828
rect 35621 18819 35679 18825
rect 35621 18816 35633 18819
rect 34572 18788 35633 18816
rect 34572 18776 34578 18788
rect 35621 18785 35633 18788
rect 35667 18785 35679 18819
rect 35621 18779 35679 18785
rect 36538 18776 36544 18828
rect 36596 18816 36602 18828
rect 36596 18788 38424 18816
rect 36596 18776 36602 18788
rect 32876 18720 34468 18748
rect 35161 18751 35219 18757
rect 35161 18717 35173 18751
rect 35207 18748 35219 18751
rect 35250 18748 35256 18760
rect 35207 18720 35256 18748
rect 35207 18717 35219 18720
rect 35161 18711 35219 18717
rect 35250 18708 35256 18720
rect 35308 18708 35314 18760
rect 38396 18757 38424 18788
rect 38562 18776 38568 18828
rect 38620 18776 38626 18828
rect 41785 18819 41843 18825
rect 41785 18816 41797 18819
rect 39776 18788 41797 18816
rect 38381 18751 38439 18757
rect 38381 18717 38393 18751
rect 38427 18717 38439 18751
rect 38381 18711 38439 18717
rect 39776 18692 39804 18788
rect 41785 18785 41797 18788
rect 41831 18785 41843 18819
rect 41785 18779 41843 18785
rect 48593 18751 48651 18757
rect 48593 18717 48605 18751
rect 48639 18748 48651 18751
rect 48774 18748 48780 18760
rect 48639 18720 48780 18748
rect 48639 18717 48651 18720
rect 48593 18711 48651 18717
rect 48774 18708 48780 18720
rect 48832 18708 48838 18760
rect 49329 18751 49387 18757
rect 49329 18717 49341 18751
rect 49375 18748 49387 18751
rect 49418 18748 49424 18760
rect 49375 18720 49424 18748
rect 49375 18717 49387 18720
rect 49329 18711 49387 18717
rect 49418 18708 49424 18720
rect 49476 18708 49482 18760
rect 35618 18680 35624 18692
rect 32140 18652 35624 18680
rect 35618 18640 35624 18652
rect 35676 18680 35682 18692
rect 35897 18683 35955 18689
rect 35897 18680 35909 18683
rect 35676 18652 35909 18680
rect 35676 18640 35682 18652
rect 35897 18649 35909 18652
rect 35943 18649 35955 18683
rect 37366 18680 37372 18692
rect 37122 18652 37372 18680
rect 35897 18643 35955 18649
rect 37366 18640 37372 18652
rect 37424 18640 37430 18692
rect 39577 18683 39635 18689
rect 39577 18680 39589 18683
rect 37660 18652 39589 18680
rect 30055 18584 30236 18612
rect 30055 18581 30067 18584
rect 30009 18575 30067 18581
rect 30466 18572 30472 18624
rect 30524 18572 30530 18624
rect 30650 18572 30656 18624
rect 30708 18612 30714 18624
rect 31113 18615 31171 18621
rect 31113 18612 31125 18615
rect 30708 18584 31125 18612
rect 30708 18572 30714 18584
rect 31113 18581 31125 18584
rect 31159 18612 31171 18615
rect 31570 18612 31576 18624
rect 31159 18584 31576 18612
rect 31159 18581 31171 18584
rect 31113 18575 31171 18581
rect 31570 18572 31576 18584
rect 31628 18572 31634 18624
rect 33045 18615 33103 18621
rect 33045 18581 33057 18615
rect 33091 18612 33103 18615
rect 33410 18612 33416 18624
rect 33091 18584 33416 18612
rect 33091 18581 33103 18584
rect 33045 18575 33103 18581
rect 33410 18572 33416 18584
rect 33468 18612 33474 18624
rect 33689 18615 33747 18621
rect 33689 18612 33701 18615
rect 33468 18584 33701 18612
rect 33468 18572 33474 18584
rect 33689 18581 33701 18584
rect 33735 18581 33747 18615
rect 33689 18575 33747 18581
rect 34238 18572 34244 18624
rect 34296 18572 34302 18624
rect 34517 18615 34575 18621
rect 34517 18581 34529 18615
rect 34563 18612 34575 18615
rect 34698 18612 34704 18624
rect 34563 18584 34704 18612
rect 34563 18581 34575 18584
rect 34517 18575 34575 18581
rect 34698 18572 34704 18584
rect 34756 18572 34762 18624
rect 34882 18572 34888 18624
rect 34940 18612 34946 18624
rect 37274 18612 37280 18624
rect 34940 18584 37280 18612
rect 34940 18572 34946 18584
rect 37274 18572 37280 18584
rect 37332 18572 37338 18624
rect 37550 18572 37556 18624
rect 37608 18612 37614 18624
rect 37660 18621 37688 18652
rect 39577 18649 39589 18652
rect 39623 18680 39635 18683
rect 39758 18680 39764 18692
rect 39623 18652 39764 18680
rect 39623 18649 39635 18652
rect 39577 18643 39635 18649
rect 39758 18640 39764 18652
rect 39816 18640 39822 18692
rect 41046 18640 41052 18692
rect 41104 18640 41110 18692
rect 41509 18683 41567 18689
rect 41509 18649 41521 18683
rect 41555 18649 41567 18683
rect 41509 18643 41567 18649
rect 37645 18615 37703 18621
rect 37645 18612 37657 18615
rect 37608 18584 37657 18612
rect 37608 18572 37614 18584
rect 37645 18581 37657 18584
rect 37691 18581 37703 18615
rect 37645 18575 37703 18581
rect 38470 18572 38476 18624
rect 38528 18572 38534 18624
rect 40037 18615 40095 18621
rect 40037 18581 40049 18615
rect 40083 18612 40095 18615
rect 40126 18612 40132 18624
rect 40083 18584 40132 18612
rect 40083 18581 40095 18584
rect 40037 18575 40095 18581
rect 40126 18572 40132 18584
rect 40184 18572 40190 18624
rect 40218 18572 40224 18624
rect 40276 18612 40282 18624
rect 41524 18612 41552 18643
rect 40276 18584 41552 18612
rect 40276 18572 40282 18584
rect 48406 18572 48412 18624
rect 48464 18572 48470 18624
rect 48498 18572 48504 18624
rect 48556 18612 48562 18624
rect 49145 18615 49203 18621
rect 49145 18612 49157 18615
rect 48556 18584 49157 18612
rect 48556 18572 48562 18584
rect 49145 18581 49157 18584
rect 49191 18581 49203 18615
rect 49145 18575 49203 18581
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 3602 18368 3608 18420
rect 3660 18368 3666 18420
rect 9858 18368 9864 18420
rect 9916 18408 9922 18420
rect 10781 18411 10839 18417
rect 10781 18408 10793 18411
rect 9916 18380 10793 18408
rect 9916 18368 9922 18380
rect 10781 18377 10793 18380
rect 10827 18377 10839 18411
rect 10781 18371 10839 18377
rect 12434 18368 12440 18420
rect 12492 18408 12498 18420
rect 17957 18411 18015 18417
rect 17957 18408 17969 18411
rect 12492 18380 17969 18408
rect 12492 18368 12498 18380
rect 17957 18377 17969 18380
rect 18003 18377 18015 18411
rect 17957 18371 18015 18377
rect 18325 18411 18383 18417
rect 18325 18377 18337 18411
rect 18371 18408 18383 18411
rect 18371 18380 18662 18408
rect 18371 18377 18383 18380
rect 18325 18371 18383 18377
rect 4154 18340 4160 18352
rect 3436 18312 4160 18340
rect 3436 18281 3464 18312
rect 4154 18300 4160 18312
rect 4212 18300 4218 18352
rect 5626 18300 5632 18352
rect 5684 18340 5690 18352
rect 7653 18343 7711 18349
rect 7653 18340 7665 18343
rect 5684 18312 7665 18340
rect 5684 18300 5690 18312
rect 7653 18309 7665 18312
rect 7699 18309 7711 18343
rect 9766 18340 9772 18352
rect 7653 18303 7711 18309
rect 7760 18312 9772 18340
rect 2961 18275 3019 18281
rect 2961 18241 2973 18275
rect 3007 18241 3019 18275
rect 2961 18235 3019 18241
rect 3421 18275 3479 18281
rect 3421 18241 3433 18275
rect 3467 18241 3479 18275
rect 3421 18235 3479 18241
rect 1762 18164 1768 18216
rect 1820 18164 1826 18216
rect 2976 18136 3004 18235
rect 4062 18232 4068 18284
rect 4120 18272 4126 18284
rect 4433 18275 4491 18281
rect 4433 18272 4445 18275
rect 4120 18244 4445 18272
rect 4120 18232 4126 18244
rect 4433 18241 4445 18244
rect 4479 18241 4491 18275
rect 4433 18235 4491 18241
rect 4157 18207 4215 18213
rect 4157 18173 4169 18207
rect 4203 18204 4215 18207
rect 4246 18204 4252 18216
rect 4203 18176 4252 18204
rect 4203 18173 4215 18176
rect 4157 18167 4215 18173
rect 4246 18164 4252 18176
rect 4304 18164 4310 18216
rect 7760 18136 7788 18312
rect 9766 18300 9772 18312
rect 9824 18300 9830 18352
rect 11238 18340 11244 18352
rect 9968 18312 11244 18340
rect 9968 18281 9996 18312
rect 11238 18300 11244 18312
rect 11296 18300 11302 18352
rect 11514 18300 11520 18352
rect 11572 18340 11578 18352
rect 11572 18312 12006 18340
rect 11572 18300 11578 18312
rect 13170 18300 13176 18352
rect 13228 18300 13234 18352
rect 13906 18300 13912 18352
rect 13964 18340 13970 18352
rect 14277 18343 14335 18349
rect 14277 18340 14289 18343
rect 13964 18312 14289 18340
rect 13964 18300 13970 18312
rect 14277 18309 14289 18312
rect 14323 18309 14335 18343
rect 14277 18303 14335 18309
rect 14369 18343 14427 18349
rect 14369 18309 14381 18343
rect 14415 18340 14427 18343
rect 16758 18340 16764 18352
rect 14415 18312 16764 18340
rect 14415 18309 14427 18312
rect 14369 18303 14427 18309
rect 16758 18300 16764 18312
rect 16816 18300 16822 18352
rect 17405 18343 17463 18349
rect 17405 18309 17417 18343
rect 17451 18340 17463 18343
rect 17451 18312 18552 18340
rect 17451 18309 17463 18312
rect 17405 18303 17463 18309
rect 7837 18275 7895 18281
rect 7837 18241 7849 18275
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 9953 18275 10011 18281
rect 9953 18241 9965 18275
rect 9999 18241 10011 18275
rect 9953 18235 10011 18241
rect 10873 18275 10931 18281
rect 10873 18241 10885 18275
rect 10919 18272 10931 18275
rect 11790 18272 11796 18284
rect 10919 18244 11796 18272
rect 10919 18241 10931 18244
rect 10873 18235 10931 18241
rect 7852 18204 7880 18235
rect 11790 18232 11796 18244
rect 11848 18232 11854 18284
rect 12158 18232 12164 18284
rect 12216 18232 12222 18284
rect 13446 18232 13452 18284
rect 13504 18232 13510 18284
rect 14826 18272 14832 18284
rect 14108 18244 14832 18272
rect 7852 18176 10824 18204
rect 2976 18108 7788 18136
rect 9769 18139 9827 18145
rect 9769 18105 9781 18139
rect 9815 18136 9827 18139
rect 10042 18136 10048 18148
rect 9815 18108 10048 18136
rect 9815 18105 9827 18108
rect 9769 18099 9827 18105
rect 10042 18096 10048 18108
rect 10100 18096 10106 18148
rect 10796 18136 10824 18176
rect 10962 18164 10968 18216
rect 11020 18164 11026 18216
rect 11701 18207 11759 18213
rect 11701 18173 11713 18207
rect 11747 18204 11759 18207
rect 12176 18204 12204 18232
rect 14108 18204 14136 18244
rect 14826 18232 14832 18244
rect 14884 18272 14890 18284
rect 15105 18275 15163 18281
rect 15105 18272 15117 18275
rect 14884 18244 15117 18272
rect 14884 18232 14890 18244
rect 15105 18241 15117 18244
rect 15151 18241 15163 18275
rect 15105 18235 15163 18241
rect 16301 18275 16359 18281
rect 16301 18241 16313 18275
rect 16347 18272 16359 18275
rect 17862 18272 17868 18284
rect 16347 18244 17868 18272
rect 16347 18241 16359 18244
rect 16301 18235 16359 18241
rect 11747 18176 12112 18204
rect 12176 18176 14136 18204
rect 11747 18173 11759 18176
rect 11701 18167 11759 18173
rect 12084 18148 12112 18176
rect 14550 18164 14556 18216
rect 14608 18164 14614 18216
rect 10796 18108 11836 18136
rect 9674 18028 9680 18080
rect 9732 18068 9738 18080
rect 10413 18071 10471 18077
rect 10413 18068 10425 18071
rect 9732 18040 10425 18068
rect 9732 18028 9738 18040
rect 10413 18037 10425 18040
rect 10459 18037 10471 18071
rect 11808 18068 11836 18108
rect 12066 18096 12072 18148
rect 12124 18096 12130 18148
rect 13722 18096 13728 18148
rect 13780 18136 13786 18148
rect 13909 18139 13967 18145
rect 13909 18136 13921 18139
rect 13780 18108 13921 18136
rect 13780 18096 13786 18108
rect 13909 18105 13921 18108
rect 13955 18105 13967 18139
rect 15120 18136 15148 18235
rect 17862 18232 17868 18244
rect 17920 18232 17926 18284
rect 15657 18207 15715 18213
rect 15657 18173 15669 18207
rect 15703 18204 15715 18207
rect 16482 18204 16488 18216
rect 15703 18176 16488 18204
rect 15703 18173 15715 18176
rect 15657 18167 15715 18173
rect 16482 18164 16488 18176
rect 16540 18164 16546 18216
rect 18417 18207 18475 18213
rect 18417 18204 18429 18207
rect 18340 18176 18429 18204
rect 15120 18108 15240 18136
rect 13909 18099 13967 18105
rect 13630 18068 13636 18080
rect 11808 18040 13636 18068
rect 10413 18031 10471 18037
rect 13630 18028 13636 18040
rect 13688 18028 13694 18080
rect 15013 18071 15071 18077
rect 15013 18037 15025 18071
rect 15059 18068 15071 18071
rect 15102 18068 15108 18080
rect 15059 18040 15108 18068
rect 15059 18037 15071 18040
rect 15013 18031 15071 18037
rect 15102 18028 15108 18040
rect 15160 18028 15166 18080
rect 15212 18068 15240 18108
rect 15286 18096 15292 18148
rect 15344 18136 15350 18148
rect 16117 18139 16175 18145
rect 16117 18136 16129 18139
rect 15344 18108 16129 18136
rect 15344 18096 15350 18108
rect 16117 18105 16129 18108
rect 16163 18105 16175 18139
rect 17221 18139 17279 18145
rect 17221 18136 17233 18139
rect 16117 18099 16175 18105
rect 16224 18108 17233 18136
rect 16224 18068 16252 18108
rect 17221 18105 17233 18108
rect 17267 18105 17279 18139
rect 17221 18099 17279 18105
rect 15212 18040 16252 18068
rect 16298 18028 16304 18080
rect 16356 18068 16362 18080
rect 16669 18071 16727 18077
rect 16669 18068 16681 18071
rect 16356 18040 16681 18068
rect 16356 18028 16362 18040
rect 16669 18037 16681 18040
rect 16715 18037 16727 18071
rect 16669 18031 16727 18037
rect 16942 18028 16948 18080
rect 17000 18028 17006 18080
rect 18340 18068 18368 18176
rect 18417 18173 18429 18176
rect 18463 18173 18475 18207
rect 18417 18167 18475 18173
rect 18524 18136 18552 18312
rect 18634 18272 18662 18380
rect 18690 18368 18696 18420
rect 18748 18408 18754 18420
rect 19061 18411 19119 18417
rect 19061 18408 19073 18411
rect 18748 18380 19073 18408
rect 18748 18368 18754 18380
rect 19061 18377 19073 18380
rect 19107 18408 19119 18411
rect 22465 18411 22523 18417
rect 19107 18380 22094 18408
rect 19107 18377 19119 18380
rect 19061 18371 19119 18377
rect 19150 18300 19156 18352
rect 19208 18340 19214 18352
rect 19889 18343 19947 18349
rect 19889 18340 19901 18343
rect 19208 18312 19901 18340
rect 19208 18300 19214 18312
rect 19889 18309 19901 18312
rect 19935 18309 19947 18343
rect 21174 18340 21180 18352
rect 21114 18312 21180 18340
rect 19889 18303 19947 18309
rect 21174 18300 21180 18312
rect 21232 18340 21238 18352
rect 21634 18340 21640 18352
rect 21232 18312 21640 18340
rect 21232 18300 21238 18312
rect 21634 18300 21640 18312
rect 21692 18300 21698 18352
rect 22066 18340 22094 18380
rect 22465 18377 22477 18411
rect 22511 18408 22523 18411
rect 25774 18408 25780 18420
rect 22511 18380 25780 18408
rect 22511 18377 22523 18380
rect 22465 18371 22523 18377
rect 25774 18368 25780 18380
rect 25832 18368 25838 18420
rect 26237 18411 26295 18417
rect 26237 18377 26249 18411
rect 26283 18408 26295 18411
rect 27246 18408 27252 18420
rect 26283 18380 27252 18408
rect 26283 18377 26295 18380
rect 26237 18371 26295 18377
rect 27246 18368 27252 18380
rect 27304 18368 27310 18420
rect 27617 18411 27675 18417
rect 27617 18377 27629 18411
rect 27663 18408 27675 18411
rect 27706 18408 27712 18420
rect 27663 18380 27712 18408
rect 27663 18377 27675 18380
rect 27617 18371 27675 18377
rect 27706 18368 27712 18380
rect 27764 18368 27770 18420
rect 28721 18411 28779 18417
rect 28721 18377 28733 18411
rect 28767 18408 28779 18411
rect 29730 18408 29736 18420
rect 28767 18380 29736 18408
rect 28767 18377 28779 18380
rect 28721 18371 28779 18377
rect 29730 18368 29736 18380
rect 29788 18368 29794 18420
rect 30837 18411 30895 18417
rect 30837 18377 30849 18411
rect 30883 18408 30895 18411
rect 31202 18408 31208 18420
rect 30883 18380 31208 18408
rect 30883 18377 30895 18380
rect 30837 18371 30895 18377
rect 31202 18368 31208 18380
rect 31260 18368 31266 18420
rect 33045 18411 33103 18417
rect 33045 18377 33057 18411
rect 33091 18408 33103 18411
rect 35526 18408 35532 18420
rect 33091 18380 35532 18408
rect 33091 18377 33103 18380
rect 33045 18371 33103 18377
rect 35526 18368 35532 18380
rect 35584 18368 35590 18420
rect 36906 18368 36912 18420
rect 36964 18368 36970 18420
rect 37366 18368 37372 18420
rect 37424 18408 37430 18420
rect 37461 18411 37519 18417
rect 37461 18408 37473 18411
rect 37424 18380 37473 18408
rect 37424 18368 37430 18380
rect 37461 18377 37473 18380
rect 37507 18377 37519 18411
rect 37461 18371 37519 18377
rect 38194 18368 38200 18420
rect 38252 18408 38258 18420
rect 40405 18411 40463 18417
rect 40405 18408 40417 18411
rect 38252 18380 40417 18408
rect 38252 18368 38258 18380
rect 40405 18377 40417 18380
rect 40451 18377 40463 18411
rect 40405 18371 40463 18377
rect 40770 18368 40776 18420
rect 40828 18408 40834 18420
rect 40865 18411 40923 18417
rect 40865 18408 40877 18411
rect 40828 18380 40877 18408
rect 40828 18368 40834 18380
rect 40865 18377 40877 18380
rect 40911 18377 40923 18411
rect 40865 18371 40923 18377
rect 48774 18368 48780 18420
rect 48832 18368 48838 18420
rect 22646 18340 22652 18352
rect 22066 18312 22652 18340
rect 22646 18300 22652 18312
rect 22704 18340 22710 18352
rect 23290 18340 23296 18352
rect 22704 18312 23296 18340
rect 22704 18300 22710 18312
rect 23290 18300 23296 18312
rect 23348 18300 23354 18352
rect 24118 18300 24124 18352
rect 24176 18300 24182 18352
rect 24762 18300 24768 18352
rect 24820 18340 24826 18352
rect 25133 18343 25191 18349
rect 25133 18340 25145 18343
rect 24820 18312 25145 18340
rect 24820 18300 24826 18312
rect 25133 18309 25145 18312
rect 25179 18309 25191 18343
rect 25133 18303 25191 18309
rect 25222 18300 25228 18352
rect 25280 18300 25286 18352
rect 28813 18343 28871 18349
rect 28813 18309 28825 18343
rect 28859 18340 28871 18343
rect 32122 18340 32128 18352
rect 28859 18312 32128 18340
rect 28859 18309 28871 18312
rect 28813 18303 28871 18309
rect 32122 18300 32128 18312
rect 32180 18300 32186 18352
rect 33594 18340 33600 18352
rect 33520 18312 33600 18340
rect 19426 18272 19432 18284
rect 18634 18244 19432 18272
rect 19426 18232 19432 18244
rect 19484 18232 19490 18284
rect 22557 18275 22615 18281
rect 22557 18241 22569 18275
rect 22603 18272 22615 18275
rect 23106 18272 23112 18284
rect 22603 18244 23112 18272
rect 22603 18241 22615 18244
rect 22557 18235 22615 18241
rect 23106 18232 23112 18244
rect 23164 18232 23170 18284
rect 25038 18232 25044 18284
rect 25096 18232 25102 18284
rect 18601 18207 18659 18213
rect 18601 18173 18613 18207
rect 18647 18204 18659 18207
rect 19150 18204 19156 18216
rect 18647 18176 19156 18204
rect 18647 18173 18659 18176
rect 18601 18167 18659 18173
rect 19150 18164 19156 18176
rect 19208 18164 19214 18216
rect 19337 18207 19395 18213
rect 19337 18173 19349 18207
rect 19383 18204 19395 18207
rect 19610 18204 19616 18216
rect 19383 18176 19616 18204
rect 19383 18173 19395 18176
rect 19337 18167 19395 18173
rect 19610 18164 19616 18176
rect 19668 18164 19674 18216
rect 21542 18204 21548 18216
rect 19720 18176 21548 18204
rect 19720 18136 19748 18176
rect 21542 18164 21548 18176
rect 21600 18164 21606 18216
rect 25240 18213 25268 18300
rect 26326 18232 26332 18284
rect 26384 18232 26390 18284
rect 27525 18275 27583 18281
rect 27525 18241 27537 18275
rect 27571 18272 27583 18275
rect 29086 18272 29092 18284
rect 27571 18244 29092 18272
rect 27571 18241 27583 18244
rect 27525 18235 27583 18241
rect 29086 18232 29092 18244
rect 29144 18232 29150 18284
rect 29362 18232 29368 18284
rect 29420 18272 29426 18284
rect 30377 18275 30435 18281
rect 30377 18272 30389 18275
rect 29420 18244 30389 18272
rect 29420 18232 29426 18244
rect 30377 18241 30389 18244
rect 30423 18241 30435 18275
rect 30377 18235 30435 18241
rect 30469 18275 30527 18281
rect 30469 18241 30481 18275
rect 30515 18272 30527 18275
rect 31297 18275 31355 18281
rect 31297 18272 31309 18275
rect 30515 18244 31309 18272
rect 30515 18241 30527 18244
rect 30469 18235 30527 18241
rect 31297 18241 31309 18244
rect 31343 18241 31355 18275
rect 32585 18275 32643 18281
rect 32585 18272 32597 18275
rect 31297 18235 31355 18241
rect 31404 18244 32597 18272
rect 22649 18207 22707 18213
rect 22649 18204 22661 18207
rect 22204 18176 22661 18204
rect 22097 18139 22155 18145
rect 22097 18136 22109 18139
rect 18524 18108 19748 18136
rect 20916 18108 22109 18136
rect 20916 18068 20944 18108
rect 22097 18105 22109 18108
rect 22143 18105 22155 18139
rect 22097 18099 22155 18105
rect 18340 18040 20944 18068
rect 21266 18028 21272 18080
rect 21324 18068 21330 18080
rect 21361 18071 21419 18077
rect 21361 18068 21373 18071
rect 21324 18040 21373 18068
rect 21324 18028 21330 18040
rect 21361 18037 21373 18040
rect 21407 18037 21419 18071
rect 21361 18031 21419 18037
rect 21450 18028 21456 18080
rect 21508 18068 21514 18080
rect 22204 18068 22232 18176
rect 22649 18173 22661 18176
rect 22695 18173 22707 18207
rect 22649 18167 22707 18173
rect 25225 18207 25283 18213
rect 25225 18173 25237 18207
rect 25271 18173 25283 18207
rect 25225 18167 25283 18173
rect 26510 18164 26516 18216
rect 26568 18164 26574 18216
rect 26602 18164 26608 18216
rect 26660 18204 26666 18216
rect 27709 18207 27767 18213
rect 27709 18204 27721 18207
rect 26660 18176 27721 18204
rect 26660 18164 26666 18176
rect 27709 18173 27721 18176
rect 27755 18173 27767 18207
rect 28905 18207 28963 18213
rect 28905 18204 28917 18207
rect 27709 18167 27767 18173
rect 28460 18176 28917 18204
rect 23750 18096 23756 18148
rect 23808 18136 23814 18148
rect 24673 18139 24731 18145
rect 24673 18136 24685 18139
rect 23808 18108 24685 18136
rect 23808 18096 23814 18108
rect 24673 18105 24685 18108
rect 24719 18105 24731 18139
rect 24673 18099 24731 18105
rect 26050 18096 26056 18148
rect 26108 18136 26114 18148
rect 28353 18139 28411 18145
rect 28353 18136 28365 18139
rect 26108 18108 28365 18136
rect 26108 18096 26114 18108
rect 28353 18105 28365 18108
rect 28399 18105 28411 18139
rect 28353 18099 28411 18105
rect 21508 18040 22232 18068
rect 21508 18028 21514 18040
rect 25038 18028 25044 18080
rect 25096 18068 25102 18080
rect 25869 18071 25927 18077
rect 25869 18068 25881 18071
rect 25096 18040 25881 18068
rect 25096 18028 25102 18040
rect 25869 18037 25881 18040
rect 25915 18037 25927 18071
rect 25869 18031 25927 18037
rect 27154 18028 27160 18080
rect 27212 18028 27218 18080
rect 27522 18028 27528 18080
rect 27580 18068 27586 18080
rect 28460 18068 28488 18176
rect 28905 18173 28917 18176
rect 28951 18173 28963 18207
rect 28905 18167 28963 18173
rect 30098 18164 30104 18216
rect 30156 18204 30162 18216
rect 30193 18207 30251 18213
rect 30193 18204 30205 18207
rect 30156 18176 30205 18204
rect 30156 18164 30162 18176
rect 30193 18173 30205 18176
rect 30239 18173 30251 18207
rect 31404 18204 31432 18244
rect 32585 18241 32597 18244
rect 32631 18241 32643 18275
rect 32585 18235 32643 18241
rect 32674 18232 32680 18284
rect 32732 18232 32738 18284
rect 30193 18167 30251 18173
rect 30300 18176 31432 18204
rect 28534 18096 28540 18148
rect 28592 18136 28598 18148
rect 30300 18136 30328 18176
rect 31938 18164 31944 18216
rect 31996 18204 32002 18216
rect 32401 18207 32459 18213
rect 32401 18204 32413 18207
rect 31996 18176 32413 18204
rect 31996 18164 32002 18176
rect 32401 18173 32413 18176
rect 32447 18204 32459 18207
rect 33520 18204 33548 18312
rect 33594 18300 33600 18312
rect 33652 18300 33658 18352
rect 34330 18300 34336 18352
rect 34388 18300 34394 18352
rect 36998 18300 37004 18352
rect 37056 18340 37062 18352
rect 37734 18340 37740 18352
rect 37056 18312 37740 18340
rect 37056 18300 37062 18312
rect 37734 18300 37740 18312
rect 37792 18300 37798 18352
rect 38746 18300 38752 18352
rect 38804 18300 38810 18352
rect 40034 18300 40040 18352
rect 40092 18340 40098 18352
rect 40129 18343 40187 18349
rect 40129 18340 40141 18343
rect 40092 18312 40141 18340
rect 40092 18300 40098 18312
rect 40129 18309 40141 18312
rect 40175 18340 40187 18343
rect 41046 18340 41052 18352
rect 40175 18312 41052 18340
rect 40175 18309 40187 18312
rect 40129 18303 40187 18309
rect 41046 18300 41052 18312
rect 41104 18300 41110 18352
rect 35710 18232 35716 18284
rect 35768 18272 35774 18284
rect 36265 18275 36323 18281
rect 36265 18272 36277 18275
rect 35768 18244 36277 18272
rect 35768 18232 35774 18244
rect 36265 18241 36277 18244
rect 36311 18241 36323 18275
rect 36265 18235 36323 18241
rect 36354 18232 36360 18284
rect 36412 18232 36418 18284
rect 37108 18244 37412 18272
rect 32447 18176 33548 18204
rect 32447 18173 32459 18176
rect 32401 18167 32459 18173
rect 33594 18164 33600 18216
rect 33652 18164 33658 18216
rect 33873 18207 33931 18213
rect 33873 18173 33885 18207
rect 33919 18204 33931 18207
rect 34606 18204 34612 18216
rect 33919 18176 34612 18204
rect 33919 18173 33931 18176
rect 33873 18167 33931 18173
rect 34606 18164 34612 18176
rect 34664 18204 34670 18216
rect 36446 18204 36452 18216
rect 34664 18176 36452 18204
rect 34664 18164 34670 18176
rect 36446 18164 36452 18176
rect 36504 18164 36510 18216
rect 36541 18207 36599 18213
rect 36541 18173 36553 18207
rect 36587 18204 36599 18207
rect 37108 18204 37136 18244
rect 36587 18176 37136 18204
rect 36587 18173 36599 18176
rect 36541 18167 36599 18173
rect 37274 18164 37280 18216
rect 37332 18164 37338 18216
rect 37384 18204 37412 18244
rect 37458 18232 37464 18284
rect 37516 18272 37522 18284
rect 38010 18272 38016 18284
rect 37516 18244 38016 18272
rect 37516 18232 37522 18244
rect 38010 18232 38016 18244
rect 38068 18232 38074 18284
rect 39758 18232 39764 18284
rect 39816 18232 39822 18284
rect 40773 18275 40831 18281
rect 40773 18241 40785 18275
rect 40819 18272 40831 18275
rect 48406 18272 48412 18284
rect 40819 18244 48412 18272
rect 40819 18241 40831 18244
rect 40773 18235 40831 18241
rect 48406 18232 48412 18244
rect 48464 18232 48470 18284
rect 48593 18275 48651 18281
rect 48593 18241 48605 18275
rect 48639 18272 48651 18275
rect 49326 18272 49332 18284
rect 48639 18244 49332 18272
rect 48639 18241 48651 18244
rect 48593 18235 48651 18241
rect 49326 18232 49332 18244
rect 49384 18232 49390 18284
rect 37734 18204 37740 18216
rect 37384 18176 37740 18204
rect 37734 18164 37740 18176
rect 37792 18164 37798 18216
rect 37826 18164 37832 18216
rect 37884 18204 37890 18216
rect 39485 18207 39543 18213
rect 39485 18204 39497 18207
rect 37884 18176 39497 18204
rect 37884 18164 37890 18176
rect 39485 18173 39497 18176
rect 39531 18204 39543 18207
rect 40957 18207 41015 18213
rect 40957 18204 40969 18207
rect 39531 18176 40969 18204
rect 39531 18173 39543 18176
rect 39485 18167 39543 18173
rect 40957 18173 40969 18176
rect 41003 18173 41015 18207
rect 40957 18167 41015 18173
rect 28592 18108 30328 18136
rect 28592 18096 28598 18108
rect 31018 18096 31024 18148
rect 31076 18136 31082 18148
rect 35897 18139 35955 18145
rect 35897 18136 35909 18139
rect 31076 18108 33732 18136
rect 31076 18096 31082 18108
rect 27580 18040 28488 18068
rect 27580 18028 27586 18040
rect 29362 18028 29368 18080
rect 29420 18068 29426 18080
rect 29733 18071 29791 18077
rect 29733 18068 29745 18071
rect 29420 18040 29745 18068
rect 29420 18028 29426 18040
rect 29733 18037 29745 18040
rect 29779 18037 29791 18071
rect 29733 18031 29791 18037
rect 30098 18028 30104 18080
rect 30156 18068 30162 18080
rect 32582 18068 32588 18080
rect 30156 18040 32588 18068
rect 30156 18028 30162 18040
rect 32582 18028 32588 18040
rect 32640 18028 32646 18080
rect 33704 18068 33732 18108
rect 34900 18108 35909 18136
rect 34900 18068 34928 18108
rect 35897 18105 35909 18108
rect 35943 18105 35955 18139
rect 35897 18099 35955 18105
rect 38010 18096 38016 18148
rect 38068 18096 38074 18148
rect 33704 18040 34928 18068
rect 35345 18071 35403 18077
rect 35345 18037 35357 18071
rect 35391 18068 35403 18071
rect 35618 18068 35624 18080
rect 35391 18040 35624 18068
rect 35391 18037 35403 18040
rect 35345 18031 35403 18037
rect 35618 18028 35624 18040
rect 35676 18028 35682 18080
rect 36354 18028 36360 18080
rect 36412 18068 36418 18080
rect 37090 18068 37096 18080
rect 36412 18040 37096 18068
rect 36412 18028 36418 18040
rect 37090 18028 37096 18040
rect 37148 18028 37154 18080
rect 37274 18028 37280 18080
rect 37332 18068 37338 18080
rect 37645 18071 37703 18077
rect 37645 18068 37657 18071
rect 37332 18040 37657 18068
rect 37332 18028 37338 18040
rect 37645 18037 37657 18040
rect 37691 18037 37703 18071
rect 38028 18068 38056 18096
rect 40218 18068 40224 18080
rect 38028 18040 40224 18068
rect 37645 18031 37703 18037
rect 40218 18028 40224 18040
rect 40276 18028 40282 18080
rect 48314 18028 48320 18080
rect 48372 18068 48378 18080
rect 49145 18071 49203 18077
rect 49145 18068 49157 18071
rect 48372 18040 49157 18068
rect 48372 18028 48378 18040
rect 49145 18037 49157 18040
rect 49191 18037 49203 18071
rect 49145 18031 49203 18037
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 10134 17824 10140 17876
rect 10192 17824 10198 17876
rect 10597 17867 10655 17873
rect 10597 17833 10609 17867
rect 10643 17864 10655 17867
rect 10962 17864 10968 17876
rect 10643 17836 10968 17864
rect 10643 17833 10655 17836
rect 10597 17827 10655 17833
rect 10962 17824 10968 17836
rect 11020 17824 11026 17876
rect 12342 17864 12348 17876
rect 11072 17836 12348 17864
rect 9858 17756 9864 17808
rect 9916 17796 9922 17808
rect 11072 17796 11100 17836
rect 12342 17824 12348 17836
rect 12400 17824 12406 17876
rect 12618 17824 12624 17876
rect 12676 17864 12682 17876
rect 12897 17867 12955 17873
rect 12897 17864 12909 17867
rect 12676 17836 12909 17864
rect 12676 17824 12682 17836
rect 12897 17833 12909 17836
rect 12943 17833 12955 17867
rect 12897 17827 12955 17833
rect 14277 17867 14335 17873
rect 14277 17833 14289 17867
rect 14323 17864 14335 17867
rect 14550 17864 14556 17876
rect 14323 17836 14556 17864
rect 14323 17833 14335 17836
rect 14277 17827 14335 17833
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 15194 17824 15200 17876
rect 15252 17864 15258 17876
rect 15746 17864 15752 17876
rect 15252 17836 15752 17864
rect 15252 17824 15258 17836
rect 15746 17824 15752 17836
rect 15804 17824 15810 17876
rect 17218 17824 17224 17876
rect 17276 17864 17282 17876
rect 17497 17867 17555 17873
rect 17497 17864 17509 17867
rect 17276 17836 17509 17864
rect 17276 17824 17282 17836
rect 17497 17833 17509 17836
rect 17543 17833 17555 17867
rect 17497 17827 17555 17833
rect 19334 17824 19340 17876
rect 19392 17864 19398 17876
rect 19429 17867 19487 17873
rect 19429 17864 19441 17867
rect 19392 17836 19441 17864
rect 19392 17824 19398 17836
rect 19429 17833 19441 17836
rect 19475 17833 19487 17867
rect 19429 17827 19487 17833
rect 19610 17824 19616 17876
rect 19668 17864 19674 17876
rect 21358 17864 21364 17876
rect 19668 17836 21364 17864
rect 19668 17824 19674 17836
rect 21358 17824 21364 17836
rect 21416 17824 21422 17876
rect 21542 17824 21548 17876
rect 21600 17864 21606 17876
rect 24581 17867 24639 17873
rect 24581 17864 24593 17867
rect 21600 17836 24593 17864
rect 21600 17824 21606 17836
rect 24581 17833 24593 17836
rect 24627 17833 24639 17867
rect 30926 17864 30932 17876
rect 24581 17827 24639 17833
rect 25976 17836 30932 17864
rect 20714 17796 20720 17808
rect 9916 17768 11100 17796
rect 16408 17768 20720 17796
rect 9916 17756 9922 17768
rect 10321 17731 10379 17737
rect 10321 17697 10333 17731
rect 10367 17728 10379 17731
rect 11422 17728 11428 17740
rect 10367 17700 11428 17728
rect 10367 17697 10379 17700
rect 10321 17691 10379 17697
rect 11422 17688 11428 17700
rect 11480 17688 11486 17740
rect 12345 17731 12403 17737
rect 12345 17697 12357 17731
rect 12391 17728 12403 17731
rect 12526 17728 12532 17740
rect 12391 17700 12532 17728
rect 12391 17697 12403 17700
rect 12345 17691 12403 17697
rect 12526 17688 12532 17700
rect 12584 17728 12590 17740
rect 13446 17728 13452 17740
rect 12584 17700 13452 17728
rect 12584 17688 12590 17700
rect 13446 17688 13452 17700
rect 13504 17688 13510 17740
rect 14734 17728 14740 17740
rect 13648 17700 14740 17728
rect 2961 17663 3019 17669
rect 2961 17629 2973 17663
rect 3007 17660 3019 17663
rect 10226 17660 10232 17672
rect 3007 17632 10232 17660
rect 3007 17629 3019 17632
rect 2961 17623 3019 17629
rect 10226 17620 10232 17632
rect 10284 17620 10290 17672
rect 13081 17663 13139 17669
rect 13081 17629 13093 17663
rect 13127 17660 13139 17663
rect 13354 17660 13360 17672
rect 13127 17632 13360 17660
rect 13127 17629 13139 17632
rect 13081 17623 13139 17629
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 934 17552 940 17604
rect 992 17592 998 17604
rect 1765 17595 1823 17601
rect 1765 17592 1777 17595
rect 992 17564 1777 17592
rect 992 17552 998 17564
rect 1765 17561 1777 17564
rect 1811 17561 1823 17595
rect 1765 17555 1823 17561
rect 10134 17552 10140 17604
rect 10192 17592 10198 17604
rect 10192 17564 10902 17592
rect 10192 17552 10198 17564
rect 10796 17524 10824 17564
rect 12066 17552 12072 17604
rect 12124 17552 12130 17604
rect 13648 17592 13676 17700
rect 13725 17663 13783 17669
rect 13725 17629 13737 17663
rect 13771 17629 13783 17663
rect 14660 17646 14688 17700
rect 14734 17688 14740 17700
rect 14792 17688 14798 17740
rect 15378 17688 15384 17740
rect 15436 17728 15442 17740
rect 16022 17728 16028 17740
rect 15436 17700 16028 17728
rect 15436 17688 15442 17700
rect 16022 17688 16028 17700
rect 16080 17688 16086 17740
rect 13725 17623 13783 17629
rect 13464 17564 13676 17592
rect 11146 17524 11152 17536
rect 10796 17496 11152 17524
rect 11146 17484 11152 17496
rect 11204 17524 11210 17536
rect 13464 17524 13492 17564
rect 11204 17496 13492 17524
rect 13541 17527 13599 17533
rect 11204 17484 11210 17496
rect 13541 17493 13553 17527
rect 13587 17524 13599 17527
rect 13630 17524 13636 17536
rect 13587 17496 13636 17524
rect 13587 17493 13599 17496
rect 13541 17487 13599 17493
rect 13630 17484 13636 17496
rect 13688 17484 13694 17536
rect 13740 17524 13768 17623
rect 15749 17595 15807 17601
rect 15749 17561 15761 17595
rect 15795 17592 15807 17595
rect 16206 17592 16212 17604
rect 15795 17564 16212 17592
rect 15795 17561 15807 17564
rect 15749 17555 15807 17561
rect 16206 17552 16212 17564
rect 16264 17552 16270 17604
rect 16408 17524 16436 17768
rect 20714 17756 20720 17768
rect 20772 17756 20778 17808
rect 22278 17756 22284 17808
rect 22336 17796 22342 17808
rect 23293 17799 23351 17805
rect 23293 17796 23305 17799
rect 22336 17768 23305 17796
rect 22336 17756 22342 17768
rect 23293 17765 23305 17768
rect 23339 17765 23351 17799
rect 23293 17759 23351 17765
rect 23566 17756 23572 17808
rect 23624 17796 23630 17808
rect 25777 17799 25835 17805
rect 25777 17796 25789 17799
rect 23624 17768 25789 17796
rect 23624 17756 23630 17768
rect 25777 17765 25789 17768
rect 25823 17765 25835 17799
rect 25777 17759 25835 17765
rect 16850 17688 16856 17740
rect 16908 17688 16914 17740
rect 16942 17688 16948 17740
rect 17000 17728 17006 17740
rect 18785 17731 18843 17737
rect 18785 17728 18797 17731
rect 17000 17700 18797 17728
rect 17000 17688 17006 17700
rect 18785 17697 18797 17700
rect 18831 17728 18843 17731
rect 19702 17728 19708 17740
rect 18831 17700 19708 17728
rect 18831 17697 18843 17700
rect 18785 17691 18843 17697
rect 19702 17688 19708 17700
rect 19760 17688 19766 17740
rect 20257 17731 20315 17737
rect 20257 17697 20269 17731
rect 20303 17728 20315 17731
rect 20346 17728 20352 17740
rect 20303 17700 20352 17728
rect 20303 17697 20315 17700
rect 20257 17691 20315 17697
rect 20346 17688 20352 17700
rect 20404 17688 20410 17740
rect 21726 17688 21732 17740
rect 21784 17688 21790 17740
rect 22005 17731 22063 17737
rect 22005 17697 22017 17731
rect 22051 17728 22063 17731
rect 22094 17728 22100 17740
rect 22051 17700 22100 17728
rect 22051 17697 22063 17700
rect 22005 17691 22063 17697
rect 22094 17688 22100 17700
rect 22152 17688 22158 17740
rect 23937 17731 23995 17737
rect 23937 17697 23949 17731
rect 23983 17728 23995 17731
rect 24946 17728 24952 17740
rect 23983 17700 24952 17728
rect 23983 17697 23995 17700
rect 23937 17691 23995 17697
rect 24946 17688 24952 17700
rect 25004 17688 25010 17740
rect 25038 17688 25044 17740
rect 25096 17688 25102 17740
rect 25133 17731 25191 17737
rect 25133 17697 25145 17731
rect 25179 17697 25191 17731
rect 25133 17691 25191 17697
rect 16482 17620 16488 17672
rect 16540 17660 16546 17672
rect 17129 17663 17187 17669
rect 17129 17660 17141 17663
rect 16540 17632 17141 17660
rect 16540 17620 16546 17632
rect 17129 17629 17141 17632
rect 17175 17629 17187 17663
rect 17129 17623 17187 17629
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17660 19671 17663
rect 19659 17632 20484 17660
rect 19659 17629 19671 17632
rect 19613 17623 19671 17629
rect 17957 17595 18015 17601
rect 17957 17561 17969 17595
rect 18003 17592 18015 17595
rect 18598 17592 18604 17604
rect 18003 17564 18604 17592
rect 18003 17561 18015 17564
rect 17957 17555 18015 17561
rect 18598 17552 18604 17564
rect 18656 17552 18662 17604
rect 13740 17496 16436 17524
rect 16482 17484 16488 17536
rect 16540 17484 16546 17536
rect 17037 17527 17095 17533
rect 17037 17493 17049 17527
rect 17083 17524 17095 17527
rect 17402 17524 17408 17536
rect 17083 17496 17408 17524
rect 17083 17493 17095 17496
rect 17037 17487 17095 17493
rect 17402 17484 17408 17496
rect 17460 17484 17466 17536
rect 18874 17484 18880 17536
rect 18932 17524 18938 17536
rect 20346 17524 20352 17536
rect 18932 17496 20352 17524
rect 18932 17484 18938 17496
rect 20346 17484 20352 17496
rect 20404 17484 20410 17536
rect 20456 17524 20484 17632
rect 23474 17620 23480 17672
rect 23532 17660 23538 17672
rect 25148 17660 25176 17691
rect 25976 17669 26004 17836
rect 30926 17824 30932 17836
rect 30984 17824 30990 17876
rect 31386 17824 31392 17876
rect 31444 17864 31450 17876
rect 33505 17867 33563 17873
rect 31444 17836 31616 17864
rect 31444 17824 31450 17836
rect 26326 17756 26332 17808
rect 26384 17756 26390 17808
rect 29641 17799 29699 17805
rect 29641 17765 29653 17799
rect 29687 17796 29699 17799
rect 29822 17796 29828 17808
rect 29687 17768 29828 17796
rect 29687 17765 29699 17768
rect 29641 17759 29699 17765
rect 29822 17756 29828 17768
rect 29880 17756 29886 17808
rect 26418 17688 26424 17740
rect 26476 17728 26482 17740
rect 31386 17728 31392 17740
rect 26476 17700 31392 17728
rect 26476 17688 26482 17700
rect 31386 17688 31392 17700
rect 31444 17688 31450 17740
rect 31478 17688 31484 17740
rect 31536 17688 31542 17740
rect 23532 17632 25176 17660
rect 25961 17663 26019 17669
rect 23532 17620 23538 17632
rect 25961 17629 25973 17663
rect 26007 17629 26019 17663
rect 25961 17623 26019 17629
rect 27430 17620 27436 17672
rect 27488 17620 27494 17672
rect 28813 17663 28871 17669
rect 28813 17629 28825 17663
rect 28859 17660 28871 17663
rect 28902 17660 28908 17672
rect 28859 17632 28908 17660
rect 28859 17629 28871 17632
rect 28813 17623 28871 17629
rect 28902 17620 28908 17632
rect 28960 17660 28966 17672
rect 31588 17660 31616 17836
rect 33505 17833 33517 17867
rect 33551 17864 33563 17867
rect 33686 17864 33692 17876
rect 33551 17836 33692 17864
rect 33551 17833 33563 17836
rect 33505 17827 33563 17833
rect 33686 17824 33692 17836
rect 33744 17824 33750 17876
rect 33870 17824 33876 17876
rect 33928 17864 33934 17876
rect 33928 17836 37504 17864
rect 33928 17824 33934 17836
rect 32858 17756 32864 17808
rect 32916 17796 32922 17808
rect 34241 17799 34299 17805
rect 34241 17796 34253 17799
rect 32916 17768 34253 17796
rect 32916 17756 32922 17768
rect 34241 17765 34253 17768
rect 34287 17796 34299 17799
rect 34330 17796 34336 17808
rect 34287 17768 34336 17796
rect 34287 17765 34299 17768
rect 34241 17759 34299 17765
rect 34330 17756 34336 17768
rect 34388 17796 34394 17808
rect 37476 17796 37504 17836
rect 38470 17824 38476 17876
rect 38528 17864 38534 17876
rect 40497 17867 40555 17873
rect 40497 17864 40509 17867
rect 38528 17836 40509 17864
rect 38528 17824 38534 17836
rect 40497 17833 40509 17836
rect 40543 17833 40555 17867
rect 40497 17827 40555 17833
rect 38749 17799 38807 17805
rect 34388 17768 36216 17796
rect 37476 17768 38654 17796
rect 34388 17756 34394 17768
rect 32950 17688 32956 17740
rect 33008 17688 33014 17740
rect 33045 17731 33103 17737
rect 33045 17697 33057 17731
rect 33091 17728 33103 17731
rect 33502 17728 33508 17740
rect 33091 17700 33508 17728
rect 33091 17697 33103 17700
rect 33045 17691 33103 17697
rect 33502 17688 33508 17700
rect 33560 17688 33566 17740
rect 34606 17688 34612 17740
rect 34664 17728 34670 17740
rect 35805 17731 35863 17737
rect 35805 17728 35817 17731
rect 34664 17700 35817 17728
rect 34664 17688 34670 17700
rect 35805 17697 35817 17700
rect 35851 17697 35863 17731
rect 35805 17691 35863 17697
rect 36188 17728 36216 17768
rect 36722 17728 36728 17740
rect 36188 17700 36728 17728
rect 31665 17663 31723 17669
rect 31665 17660 31677 17663
rect 28960 17632 30788 17660
rect 31588 17632 31677 17660
rect 28960 17620 28966 17632
rect 21634 17592 21640 17604
rect 21298 17564 21640 17592
rect 21634 17552 21640 17564
rect 21692 17552 21698 17604
rect 21818 17552 21824 17604
rect 21876 17592 21882 17604
rect 22281 17595 22339 17601
rect 22281 17592 22293 17595
rect 21876 17564 22293 17592
rect 21876 17552 21882 17564
rect 22281 17561 22293 17564
rect 22327 17561 22339 17595
rect 22281 17555 22339 17561
rect 22833 17595 22891 17601
rect 22833 17561 22845 17595
rect 22879 17592 22891 17595
rect 23661 17595 23719 17601
rect 23661 17592 23673 17595
rect 22879 17564 23673 17592
rect 22879 17561 22891 17564
rect 22833 17555 22891 17561
rect 23661 17561 23673 17564
rect 23707 17561 23719 17595
rect 23661 17555 23719 17561
rect 24486 17552 24492 17604
rect 24544 17592 24550 17604
rect 26510 17592 26516 17604
rect 24544 17564 26516 17592
rect 24544 17552 24550 17564
rect 26510 17552 26516 17564
rect 26568 17552 26574 17604
rect 28537 17595 28595 17601
rect 28537 17561 28549 17595
rect 28583 17561 28595 17595
rect 28537 17555 28595 17561
rect 22186 17524 22192 17536
rect 20456 17496 22192 17524
rect 22186 17484 22192 17496
rect 22244 17484 22250 17536
rect 23750 17484 23756 17536
rect 23808 17484 23814 17536
rect 24670 17484 24676 17536
rect 24728 17524 24734 17536
rect 24949 17527 25007 17533
rect 24949 17524 24961 17527
rect 24728 17496 24961 17524
rect 24728 17484 24734 17496
rect 24949 17493 24961 17496
rect 24995 17493 25007 17527
rect 24949 17487 25007 17493
rect 25038 17484 25044 17536
rect 25096 17524 25102 17536
rect 26421 17527 26479 17533
rect 26421 17524 26433 17527
rect 25096 17496 26433 17524
rect 25096 17484 25102 17496
rect 26421 17493 26433 17496
rect 26467 17524 26479 17527
rect 26970 17524 26976 17536
rect 26467 17496 26976 17524
rect 26467 17493 26479 17496
rect 26421 17487 26479 17493
rect 26970 17484 26976 17496
rect 27028 17484 27034 17536
rect 27062 17484 27068 17536
rect 27120 17524 27126 17536
rect 27522 17524 27528 17536
rect 27120 17496 27528 17524
rect 27120 17484 27126 17496
rect 27522 17484 27528 17496
rect 27580 17484 27586 17536
rect 28552 17524 28580 17555
rect 28626 17552 28632 17604
rect 28684 17592 28690 17604
rect 29365 17595 29423 17601
rect 29365 17592 29377 17595
rect 28684 17564 29377 17592
rect 28684 17552 28690 17564
rect 29365 17561 29377 17564
rect 29411 17592 29423 17595
rect 29914 17592 29920 17604
rect 29411 17564 29920 17592
rect 29411 17561 29423 17564
rect 29365 17555 29423 17561
rect 29914 17552 29920 17564
rect 29972 17552 29978 17604
rect 30760 17601 30788 17632
rect 31665 17629 31677 17632
rect 31711 17629 31723 17663
rect 33870 17660 33876 17672
rect 31665 17623 31723 17629
rect 32876 17632 33876 17660
rect 30745 17595 30803 17601
rect 30745 17561 30757 17595
rect 30791 17592 30803 17595
rect 31478 17592 31484 17604
rect 30791 17564 31484 17592
rect 30791 17561 30803 17564
rect 30745 17555 30803 17561
rect 31478 17552 31484 17564
rect 31536 17552 31542 17604
rect 32876 17592 32904 17632
rect 33870 17620 33876 17632
rect 33928 17620 33934 17672
rect 34057 17663 34115 17669
rect 34057 17629 34069 17663
rect 34103 17660 34115 17663
rect 35066 17660 35072 17672
rect 34103 17632 35072 17660
rect 34103 17629 34115 17632
rect 34057 17623 34115 17629
rect 31956 17564 32904 17592
rect 28994 17524 29000 17536
rect 28552 17496 29000 17524
rect 28994 17484 29000 17496
rect 29052 17484 29058 17536
rect 29178 17484 29184 17536
rect 29236 17484 29242 17536
rect 30006 17484 30012 17536
rect 30064 17524 30070 17536
rect 31573 17527 31631 17533
rect 31573 17524 31585 17527
rect 30064 17496 31585 17524
rect 30064 17484 30070 17496
rect 31573 17493 31585 17496
rect 31619 17524 31631 17527
rect 31956 17524 31984 17564
rect 33226 17552 33232 17604
rect 33284 17592 33290 17604
rect 34072 17592 34100 17623
rect 35066 17620 35072 17632
rect 35124 17660 35130 17672
rect 35250 17660 35256 17672
rect 35124 17632 35256 17660
rect 35124 17620 35130 17632
rect 35250 17620 35256 17632
rect 35308 17620 35314 17672
rect 36188 17646 36216 17700
rect 36722 17688 36728 17700
rect 36780 17688 36786 17740
rect 37274 17688 37280 17740
rect 37332 17728 37338 17740
rect 38105 17731 38163 17737
rect 38105 17728 38117 17731
rect 37332 17700 38117 17728
rect 37332 17688 37338 17700
rect 38105 17697 38117 17700
rect 38151 17697 38163 17731
rect 38105 17691 38163 17697
rect 37550 17620 37556 17672
rect 37608 17620 37614 17672
rect 38626 17660 38654 17768
rect 38749 17765 38761 17799
rect 38795 17796 38807 17799
rect 40862 17796 40868 17808
rect 38795 17768 40868 17796
rect 38795 17765 38807 17768
rect 38749 17759 38807 17765
rect 40862 17756 40868 17768
rect 40920 17756 40926 17808
rect 43438 17796 43444 17808
rect 41386 17768 43444 17796
rect 40678 17688 40684 17740
rect 40736 17728 40742 17740
rect 40957 17731 41015 17737
rect 40957 17728 40969 17731
rect 40736 17700 40969 17728
rect 40736 17688 40742 17700
rect 40957 17697 40969 17700
rect 41003 17697 41015 17731
rect 40957 17691 41015 17697
rect 41046 17688 41052 17740
rect 41104 17688 41110 17740
rect 41386 17660 41414 17768
rect 43438 17756 43444 17768
rect 43496 17756 43502 17808
rect 38626 17632 41414 17660
rect 48593 17663 48651 17669
rect 48593 17629 48605 17663
rect 48639 17660 48651 17663
rect 49326 17660 49332 17672
rect 48639 17632 49332 17660
rect 48639 17629 48651 17632
rect 48593 17623 48651 17629
rect 49326 17620 49332 17632
rect 49384 17620 49390 17672
rect 33284 17564 34100 17592
rect 33284 17552 33290 17564
rect 36998 17552 37004 17604
rect 37056 17592 37062 17604
rect 37277 17595 37335 17601
rect 37277 17592 37289 17595
rect 37056 17564 37289 17592
rect 37056 17552 37062 17564
rect 37277 17561 37289 17564
rect 37323 17561 37335 17595
rect 37277 17555 37335 17561
rect 37366 17552 37372 17604
rect 37424 17592 37430 17604
rect 38381 17595 38439 17601
rect 38381 17592 38393 17595
rect 37424 17564 38393 17592
rect 37424 17552 37430 17564
rect 38381 17561 38393 17564
rect 38427 17561 38439 17595
rect 38381 17555 38439 17561
rect 40865 17595 40923 17601
rect 40865 17561 40877 17595
rect 40911 17592 40923 17595
rect 48406 17592 48412 17604
rect 40911 17564 48412 17592
rect 40911 17561 40923 17564
rect 40865 17555 40923 17561
rect 48406 17552 48412 17564
rect 48464 17552 48470 17604
rect 31619 17496 31984 17524
rect 32033 17527 32091 17533
rect 31619 17493 31631 17496
rect 31573 17487 31631 17493
rect 32033 17493 32045 17527
rect 32079 17524 32091 17527
rect 32122 17524 32128 17536
rect 32079 17496 32128 17524
rect 32079 17493 32091 17496
rect 32033 17487 32091 17493
rect 32122 17484 32128 17496
rect 32180 17484 32186 17536
rect 32306 17484 32312 17536
rect 32364 17524 32370 17536
rect 32401 17527 32459 17533
rect 32401 17524 32413 17527
rect 32364 17496 32413 17524
rect 32364 17484 32370 17496
rect 32401 17493 32413 17496
rect 32447 17524 32459 17527
rect 32674 17524 32680 17536
rect 32447 17496 32680 17524
rect 32447 17493 32459 17496
rect 32401 17487 32459 17493
rect 32674 17484 32680 17496
rect 32732 17484 32738 17536
rect 33137 17527 33195 17533
rect 33137 17493 33149 17527
rect 33183 17524 33195 17527
rect 33318 17524 33324 17536
rect 33183 17496 33324 17524
rect 33183 17493 33195 17496
rect 33137 17487 33195 17493
rect 33318 17484 33324 17496
rect 33376 17484 33382 17536
rect 34514 17484 34520 17536
rect 34572 17484 34578 17536
rect 35066 17484 35072 17536
rect 35124 17484 35130 17536
rect 35437 17527 35495 17533
rect 35437 17493 35449 17527
rect 35483 17524 35495 17527
rect 35526 17524 35532 17536
rect 35483 17496 35532 17524
rect 35483 17493 35495 17496
rect 35437 17487 35495 17493
rect 35526 17484 35532 17496
rect 35584 17484 35590 17536
rect 36630 17484 36636 17536
rect 36688 17524 36694 17536
rect 38289 17527 38347 17533
rect 38289 17524 38301 17527
rect 36688 17496 38301 17524
rect 36688 17484 36694 17496
rect 38289 17493 38301 17496
rect 38335 17493 38347 17527
rect 38289 17487 38347 17493
rect 38930 17484 38936 17536
rect 38988 17524 38994 17536
rect 39025 17527 39083 17533
rect 39025 17524 39037 17527
rect 38988 17496 39037 17524
rect 38988 17484 38994 17496
rect 39025 17493 39037 17496
rect 39071 17493 39083 17527
rect 39025 17487 39083 17493
rect 39301 17527 39359 17533
rect 39301 17493 39313 17527
rect 39347 17524 39359 17527
rect 40034 17524 40040 17536
rect 39347 17496 40040 17524
rect 39347 17493 39359 17496
rect 39301 17487 39359 17493
rect 40034 17484 40040 17496
rect 40092 17484 40098 17536
rect 48682 17484 48688 17536
rect 48740 17484 48746 17536
rect 49142 17484 49148 17536
rect 49200 17484 49206 17536
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 13814 17320 13820 17332
rect 2746 17292 13820 17320
rect 1026 17076 1032 17128
rect 1084 17116 1090 17128
rect 1765 17119 1823 17125
rect 1765 17116 1777 17119
rect 1084 17088 1777 17116
rect 1084 17076 1090 17088
rect 1765 17085 1777 17088
rect 1811 17085 1823 17119
rect 1765 17079 1823 17085
rect 2130 17008 2136 17060
rect 2188 17048 2194 17060
rect 2746 17048 2774 17292
rect 13814 17280 13820 17292
rect 13872 17280 13878 17332
rect 13998 17280 14004 17332
rect 14056 17320 14062 17332
rect 14921 17323 14979 17329
rect 14921 17320 14933 17323
rect 14056 17292 14933 17320
rect 14056 17280 14062 17292
rect 14921 17289 14933 17292
rect 14967 17289 14979 17323
rect 14921 17283 14979 17289
rect 15562 17280 15568 17332
rect 15620 17280 15626 17332
rect 15672 17292 18828 17320
rect 10410 17212 10416 17264
rect 10468 17252 10474 17264
rect 10468 17224 10916 17252
rect 10468 17212 10474 17224
rect 2961 17187 3019 17193
rect 2961 17153 2973 17187
rect 3007 17184 3019 17187
rect 4338 17184 4344 17196
rect 3007 17156 4344 17184
rect 3007 17153 3019 17156
rect 2961 17147 3019 17153
rect 4338 17144 4344 17156
rect 4396 17144 4402 17196
rect 5902 17144 5908 17196
rect 5960 17184 5966 17196
rect 9858 17184 9864 17196
rect 5960 17156 9864 17184
rect 5960 17144 5966 17156
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 9950 17144 9956 17196
rect 10008 17184 10014 17196
rect 10781 17187 10839 17193
rect 10781 17184 10793 17187
rect 10008 17156 10793 17184
rect 10008 17144 10014 17156
rect 10781 17153 10793 17156
rect 10827 17153 10839 17187
rect 10888 17184 10916 17224
rect 11422 17212 11428 17264
rect 11480 17252 11486 17264
rect 11882 17252 11888 17264
rect 11480 17224 11888 17252
rect 11480 17212 11486 17224
rect 11882 17212 11888 17224
rect 11940 17212 11946 17264
rect 12342 17212 12348 17264
rect 12400 17252 12406 17264
rect 12989 17255 13047 17261
rect 12989 17252 13001 17255
rect 12400 17224 13001 17252
rect 12400 17212 12406 17224
rect 12989 17221 13001 17224
rect 13035 17221 13047 17255
rect 12989 17215 13047 17221
rect 13081 17255 13139 17261
rect 13081 17221 13093 17255
rect 13127 17252 13139 17255
rect 13262 17252 13268 17264
rect 13127 17224 13268 17252
rect 13127 17221 13139 17224
rect 13081 17215 13139 17221
rect 13262 17212 13268 17224
rect 13320 17212 13326 17264
rect 14090 17212 14096 17264
rect 14148 17252 14154 17264
rect 14277 17255 14335 17261
rect 14277 17252 14289 17255
rect 14148 17224 14289 17252
rect 14148 17212 14154 17224
rect 14277 17221 14289 17224
rect 14323 17221 14335 17255
rect 14277 17215 14335 17221
rect 14734 17212 14740 17264
rect 14792 17252 14798 17264
rect 15672 17252 15700 17292
rect 14792 17224 15700 17252
rect 14792 17212 14798 17224
rect 15746 17212 15752 17264
rect 15804 17252 15810 17264
rect 15933 17255 15991 17261
rect 15933 17252 15945 17255
rect 15804 17224 15945 17252
rect 15804 17212 15810 17224
rect 15933 17221 15945 17224
rect 15979 17221 15991 17255
rect 15933 17215 15991 17221
rect 16022 17212 16028 17264
rect 16080 17252 16086 17264
rect 17954 17252 17960 17264
rect 16080 17224 17960 17252
rect 16080 17212 16086 17224
rect 17954 17212 17960 17224
rect 18012 17212 18018 17264
rect 18690 17212 18696 17264
rect 18748 17212 18754 17264
rect 18800 17252 18828 17292
rect 19150 17280 19156 17332
rect 19208 17280 19214 17332
rect 20254 17320 20260 17332
rect 19260 17292 20260 17320
rect 19260 17252 19288 17292
rect 20254 17280 20260 17292
rect 20312 17280 20318 17332
rect 21726 17280 21732 17332
rect 21784 17320 21790 17332
rect 22002 17320 22008 17332
rect 21784 17292 22008 17320
rect 21784 17280 21790 17292
rect 22002 17280 22008 17292
rect 22060 17280 22066 17332
rect 22649 17323 22707 17329
rect 22649 17289 22661 17323
rect 22695 17320 22707 17323
rect 23474 17320 23480 17332
rect 22695 17292 23480 17320
rect 22695 17289 22707 17292
rect 22649 17283 22707 17289
rect 23474 17280 23480 17292
rect 23532 17280 23538 17332
rect 24026 17280 24032 17332
rect 24084 17320 24090 17332
rect 24857 17323 24915 17329
rect 24857 17320 24869 17323
rect 24084 17292 24869 17320
rect 24084 17280 24090 17292
rect 24857 17289 24869 17292
rect 24903 17289 24915 17323
rect 24857 17283 24915 17289
rect 25317 17323 25375 17329
rect 25317 17289 25329 17323
rect 25363 17320 25375 17323
rect 27341 17323 27399 17329
rect 27341 17320 27353 17323
rect 25363 17292 27353 17320
rect 25363 17289 25375 17292
rect 25317 17283 25375 17289
rect 27341 17289 27353 17292
rect 27387 17289 27399 17323
rect 27341 17283 27399 17289
rect 27706 17280 27712 17332
rect 27764 17280 27770 17332
rect 27798 17280 27804 17332
rect 27856 17320 27862 17332
rect 28997 17323 29055 17329
rect 28997 17320 29009 17323
rect 27856 17292 29009 17320
rect 27856 17280 27862 17292
rect 28997 17289 29009 17292
rect 29043 17289 29055 17323
rect 28997 17283 29055 17289
rect 30193 17323 30251 17329
rect 30193 17289 30205 17323
rect 30239 17320 30251 17323
rect 32306 17320 32312 17332
rect 30239 17292 32312 17320
rect 30239 17289 30251 17292
rect 30193 17283 30251 17289
rect 32306 17280 32312 17292
rect 32364 17280 32370 17332
rect 33594 17320 33600 17332
rect 32416 17292 33600 17320
rect 20530 17252 20536 17264
rect 18800 17224 19288 17252
rect 20194 17224 20536 17252
rect 20530 17212 20536 17224
rect 20588 17212 20594 17264
rect 20625 17255 20683 17261
rect 20625 17221 20637 17255
rect 20671 17252 20683 17255
rect 20990 17252 20996 17264
rect 20671 17224 20996 17252
rect 20671 17221 20683 17224
rect 20625 17215 20683 17221
rect 20990 17212 20996 17224
rect 21048 17252 21054 17264
rect 21450 17252 21456 17264
rect 21048 17224 21456 17252
rect 21048 17212 21054 17224
rect 21450 17212 21456 17224
rect 21508 17212 21514 17264
rect 23658 17212 23664 17264
rect 23716 17212 23722 17264
rect 24118 17212 24124 17264
rect 24176 17252 24182 17264
rect 24176 17224 24440 17252
rect 24176 17212 24182 17224
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 10888 17156 11713 17184
rect 10781 17147 10839 17153
rect 11701 17153 11713 17156
rect 11747 17153 11759 17187
rect 11701 17147 11759 17153
rect 11974 17144 11980 17196
rect 12032 17184 12038 17196
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 12032 17156 12449 17184
rect 12032 17144 12038 17156
rect 12437 17153 12449 17156
rect 12483 17184 12495 17187
rect 14752 17184 14780 17212
rect 12483 17156 14780 17184
rect 12483 17153 12495 17156
rect 12437 17147 12495 17153
rect 10505 17119 10563 17125
rect 10505 17085 10517 17119
rect 10551 17085 10563 17119
rect 10505 17079 10563 17085
rect 2188 17020 2774 17048
rect 9769 17051 9827 17057
rect 2188 17008 2194 17020
rect 9769 17017 9781 17051
rect 9815 17048 9827 17051
rect 10045 17051 10103 17057
rect 10045 17048 10057 17051
rect 9815 17020 10057 17048
rect 9815 17017 9827 17020
rect 9769 17011 9827 17017
rect 10045 17017 10057 17020
rect 10091 17048 10103 17051
rect 10520 17048 10548 17079
rect 10594 17076 10600 17128
rect 10652 17116 10658 17128
rect 10689 17119 10747 17125
rect 10689 17116 10701 17119
rect 10652 17088 10701 17116
rect 10652 17076 10658 17088
rect 10689 17085 10701 17088
rect 10735 17085 10747 17119
rect 12342 17116 12348 17128
rect 10689 17079 10747 17085
rect 11072 17088 12348 17116
rect 11072 17048 11100 17088
rect 12342 17076 12348 17088
rect 12400 17116 12406 17128
rect 12805 17119 12863 17125
rect 12805 17116 12817 17119
rect 12400 17088 12817 17116
rect 12400 17076 12406 17088
rect 12805 17085 12817 17088
rect 12851 17085 12863 17119
rect 12805 17079 12863 17085
rect 10091 17020 11100 17048
rect 11149 17051 11207 17057
rect 10091 17017 10103 17020
rect 10045 17011 10103 17017
rect 11149 17017 11161 17051
rect 11195 17048 11207 17051
rect 12710 17048 12716 17060
rect 11195 17020 12716 17048
rect 11195 17017 11207 17020
rect 11149 17011 11207 17017
rect 12710 17008 12716 17020
rect 12768 17008 12774 17060
rect 9490 16940 9496 16992
rect 9548 16980 9554 16992
rect 10502 16980 10508 16992
rect 9548 16952 10508 16980
rect 9548 16940 9554 16952
rect 10502 16940 10508 16952
rect 10560 16940 10566 16992
rect 10594 16940 10600 16992
rect 10652 16980 10658 16992
rect 11974 16980 11980 16992
rect 10652 16952 11980 16980
rect 10652 16940 10658 16952
rect 11974 16940 11980 16952
rect 12032 16940 12038 16992
rect 12802 16940 12808 16992
rect 12860 16980 12866 16992
rect 12912 16980 12940 17156
rect 15102 17144 15108 17196
rect 15160 17144 15166 17196
rect 16850 17184 16856 17196
rect 15948 17156 16856 17184
rect 14274 17076 14280 17128
rect 14332 17116 14338 17128
rect 15948 17116 15976 17156
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 17037 17187 17095 17193
rect 17037 17153 17049 17187
rect 17083 17184 17095 17187
rect 19334 17184 19340 17196
rect 17083 17156 19340 17184
rect 17083 17153 17095 17156
rect 17037 17147 17095 17153
rect 19334 17144 19340 17156
rect 19392 17144 19398 17196
rect 20901 17187 20959 17193
rect 20901 17153 20913 17187
rect 20947 17184 20959 17187
rect 22094 17184 22100 17196
rect 20947 17156 22100 17184
rect 20947 17153 20959 17156
rect 20901 17147 20959 17153
rect 22094 17144 22100 17156
rect 22152 17184 22158 17196
rect 22738 17184 22744 17196
rect 22152 17156 22744 17184
rect 22152 17144 22158 17156
rect 22738 17144 22744 17156
rect 22796 17144 22802 17196
rect 24412 17193 24440 17224
rect 25774 17212 25780 17264
rect 25832 17252 25838 17264
rect 25869 17255 25927 17261
rect 25869 17252 25881 17255
rect 25832 17224 25881 17252
rect 25832 17212 25838 17224
rect 25869 17221 25881 17224
rect 25915 17252 25927 17255
rect 25958 17252 25964 17264
rect 25915 17224 25964 17252
rect 25915 17221 25927 17224
rect 25869 17215 25927 17221
rect 25958 17212 25964 17224
rect 26016 17212 26022 17264
rect 26142 17212 26148 17264
rect 26200 17252 26206 17264
rect 27614 17252 27620 17264
rect 26200 17224 27620 17252
rect 26200 17212 26206 17224
rect 27614 17212 27620 17224
rect 27672 17212 27678 17264
rect 28810 17252 28816 17264
rect 27816 17224 28816 17252
rect 24397 17187 24455 17193
rect 24397 17153 24409 17187
rect 24443 17153 24455 17187
rect 24397 17147 24455 17153
rect 25225 17187 25283 17193
rect 25225 17153 25237 17187
rect 25271 17184 25283 17187
rect 25590 17184 25596 17196
rect 25271 17156 25596 17184
rect 25271 17153 25283 17156
rect 25225 17147 25283 17153
rect 25590 17144 25596 17156
rect 25648 17144 25654 17196
rect 26326 17144 26332 17196
rect 26384 17184 26390 17196
rect 27706 17184 27712 17196
rect 26384 17156 27712 17184
rect 26384 17144 26390 17156
rect 27706 17144 27712 17156
rect 27764 17144 27770 17196
rect 27816 17193 27844 17224
rect 28810 17212 28816 17224
rect 28868 17212 28874 17264
rect 28905 17255 28963 17261
rect 28905 17221 28917 17255
rect 28951 17252 28963 17255
rect 29822 17252 29828 17264
rect 28951 17224 29828 17252
rect 28951 17221 28963 17224
rect 28905 17215 28963 17221
rect 29822 17212 29828 17224
rect 29880 17212 29886 17264
rect 30101 17255 30159 17261
rect 30101 17252 30113 17255
rect 29932 17224 30113 17252
rect 27801 17187 27859 17193
rect 27801 17153 27813 17187
rect 27847 17153 27859 17187
rect 27801 17147 27859 17153
rect 14332 17088 15976 17116
rect 16025 17119 16083 17125
rect 14332 17076 14338 17088
rect 16025 17085 16037 17119
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 16040 17048 16068 17079
rect 16114 17076 16120 17128
rect 16172 17076 16178 17128
rect 16390 17076 16396 17128
rect 16448 17116 16454 17128
rect 21174 17116 21180 17128
rect 16448 17088 21180 17116
rect 16448 17076 16454 17088
rect 21174 17076 21180 17088
rect 21232 17076 21238 17128
rect 21269 17119 21327 17125
rect 21269 17085 21281 17119
rect 21315 17116 21327 17119
rect 21634 17116 21640 17128
rect 21315 17088 21640 17116
rect 21315 17085 21327 17088
rect 21269 17079 21327 17085
rect 21634 17076 21640 17088
rect 21692 17116 21698 17128
rect 22002 17116 22008 17128
rect 21692 17088 22008 17116
rect 21692 17076 21698 17088
rect 22002 17076 22008 17088
rect 22060 17116 22066 17128
rect 22189 17119 22247 17125
rect 22189 17116 22201 17119
rect 22060 17088 22201 17116
rect 22060 17076 22066 17088
rect 22189 17085 22201 17088
rect 22235 17116 22247 17119
rect 23382 17116 23388 17128
rect 22235 17088 23388 17116
rect 22235 17085 22247 17088
rect 22189 17079 22247 17085
rect 23382 17076 23388 17088
rect 23440 17076 23446 17128
rect 24121 17119 24179 17125
rect 24121 17085 24133 17119
rect 24167 17116 24179 17119
rect 24486 17116 24492 17128
rect 24167 17088 24492 17116
rect 24167 17085 24179 17088
rect 24121 17079 24179 17085
rect 24486 17076 24492 17088
rect 24544 17076 24550 17128
rect 25498 17076 25504 17128
rect 25556 17076 25562 17128
rect 27816 17116 27844 17147
rect 28442 17144 28448 17196
rect 28500 17184 28506 17196
rect 29270 17184 29276 17196
rect 28500 17156 29276 17184
rect 28500 17144 28506 17156
rect 29270 17144 29276 17156
rect 29328 17184 29334 17196
rect 29932 17184 29960 17224
rect 30101 17221 30113 17224
rect 30147 17221 30159 17255
rect 30101 17215 30159 17221
rect 30282 17212 30288 17264
rect 30340 17252 30346 17264
rect 31297 17255 31355 17261
rect 31297 17252 31309 17255
rect 30340 17224 31309 17252
rect 30340 17212 30346 17224
rect 31297 17221 31309 17224
rect 31343 17221 31355 17255
rect 32416 17252 32444 17292
rect 33594 17280 33600 17292
rect 33652 17280 33658 17332
rect 35066 17280 35072 17332
rect 35124 17320 35130 17332
rect 37829 17323 37887 17329
rect 37829 17320 37841 17323
rect 35124 17292 37841 17320
rect 35124 17280 35130 17292
rect 37829 17289 37841 17292
rect 37875 17289 37887 17323
rect 48314 17320 48320 17332
rect 37829 17283 37887 17289
rect 37936 17292 48320 17320
rect 31297 17215 31355 17221
rect 32324 17224 32444 17252
rect 30558 17184 30564 17196
rect 29328 17156 29960 17184
rect 30024 17156 30564 17184
rect 29328 17144 29334 17156
rect 27448 17088 27844 17116
rect 27893 17119 27951 17125
rect 16482 17048 16488 17060
rect 16040 17020 16488 17048
rect 16482 17008 16488 17020
rect 16540 17048 16546 17060
rect 16540 17020 17540 17048
rect 16540 17008 16546 17020
rect 12860 16952 12940 16980
rect 12860 16940 12866 16952
rect 13446 16940 13452 16992
rect 13504 16940 13510 16992
rect 14182 16940 14188 16992
rect 14240 16940 14246 16992
rect 15930 16940 15936 16992
rect 15988 16980 15994 16992
rect 16945 16983 17003 16989
rect 16945 16980 16957 16983
rect 15988 16952 16957 16980
rect 15988 16940 15994 16952
rect 16945 16949 16957 16952
rect 16991 16949 17003 16983
rect 16945 16943 17003 16949
rect 17402 16940 17408 16992
rect 17460 16940 17466 16992
rect 17512 16980 17540 17020
rect 20824 17020 22094 17048
rect 20824 16980 20852 17020
rect 17512 16952 20852 16980
rect 21634 16940 21640 16992
rect 21692 16980 21698 16992
rect 21913 16983 21971 16989
rect 21913 16980 21925 16983
rect 21692 16952 21925 16980
rect 21692 16940 21698 16952
rect 21913 16949 21925 16952
rect 21959 16949 21971 16983
rect 22066 16980 22094 17020
rect 25130 17008 25136 17060
rect 25188 17048 25194 17060
rect 26510 17048 26516 17060
rect 25188 17020 26516 17048
rect 25188 17008 25194 17020
rect 26510 17008 26516 17020
rect 26568 17008 26574 17060
rect 27448 16980 27476 17088
rect 27893 17085 27905 17119
rect 27939 17085 27951 17119
rect 27893 17079 27951 17085
rect 28813 17119 28871 17125
rect 28813 17085 28825 17119
rect 28859 17085 28871 17119
rect 28813 17079 28871 17085
rect 27522 17008 27528 17060
rect 27580 17048 27586 17060
rect 27908 17048 27936 17079
rect 27580 17020 27936 17048
rect 28828 17048 28856 17079
rect 28994 17076 29000 17128
rect 29052 17116 29058 17128
rect 29454 17116 29460 17128
rect 29052 17088 29460 17116
rect 29052 17076 29058 17088
rect 29454 17076 29460 17088
rect 29512 17076 29518 17128
rect 30024 17125 30052 17156
rect 30300 17128 30328 17156
rect 30558 17144 30564 17156
rect 30616 17144 30622 17196
rect 31386 17144 31392 17196
rect 31444 17144 31450 17196
rect 31478 17144 31484 17196
rect 31536 17184 31542 17196
rect 32214 17184 32220 17196
rect 31536 17156 32220 17184
rect 31536 17144 31542 17156
rect 32214 17144 32220 17156
rect 32272 17184 32278 17196
rect 32324 17193 32352 17224
rect 33042 17212 33048 17264
rect 33100 17212 33106 17264
rect 35526 17212 35532 17264
rect 35584 17252 35590 17264
rect 37001 17255 37059 17261
rect 37001 17252 37013 17255
rect 35584 17224 37013 17252
rect 35584 17212 35590 17224
rect 37001 17221 37013 17224
rect 37047 17221 37059 17255
rect 37936 17252 37964 17292
rect 48314 17280 48320 17292
rect 48372 17280 48378 17332
rect 48406 17280 48412 17332
rect 48464 17280 48470 17332
rect 37001 17215 37059 17221
rect 37108 17224 37964 17252
rect 32309 17187 32367 17193
rect 32309 17184 32321 17187
rect 32272 17156 32321 17184
rect 32272 17144 32278 17156
rect 32309 17153 32321 17156
rect 32355 17153 32367 17187
rect 32309 17147 32367 17153
rect 35158 17144 35164 17196
rect 35216 17184 35222 17196
rect 36265 17187 36323 17193
rect 36265 17184 36277 17187
rect 35216 17156 36277 17184
rect 35216 17144 35222 17156
rect 36265 17153 36277 17156
rect 36311 17153 36323 17187
rect 36265 17147 36323 17153
rect 36354 17144 36360 17196
rect 36412 17144 36418 17196
rect 30009 17119 30067 17125
rect 30009 17085 30021 17119
rect 30055 17085 30067 17119
rect 30009 17079 30067 17085
rect 30282 17076 30288 17128
rect 30340 17076 30346 17128
rect 30742 17076 30748 17128
rect 30800 17116 30806 17128
rect 31113 17119 31171 17125
rect 31113 17116 31125 17119
rect 30800 17088 31125 17116
rect 30800 17076 30806 17088
rect 31113 17085 31125 17088
rect 31159 17085 31171 17119
rect 31113 17079 31171 17085
rect 32582 17076 32588 17128
rect 32640 17076 32646 17128
rect 32950 17076 32956 17128
rect 33008 17116 33014 17128
rect 34057 17119 34115 17125
rect 34057 17116 34069 17119
rect 33008 17088 34069 17116
rect 33008 17076 33014 17088
rect 34057 17085 34069 17088
rect 34103 17085 34115 17119
rect 34057 17079 34115 17085
rect 34790 17076 34796 17128
rect 34848 17076 34854 17128
rect 36170 17076 36176 17128
rect 36228 17076 36234 17128
rect 29365 17051 29423 17057
rect 28828 17020 29040 17048
rect 27580 17008 27586 17020
rect 22066 16952 27476 16980
rect 29012 16980 29040 17020
rect 29365 17017 29377 17051
rect 29411 17048 29423 17051
rect 32306 17048 32312 17060
rect 29411 17020 32312 17048
rect 29411 17017 29423 17020
rect 29365 17011 29423 17017
rect 32306 17008 32312 17020
rect 32364 17008 32370 17060
rect 33686 17008 33692 17060
rect 33744 17048 33750 17060
rect 36078 17048 36084 17060
rect 33744 17020 36084 17048
rect 33744 17008 33750 17020
rect 36078 17008 36084 17020
rect 36136 17008 36142 17060
rect 37108 17048 37136 17224
rect 39942 17212 39948 17264
rect 40000 17212 40006 17264
rect 40126 17212 40132 17264
rect 40184 17252 40190 17264
rect 40405 17255 40463 17261
rect 40405 17252 40417 17255
rect 40184 17224 40417 17252
rect 40184 17212 40190 17224
rect 40405 17221 40417 17224
rect 40451 17221 40463 17255
rect 40405 17215 40463 17221
rect 40954 17212 40960 17264
rect 41012 17212 41018 17264
rect 48222 17212 48228 17264
rect 48280 17252 48286 17264
rect 48682 17252 48688 17264
rect 48280 17224 48688 17252
rect 48280 17212 48286 17224
rect 48682 17212 48688 17224
rect 48740 17252 48746 17264
rect 49237 17255 49295 17261
rect 49237 17252 49249 17255
rect 48740 17224 49249 17252
rect 48740 17212 48746 17224
rect 49237 17221 49249 17224
rect 49283 17221 49295 17255
rect 49237 17215 49295 17221
rect 37921 17187 37979 17193
rect 37921 17153 37933 17187
rect 37967 17184 37979 17187
rect 38930 17184 38936 17196
rect 37967 17156 38936 17184
rect 37967 17153 37979 17156
rect 37921 17147 37979 17153
rect 38930 17144 38936 17156
rect 38988 17144 38994 17196
rect 48593 17187 48651 17193
rect 48593 17153 48605 17187
rect 48639 17184 48651 17187
rect 48774 17184 48780 17196
rect 48639 17156 48780 17184
rect 48639 17153 48651 17156
rect 48593 17147 48651 17153
rect 48774 17144 48780 17156
rect 48832 17144 48838 17196
rect 37826 17076 37832 17128
rect 37884 17116 37890 17128
rect 38013 17119 38071 17125
rect 38013 17116 38025 17119
rect 37884 17088 38025 17116
rect 37884 17076 37890 17088
rect 38013 17085 38025 17088
rect 38059 17085 38071 17119
rect 38013 17079 38071 17085
rect 40678 17076 40684 17128
rect 40736 17076 40742 17128
rect 49050 17076 49056 17128
rect 49108 17076 49114 17128
rect 36372 17020 37136 17048
rect 29454 16980 29460 16992
rect 29012 16952 29460 16980
rect 21913 16943 21971 16949
rect 29454 16940 29460 16952
rect 29512 16940 29518 16992
rect 30558 16940 30564 16992
rect 30616 16940 30622 16992
rect 31757 16983 31815 16989
rect 31757 16949 31769 16983
rect 31803 16980 31815 16983
rect 33778 16980 33784 16992
rect 31803 16952 33784 16980
rect 31803 16949 31815 16952
rect 31757 16943 31815 16949
rect 33778 16940 33784 16952
rect 33836 16940 33842 16992
rect 35618 16940 35624 16992
rect 35676 16980 35682 16992
rect 36372 16980 36400 17020
rect 37182 17008 37188 17060
rect 37240 17048 37246 17060
rect 37461 17051 37519 17057
rect 37461 17048 37473 17051
rect 37240 17020 37473 17048
rect 37240 17008 37246 17020
rect 37461 17017 37473 17020
rect 37507 17017 37519 17051
rect 41046 17048 41052 17060
rect 37461 17011 37519 17017
rect 40880 17020 41052 17048
rect 35676 16952 36400 16980
rect 35676 16940 35682 16952
rect 36722 16940 36728 16992
rect 36780 16940 36786 16992
rect 38565 16983 38623 16989
rect 38565 16949 38577 16983
rect 38611 16980 38623 16983
rect 38746 16980 38752 16992
rect 38611 16952 38752 16980
rect 38611 16949 38623 16952
rect 38565 16943 38623 16949
rect 38746 16940 38752 16952
rect 38804 16940 38810 16992
rect 38838 16940 38844 16992
rect 38896 16980 38902 16992
rect 38933 16983 38991 16989
rect 38933 16980 38945 16983
rect 38896 16952 38945 16980
rect 38896 16940 38902 16952
rect 38933 16949 38945 16952
rect 38979 16980 38991 16983
rect 40880 16980 40908 17020
rect 41046 17008 41052 17020
rect 41104 17008 41110 17060
rect 38979 16952 40908 16980
rect 38979 16949 38991 16952
rect 38933 16943 38991 16949
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 14182 16776 14188 16788
rect 2976 16748 14188 16776
rect 2976 16581 3004 16748
rect 14182 16736 14188 16748
rect 14240 16736 14246 16788
rect 14642 16736 14648 16788
rect 14700 16776 14706 16788
rect 18619 16779 18677 16785
rect 14700 16748 17356 16776
rect 14700 16736 14706 16748
rect 4430 16668 4436 16720
rect 4488 16708 4494 16720
rect 5442 16708 5448 16720
rect 4488 16680 5448 16708
rect 4488 16668 4494 16680
rect 5442 16668 5448 16680
rect 5500 16708 5506 16720
rect 5500 16680 8064 16708
rect 5500 16668 5506 16680
rect 8036 16649 8064 16680
rect 10226 16668 10232 16720
rect 10284 16708 10290 16720
rect 10321 16711 10379 16717
rect 10321 16708 10333 16711
rect 10284 16680 10333 16708
rect 10284 16668 10290 16680
rect 10321 16677 10333 16680
rect 10367 16677 10379 16711
rect 10321 16671 10379 16677
rect 12434 16668 12440 16720
rect 12492 16708 12498 16720
rect 12529 16711 12587 16717
rect 12529 16708 12541 16711
rect 12492 16680 12541 16708
rect 12492 16668 12498 16680
rect 12529 16677 12541 16680
rect 12575 16677 12587 16711
rect 12529 16671 12587 16677
rect 13814 16668 13820 16720
rect 13872 16708 13878 16720
rect 16666 16708 16672 16720
rect 13872 16680 16672 16708
rect 13872 16668 13878 16680
rect 7929 16643 7987 16649
rect 7929 16609 7941 16643
rect 7975 16609 7987 16643
rect 7929 16603 7987 16609
rect 8021 16643 8079 16649
rect 8021 16609 8033 16643
rect 8067 16609 8079 16643
rect 8021 16603 8079 16609
rect 2961 16575 3019 16581
rect 2961 16541 2973 16575
rect 3007 16541 3019 16575
rect 7944 16572 7972 16603
rect 10870 16600 10876 16652
rect 10928 16640 10934 16652
rect 11149 16643 11207 16649
rect 11149 16640 11161 16643
rect 10928 16612 11161 16640
rect 10928 16600 10934 16612
rect 11149 16609 11161 16612
rect 11195 16609 11207 16643
rect 11149 16603 11207 16609
rect 13173 16643 13231 16649
rect 13173 16609 13185 16643
rect 13219 16640 13231 16643
rect 14645 16643 14703 16649
rect 13219 16612 14596 16640
rect 13219 16609 13231 16612
rect 13173 16603 13231 16609
rect 9030 16572 9036 16584
rect 7944 16544 9036 16572
rect 2961 16535 3019 16541
rect 9030 16532 9036 16544
rect 9088 16532 9094 16584
rect 12345 16575 12403 16581
rect 12345 16541 12357 16575
rect 12391 16572 12403 16575
rect 12391 16544 12756 16572
rect 12391 16541 12403 16544
rect 12345 16535 12403 16541
rect 1026 16464 1032 16516
rect 1084 16504 1090 16516
rect 1765 16507 1823 16513
rect 1765 16504 1777 16507
rect 1084 16476 1777 16504
rect 1084 16464 1090 16476
rect 1765 16473 1777 16476
rect 1811 16473 1823 16507
rect 1765 16467 1823 16473
rect 7834 16464 7840 16516
rect 7892 16504 7898 16516
rect 8113 16507 8171 16513
rect 8113 16504 8125 16507
rect 7892 16476 8125 16504
rect 7892 16464 7898 16476
rect 8113 16473 8125 16476
rect 8159 16473 8171 16507
rect 9674 16504 9680 16516
rect 8113 16467 8171 16473
rect 8496 16476 9680 16504
rect 8496 16445 8524 16476
rect 9674 16464 9680 16476
rect 9732 16464 9738 16516
rect 10045 16507 10103 16513
rect 10045 16473 10057 16507
rect 10091 16504 10103 16507
rect 10502 16504 10508 16516
rect 10091 16476 10508 16504
rect 10091 16473 10103 16476
rect 10045 16467 10103 16473
rect 10502 16464 10508 16476
rect 10560 16464 10566 16516
rect 11425 16507 11483 16513
rect 11425 16473 11437 16507
rect 11471 16504 11483 16507
rect 12618 16504 12624 16516
rect 11471 16476 12624 16504
rect 11471 16473 11483 16476
rect 11425 16467 11483 16473
rect 12618 16464 12624 16476
rect 12676 16464 12682 16516
rect 12728 16504 12756 16544
rect 12802 16532 12808 16584
rect 12860 16572 12866 16584
rect 13538 16572 13544 16584
rect 12860 16544 13544 16572
rect 12860 16532 12866 16544
rect 13538 16532 13544 16544
rect 13596 16532 13602 16584
rect 14568 16572 14596 16612
rect 14645 16609 14657 16643
rect 14691 16640 14703 16643
rect 15378 16640 15384 16652
rect 14691 16612 15384 16640
rect 14691 16609 14703 16612
rect 14645 16603 14703 16609
rect 15378 16600 15384 16612
rect 15436 16600 15442 16652
rect 16132 16649 16160 16680
rect 16666 16668 16672 16680
rect 16724 16668 16730 16720
rect 16117 16643 16175 16649
rect 16117 16609 16129 16643
rect 16163 16609 16175 16643
rect 16117 16603 16175 16609
rect 16209 16643 16267 16649
rect 16209 16609 16221 16643
rect 16255 16609 16267 16643
rect 16209 16603 16267 16609
rect 14918 16572 14924 16584
rect 14568 16544 14924 16572
rect 14918 16532 14924 16544
rect 14976 16572 14982 16584
rect 16224 16572 16252 16603
rect 14976 16544 16252 16572
rect 14976 16532 14982 16544
rect 16666 16532 16672 16584
rect 16724 16532 16730 16584
rect 16684 16504 16712 16532
rect 12728 16476 16712 16504
rect 8481 16439 8539 16445
rect 8481 16405 8493 16439
rect 8527 16405 8539 16439
rect 8481 16399 8539 16405
rect 9030 16396 9036 16448
rect 9088 16396 9094 16448
rect 11330 16396 11336 16448
rect 11388 16396 11394 16448
rect 11793 16439 11851 16445
rect 11793 16405 11805 16439
rect 11839 16436 11851 16439
rect 11974 16436 11980 16448
rect 11839 16408 11980 16436
rect 11839 16405 11851 16408
rect 11793 16399 11851 16405
rect 11974 16396 11980 16408
rect 12032 16396 12038 16448
rect 12894 16396 12900 16448
rect 12952 16436 12958 16448
rect 13265 16439 13323 16445
rect 13265 16436 13277 16439
rect 12952 16408 13277 16436
rect 12952 16396 12958 16408
rect 13265 16405 13277 16408
rect 13311 16405 13323 16439
rect 13265 16399 13323 16405
rect 13357 16439 13415 16445
rect 13357 16405 13369 16439
rect 13403 16436 13415 16439
rect 13538 16436 13544 16448
rect 13403 16408 13544 16436
rect 13403 16405 13415 16408
rect 13357 16399 13415 16405
rect 13538 16396 13544 16408
rect 13596 16396 13602 16448
rect 13630 16396 13636 16448
rect 13688 16436 13694 16448
rect 13725 16439 13783 16445
rect 13725 16436 13737 16439
rect 13688 16408 13737 16436
rect 13688 16396 13694 16408
rect 13725 16405 13737 16408
rect 13771 16405 13783 16439
rect 13725 16399 13783 16405
rect 14182 16396 14188 16448
rect 14240 16396 14246 16448
rect 14734 16396 14740 16448
rect 14792 16396 14798 16448
rect 14826 16396 14832 16448
rect 14884 16396 14890 16448
rect 15197 16439 15255 16445
rect 15197 16405 15209 16439
rect 15243 16436 15255 16439
rect 15470 16436 15476 16448
rect 15243 16408 15476 16436
rect 15243 16405 15255 16408
rect 15197 16399 15255 16405
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 15654 16396 15660 16448
rect 15712 16396 15718 16448
rect 16025 16439 16083 16445
rect 16025 16405 16037 16439
rect 16071 16436 16083 16439
rect 16390 16436 16396 16448
rect 16071 16408 16396 16436
rect 16071 16405 16083 16408
rect 16025 16399 16083 16405
rect 16390 16396 16396 16408
rect 16448 16436 16454 16448
rect 16669 16439 16727 16445
rect 16669 16436 16681 16439
rect 16448 16408 16681 16436
rect 16448 16396 16454 16408
rect 16669 16405 16681 16408
rect 16715 16405 16727 16439
rect 16669 16399 16727 16405
rect 17126 16396 17132 16448
rect 17184 16396 17190 16448
rect 17328 16436 17356 16748
rect 18619 16745 18631 16779
rect 18665 16776 18677 16779
rect 18874 16776 18880 16788
rect 18665 16748 18880 16776
rect 18665 16745 18677 16748
rect 18619 16739 18677 16745
rect 18874 16736 18880 16748
rect 18932 16736 18938 16788
rect 20990 16736 20996 16788
rect 21048 16736 21054 16788
rect 21174 16736 21180 16788
rect 21232 16776 21238 16788
rect 21232 16748 23244 16776
rect 21232 16736 21238 16748
rect 20162 16668 20168 16720
rect 20220 16708 20226 16720
rect 21008 16708 21036 16736
rect 22830 16708 22836 16720
rect 20220 16680 21036 16708
rect 22664 16680 22836 16708
rect 20220 16668 20226 16680
rect 17954 16600 17960 16652
rect 18012 16640 18018 16652
rect 18877 16643 18935 16649
rect 18877 16640 18889 16643
rect 18012 16612 18889 16640
rect 18012 16600 18018 16612
rect 18877 16609 18889 16612
rect 18923 16640 18935 16643
rect 19150 16640 19156 16652
rect 18923 16612 19156 16640
rect 18923 16609 18935 16612
rect 18877 16603 18935 16609
rect 19150 16600 19156 16612
rect 19208 16600 19214 16652
rect 20622 16600 20628 16652
rect 20680 16640 20686 16652
rect 22370 16640 22376 16652
rect 20680 16612 22376 16640
rect 20680 16600 20686 16612
rect 22370 16600 22376 16612
rect 22428 16600 22434 16652
rect 22465 16643 22523 16649
rect 22465 16609 22477 16643
rect 22511 16640 22523 16643
rect 22664 16640 22692 16680
rect 22830 16668 22836 16680
rect 22888 16668 22894 16720
rect 23216 16708 23244 16748
rect 23290 16736 23296 16788
rect 23348 16776 23354 16788
rect 24673 16779 24731 16785
rect 24673 16776 24685 16779
rect 23348 16748 24685 16776
rect 23348 16736 23354 16748
rect 24673 16745 24685 16748
rect 24719 16776 24731 16779
rect 27614 16776 27620 16788
rect 24719 16748 27620 16776
rect 24719 16745 24731 16748
rect 24673 16739 24731 16745
rect 27614 16736 27620 16748
rect 27672 16776 27678 16788
rect 28626 16776 28632 16788
rect 27672 16748 28632 16776
rect 27672 16736 27678 16748
rect 28626 16736 28632 16748
rect 28684 16736 28690 16788
rect 28810 16736 28816 16788
rect 28868 16736 28874 16788
rect 31110 16776 31116 16788
rect 28920 16748 31116 16776
rect 26050 16708 26056 16720
rect 23216 16680 23704 16708
rect 22511 16612 22692 16640
rect 22511 16609 22523 16612
rect 22465 16603 22523 16609
rect 22738 16600 22744 16652
rect 22796 16600 22802 16652
rect 17494 16532 17500 16584
rect 17552 16532 17558 16584
rect 20257 16575 20315 16581
rect 20257 16541 20269 16575
rect 20303 16541 20315 16575
rect 23676 16572 23704 16680
rect 23768 16680 26056 16708
rect 23768 16649 23796 16680
rect 26050 16668 26056 16680
rect 26108 16668 26114 16720
rect 27709 16711 27767 16717
rect 27709 16677 27721 16711
rect 27755 16708 27767 16711
rect 27798 16708 27804 16720
rect 27755 16680 27804 16708
rect 27755 16677 27767 16680
rect 27709 16671 27767 16677
rect 27798 16668 27804 16680
rect 27856 16668 27862 16720
rect 28920 16708 28948 16748
rect 31110 16736 31116 16748
rect 31168 16736 31174 16788
rect 34606 16776 34612 16788
rect 31726 16748 34612 16776
rect 28092 16680 28948 16708
rect 29181 16711 29239 16717
rect 23753 16643 23811 16649
rect 23753 16609 23765 16643
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 23937 16643 23995 16649
rect 23937 16609 23949 16643
rect 23983 16640 23995 16643
rect 25593 16643 25651 16649
rect 25593 16640 25605 16643
rect 23983 16612 25605 16640
rect 23983 16609 23995 16612
rect 23937 16603 23995 16609
rect 25593 16609 25605 16612
rect 25639 16640 25651 16643
rect 25866 16640 25872 16652
rect 25639 16612 25872 16640
rect 25639 16609 25651 16612
rect 25593 16603 25651 16609
rect 25866 16600 25872 16612
rect 25924 16600 25930 16652
rect 26418 16600 26424 16652
rect 26476 16640 26482 16652
rect 27062 16640 27068 16652
rect 26476 16612 27068 16640
rect 26476 16600 26482 16612
rect 27062 16600 27068 16612
rect 27120 16600 27126 16652
rect 27430 16600 27436 16652
rect 27488 16640 27494 16652
rect 27982 16640 27988 16652
rect 27488 16612 27988 16640
rect 27488 16600 27494 16612
rect 27982 16600 27988 16612
rect 28040 16600 28046 16652
rect 27341 16575 27399 16581
rect 23676 16544 25176 16572
rect 20257 16535 20315 16541
rect 20272 16504 20300 16535
rect 18248 16476 20116 16504
rect 20272 16476 21220 16504
rect 18248 16436 18276 16476
rect 17328 16408 18276 16436
rect 18782 16396 18788 16448
rect 18840 16436 18846 16448
rect 20088 16445 20116 16476
rect 19429 16439 19487 16445
rect 19429 16436 19441 16439
rect 18840 16408 19441 16436
rect 18840 16396 18846 16408
rect 19429 16405 19441 16408
rect 19475 16405 19487 16439
rect 19429 16399 19487 16405
rect 20073 16439 20131 16445
rect 20073 16405 20085 16439
rect 20119 16405 20131 16439
rect 20073 16399 20131 16405
rect 20530 16396 20536 16448
rect 20588 16436 20594 16448
rect 20625 16439 20683 16445
rect 20625 16436 20637 16439
rect 20588 16408 20637 16436
rect 20588 16396 20594 16408
rect 20625 16405 20637 16408
rect 20671 16436 20683 16439
rect 20806 16436 20812 16448
rect 20671 16408 20812 16436
rect 20671 16405 20683 16408
rect 20625 16399 20683 16405
rect 20806 16396 20812 16408
rect 20864 16396 20870 16448
rect 21192 16436 21220 16476
rect 22002 16464 22008 16516
rect 22060 16464 22066 16516
rect 24578 16464 24584 16516
rect 24636 16464 24642 16516
rect 25148 16448 25176 16544
rect 27341 16541 27353 16575
rect 27387 16572 27399 16575
rect 27798 16572 27804 16584
rect 27387 16544 27804 16572
rect 27387 16541 27399 16544
rect 27341 16535 27399 16541
rect 27798 16532 27804 16544
rect 27856 16532 27862 16584
rect 26786 16504 26792 16516
rect 26634 16476 26792 16504
rect 26786 16464 26792 16476
rect 26844 16464 26850 16516
rect 22830 16436 22836 16448
rect 21192 16408 22836 16436
rect 22830 16396 22836 16408
rect 22888 16396 22894 16448
rect 22922 16396 22928 16448
rect 22980 16436 22986 16448
rect 23293 16439 23351 16445
rect 23293 16436 23305 16439
rect 22980 16408 23305 16436
rect 22980 16396 22986 16408
rect 23293 16405 23305 16408
rect 23339 16405 23351 16439
rect 23293 16399 23351 16405
rect 23658 16396 23664 16448
rect 23716 16396 23722 16448
rect 25130 16396 25136 16448
rect 25188 16436 25194 16448
rect 28092 16436 28120 16680
rect 29181 16677 29193 16711
rect 29227 16708 29239 16711
rect 29227 16680 30236 16708
rect 29227 16677 29239 16680
rect 29181 16671 29239 16677
rect 30208 16652 30236 16680
rect 28258 16600 28264 16652
rect 28316 16640 28322 16652
rect 28537 16643 28595 16649
rect 28537 16640 28549 16643
rect 28316 16612 28549 16640
rect 28316 16600 28322 16612
rect 28537 16609 28549 16612
rect 28583 16609 28595 16643
rect 28537 16603 28595 16609
rect 29270 16600 29276 16652
rect 29328 16600 29334 16652
rect 29917 16643 29975 16649
rect 29917 16609 29929 16643
rect 29963 16640 29975 16643
rect 30098 16640 30104 16652
rect 29963 16612 30104 16640
rect 29963 16609 29975 16612
rect 29917 16603 29975 16609
rect 30098 16600 30104 16612
rect 30156 16600 30162 16652
rect 30190 16600 30196 16652
rect 30248 16600 30254 16652
rect 31113 16643 31171 16649
rect 31113 16609 31125 16643
rect 31159 16640 31171 16643
rect 31726 16640 31754 16748
rect 34606 16736 34612 16748
rect 34664 16736 34670 16788
rect 36265 16779 36323 16785
rect 36265 16745 36277 16779
rect 36311 16776 36323 16779
rect 36354 16776 36360 16788
rect 36311 16748 36360 16776
rect 36311 16745 36323 16748
rect 36265 16739 36323 16745
rect 36354 16736 36360 16748
rect 36412 16736 36418 16788
rect 36446 16736 36452 16788
rect 36504 16776 36510 16788
rect 36630 16776 36636 16788
rect 36504 16748 36636 16776
rect 36504 16736 36510 16748
rect 36630 16736 36636 16748
rect 36688 16736 36694 16788
rect 37182 16736 37188 16788
rect 37240 16776 37246 16788
rect 37458 16776 37464 16788
rect 37240 16748 37464 16776
rect 37240 16736 37246 16748
rect 37458 16736 37464 16748
rect 37516 16736 37522 16788
rect 40218 16736 40224 16788
rect 40276 16736 40282 16788
rect 40954 16736 40960 16788
rect 41012 16776 41018 16788
rect 41049 16779 41107 16785
rect 41049 16776 41061 16779
rect 41012 16748 41061 16776
rect 41012 16736 41018 16748
rect 41049 16745 41061 16748
rect 41095 16776 41107 16779
rect 41322 16776 41328 16788
rect 41095 16748 41328 16776
rect 41095 16745 41107 16748
rect 41049 16739 41107 16745
rect 41322 16736 41328 16748
rect 41380 16736 41386 16788
rect 41509 16779 41567 16785
rect 41509 16745 41521 16779
rect 41555 16776 41567 16779
rect 46014 16776 46020 16788
rect 41555 16748 46020 16776
rect 41555 16745 41567 16748
rect 41509 16739 41567 16745
rect 34054 16668 34060 16720
rect 34112 16708 34118 16720
rect 34241 16711 34299 16717
rect 34241 16708 34253 16711
rect 34112 16680 34253 16708
rect 34112 16668 34118 16680
rect 34241 16677 34253 16680
rect 34287 16677 34299 16711
rect 37550 16708 37556 16720
rect 34241 16671 34299 16677
rect 35084 16680 37556 16708
rect 31159 16612 31754 16640
rect 31159 16609 31171 16612
rect 31113 16603 31171 16609
rect 31938 16600 31944 16652
rect 31996 16600 32002 16652
rect 32214 16600 32220 16652
rect 32272 16600 32278 16652
rect 33686 16600 33692 16652
rect 33744 16640 33750 16652
rect 35084 16649 35112 16680
rect 37550 16668 37556 16680
rect 37608 16668 37614 16720
rect 40236 16708 40264 16736
rect 40236 16680 41184 16708
rect 34425 16643 34483 16649
rect 34425 16640 34437 16643
rect 33744 16612 34437 16640
rect 33744 16600 33750 16612
rect 34425 16609 34437 16612
rect 34471 16609 34483 16643
rect 34425 16603 34483 16609
rect 35069 16643 35127 16649
rect 35069 16609 35081 16643
rect 35115 16609 35127 16643
rect 35069 16603 35127 16609
rect 35342 16600 35348 16652
rect 35400 16640 35406 16652
rect 36725 16643 36783 16649
rect 36725 16640 36737 16643
rect 35400 16612 36737 16640
rect 35400 16600 35406 16612
rect 36725 16609 36737 16612
rect 36771 16609 36783 16643
rect 36725 16603 36783 16609
rect 28350 16532 28356 16584
rect 28408 16532 28414 16584
rect 30009 16575 30067 16581
rect 30009 16541 30021 16575
rect 30055 16572 30067 16575
rect 30208 16572 30236 16600
rect 31956 16572 31984 16600
rect 30055 16544 30236 16572
rect 30392 16544 32260 16572
rect 30055 16541 30067 16544
rect 30009 16535 30067 16541
rect 28261 16507 28319 16513
rect 28261 16473 28273 16507
rect 28307 16504 28319 16507
rect 28626 16504 28632 16516
rect 28307 16476 28632 16504
rect 28307 16473 28319 16476
rect 28261 16467 28319 16473
rect 28626 16464 28632 16476
rect 28684 16504 28690 16516
rect 28994 16504 29000 16516
rect 28684 16476 29000 16504
rect 28684 16464 28690 16476
rect 28994 16464 29000 16476
rect 29052 16464 29058 16516
rect 29086 16464 29092 16516
rect 29144 16504 29150 16516
rect 30101 16507 30159 16513
rect 30101 16504 30113 16507
rect 29144 16476 30113 16504
rect 29144 16464 29150 16476
rect 30101 16473 30113 16476
rect 30147 16473 30159 16507
rect 30101 16467 30159 16473
rect 25188 16408 28120 16436
rect 25188 16396 25194 16408
rect 29730 16396 29736 16448
rect 29788 16436 29794 16448
rect 30392 16436 30420 16544
rect 31938 16504 31944 16516
rect 30484 16476 31944 16504
rect 30484 16445 30512 16476
rect 31938 16464 31944 16476
rect 31996 16464 32002 16516
rect 32232 16504 32260 16544
rect 35526 16532 35532 16584
rect 35584 16572 35590 16584
rect 35805 16575 35863 16581
rect 35805 16572 35817 16575
rect 35584 16544 35817 16572
rect 35584 16532 35590 16544
rect 35805 16541 35817 16544
rect 35851 16541 35863 16575
rect 36740 16572 36768 16603
rect 36814 16600 36820 16652
rect 36872 16600 36878 16652
rect 37458 16600 37464 16652
rect 37516 16640 37522 16652
rect 38838 16640 38844 16652
rect 37516 16612 38844 16640
rect 37516 16600 37522 16612
rect 38838 16600 38844 16612
rect 38896 16640 38902 16652
rect 39209 16643 39267 16649
rect 39209 16640 39221 16643
rect 38896 16612 39221 16640
rect 38896 16600 38902 16612
rect 39209 16609 39221 16612
rect 39255 16609 39267 16643
rect 39209 16603 39267 16609
rect 40221 16643 40279 16649
rect 40221 16609 40233 16643
rect 40267 16640 40279 16643
rect 40310 16640 40316 16652
rect 40267 16612 40316 16640
rect 40267 16609 40279 16612
rect 40221 16603 40279 16609
rect 40310 16600 40316 16612
rect 40368 16600 40374 16652
rect 41156 16640 41184 16680
rect 41230 16668 41236 16720
rect 41288 16668 41294 16720
rect 41524 16708 41552 16739
rect 46014 16736 46020 16748
rect 46072 16736 46078 16788
rect 48774 16736 48780 16788
rect 48832 16736 48838 16788
rect 41386 16680 41552 16708
rect 41386 16640 41414 16680
rect 41156 16612 41414 16640
rect 37277 16575 37335 16581
rect 37277 16572 37289 16575
rect 36740 16544 37289 16572
rect 35805 16535 35863 16541
rect 37277 16541 37289 16544
rect 37323 16541 37335 16575
rect 37277 16535 37335 16541
rect 39482 16532 39488 16584
rect 39540 16572 39546 16584
rect 40678 16572 40684 16584
rect 39540 16544 40684 16572
rect 39540 16532 39546 16544
rect 40678 16532 40684 16544
rect 40736 16532 40742 16584
rect 48593 16575 48651 16581
rect 48593 16541 48605 16575
rect 48639 16572 48651 16575
rect 49329 16575 49387 16581
rect 49329 16572 49341 16575
rect 48639 16544 49341 16572
rect 48639 16541 48651 16544
rect 48593 16535 48651 16541
rect 49329 16541 49341 16544
rect 49375 16572 49387 16575
rect 49418 16572 49424 16584
rect 49375 16544 49424 16572
rect 49375 16541 49387 16544
rect 49329 16535 49387 16541
rect 49418 16532 49424 16544
rect 49476 16532 49482 16584
rect 32493 16507 32551 16513
rect 32493 16504 32505 16507
rect 32232 16476 32505 16504
rect 32493 16473 32505 16476
rect 32539 16504 32551 16507
rect 32766 16504 32772 16516
rect 32539 16476 32772 16504
rect 32539 16473 32551 16476
rect 32493 16467 32551 16473
rect 32766 16464 32772 16476
rect 32824 16464 32830 16516
rect 32950 16464 32956 16516
rect 33008 16464 33014 16516
rect 35894 16504 35900 16516
rect 33980 16476 35900 16504
rect 33980 16448 34008 16476
rect 35894 16464 35900 16476
rect 35952 16464 35958 16516
rect 36078 16464 36084 16516
rect 36136 16504 36142 16516
rect 36814 16504 36820 16516
rect 36136 16476 36820 16504
rect 36136 16464 36142 16476
rect 36814 16464 36820 16476
rect 36872 16464 36878 16516
rect 38746 16464 38752 16516
rect 38804 16504 38810 16516
rect 39942 16504 39948 16516
rect 38804 16476 39948 16504
rect 38804 16464 38810 16476
rect 39942 16464 39948 16476
rect 40000 16464 40006 16516
rect 40218 16464 40224 16516
rect 40276 16504 40282 16516
rect 40313 16507 40371 16513
rect 40313 16504 40325 16507
rect 40276 16476 40325 16504
rect 40276 16464 40282 16476
rect 40313 16473 40325 16476
rect 40359 16473 40371 16507
rect 40313 16467 40371 16473
rect 40405 16507 40463 16513
rect 40405 16473 40417 16507
rect 40451 16504 40463 16507
rect 41230 16504 41236 16516
rect 40451 16476 41236 16504
rect 40451 16473 40463 16476
rect 40405 16467 40463 16473
rect 41230 16464 41236 16476
rect 41288 16464 41294 16516
rect 29788 16408 30420 16436
rect 30469 16439 30527 16445
rect 29788 16396 29794 16408
rect 30469 16405 30481 16439
rect 30515 16405 30527 16439
rect 30469 16399 30527 16405
rect 31202 16396 31208 16448
rect 31260 16396 31266 16448
rect 31294 16396 31300 16448
rect 31352 16396 31358 16448
rect 31662 16396 31668 16448
rect 31720 16396 31726 16448
rect 32674 16396 32680 16448
rect 32732 16436 32738 16448
rect 33410 16436 33416 16448
rect 32732 16408 33416 16436
rect 32732 16396 32738 16408
rect 33410 16396 33416 16408
rect 33468 16396 33474 16448
rect 33962 16396 33968 16448
rect 34020 16396 34026 16448
rect 34606 16396 34612 16448
rect 34664 16436 34670 16448
rect 35802 16436 35808 16448
rect 34664 16408 35808 16436
rect 34664 16396 34670 16408
rect 35802 16396 35808 16408
rect 35860 16396 35866 16448
rect 36633 16439 36691 16445
rect 36633 16405 36645 16439
rect 36679 16436 36691 16439
rect 37182 16436 37188 16448
rect 36679 16408 37188 16436
rect 36679 16405 36691 16408
rect 36633 16399 36691 16405
rect 37182 16396 37188 16408
rect 37240 16396 37246 16448
rect 37737 16439 37795 16445
rect 37737 16405 37749 16439
rect 37783 16436 37795 16439
rect 38562 16436 38568 16448
rect 37783 16408 38568 16436
rect 37783 16405 37795 16408
rect 37737 16399 37795 16405
rect 38562 16396 38568 16408
rect 38620 16396 38626 16448
rect 40773 16439 40831 16445
rect 40773 16405 40785 16439
rect 40819 16436 40831 16439
rect 40954 16436 40960 16448
rect 40819 16408 40960 16436
rect 40819 16405 40831 16408
rect 40773 16399 40831 16405
rect 40954 16396 40960 16408
rect 41012 16396 41018 16448
rect 49142 16396 49148 16448
rect 49200 16396 49206 16448
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 8294 16192 8300 16244
rect 8352 16192 8358 16244
rect 9214 16192 9220 16244
rect 9272 16192 9278 16244
rect 9766 16192 9772 16244
rect 9824 16232 9830 16244
rect 10965 16235 11023 16241
rect 10965 16232 10977 16235
rect 9824 16204 10977 16232
rect 9824 16192 9830 16204
rect 10965 16201 10977 16204
rect 11011 16201 11023 16235
rect 10965 16195 11023 16201
rect 11054 16192 11060 16244
rect 11112 16192 11118 16244
rect 11330 16192 11336 16244
rect 11388 16232 11394 16244
rect 11977 16235 12035 16241
rect 11977 16232 11989 16235
rect 11388 16204 11989 16232
rect 11388 16192 11394 16204
rect 11977 16201 11989 16204
rect 12023 16201 12035 16235
rect 11977 16195 12035 16201
rect 12437 16235 12495 16241
rect 12437 16201 12449 16235
rect 12483 16232 12495 16235
rect 13173 16235 13231 16241
rect 13173 16232 13185 16235
rect 12483 16204 13185 16232
rect 12483 16201 12495 16204
rect 12437 16195 12495 16201
rect 13173 16201 13185 16204
rect 13219 16201 13231 16235
rect 13173 16195 13231 16201
rect 13630 16192 13636 16244
rect 13688 16192 13694 16244
rect 14369 16235 14427 16241
rect 14369 16201 14381 16235
rect 14415 16201 14427 16235
rect 14369 16195 14427 16201
rect 10870 16164 10876 16176
rect 2976 16136 10876 16164
rect 2976 16105 3004 16136
rect 10870 16124 10876 16136
rect 10928 16124 10934 16176
rect 11072 16164 11100 16192
rect 13541 16167 13599 16173
rect 11072 16136 12296 16164
rect 2961 16099 3019 16105
rect 2961 16065 2973 16099
rect 3007 16065 3019 16099
rect 2961 16059 3019 16065
rect 4246 16056 4252 16108
rect 4304 16096 4310 16108
rect 8205 16099 8263 16105
rect 8205 16096 8217 16099
rect 4304 16068 8217 16096
rect 4304 16056 4310 16068
rect 8205 16065 8217 16068
rect 8251 16065 8263 16099
rect 8205 16059 8263 16065
rect 9309 16099 9367 16105
rect 9309 16065 9321 16099
rect 9355 16065 9367 16099
rect 9309 16059 9367 16065
rect 10413 16099 10471 16105
rect 10413 16065 10425 16099
rect 10459 16096 10471 16099
rect 11057 16099 11115 16105
rect 11057 16096 11069 16099
rect 10459 16068 11069 16096
rect 10459 16065 10471 16068
rect 10413 16059 10471 16065
rect 11057 16065 11069 16068
rect 11103 16096 11115 16099
rect 12158 16096 12164 16108
rect 11103 16068 12164 16096
rect 11103 16065 11115 16068
rect 11057 16059 11115 16065
rect 1026 15988 1032 16040
rect 1084 16028 1090 16040
rect 1765 16031 1823 16037
rect 1765 16028 1777 16031
rect 1084 16000 1777 16028
rect 1084 15988 1090 16000
rect 1765 15997 1777 16000
rect 1811 15997 1823 16031
rect 1765 15991 1823 15997
rect 8113 16031 8171 16037
rect 8113 15997 8125 16031
rect 8159 16028 8171 16031
rect 9030 16028 9036 16040
rect 8159 16000 9036 16028
rect 8159 15997 8171 16000
rect 8113 15991 8171 15997
rect 9030 15988 9036 16000
rect 9088 15988 9094 16040
rect 9324 16028 9352 16059
rect 12158 16056 12164 16068
rect 12216 16056 12222 16108
rect 12268 16028 12296 16136
rect 13541 16133 13553 16167
rect 13587 16164 13599 16167
rect 14384 16164 14412 16195
rect 15838 16192 15844 16244
rect 15896 16232 15902 16244
rect 15933 16235 15991 16241
rect 15933 16232 15945 16235
rect 15896 16204 15945 16232
rect 15896 16192 15902 16204
rect 15933 16201 15945 16204
rect 15979 16201 15991 16235
rect 17405 16235 17463 16241
rect 17405 16232 17417 16235
rect 15933 16195 15991 16201
rect 16040 16204 17417 16232
rect 13587 16136 14412 16164
rect 13587 16133 13599 16136
rect 13541 16127 13599 16133
rect 15010 16124 15016 16176
rect 15068 16164 15074 16176
rect 16040 16164 16068 16204
rect 17405 16201 17417 16204
rect 17451 16201 17463 16235
rect 17405 16195 17463 16201
rect 17773 16235 17831 16241
rect 17773 16201 17785 16235
rect 17819 16232 17831 16235
rect 18322 16232 18328 16244
rect 17819 16204 18328 16232
rect 17819 16201 17831 16204
rect 17773 16195 17831 16201
rect 18322 16192 18328 16204
rect 18380 16192 18386 16244
rect 18690 16192 18696 16244
rect 18748 16232 18754 16244
rect 18785 16235 18843 16241
rect 18785 16232 18797 16235
rect 18748 16204 18797 16232
rect 18748 16192 18754 16204
rect 18785 16201 18797 16204
rect 18831 16201 18843 16235
rect 18785 16195 18843 16201
rect 21266 16192 21272 16244
rect 21324 16232 21330 16244
rect 21450 16232 21456 16244
rect 21324 16204 21456 16232
rect 21324 16192 21330 16204
rect 21450 16192 21456 16204
rect 21508 16192 21514 16244
rect 22646 16192 22652 16244
rect 22704 16232 22710 16244
rect 22833 16235 22891 16241
rect 22833 16232 22845 16235
rect 22704 16204 22845 16232
rect 22704 16192 22710 16204
rect 22833 16201 22845 16204
rect 22879 16232 22891 16235
rect 23382 16232 23388 16244
rect 22879 16204 23388 16232
rect 22879 16201 22891 16204
rect 22833 16195 22891 16201
rect 23382 16192 23388 16204
rect 23440 16192 23446 16244
rect 23845 16235 23903 16241
rect 23845 16201 23857 16235
rect 23891 16232 23903 16235
rect 24670 16232 24676 16244
rect 23891 16204 24676 16232
rect 23891 16201 23903 16204
rect 23845 16195 23903 16201
rect 24670 16192 24676 16204
rect 24728 16192 24734 16244
rect 24762 16192 24768 16244
rect 24820 16232 24826 16244
rect 26602 16232 26608 16244
rect 24820 16204 26608 16232
rect 24820 16192 24826 16204
rect 26602 16192 26608 16204
rect 26660 16192 26666 16244
rect 26697 16235 26755 16241
rect 26697 16201 26709 16235
rect 26743 16232 26755 16235
rect 26786 16232 26792 16244
rect 26743 16204 26792 16232
rect 26743 16201 26755 16204
rect 26697 16195 26755 16201
rect 26786 16192 26792 16204
rect 26844 16192 26850 16244
rect 26970 16192 26976 16244
rect 27028 16232 27034 16244
rect 27430 16232 27436 16244
rect 27028 16204 27436 16232
rect 27028 16192 27034 16204
rect 27430 16192 27436 16204
rect 27488 16232 27494 16244
rect 27525 16235 27583 16241
rect 27525 16232 27537 16235
rect 27488 16204 27537 16232
rect 27488 16192 27494 16204
rect 27525 16201 27537 16204
rect 27571 16201 27583 16235
rect 27525 16195 27583 16201
rect 27617 16235 27675 16241
rect 27617 16201 27629 16235
rect 27663 16232 27675 16235
rect 28350 16232 28356 16244
rect 27663 16204 28356 16232
rect 27663 16201 27675 16204
rect 27617 16195 27675 16201
rect 28350 16192 28356 16204
rect 28408 16192 28414 16244
rect 30558 16192 30564 16244
rect 30616 16232 30622 16244
rect 30929 16235 30987 16241
rect 30929 16232 30941 16235
rect 30616 16204 30941 16232
rect 30616 16192 30622 16204
rect 30929 16201 30941 16204
rect 30975 16201 30987 16235
rect 30929 16195 30987 16201
rect 32030 16192 32036 16244
rect 32088 16232 32094 16244
rect 32950 16232 32956 16244
rect 32088 16204 32956 16232
rect 32088 16192 32094 16204
rect 32950 16192 32956 16204
rect 33008 16232 33014 16244
rect 33686 16232 33692 16244
rect 33008 16204 33692 16232
rect 33008 16192 33014 16204
rect 33686 16192 33692 16204
rect 33744 16192 33750 16244
rect 33778 16192 33784 16244
rect 33836 16192 33842 16244
rect 34790 16192 34796 16244
rect 34848 16232 34854 16244
rect 34848 16204 36952 16232
rect 34848 16192 34854 16204
rect 15068 16136 16068 16164
rect 15068 16124 15074 16136
rect 17126 16124 17132 16176
rect 17184 16164 17190 16176
rect 19429 16167 19487 16173
rect 19429 16164 19441 16167
rect 17184 16136 19441 16164
rect 17184 16124 17190 16136
rect 12345 16099 12403 16105
rect 12345 16065 12357 16099
rect 12391 16096 12403 16099
rect 14458 16096 14464 16108
rect 12391 16068 14464 16096
rect 12391 16065 12403 16068
rect 12345 16059 12403 16065
rect 14458 16056 14464 16068
rect 14516 16056 14522 16108
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16065 14795 16099
rect 14737 16059 14795 16065
rect 14829 16099 14887 16105
rect 14829 16065 14841 16099
rect 14875 16096 14887 16099
rect 15286 16096 15292 16108
rect 14875 16068 15292 16096
rect 14875 16065 14887 16068
rect 14829 16059 14887 16065
rect 12621 16031 12679 16037
rect 12621 16028 12633 16031
rect 9324 16000 11836 16028
rect 12268 16000 12633 16028
rect 8665 15963 8723 15969
rect 8665 15929 8677 15963
rect 8711 15960 8723 15963
rect 9766 15960 9772 15972
rect 8711 15932 9772 15960
rect 8711 15929 8723 15932
rect 8665 15923 8723 15929
rect 9766 15920 9772 15932
rect 9824 15920 9830 15972
rect 9858 15852 9864 15904
rect 9916 15892 9922 15904
rect 10505 15895 10563 15901
rect 10505 15892 10517 15895
rect 9916 15864 10517 15892
rect 9916 15852 9922 15864
rect 10505 15861 10517 15864
rect 10551 15892 10563 15895
rect 10594 15892 10600 15904
rect 10551 15864 10600 15892
rect 10551 15861 10563 15864
rect 10505 15855 10563 15861
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 11514 15852 11520 15904
rect 11572 15892 11578 15904
rect 11609 15895 11667 15901
rect 11609 15892 11621 15895
rect 11572 15864 11621 15892
rect 11572 15852 11578 15864
rect 11609 15861 11621 15864
rect 11655 15861 11667 15895
rect 11808 15892 11836 16000
rect 12621 15997 12633 16000
rect 12667 16028 12679 16031
rect 13630 16028 13636 16040
rect 12667 16000 13636 16028
rect 12667 15997 12679 16000
rect 12621 15991 12679 15997
rect 13630 15988 13636 16000
rect 13688 15988 13694 16040
rect 13817 16031 13875 16037
rect 13817 15997 13829 16031
rect 13863 16028 13875 16031
rect 14274 16028 14280 16040
rect 13863 16000 14280 16028
rect 13863 15997 13875 16000
rect 13817 15991 13875 15997
rect 14274 15988 14280 16000
rect 14332 15988 14338 16040
rect 13538 15920 13544 15972
rect 13596 15960 13602 15972
rect 14752 15960 14780 16059
rect 15286 16056 15292 16068
rect 15344 16056 15350 16108
rect 15378 16056 15384 16108
rect 15436 16096 15442 16108
rect 16114 16096 16120 16108
rect 15436 16068 16120 16096
rect 15436 16056 15442 16068
rect 14918 15988 14924 16040
rect 14976 15988 14982 16040
rect 15764 16037 15792 16068
rect 16114 16056 16120 16068
rect 16172 16096 16178 16108
rect 16172 16068 17724 16096
rect 16172 16056 16178 16068
rect 15749 16031 15807 16037
rect 15749 15997 15761 16031
rect 15795 15997 15807 16031
rect 15749 15991 15807 15997
rect 15838 15988 15844 16040
rect 15896 15988 15902 16040
rect 16761 16031 16819 16037
rect 16761 15997 16773 16031
rect 16807 16028 16819 16031
rect 17126 16028 17132 16040
rect 16807 16000 17132 16028
rect 16807 15997 16819 16000
rect 16761 15991 16819 15997
rect 17126 15988 17132 16000
rect 17184 15988 17190 16040
rect 15930 15960 15936 15972
rect 13596 15932 15936 15960
rect 13596 15920 13602 15932
rect 15930 15920 15936 15932
rect 15988 15920 15994 15972
rect 16301 15963 16359 15969
rect 16301 15929 16313 15963
rect 16347 15960 16359 15963
rect 17586 15960 17592 15972
rect 16347 15932 17592 15960
rect 16347 15929 16359 15932
rect 16301 15923 16359 15929
rect 17586 15920 17592 15932
rect 17644 15920 17650 15972
rect 16390 15892 16396 15904
rect 11808 15864 16396 15892
rect 11609 15855 11667 15861
rect 16390 15852 16396 15864
rect 16448 15852 16454 15904
rect 16942 15852 16948 15904
rect 17000 15852 17006 15904
rect 17129 15895 17187 15901
rect 17129 15861 17141 15895
rect 17175 15892 17187 15895
rect 17218 15892 17224 15904
rect 17175 15864 17224 15892
rect 17175 15861 17187 15864
rect 17129 15855 17187 15861
rect 17218 15852 17224 15864
rect 17276 15852 17282 15904
rect 17696 15892 17724 16068
rect 17972 16037 18000 16136
rect 19429 16133 19441 16136
rect 19475 16133 19487 16167
rect 20806 16164 20812 16176
rect 20654 16136 20812 16164
rect 19429 16127 19487 16133
rect 20806 16124 20812 16136
rect 20864 16124 20870 16176
rect 20898 16124 20904 16176
rect 20956 16164 20962 16176
rect 20956 16136 21404 16164
rect 20956 16124 20962 16136
rect 19150 16056 19156 16108
rect 19208 16056 19214 16108
rect 21376 16096 21404 16136
rect 21542 16124 21548 16176
rect 21600 16164 21606 16176
rect 21910 16164 21916 16176
rect 21600 16136 21916 16164
rect 21600 16124 21606 16136
rect 21910 16124 21916 16136
rect 21968 16124 21974 16176
rect 25774 16164 25780 16176
rect 25622 16136 25780 16164
rect 25774 16124 25780 16136
rect 25832 16124 25838 16176
rect 27798 16124 27804 16176
rect 27856 16164 27862 16176
rect 28902 16164 28908 16176
rect 27856 16136 28908 16164
rect 27856 16124 27862 16136
rect 22922 16096 22928 16108
rect 21376 16068 22928 16096
rect 22922 16056 22928 16068
rect 22980 16056 22986 16108
rect 23474 16056 23480 16108
rect 23532 16056 23538 16108
rect 26329 16099 26387 16105
rect 26329 16065 26341 16099
rect 26375 16096 26387 16099
rect 27816 16096 27844 16124
rect 28368 16105 28396 16136
rect 28902 16124 28908 16136
rect 28960 16124 28966 16176
rect 29178 16124 29184 16176
rect 29236 16124 29242 16176
rect 29914 16124 29920 16176
rect 29972 16164 29978 16176
rect 30650 16164 30656 16176
rect 29972 16136 30656 16164
rect 29972 16124 29978 16136
rect 30650 16124 30656 16136
rect 30708 16124 30714 16176
rect 30834 16124 30840 16176
rect 30892 16124 30898 16176
rect 31662 16124 31668 16176
rect 31720 16164 31726 16176
rect 33873 16167 33931 16173
rect 33873 16164 33885 16167
rect 31720 16136 33885 16164
rect 31720 16124 31726 16136
rect 33873 16133 33885 16136
rect 33919 16133 33931 16167
rect 33873 16127 33931 16133
rect 26375 16068 27844 16096
rect 28353 16099 28411 16105
rect 26375 16065 26387 16068
rect 26329 16059 26387 16065
rect 28353 16065 28365 16099
rect 28399 16065 28411 16099
rect 32677 16099 32735 16105
rect 28353 16059 28411 16065
rect 30760 16068 32628 16096
rect 17865 16031 17923 16037
rect 17865 15997 17877 16031
rect 17911 15997 17923 16031
rect 17865 15991 17923 15997
rect 17957 16031 18015 16037
rect 17957 15997 17969 16031
rect 18003 15997 18015 16031
rect 19978 16028 19984 16040
rect 17957 15991 18015 15997
rect 18064 16000 19984 16028
rect 17880 15960 17908 15991
rect 18064 15960 18092 16000
rect 19978 15988 19984 16000
rect 20036 15988 20042 16040
rect 20901 16031 20959 16037
rect 20901 15997 20913 16031
rect 20947 16028 20959 16031
rect 20990 16028 20996 16040
rect 20947 16000 20996 16028
rect 20947 15997 20959 16000
rect 20901 15991 20959 15997
rect 20990 15988 20996 16000
rect 21048 16028 21054 16040
rect 21910 16028 21916 16040
rect 21048 16000 21916 16028
rect 21048 15988 21054 16000
rect 21910 15988 21916 16000
rect 21968 15988 21974 16040
rect 23293 16031 23351 16037
rect 23293 15997 23305 16031
rect 23339 15997 23351 16031
rect 23293 15991 23351 15997
rect 17880 15932 18092 15960
rect 20438 15920 20444 15972
rect 20496 15960 20502 15972
rect 22094 15960 22100 15972
rect 20496 15932 22100 15960
rect 20496 15920 20502 15932
rect 22094 15920 22100 15932
rect 22152 15920 22158 15972
rect 23308 15960 23336 15991
rect 23382 15988 23388 16040
rect 23440 15988 23446 16040
rect 24486 15988 24492 16040
rect 24544 16028 24550 16040
rect 24581 16031 24639 16037
rect 24581 16028 24593 16031
rect 24544 16000 24593 16028
rect 24544 15988 24550 16000
rect 24581 15997 24593 16000
rect 24627 15997 24639 16031
rect 24581 15991 24639 15997
rect 26050 15988 26056 16040
rect 26108 15988 26114 16040
rect 26878 15988 26884 16040
rect 26936 16028 26942 16040
rect 27709 16031 27767 16037
rect 27709 16028 27721 16031
rect 26936 16000 27721 16028
rect 26936 15988 26942 16000
rect 27709 15997 27721 16000
rect 27755 15997 27767 16031
rect 27709 15991 27767 15997
rect 28626 15988 28632 16040
rect 28684 15988 28690 16040
rect 29822 15988 29828 16040
rect 29880 16028 29886 16040
rect 30653 16031 30711 16037
rect 30653 16028 30665 16031
rect 29880 16000 30665 16028
rect 29880 15988 29886 16000
rect 30653 15997 30665 16000
rect 30699 15997 30711 16031
rect 30653 15991 30711 15997
rect 24504 15960 24532 15988
rect 30760 15960 30788 16068
rect 31202 15988 31208 16040
rect 31260 16028 31266 16040
rect 31260 16000 32168 16028
rect 31260 15988 31266 16000
rect 31573 15963 31631 15969
rect 31573 15960 31585 15963
rect 23308 15932 24532 15960
rect 29656 15932 30788 15960
rect 31220 15932 31585 15960
rect 18414 15892 18420 15904
rect 17696 15864 18420 15892
rect 18414 15852 18420 15864
rect 18472 15852 18478 15904
rect 20806 15852 20812 15904
rect 20864 15892 20870 15904
rect 21361 15895 21419 15901
rect 21361 15892 21373 15895
rect 20864 15864 21373 15892
rect 20864 15852 20870 15864
rect 21361 15861 21373 15864
rect 21407 15892 21419 15895
rect 22002 15892 22008 15904
rect 21407 15864 22008 15892
rect 21407 15861 21419 15864
rect 21361 15855 21419 15861
rect 22002 15852 22008 15864
rect 22060 15852 22066 15904
rect 26694 15852 26700 15904
rect 26752 15892 26758 15904
rect 27157 15895 27215 15901
rect 27157 15892 27169 15895
rect 26752 15864 27169 15892
rect 26752 15852 26758 15864
rect 27157 15861 27169 15864
rect 27203 15861 27215 15895
rect 27157 15855 27215 15861
rect 27246 15852 27252 15904
rect 27304 15892 27310 15904
rect 29656 15892 29684 15932
rect 31220 15904 31248 15932
rect 31573 15929 31585 15932
rect 31619 15960 31631 15963
rect 32030 15960 32036 15972
rect 31619 15932 32036 15960
rect 31619 15929 31631 15932
rect 31573 15923 31631 15929
rect 32030 15920 32036 15932
rect 32088 15920 32094 15972
rect 27304 15864 29684 15892
rect 30101 15895 30159 15901
rect 27304 15852 27310 15864
rect 30101 15861 30113 15895
rect 30147 15892 30159 15895
rect 30742 15892 30748 15904
rect 30147 15864 30748 15892
rect 30147 15861 30159 15864
rect 30101 15855 30159 15861
rect 30742 15852 30748 15864
rect 30800 15852 30806 15904
rect 31202 15852 31208 15904
rect 31260 15852 31266 15904
rect 31297 15895 31355 15901
rect 31297 15861 31309 15895
rect 31343 15892 31355 15895
rect 31478 15892 31484 15904
rect 31343 15864 31484 15892
rect 31343 15861 31355 15864
rect 31297 15855 31355 15861
rect 31478 15852 31484 15864
rect 31536 15852 31542 15904
rect 31849 15895 31907 15901
rect 31849 15861 31861 15895
rect 31895 15892 31907 15895
rect 32140 15892 32168 16000
rect 32398 15988 32404 16040
rect 32456 15988 32462 16040
rect 32600 16037 32628 16068
rect 32677 16065 32689 16099
rect 32723 16096 32735 16099
rect 33318 16096 33324 16108
rect 32723 16068 33324 16096
rect 32723 16065 32735 16068
rect 32677 16059 32735 16065
rect 33318 16056 33324 16068
rect 33376 16096 33382 16108
rect 33376 16068 34468 16096
rect 33376 16056 33382 16068
rect 34440 16040 34468 16068
rect 35526 16056 35532 16108
rect 35584 16056 35590 16108
rect 36924 16105 36952 16204
rect 37090 16192 37096 16244
rect 37148 16232 37154 16244
rect 40497 16235 40555 16241
rect 40497 16232 40509 16235
rect 37148 16204 40509 16232
rect 37148 16192 37154 16204
rect 40497 16201 40509 16204
rect 40543 16201 40555 16235
rect 40497 16195 40555 16201
rect 40954 16192 40960 16244
rect 41012 16192 41018 16244
rect 41414 16192 41420 16244
rect 41472 16232 41478 16244
rect 41509 16235 41567 16241
rect 41509 16232 41521 16235
rect 41472 16204 41521 16232
rect 41472 16192 41478 16204
rect 41509 16201 41521 16204
rect 41555 16201 41567 16235
rect 41509 16195 41567 16201
rect 38473 16167 38531 16173
rect 38473 16133 38485 16167
rect 38519 16164 38531 16167
rect 38562 16164 38568 16176
rect 38519 16136 38568 16164
rect 38519 16133 38531 16136
rect 38473 16127 38531 16133
rect 38562 16124 38568 16136
rect 38620 16124 38626 16176
rect 39942 16164 39948 16176
rect 39698 16136 39948 16164
rect 39942 16124 39948 16136
rect 40000 16124 40006 16176
rect 36909 16099 36967 16105
rect 36909 16065 36921 16099
rect 36955 16096 36967 16099
rect 37366 16096 37372 16108
rect 36955 16068 37372 16096
rect 36955 16065 36967 16068
rect 36909 16059 36967 16065
rect 37366 16056 37372 16068
rect 37424 16096 37430 16108
rect 38197 16099 38255 16105
rect 38197 16096 38209 16099
rect 37424 16068 38209 16096
rect 37424 16056 37430 16068
rect 38197 16065 38209 16068
rect 38243 16065 38255 16099
rect 38197 16059 38255 16065
rect 40865 16099 40923 16105
rect 40865 16065 40877 16099
rect 40911 16096 40923 16099
rect 48682 16096 48688 16108
rect 40911 16068 48688 16096
rect 40911 16065 40923 16068
rect 40865 16059 40923 16065
rect 48682 16056 48688 16068
rect 48740 16056 48746 16108
rect 48777 16099 48835 16105
rect 48777 16065 48789 16099
rect 48823 16096 48835 16099
rect 49326 16096 49332 16108
rect 48823 16068 49332 16096
rect 48823 16065 48835 16068
rect 48777 16059 48835 16065
rect 49326 16056 49332 16068
rect 49384 16056 49390 16108
rect 32585 16031 32643 16037
rect 32585 15997 32597 16031
rect 32631 15997 32643 16031
rect 32585 15991 32643 15997
rect 32600 15960 32628 15991
rect 32766 15988 32772 16040
rect 32824 16028 32830 16040
rect 33597 16031 33655 16037
rect 33597 16028 33609 16031
rect 32824 16000 33609 16028
rect 32824 15988 32830 16000
rect 33597 15997 33609 16000
rect 33643 15997 33655 16031
rect 33597 15991 33655 15997
rect 34422 15988 34428 16040
rect 34480 16028 34486 16040
rect 34701 16031 34759 16037
rect 34701 16028 34713 16031
rect 34480 16000 34713 16028
rect 34480 15988 34486 16000
rect 34701 15997 34713 16000
rect 34747 15997 34759 16031
rect 34701 15991 34759 15997
rect 35158 15988 35164 16040
rect 35216 16028 35222 16040
rect 36078 16028 36084 16040
rect 35216 16000 36084 16028
rect 35216 15988 35222 16000
rect 36078 15988 36084 16000
rect 36136 15988 36142 16040
rect 36633 16031 36691 16037
rect 36633 15997 36645 16031
rect 36679 16028 36691 16031
rect 36679 16000 36952 16028
rect 36679 15997 36691 16000
rect 36633 15991 36691 15997
rect 34517 15963 34575 15969
rect 34517 15960 34529 15963
rect 32600 15932 34529 15960
rect 34517 15929 34529 15932
rect 34563 15929 34575 15963
rect 36924 15960 36952 16000
rect 36998 15988 37004 16040
rect 37056 16028 37062 16040
rect 37461 16031 37519 16037
rect 37461 16028 37473 16031
rect 37056 16000 37473 16028
rect 37056 15988 37062 16000
rect 37461 15997 37473 16000
rect 37507 15997 37519 16031
rect 37461 15991 37519 15997
rect 39206 15988 39212 16040
rect 39264 16028 39270 16040
rect 41049 16031 41107 16037
rect 41049 16028 41061 16031
rect 39264 16000 41061 16028
rect 39264 15988 39270 16000
rect 41049 15997 41061 16000
rect 41095 16028 41107 16031
rect 41782 16028 41788 16040
rect 41095 16000 41788 16028
rect 41095 15997 41107 16000
rect 41049 15991 41107 15997
rect 41782 15988 41788 16000
rect 41840 15988 41846 16040
rect 37274 15960 37280 15972
rect 34517 15923 34575 15929
rect 34624 15932 35664 15960
rect 36924 15932 37280 15960
rect 32766 15892 32772 15904
rect 31895 15864 32772 15892
rect 31895 15861 31907 15864
rect 31849 15855 31907 15861
rect 32766 15852 32772 15864
rect 32824 15852 32830 15904
rect 32858 15852 32864 15904
rect 32916 15892 32922 15904
rect 33045 15895 33103 15901
rect 33045 15892 33057 15895
rect 32916 15864 33057 15892
rect 32916 15852 32922 15864
rect 33045 15861 33057 15864
rect 33091 15861 33103 15895
rect 33045 15855 33103 15861
rect 34241 15895 34299 15901
rect 34241 15861 34253 15895
rect 34287 15892 34299 15895
rect 34624 15892 34652 15932
rect 34287 15864 34652 15892
rect 35636 15892 35664 15932
rect 37274 15920 37280 15932
rect 37332 15920 37338 15972
rect 49142 15920 49148 15972
rect 49200 15920 49206 15972
rect 38562 15892 38568 15904
rect 35636 15864 38568 15892
rect 34287 15861 34299 15864
rect 34241 15855 34299 15861
rect 38562 15852 38568 15864
rect 38620 15852 38626 15904
rect 39945 15895 40003 15901
rect 39945 15861 39957 15895
rect 39991 15892 40003 15895
rect 40310 15892 40316 15904
rect 39991 15864 40316 15892
rect 39991 15861 40003 15864
rect 39945 15855 40003 15861
rect 40310 15852 40316 15864
rect 40368 15852 40374 15904
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 10686 15648 10692 15700
rect 10744 15688 10750 15700
rect 10781 15691 10839 15697
rect 10781 15688 10793 15691
rect 10744 15660 10793 15688
rect 10744 15648 10750 15660
rect 10781 15657 10793 15660
rect 10827 15657 10839 15691
rect 10781 15651 10839 15657
rect 11514 15648 11520 15700
rect 11572 15688 11578 15700
rect 15286 15688 15292 15700
rect 11572 15660 15292 15688
rect 11572 15648 11578 15660
rect 15286 15648 15292 15660
rect 15344 15648 15350 15700
rect 16758 15648 16764 15700
rect 16816 15648 16822 15700
rect 17310 15648 17316 15700
rect 17368 15688 17374 15700
rect 17865 15691 17923 15697
rect 17865 15688 17877 15691
rect 17368 15660 17877 15688
rect 17368 15648 17374 15660
rect 17865 15657 17877 15660
rect 17911 15688 17923 15691
rect 20806 15688 20812 15700
rect 17911 15660 20812 15688
rect 17911 15657 17923 15660
rect 17865 15651 17923 15657
rect 20806 15648 20812 15660
rect 20864 15648 20870 15700
rect 22462 15648 22468 15700
rect 22520 15648 22526 15700
rect 22554 15648 22560 15700
rect 22612 15688 22618 15700
rect 32217 15691 32275 15697
rect 22612 15660 31800 15688
rect 22612 15648 22618 15660
rect 14274 15620 14280 15632
rect 12452 15592 14280 15620
rect 10505 15555 10563 15561
rect 10505 15521 10517 15555
rect 10551 15552 10563 15555
rect 11054 15552 11060 15564
rect 10551 15524 11060 15552
rect 10551 15521 10563 15524
rect 10505 15515 10563 15521
rect 11054 15512 11060 15524
rect 11112 15512 11118 15564
rect 12253 15555 12311 15561
rect 12253 15521 12265 15555
rect 12299 15552 12311 15555
rect 12452 15552 12480 15592
rect 14274 15580 14280 15592
rect 14332 15580 14338 15632
rect 17494 15580 17500 15632
rect 17552 15620 17558 15632
rect 18049 15623 18107 15629
rect 18049 15620 18061 15623
rect 17552 15592 18061 15620
rect 17552 15580 17558 15592
rect 18049 15589 18061 15592
rect 18095 15620 18107 15623
rect 18598 15620 18604 15632
rect 18095 15592 18604 15620
rect 18095 15589 18107 15592
rect 18049 15583 18107 15589
rect 18598 15580 18604 15592
rect 18656 15580 18662 15632
rect 18966 15580 18972 15632
rect 19024 15580 19030 15632
rect 19334 15580 19340 15632
rect 19392 15620 19398 15632
rect 19889 15623 19947 15629
rect 19889 15620 19901 15623
rect 19392 15592 19901 15620
rect 19392 15580 19398 15592
rect 19889 15589 19901 15592
rect 19935 15589 19947 15623
rect 22094 15620 22100 15632
rect 19889 15583 19947 15589
rect 20364 15592 22100 15620
rect 12299 15524 12480 15552
rect 12299 15521 12311 15524
rect 12253 15515 12311 15521
rect 12526 15512 12532 15564
rect 12584 15512 12590 15564
rect 13173 15555 13231 15561
rect 13173 15521 13185 15555
rect 13219 15552 13231 15555
rect 14090 15552 14096 15564
rect 13219 15524 14096 15552
rect 13219 15521 13231 15524
rect 13173 15515 13231 15521
rect 14090 15512 14096 15524
rect 14148 15512 14154 15564
rect 14918 15512 14924 15564
rect 14976 15512 14982 15564
rect 16114 15512 16120 15564
rect 16172 15512 16178 15564
rect 16206 15512 16212 15564
rect 16264 15552 16270 15564
rect 16482 15552 16488 15564
rect 16264 15524 16488 15552
rect 16264 15512 16270 15524
rect 16482 15512 16488 15524
rect 16540 15552 16546 15564
rect 17313 15555 17371 15561
rect 17313 15552 17325 15555
rect 16540 15524 17325 15552
rect 16540 15512 16546 15524
rect 17313 15521 17325 15524
rect 17359 15521 17371 15555
rect 17313 15515 17371 15521
rect 19245 15555 19303 15561
rect 19245 15521 19257 15555
rect 19291 15552 19303 15555
rect 19518 15552 19524 15564
rect 19291 15524 19524 15552
rect 19291 15521 19303 15524
rect 19245 15515 19303 15521
rect 19518 15512 19524 15524
rect 19576 15512 19582 15564
rect 20364 15561 20392 15592
rect 22094 15580 22100 15592
rect 22152 15580 22158 15632
rect 24026 15580 24032 15632
rect 24084 15620 24090 15632
rect 27433 15623 27491 15629
rect 27433 15620 27445 15623
rect 24084 15592 27445 15620
rect 24084 15580 24090 15592
rect 27433 15589 27445 15592
rect 27479 15589 27491 15623
rect 27433 15583 27491 15589
rect 29178 15580 29184 15632
rect 29236 15620 29242 15632
rect 29273 15623 29331 15629
rect 29273 15620 29285 15623
rect 29236 15592 29285 15620
rect 29236 15580 29242 15592
rect 29273 15589 29285 15592
rect 29319 15589 29331 15623
rect 29273 15583 29331 15589
rect 20349 15555 20407 15561
rect 20349 15521 20361 15555
rect 20395 15521 20407 15555
rect 20349 15515 20407 15521
rect 20533 15555 20591 15561
rect 20533 15521 20545 15555
rect 20579 15552 20591 15555
rect 21266 15552 21272 15564
rect 20579 15524 21272 15552
rect 20579 15521 20591 15524
rect 20533 15515 20591 15521
rect 21266 15512 21272 15524
rect 21324 15512 21330 15564
rect 21450 15512 21456 15564
rect 21508 15552 21514 15564
rect 21729 15555 21787 15561
rect 21729 15552 21741 15555
rect 21508 15524 21741 15552
rect 21508 15512 21514 15524
rect 21729 15521 21741 15524
rect 21775 15521 21787 15555
rect 21729 15515 21787 15521
rect 22002 15512 22008 15564
rect 22060 15552 22066 15564
rect 23661 15555 23719 15561
rect 23661 15552 23673 15555
rect 22060 15524 23673 15552
rect 22060 15512 22066 15524
rect 23661 15521 23673 15524
rect 23707 15521 23719 15555
rect 23661 15515 23719 15521
rect 24762 15512 24768 15564
rect 24820 15552 24826 15564
rect 25225 15555 25283 15561
rect 25225 15552 25237 15555
rect 24820 15524 25237 15552
rect 24820 15512 24826 15524
rect 25225 15521 25237 15524
rect 25271 15521 25283 15555
rect 25225 15515 25283 15521
rect 25314 15512 25320 15564
rect 25372 15552 25378 15564
rect 26421 15555 26479 15561
rect 26421 15552 26433 15555
rect 25372 15524 26433 15552
rect 25372 15512 25378 15524
rect 26421 15521 26433 15524
rect 26467 15521 26479 15555
rect 26421 15515 26479 15521
rect 26602 15512 26608 15564
rect 26660 15552 26666 15564
rect 27985 15555 28043 15561
rect 27985 15552 27997 15555
rect 26660 15524 27997 15552
rect 26660 15512 26666 15524
rect 27985 15521 27997 15524
rect 28031 15521 28043 15555
rect 27985 15515 28043 15521
rect 28718 15512 28724 15564
rect 28776 15512 28782 15564
rect 30469 15555 30527 15561
rect 30469 15521 30481 15555
rect 30515 15552 30527 15555
rect 31110 15552 31116 15564
rect 30515 15524 31116 15552
rect 30515 15521 30527 15524
rect 30469 15515 30527 15521
rect 31110 15512 31116 15524
rect 31168 15512 31174 15564
rect 31772 15552 31800 15660
rect 32217 15657 32229 15691
rect 32263 15688 32275 15691
rect 32582 15688 32588 15700
rect 32263 15660 32588 15688
rect 32263 15657 32275 15660
rect 32217 15651 32275 15657
rect 32582 15648 32588 15660
rect 32640 15648 32646 15700
rect 33686 15648 33692 15700
rect 33744 15688 33750 15700
rect 34333 15691 34391 15697
rect 34333 15688 34345 15691
rect 33744 15660 34345 15688
rect 33744 15648 33750 15660
rect 34333 15657 34345 15660
rect 34379 15688 34391 15691
rect 35526 15688 35532 15700
rect 34379 15660 35532 15688
rect 34379 15657 34391 15660
rect 34333 15651 34391 15657
rect 35526 15648 35532 15660
rect 35584 15648 35590 15700
rect 36633 15691 36691 15697
rect 36633 15657 36645 15691
rect 36679 15688 36691 15691
rect 37274 15688 37280 15700
rect 36679 15660 37280 15688
rect 36679 15657 36691 15660
rect 36633 15651 36691 15657
rect 37274 15648 37280 15660
rect 37332 15648 37338 15700
rect 37734 15648 37740 15700
rect 37792 15648 37798 15700
rect 41414 15648 41420 15700
rect 41472 15688 41478 15700
rect 42061 15691 42119 15697
rect 42061 15688 42073 15691
rect 41472 15660 42073 15688
rect 41472 15648 41478 15660
rect 42061 15657 42073 15660
rect 42107 15657 42119 15691
rect 42061 15651 42119 15657
rect 48682 15648 48688 15700
rect 48740 15688 48746 15700
rect 49145 15691 49203 15697
rect 49145 15688 49157 15691
rect 48740 15660 49157 15688
rect 48740 15648 48746 15660
rect 49145 15657 49157 15660
rect 49191 15657 49203 15691
rect 49145 15651 49203 15657
rect 31846 15580 31852 15632
rect 31904 15620 31910 15632
rect 31904 15592 32996 15620
rect 31904 15580 31910 15592
rect 32968 15561 32996 15592
rect 41782 15580 41788 15632
rect 41840 15580 41846 15632
rect 32861 15555 32919 15561
rect 31772 15524 32812 15552
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 10226 15484 10232 15496
rect 3007 15456 10232 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 10226 15444 10232 15456
rect 10284 15444 10290 15496
rect 11146 15444 11152 15496
rect 11204 15444 11210 15496
rect 12710 15444 12716 15496
rect 12768 15484 12774 15496
rect 13265 15487 13323 15493
rect 13265 15484 13277 15487
rect 12768 15456 13277 15484
rect 12768 15444 12774 15456
rect 13265 15453 13277 15456
rect 13311 15453 13323 15487
rect 13265 15447 13323 15453
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15484 13415 15487
rect 13446 15484 13452 15496
rect 13403 15456 13452 15484
rect 13403 15453 13415 15456
rect 13357 15447 13415 15453
rect 13446 15444 13452 15456
rect 13504 15444 13510 15496
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15484 14795 15487
rect 18414 15484 18420 15496
rect 14783 15456 18420 15484
rect 14783 15453 14795 15456
rect 14737 15447 14795 15453
rect 18414 15444 18420 15456
rect 18472 15444 18478 15496
rect 18601 15487 18659 15493
rect 18601 15453 18613 15487
rect 18647 15484 18659 15487
rect 20898 15484 20904 15496
rect 18647 15456 20904 15484
rect 18647 15453 18659 15456
rect 18601 15447 18659 15453
rect 20898 15444 20904 15456
rect 20956 15444 20962 15496
rect 21174 15444 21180 15496
rect 21232 15484 21238 15496
rect 21637 15487 21695 15493
rect 21637 15484 21649 15487
rect 21232 15456 21649 15484
rect 21232 15444 21238 15456
rect 21637 15453 21649 15456
rect 21683 15484 21695 15487
rect 22462 15484 22468 15496
rect 21683 15456 22468 15484
rect 21683 15453 21695 15456
rect 21637 15447 21695 15453
rect 22462 15444 22468 15456
rect 22520 15444 22526 15496
rect 23569 15487 23627 15493
rect 23569 15453 23581 15487
rect 23615 15484 23627 15487
rect 27338 15484 27344 15496
rect 23615 15456 27344 15484
rect 23615 15453 23627 15456
rect 23569 15447 23627 15453
rect 27338 15444 27344 15456
rect 27396 15444 27402 15496
rect 27706 15444 27712 15496
rect 27764 15484 27770 15496
rect 27801 15487 27859 15493
rect 27801 15484 27813 15487
rect 27764 15456 27813 15484
rect 27764 15444 27770 15456
rect 27801 15453 27813 15456
rect 27847 15484 27859 15487
rect 28445 15487 28503 15493
rect 28445 15484 28457 15487
rect 27847 15456 28457 15484
rect 27847 15453 27859 15456
rect 27801 15447 27859 15453
rect 28445 15453 28457 15456
rect 28491 15453 28503 15487
rect 28445 15447 28503 15453
rect 934 15376 940 15428
rect 992 15416 998 15428
rect 1765 15419 1823 15425
rect 1765 15416 1777 15419
rect 992 15388 1777 15416
rect 992 15376 998 15388
rect 1765 15385 1777 15388
rect 1811 15385 1823 15419
rect 1765 15379 1823 15385
rect 4154 15376 4160 15428
rect 4212 15416 4218 15428
rect 6365 15419 6423 15425
rect 6365 15416 6377 15419
rect 4212 15388 6377 15416
rect 4212 15376 4218 15388
rect 6365 15385 6377 15388
rect 6411 15385 6423 15419
rect 6365 15379 6423 15385
rect 6549 15419 6607 15425
rect 6549 15385 6561 15419
rect 6595 15416 6607 15419
rect 6595 15388 10916 15416
rect 6595 15385 6607 15388
rect 6549 15379 6607 15385
rect 9030 15308 9036 15360
rect 9088 15308 9094 15360
rect 10888 15348 10916 15388
rect 15930 15376 15936 15428
rect 15988 15376 15994 15428
rect 16390 15376 16396 15428
rect 16448 15416 16454 15428
rect 16448 15388 18460 15416
rect 16448 15376 16454 15388
rect 11882 15348 11888 15360
rect 10888 15320 11888 15348
rect 11882 15308 11888 15320
rect 11940 15348 11946 15360
rect 12802 15348 12808 15360
rect 11940 15320 12808 15348
rect 11940 15308 11946 15320
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 13538 15308 13544 15360
rect 13596 15348 13602 15360
rect 13725 15351 13783 15357
rect 13725 15348 13737 15351
rect 13596 15320 13737 15348
rect 13596 15308 13602 15320
rect 13725 15317 13737 15320
rect 13771 15317 13783 15351
rect 13725 15311 13783 15317
rect 13906 15308 13912 15360
rect 13964 15348 13970 15360
rect 14277 15351 14335 15357
rect 14277 15348 14289 15351
rect 13964 15320 14289 15348
rect 13964 15308 13970 15320
rect 14277 15317 14289 15320
rect 14323 15317 14335 15351
rect 14277 15311 14335 15317
rect 14642 15308 14648 15360
rect 14700 15308 14706 15360
rect 15562 15308 15568 15360
rect 15620 15308 15626 15360
rect 16025 15351 16083 15357
rect 16025 15317 16037 15351
rect 16071 15348 16083 15351
rect 16114 15348 16120 15360
rect 16071 15320 16120 15348
rect 16071 15317 16083 15320
rect 16025 15311 16083 15317
rect 16114 15308 16120 15320
rect 16172 15308 16178 15360
rect 17126 15308 17132 15360
rect 17184 15308 17190 15360
rect 17221 15351 17279 15357
rect 17221 15317 17233 15351
rect 17267 15348 17279 15351
rect 17310 15348 17316 15360
rect 17267 15320 17316 15348
rect 17267 15317 17279 15320
rect 17221 15311 17279 15317
rect 17310 15308 17316 15320
rect 17368 15308 17374 15360
rect 18432 15357 18460 15388
rect 18506 15376 18512 15428
rect 18564 15416 18570 15428
rect 21450 15416 21456 15428
rect 18564 15388 21456 15416
rect 18564 15376 18570 15388
rect 21450 15376 21456 15388
rect 21508 15376 21514 15428
rect 21545 15419 21603 15425
rect 21545 15385 21557 15419
rect 21591 15416 21603 15419
rect 21591 15388 21772 15416
rect 21591 15385 21603 15388
rect 21545 15379 21603 15385
rect 18417 15351 18475 15357
rect 18417 15317 18429 15351
rect 18463 15317 18475 15351
rect 18417 15311 18475 15317
rect 19521 15351 19579 15357
rect 19521 15317 19533 15351
rect 19567 15348 19579 15351
rect 19794 15348 19800 15360
rect 19567 15320 19800 15348
rect 19567 15317 19579 15320
rect 19521 15311 19579 15317
rect 19794 15308 19800 15320
rect 19852 15308 19858 15360
rect 20254 15308 20260 15360
rect 20312 15308 20318 15360
rect 21082 15308 21088 15360
rect 21140 15348 21146 15360
rect 21177 15351 21235 15357
rect 21177 15348 21189 15351
rect 21140 15320 21189 15348
rect 21140 15308 21146 15320
rect 21177 15317 21189 15320
rect 21223 15317 21235 15351
rect 21744 15348 21772 15388
rect 22094 15376 22100 15428
rect 22152 15416 22158 15428
rect 23477 15419 23535 15425
rect 22152 15388 23152 15416
rect 22152 15376 22158 15388
rect 22278 15348 22284 15360
rect 21744 15320 22284 15348
rect 21177 15311 21235 15317
rect 22278 15308 22284 15320
rect 22336 15308 22342 15360
rect 23124 15357 23152 15388
rect 23477 15385 23489 15419
rect 23523 15416 23535 15419
rect 25041 15419 25099 15425
rect 23523 15388 24716 15416
rect 23523 15385 23535 15388
rect 23477 15379 23535 15385
rect 24688 15357 24716 15388
rect 25041 15385 25053 15419
rect 25087 15416 25099 15419
rect 25682 15416 25688 15428
rect 25087 15388 25688 15416
rect 25087 15385 25099 15388
rect 25041 15379 25099 15385
rect 25682 15376 25688 15388
rect 25740 15376 25746 15428
rect 26326 15376 26332 15428
rect 26384 15416 26390 15428
rect 26970 15416 26976 15428
rect 26384 15388 26976 15416
rect 26384 15376 26390 15388
rect 26970 15376 26976 15388
rect 27028 15376 27034 15428
rect 27893 15419 27951 15425
rect 27893 15385 27905 15419
rect 27939 15416 27951 15419
rect 28736 15416 28764 15512
rect 27939 15388 28764 15416
rect 29181 15419 29239 15425
rect 27939 15385 27951 15388
rect 27893 15379 27951 15385
rect 29181 15385 29193 15419
rect 29227 15416 29239 15419
rect 30282 15416 30288 15428
rect 29227 15388 30288 15416
rect 29227 15385 29239 15388
rect 29181 15379 29239 15385
rect 30282 15376 30288 15388
rect 30340 15376 30346 15428
rect 30742 15376 30748 15428
rect 30800 15376 30806 15428
rect 31202 15376 31208 15428
rect 31260 15376 31266 15428
rect 32784 15416 32812 15524
rect 32861 15521 32873 15555
rect 32907 15521 32919 15555
rect 32861 15515 32919 15521
rect 32953 15555 33011 15561
rect 32953 15521 32965 15555
rect 32999 15521 33011 15555
rect 32953 15515 33011 15521
rect 32876 15484 32904 15515
rect 34790 15512 34796 15564
rect 34848 15552 34854 15564
rect 34885 15555 34943 15561
rect 34885 15552 34897 15555
rect 34848 15524 34897 15552
rect 34848 15512 34854 15524
rect 34885 15521 34897 15524
rect 34931 15521 34943 15555
rect 34885 15515 34943 15521
rect 35161 15555 35219 15561
rect 35161 15521 35173 15555
rect 35207 15552 35219 15555
rect 35894 15552 35900 15564
rect 35207 15524 35900 15552
rect 35207 15521 35219 15524
rect 35161 15515 35219 15521
rect 35894 15512 35900 15524
rect 35952 15512 35958 15564
rect 37366 15512 37372 15564
rect 37424 15552 37430 15564
rect 39482 15552 39488 15564
rect 37424 15524 39488 15552
rect 37424 15512 37430 15524
rect 39482 15512 39488 15524
rect 39540 15552 39546 15564
rect 40037 15555 40095 15561
rect 40037 15552 40049 15555
rect 39540 15524 40049 15552
rect 39540 15512 39546 15524
rect 40037 15521 40049 15524
rect 40083 15521 40095 15555
rect 40037 15515 40095 15521
rect 40310 15512 40316 15564
rect 40368 15512 40374 15564
rect 34054 15484 34060 15496
rect 32876 15456 34060 15484
rect 34054 15444 34060 15456
rect 34112 15444 34118 15496
rect 48869 15487 48927 15493
rect 48869 15453 48881 15487
rect 48915 15484 48927 15487
rect 49326 15484 49332 15496
rect 48915 15456 49332 15484
rect 48915 15453 48927 15456
rect 48869 15447 48927 15453
rect 49326 15444 49332 15456
rect 49384 15444 49390 15496
rect 34606 15416 34612 15428
rect 32784 15388 34612 15416
rect 34606 15376 34612 15388
rect 34664 15376 34670 15428
rect 35618 15376 35624 15428
rect 35676 15376 35682 15428
rect 38746 15376 38752 15428
rect 38804 15376 38810 15428
rect 39206 15376 39212 15428
rect 39264 15376 39270 15428
rect 39942 15376 39948 15428
rect 40000 15416 40006 15428
rect 40000 15388 40802 15416
rect 40000 15376 40006 15388
rect 23109 15351 23167 15357
rect 23109 15317 23121 15351
rect 23155 15317 23167 15351
rect 23109 15311 23167 15317
rect 24673 15351 24731 15357
rect 24673 15317 24685 15351
rect 24719 15317 24731 15351
rect 24673 15311 24731 15317
rect 25130 15308 25136 15360
rect 25188 15308 25194 15360
rect 25866 15308 25872 15360
rect 25924 15308 25930 15360
rect 26234 15308 26240 15360
rect 26292 15348 26298 15360
rect 26786 15348 26792 15360
rect 26292 15320 26792 15348
rect 26292 15308 26298 15320
rect 26786 15308 26792 15320
rect 26844 15348 26850 15360
rect 26881 15351 26939 15357
rect 26881 15348 26893 15351
rect 26844 15320 26893 15348
rect 26844 15308 26850 15320
rect 26881 15317 26893 15320
rect 26927 15317 26939 15351
rect 26881 15311 26939 15317
rect 27154 15308 27160 15360
rect 27212 15308 27218 15360
rect 28994 15308 29000 15360
rect 29052 15308 29058 15360
rect 30009 15351 30067 15357
rect 30009 15317 30021 15351
rect 30055 15348 30067 15351
rect 31018 15348 31024 15360
rect 30055 15320 31024 15348
rect 30055 15317 30067 15320
rect 30009 15311 30067 15317
rect 31018 15308 31024 15320
rect 31076 15308 31082 15360
rect 32306 15308 32312 15360
rect 32364 15348 32370 15360
rect 32674 15348 32680 15360
rect 32364 15320 32680 15348
rect 32364 15308 32370 15320
rect 32674 15308 32680 15320
rect 32732 15308 32738 15360
rect 33045 15351 33103 15357
rect 33045 15317 33057 15351
rect 33091 15348 33103 15351
rect 33318 15348 33324 15360
rect 33091 15320 33324 15348
rect 33091 15317 33103 15320
rect 33045 15311 33103 15317
rect 33318 15308 33324 15320
rect 33376 15308 33382 15360
rect 33413 15351 33471 15357
rect 33413 15317 33425 15351
rect 33459 15348 33471 15351
rect 33686 15348 33692 15360
rect 33459 15320 33692 15348
rect 33459 15317 33471 15320
rect 33413 15311 33471 15317
rect 33686 15308 33692 15320
rect 33744 15308 33750 15360
rect 33870 15308 33876 15360
rect 33928 15308 33934 15360
rect 36446 15308 36452 15360
rect 36504 15348 36510 15360
rect 37093 15351 37151 15357
rect 37093 15348 37105 15351
rect 36504 15320 37105 15348
rect 36504 15308 36510 15320
rect 37093 15317 37105 15320
rect 37139 15317 37151 15351
rect 37093 15311 37151 15317
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 9674 15104 9680 15156
rect 9732 15104 9738 15156
rect 9766 15104 9772 15156
rect 9824 15104 9830 15156
rect 10137 15147 10195 15153
rect 10137 15113 10149 15147
rect 10183 15144 10195 15147
rect 11330 15144 11336 15156
rect 10183 15116 11336 15144
rect 10183 15113 10195 15116
rect 10137 15107 10195 15113
rect 11330 15104 11336 15116
rect 11388 15104 11394 15156
rect 11790 15104 11796 15156
rect 11848 15144 11854 15156
rect 11885 15147 11943 15153
rect 11885 15144 11897 15147
rect 11848 15116 11897 15144
rect 11848 15104 11854 15116
rect 11885 15113 11897 15116
rect 11931 15113 11943 15147
rect 15933 15147 15991 15153
rect 11885 15107 11943 15113
rect 12912 15116 13768 15144
rect 10870 15036 10876 15088
rect 10928 15036 10934 15088
rect 11054 15036 11060 15088
rect 11112 15036 11118 15088
rect 11146 15036 11152 15088
rect 11204 15076 11210 15088
rect 12912 15085 12940 15116
rect 12897 15079 12955 15085
rect 12897 15076 12909 15079
rect 11204 15048 12909 15076
rect 11204 15036 11210 15048
rect 12897 15045 12909 15048
rect 12943 15045 12955 15079
rect 12897 15039 12955 15045
rect 13740 15020 13768 15116
rect 15933 15113 15945 15147
rect 15979 15144 15991 15147
rect 18325 15147 18383 15153
rect 18325 15144 18337 15147
rect 15979 15116 18337 15144
rect 15979 15113 15991 15116
rect 15933 15107 15991 15113
rect 18325 15113 18337 15116
rect 18371 15113 18383 15147
rect 18325 15107 18383 15113
rect 18693 15147 18751 15153
rect 18693 15113 18705 15147
rect 18739 15144 18751 15147
rect 19334 15144 19340 15156
rect 18739 15116 19340 15144
rect 18739 15113 18751 15116
rect 18693 15107 18751 15113
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 19426 15104 19432 15156
rect 19484 15144 19490 15156
rect 19521 15147 19579 15153
rect 19521 15144 19533 15147
rect 19484 15116 19533 15144
rect 19484 15104 19490 15116
rect 19521 15113 19533 15116
rect 19567 15113 19579 15147
rect 21542 15144 21548 15156
rect 19521 15107 19579 15113
rect 19628 15116 21548 15144
rect 14826 15036 14832 15088
rect 14884 15036 14890 15088
rect 15654 15036 15660 15088
rect 15712 15076 15718 15088
rect 16025 15079 16083 15085
rect 16025 15076 16037 15079
rect 15712 15048 16037 15076
rect 15712 15036 15718 15048
rect 16025 15045 16037 15048
rect 16071 15045 16083 15079
rect 16025 15039 16083 15045
rect 16114 15036 16120 15088
rect 16172 15076 16178 15088
rect 19628 15076 19656 15116
rect 21542 15104 21548 15116
rect 21600 15104 21606 15156
rect 22830 15104 22836 15156
rect 22888 15144 22894 15156
rect 22925 15147 22983 15153
rect 22925 15144 22937 15147
rect 22888 15116 22937 15144
rect 22888 15104 22894 15116
rect 22925 15113 22937 15116
rect 22971 15113 22983 15147
rect 22925 15107 22983 15113
rect 23750 15104 23756 15156
rect 23808 15144 23814 15156
rect 24121 15147 24179 15153
rect 24121 15144 24133 15147
rect 23808 15116 24133 15144
rect 23808 15104 23814 15116
rect 24121 15113 24133 15116
rect 24167 15113 24179 15147
rect 24121 15107 24179 15113
rect 24581 15147 24639 15153
rect 24581 15113 24593 15147
rect 24627 15144 24639 15147
rect 24670 15144 24676 15156
rect 24627 15116 24676 15144
rect 24627 15113 24639 15116
rect 24581 15107 24639 15113
rect 24670 15104 24676 15116
rect 24728 15144 24734 15156
rect 26329 15147 26387 15153
rect 24728 15116 26280 15144
rect 24728 15104 24734 15116
rect 16172 15048 19656 15076
rect 19889 15079 19947 15085
rect 16172 15036 16178 15048
rect 19889 15045 19901 15079
rect 19935 15076 19947 15079
rect 20806 15076 20812 15088
rect 19935 15048 20812 15076
rect 19935 15045 19947 15048
rect 19889 15039 19947 15045
rect 20806 15036 20812 15048
rect 20864 15036 20870 15088
rect 21085 15079 21143 15085
rect 21085 15045 21097 15079
rect 21131 15076 21143 15079
rect 21634 15076 21640 15088
rect 21131 15048 21640 15076
rect 21131 15045 21143 15048
rect 21085 15039 21143 15045
rect 21634 15036 21640 15048
rect 21692 15076 21698 15088
rect 21821 15079 21879 15085
rect 21821 15076 21833 15079
rect 21692 15048 21833 15076
rect 21692 15036 21698 15048
rect 21821 15045 21833 15048
rect 21867 15045 21879 15079
rect 21821 15039 21879 15045
rect 23385 15079 23443 15085
rect 23385 15045 23397 15079
rect 23431 15076 23443 15079
rect 25866 15076 25872 15088
rect 23431 15048 25872 15076
rect 23431 15045 23443 15048
rect 23385 15039 23443 15045
rect 25866 15036 25872 15048
rect 25924 15036 25930 15088
rect 934 14968 940 15020
rect 992 15008 998 15020
rect 1765 15011 1823 15017
rect 1765 15008 1777 15011
rect 992 14980 1777 15008
rect 992 14968 998 14980
rect 1765 14977 1777 14980
rect 1811 14977 1823 15011
rect 1765 14971 1823 14977
rect 2961 15011 3019 15017
rect 2961 14977 2973 15011
rect 3007 15008 3019 15011
rect 4154 15008 4160 15020
rect 3007 14980 4160 15008
rect 3007 14977 3019 14980
rect 2961 14971 3019 14977
rect 4154 14968 4160 14980
rect 4212 14968 4218 15020
rect 12250 14968 12256 15020
rect 12308 14968 12314 15020
rect 13722 14968 13728 15020
rect 13780 14968 13786 15020
rect 15102 14968 15108 15020
rect 15160 14968 15166 15020
rect 15286 14968 15292 15020
rect 15344 15008 15350 15020
rect 16132 15008 16160 15036
rect 15344 14980 16160 15008
rect 17221 15011 17279 15017
rect 15344 14968 15350 14980
rect 17221 14977 17233 15011
rect 17267 15008 17279 15011
rect 17494 15008 17500 15020
rect 17267 14980 17500 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 17494 14968 17500 14980
rect 17552 14968 17558 15020
rect 18506 14968 18512 15020
rect 18564 15008 18570 15020
rect 19981 15011 20039 15017
rect 18564 14980 18920 15008
rect 18564 14968 18570 14980
rect 9585 14943 9643 14949
rect 9585 14909 9597 14943
rect 9631 14940 9643 14943
rect 9766 14940 9772 14952
rect 9631 14912 9772 14940
rect 9631 14909 9643 14912
rect 9585 14903 9643 14909
rect 9766 14900 9772 14912
rect 9824 14900 9830 14952
rect 11609 14943 11667 14949
rect 11609 14909 11621 14943
rect 11655 14940 11667 14943
rect 12342 14940 12348 14952
rect 11655 14912 12348 14940
rect 11655 14909 11667 14912
rect 11609 14903 11667 14909
rect 12342 14900 12348 14912
rect 12400 14900 12406 14952
rect 12437 14943 12495 14949
rect 12437 14909 12449 14943
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 11054 14832 11060 14884
rect 11112 14872 11118 14884
rect 11112 14844 12020 14872
rect 11112 14832 11118 14844
rect 10597 14807 10655 14813
rect 10597 14773 10609 14807
rect 10643 14804 10655 14807
rect 10686 14804 10692 14816
rect 10643 14776 10692 14804
rect 10643 14773 10655 14776
rect 10597 14767 10655 14773
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 11992 14804 12020 14844
rect 12066 14832 12072 14884
rect 12124 14872 12130 14884
rect 12452 14872 12480 14903
rect 13814 14900 13820 14952
rect 13872 14940 13878 14952
rect 14182 14940 14188 14952
rect 13872 14912 14188 14940
rect 13872 14900 13878 14912
rect 14182 14900 14188 14912
rect 14240 14900 14246 14952
rect 14274 14900 14280 14952
rect 14332 14940 14338 14952
rect 14332 14912 15056 14940
rect 14332 14900 14338 14912
rect 12124 14844 12480 14872
rect 15028 14872 15056 14912
rect 15378 14900 15384 14952
rect 15436 14940 15442 14952
rect 16117 14943 16175 14949
rect 16117 14940 16129 14943
rect 15436 14912 16129 14940
rect 15436 14900 15442 14912
rect 16117 14909 16129 14912
rect 16163 14909 16175 14943
rect 16117 14903 16175 14909
rect 17310 14900 17316 14952
rect 17368 14900 17374 14952
rect 17402 14900 17408 14952
rect 17460 14900 17466 14952
rect 18046 14900 18052 14952
rect 18104 14940 18110 14952
rect 18892 14949 18920 14980
rect 19981 14977 19993 15011
rect 20027 15008 20039 15011
rect 20898 15008 20904 15020
rect 20027 14980 20904 15008
rect 20027 14977 20039 14980
rect 19981 14971 20039 14977
rect 20898 14968 20904 14980
rect 20956 14968 20962 15020
rect 21450 15008 21456 15020
rect 21284 14980 21456 15008
rect 18785 14943 18843 14949
rect 18785 14940 18797 14943
rect 18104 14912 18797 14940
rect 18104 14900 18110 14912
rect 18785 14909 18797 14912
rect 18831 14909 18843 14943
rect 18785 14903 18843 14909
rect 18877 14943 18935 14949
rect 18877 14909 18889 14943
rect 18923 14909 18935 14943
rect 18877 14903 18935 14909
rect 20162 14900 20168 14952
rect 20220 14900 20226 14952
rect 20530 14900 20536 14952
rect 20588 14940 20594 14952
rect 21284 14949 21312 14980
rect 21450 14968 21456 14980
rect 21508 14968 21514 15020
rect 23290 14968 23296 15020
rect 23348 14968 23354 15020
rect 24489 15011 24547 15017
rect 24489 14977 24501 15011
rect 24535 15008 24547 15011
rect 25038 15008 25044 15020
rect 24535 14980 25044 15008
rect 24535 14977 24547 14980
rect 24489 14971 24547 14977
rect 25038 14968 25044 14980
rect 25096 14968 25102 15020
rect 25130 14968 25136 15020
rect 25188 15008 25194 15020
rect 25317 15011 25375 15017
rect 25317 15008 25329 15011
rect 25188 14980 25329 15008
rect 25188 14968 25194 14980
rect 25317 14977 25329 14980
rect 25363 14977 25375 15011
rect 25317 14971 25375 14977
rect 25406 14968 25412 15020
rect 25464 15008 25470 15020
rect 25593 15011 25651 15017
rect 25593 15008 25605 15011
rect 25464 14980 25605 15008
rect 25464 14968 25470 14980
rect 25593 14977 25605 14980
rect 25639 15008 25651 15011
rect 25682 15008 25688 15020
rect 25639 14980 25688 15008
rect 25639 14977 25651 14980
rect 25593 14971 25651 14977
rect 25682 14968 25688 14980
rect 25740 14968 25746 15020
rect 26252 15017 26280 15116
rect 26329 15113 26341 15147
rect 26375 15144 26387 15147
rect 27433 15147 27491 15153
rect 27433 15144 27445 15147
rect 26375 15116 27445 15144
rect 26375 15113 26387 15116
rect 26329 15107 26387 15113
rect 27433 15113 27445 15116
rect 27479 15144 27491 15147
rect 29638 15144 29644 15156
rect 27479 15116 29644 15144
rect 27479 15113 27491 15116
rect 27433 15107 27491 15113
rect 29638 15104 29644 15116
rect 29696 15104 29702 15156
rect 31294 15104 31300 15156
rect 31352 15144 31358 15156
rect 31389 15147 31447 15153
rect 31389 15144 31401 15147
rect 31352 15116 31401 15144
rect 31352 15104 31358 15116
rect 31389 15113 31401 15116
rect 31435 15113 31447 15147
rect 32309 15147 32367 15153
rect 32309 15144 32321 15147
rect 31389 15107 31447 15113
rect 31496 15116 32321 15144
rect 27062 15036 27068 15088
rect 27120 15036 27126 15088
rect 27890 15036 27896 15088
rect 27948 15076 27954 15088
rect 28534 15076 28540 15088
rect 27948 15048 28540 15076
rect 27948 15036 27954 15048
rect 28534 15036 28540 15048
rect 28592 15036 28598 15088
rect 29270 15036 29276 15088
rect 29328 15036 29334 15088
rect 29546 15036 29552 15088
rect 29604 15076 29610 15088
rect 29604 15048 30788 15076
rect 29604 15036 29610 15048
rect 26237 15011 26295 15017
rect 26237 14977 26249 15011
rect 26283 15008 26295 15011
rect 27246 15008 27252 15020
rect 26283 14980 27252 15008
rect 26283 14977 26295 14980
rect 26237 14971 26295 14977
rect 27246 14968 27252 14980
rect 27304 14968 27310 15020
rect 27798 14968 27804 15020
rect 27856 15008 27862 15020
rect 27985 15011 28043 15017
rect 27985 15008 27997 15011
rect 27856 14980 27997 15008
rect 27856 14968 27862 14980
rect 27985 14977 27997 14980
rect 28031 14977 28043 15011
rect 30190 15008 30196 15020
rect 27985 14971 28043 14977
rect 29564 14980 30196 15008
rect 21177 14943 21235 14949
rect 21177 14940 21189 14943
rect 20588 14912 21189 14940
rect 20588 14900 20594 14912
rect 21177 14909 21189 14912
rect 21223 14909 21235 14943
rect 21177 14903 21235 14909
rect 21269 14943 21327 14949
rect 21269 14909 21281 14943
rect 21315 14909 21327 14943
rect 21269 14903 21327 14909
rect 21358 14900 21364 14952
rect 21416 14940 21422 14952
rect 22005 14943 22063 14949
rect 22005 14940 22017 14943
rect 21416 14912 22017 14940
rect 21416 14900 21422 14912
rect 22005 14909 22017 14912
rect 22051 14909 22063 14943
rect 22005 14903 22063 14909
rect 23566 14900 23572 14952
rect 23624 14900 23630 14952
rect 24210 14900 24216 14952
rect 24268 14940 24274 14952
rect 24673 14943 24731 14949
rect 24673 14940 24685 14943
rect 24268 14912 24685 14940
rect 24268 14900 24274 14912
rect 24673 14909 24685 14912
rect 24719 14909 24731 14943
rect 24673 14903 24731 14909
rect 24762 14900 24768 14952
rect 24820 14940 24826 14952
rect 26421 14943 26479 14949
rect 26421 14940 26433 14943
rect 24820 14912 26433 14940
rect 24820 14900 24826 14912
rect 26421 14909 26433 14912
rect 26467 14909 26479 14943
rect 26421 14903 26479 14909
rect 27338 14900 27344 14952
rect 27396 14940 27402 14952
rect 28261 14943 28319 14949
rect 28261 14940 28273 14943
rect 27396 14912 28273 14940
rect 27396 14900 27402 14912
rect 28261 14909 28273 14912
rect 28307 14940 28319 14943
rect 29564 14940 29592 14980
rect 30190 14968 30196 14980
rect 30248 14968 30254 15020
rect 30558 14968 30564 15020
rect 30616 14968 30622 15020
rect 28307 14912 29592 14940
rect 29733 14943 29791 14949
rect 28307 14909 28319 14912
rect 28261 14903 28319 14909
rect 29733 14909 29745 14943
rect 29779 14940 29791 14943
rect 29822 14940 29828 14952
rect 29779 14912 29828 14940
rect 29779 14909 29791 14912
rect 29733 14903 29791 14909
rect 29822 14900 29828 14912
rect 29880 14900 29886 14952
rect 30006 14900 30012 14952
rect 30064 14940 30070 14952
rect 30650 14940 30656 14952
rect 30064 14912 30656 14940
rect 30064 14900 30070 14912
rect 30650 14900 30656 14912
rect 30708 14900 30714 14952
rect 30760 14949 30788 15048
rect 30926 15036 30932 15088
rect 30984 15076 30990 15088
rect 31496 15076 31524 15116
rect 32309 15113 32321 15116
rect 32355 15113 32367 15147
rect 32309 15107 32367 15113
rect 33870 15104 33876 15156
rect 33928 15104 33934 15156
rect 35069 15147 35127 15153
rect 35069 15113 35081 15147
rect 35115 15144 35127 15147
rect 36998 15144 37004 15156
rect 35115 15116 37004 15144
rect 35115 15113 35127 15116
rect 35069 15107 35127 15113
rect 36998 15104 37004 15116
rect 37056 15104 37062 15156
rect 37642 15104 37648 15156
rect 37700 15144 37706 15156
rect 39209 15147 39267 15153
rect 39209 15144 39221 15147
rect 37700 15116 39221 15144
rect 37700 15104 37706 15116
rect 39209 15113 39221 15116
rect 39255 15113 39267 15147
rect 39209 15107 39267 15113
rect 40126 15104 40132 15156
rect 40184 15104 40190 15156
rect 30984 15048 31524 15076
rect 30984 15036 30990 15048
rect 35986 15036 35992 15088
rect 36044 15076 36050 15088
rect 36173 15079 36231 15085
rect 36173 15076 36185 15079
rect 36044 15048 36185 15076
rect 36044 15036 36050 15048
rect 36173 15045 36185 15048
rect 36219 15045 36231 15079
rect 36173 15039 36231 15045
rect 36262 15036 36268 15088
rect 36320 15036 36326 15088
rect 37734 15036 37740 15088
rect 37792 15036 37798 15088
rect 38746 15036 38752 15088
rect 38804 15036 38810 15088
rect 40037 15079 40095 15085
rect 40037 15045 40049 15079
rect 40083 15076 40095 15079
rect 48406 15076 48412 15088
rect 40083 15048 48412 15076
rect 40083 15045 40095 15048
rect 40037 15039 40095 15045
rect 48406 15036 48412 15048
rect 48464 15036 48470 15088
rect 31754 14968 31760 15020
rect 31812 15008 31818 15020
rect 32677 15011 32735 15017
rect 32677 15008 32689 15011
rect 31812 14980 32689 15008
rect 31812 14968 31818 14980
rect 32677 14977 32689 14980
rect 32723 14977 32735 15011
rect 32677 14971 32735 14977
rect 32769 15011 32827 15017
rect 32769 14977 32781 15011
rect 32815 15008 32827 15011
rect 35894 15008 35900 15020
rect 32815 14980 35900 15008
rect 32815 14977 32827 14980
rect 32769 14971 32827 14977
rect 35894 14968 35900 14980
rect 35952 14968 35958 15020
rect 36909 15011 36967 15017
rect 36909 15008 36921 15011
rect 36004 14980 36921 15008
rect 30745 14943 30803 14949
rect 30745 14909 30757 14943
rect 30791 14909 30803 14943
rect 30745 14903 30803 14909
rect 31846 14900 31852 14952
rect 31904 14900 31910 14952
rect 32306 14900 32312 14952
rect 32364 14940 32370 14952
rect 32861 14943 32919 14949
rect 32861 14940 32873 14943
rect 32364 14912 32873 14940
rect 32364 14900 32370 14912
rect 32861 14909 32873 14912
rect 32907 14909 32919 14943
rect 32861 14903 32919 14909
rect 33689 14943 33747 14949
rect 33689 14909 33701 14943
rect 33735 14909 33747 14943
rect 33689 14903 33747 14909
rect 15396 14872 15424 14900
rect 15028 14844 15424 14872
rect 12124 14832 12130 14844
rect 17954 14832 17960 14884
rect 18012 14872 18018 14884
rect 20717 14875 20775 14881
rect 20717 14872 20729 14875
rect 18012 14844 20729 14872
rect 18012 14832 18018 14844
rect 20717 14841 20729 14844
rect 20763 14841 20775 14875
rect 27617 14875 27675 14881
rect 20717 14835 20775 14841
rect 22480 14844 26004 14872
rect 12802 14804 12808 14816
rect 11992 14776 12808 14804
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 13357 14807 13415 14813
rect 13357 14773 13369 14807
rect 13403 14804 13415 14807
rect 14274 14804 14280 14816
rect 13403 14776 14280 14804
rect 13403 14773 13415 14776
rect 13357 14767 13415 14773
rect 14274 14764 14280 14776
rect 14332 14764 14338 14816
rect 14458 14764 14464 14816
rect 14516 14804 14522 14816
rect 15565 14807 15623 14813
rect 15565 14804 15577 14807
rect 14516 14776 15577 14804
rect 14516 14764 14522 14776
rect 15565 14773 15577 14776
rect 15611 14773 15623 14807
rect 15565 14767 15623 14773
rect 15930 14764 15936 14816
rect 15988 14804 15994 14816
rect 16853 14807 16911 14813
rect 16853 14804 16865 14807
rect 15988 14776 16865 14804
rect 15988 14764 15994 14776
rect 16853 14773 16865 14776
rect 16899 14773 16911 14807
rect 16853 14767 16911 14773
rect 18598 14764 18604 14816
rect 18656 14804 18662 14816
rect 22480 14804 22508 14844
rect 18656 14776 22508 14804
rect 18656 14764 18662 14776
rect 25038 14764 25044 14816
rect 25096 14804 25102 14816
rect 25133 14807 25191 14813
rect 25133 14804 25145 14807
rect 25096 14776 25145 14804
rect 25096 14764 25102 14776
rect 25133 14773 25145 14776
rect 25179 14773 25191 14807
rect 25133 14767 25191 14773
rect 25682 14764 25688 14816
rect 25740 14804 25746 14816
rect 25869 14807 25927 14813
rect 25869 14804 25881 14807
rect 25740 14776 25881 14804
rect 25740 14764 25746 14776
rect 25869 14773 25881 14776
rect 25915 14773 25927 14807
rect 25976 14804 26004 14844
rect 27617 14841 27629 14875
rect 27663 14872 27675 14875
rect 27706 14872 27712 14884
rect 27663 14844 27712 14872
rect 27663 14841 27675 14844
rect 27617 14835 27675 14841
rect 27706 14832 27712 14844
rect 27764 14832 27770 14884
rect 33704 14872 33732 14903
rect 33778 14900 33784 14952
rect 33836 14900 33842 14952
rect 34882 14900 34888 14952
rect 34940 14900 34946 14952
rect 34977 14943 35035 14949
rect 34977 14909 34989 14943
rect 35023 14940 35035 14943
rect 36004 14940 36032 14980
rect 36280 14952 36308 14980
rect 36909 14977 36921 14980
rect 36955 14977 36967 15011
rect 36909 14971 36967 14977
rect 37366 14968 37372 15020
rect 37424 15008 37430 15020
rect 37461 15011 37519 15017
rect 37461 15008 37473 15011
rect 37424 14980 37473 15008
rect 37424 14968 37430 14980
rect 37461 14977 37473 14980
rect 37507 14977 37519 15011
rect 37461 14971 37519 14977
rect 40862 14968 40868 15020
rect 40920 14968 40926 15020
rect 48777 15011 48835 15017
rect 48777 14977 48789 15011
rect 48823 15008 48835 15011
rect 49326 15008 49332 15020
rect 48823 14980 49332 15008
rect 48823 14977 48835 14980
rect 48777 14971 48835 14977
rect 49326 14968 49332 14980
rect 49384 14968 49390 15020
rect 35023 14912 36032 14940
rect 35023 14909 35035 14912
rect 34977 14903 35035 14909
rect 36078 14900 36084 14952
rect 36136 14900 36142 14952
rect 36262 14900 36268 14952
rect 36320 14900 36326 14952
rect 37090 14900 37096 14952
rect 37148 14940 37154 14952
rect 40221 14943 40279 14949
rect 40221 14940 40233 14943
rect 37148 14912 40233 14940
rect 37148 14900 37154 14912
rect 40221 14909 40233 14912
rect 40267 14909 40279 14943
rect 40221 14903 40279 14909
rect 33962 14872 33968 14884
rect 29288 14844 30328 14872
rect 33704 14844 33968 14872
rect 29288 14804 29316 14844
rect 25976 14776 29316 14804
rect 25869 14767 25927 14773
rect 30190 14764 30196 14816
rect 30248 14764 30254 14816
rect 30300 14804 30328 14844
rect 33962 14832 33968 14844
rect 34020 14832 34026 14884
rect 35437 14875 35495 14881
rect 35437 14841 35449 14875
rect 35483 14872 35495 14875
rect 36538 14872 36544 14884
rect 35483 14844 36544 14872
rect 35483 14841 35495 14844
rect 35437 14835 35495 14841
rect 36538 14832 36544 14844
rect 36596 14832 36602 14884
rect 36633 14875 36691 14881
rect 36633 14841 36645 14875
rect 36679 14872 36691 14875
rect 36679 14844 37596 14872
rect 36679 14841 36691 14844
rect 36633 14835 36691 14841
rect 33318 14804 33324 14816
rect 30300 14776 33324 14804
rect 33318 14764 33324 14776
rect 33376 14804 33382 14816
rect 33502 14804 33508 14816
rect 33376 14776 33508 14804
rect 33376 14764 33382 14776
rect 33502 14764 33508 14776
rect 33560 14764 33566 14816
rect 34241 14807 34299 14813
rect 34241 14773 34253 14807
rect 34287 14804 34299 14807
rect 37458 14804 37464 14816
rect 34287 14776 37464 14804
rect 34287 14773 34299 14776
rect 34241 14767 34299 14773
rect 37458 14764 37464 14776
rect 37516 14764 37522 14816
rect 37568 14804 37596 14844
rect 39666 14832 39672 14884
rect 39724 14832 39730 14884
rect 39758 14832 39764 14884
rect 39816 14872 39822 14884
rect 49145 14875 49203 14881
rect 49145 14872 49157 14875
rect 39816 14844 49157 14872
rect 39816 14832 39822 14844
rect 49145 14841 49157 14844
rect 49191 14841 49203 14875
rect 49145 14835 49203 14841
rect 38746 14804 38752 14816
rect 37568 14776 38752 14804
rect 38746 14764 38752 14776
rect 38804 14764 38810 14816
rect 41049 14807 41107 14813
rect 41049 14773 41061 14807
rect 41095 14804 41107 14807
rect 45646 14804 45652 14816
rect 41095 14776 45652 14804
rect 41095 14773 41107 14776
rect 41049 14767 41107 14773
rect 45646 14764 45652 14776
rect 45704 14764 45710 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 11238 14560 11244 14612
rect 11296 14600 11302 14612
rect 11793 14603 11851 14609
rect 11793 14600 11805 14603
rect 11296 14572 11805 14600
rect 11296 14560 11302 14572
rect 11793 14569 11805 14572
rect 11839 14569 11851 14603
rect 11793 14563 11851 14569
rect 12618 14560 12624 14612
rect 12676 14600 12682 14612
rect 12989 14603 13047 14609
rect 12989 14600 13001 14603
rect 12676 14572 13001 14600
rect 12676 14560 12682 14572
rect 12989 14569 13001 14572
rect 13035 14569 13047 14603
rect 12989 14563 13047 14569
rect 13998 14560 14004 14612
rect 14056 14600 14062 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 14056 14572 14105 14600
rect 14056 14560 14062 14572
rect 14093 14569 14105 14572
rect 14139 14569 14151 14603
rect 14093 14563 14151 14569
rect 14461 14603 14519 14609
rect 14461 14569 14473 14603
rect 14507 14600 14519 14603
rect 14642 14600 14648 14612
rect 14507 14572 14648 14600
rect 14507 14569 14519 14572
rect 14461 14563 14519 14569
rect 14642 14560 14648 14572
rect 14700 14560 14706 14612
rect 16758 14560 16764 14612
rect 16816 14600 16822 14612
rect 17402 14600 17408 14612
rect 16816 14572 17408 14600
rect 16816 14560 16822 14572
rect 17402 14560 17408 14572
rect 17460 14600 17466 14612
rect 17589 14603 17647 14609
rect 17589 14600 17601 14603
rect 17460 14572 17601 14600
rect 17460 14560 17466 14572
rect 17589 14569 17601 14572
rect 17635 14569 17647 14603
rect 17589 14563 17647 14569
rect 18141 14603 18199 14609
rect 18141 14569 18153 14603
rect 18187 14600 18199 14603
rect 18414 14600 18420 14612
rect 18187 14572 18420 14600
rect 18187 14569 18199 14572
rect 18141 14563 18199 14569
rect 18414 14560 18420 14572
rect 18472 14560 18478 14612
rect 18506 14560 18512 14612
rect 18564 14600 18570 14612
rect 18564 14572 25452 14600
rect 18564 14560 18570 14572
rect 10226 14492 10232 14544
rect 10284 14492 10290 14544
rect 10612 14504 15332 14532
rect 934 14424 940 14476
rect 992 14464 998 14476
rect 1765 14467 1823 14473
rect 1765 14464 1777 14467
rect 992 14436 1777 14464
rect 992 14424 998 14436
rect 1765 14433 1777 14436
rect 1811 14433 1823 14467
rect 1765 14427 1823 14433
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14396 3019 14399
rect 9493 14399 9551 14405
rect 9493 14396 9505 14399
rect 3007 14368 9505 14396
rect 3007 14365 3019 14368
rect 2961 14359 3019 14365
rect 9493 14365 9505 14368
rect 9539 14365 9551 14399
rect 9493 14359 9551 14365
rect 10410 14356 10416 14408
rect 10468 14356 10474 14408
rect 9677 14331 9735 14337
rect 9677 14297 9689 14331
rect 9723 14328 9735 14331
rect 9950 14328 9956 14340
rect 9723 14300 9956 14328
rect 9723 14297 9735 14300
rect 9677 14291 9735 14297
rect 9950 14288 9956 14300
rect 10008 14328 10014 14340
rect 10612 14328 10640 14504
rect 10686 14424 10692 14476
rect 10744 14464 10750 14476
rect 12250 14464 12256 14476
rect 10744 14436 12256 14464
rect 10744 14424 10750 14436
rect 12250 14424 12256 14436
rect 12308 14424 12314 14476
rect 12437 14467 12495 14473
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 13262 14464 13268 14476
rect 12483 14436 13268 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 13262 14424 13268 14436
rect 13320 14424 13326 14476
rect 13630 14424 13636 14476
rect 13688 14424 13694 14476
rect 14826 14424 14832 14476
rect 14884 14464 14890 14476
rect 15013 14467 15071 14473
rect 15013 14464 15025 14467
rect 14884 14436 15025 14464
rect 14884 14424 14890 14436
rect 15013 14433 15025 14436
rect 15059 14433 15071 14467
rect 15013 14427 15071 14433
rect 13814 14356 13820 14408
rect 13872 14396 13878 14408
rect 14921 14399 14979 14405
rect 14921 14396 14933 14399
rect 13872 14368 14933 14396
rect 13872 14356 13878 14368
rect 14921 14365 14933 14368
rect 14967 14365 14979 14399
rect 15304 14396 15332 14504
rect 20714 14492 20720 14544
rect 20772 14492 20778 14544
rect 22738 14492 22744 14544
rect 22796 14532 22802 14544
rect 22833 14535 22891 14541
rect 22833 14532 22845 14535
rect 22796 14504 22845 14532
rect 22796 14492 22802 14504
rect 22833 14501 22845 14504
rect 22879 14501 22891 14535
rect 22833 14495 22891 14501
rect 24670 14492 24676 14544
rect 24728 14492 24734 14544
rect 25424 14532 25452 14572
rect 25498 14560 25504 14612
rect 25556 14600 25562 14612
rect 25593 14603 25651 14609
rect 25593 14600 25605 14603
rect 25556 14572 25605 14600
rect 25556 14560 25562 14572
rect 25593 14569 25605 14572
rect 25639 14569 25651 14603
rect 26326 14600 26332 14612
rect 25593 14563 25651 14569
rect 25700 14572 26332 14600
rect 25700 14532 25728 14572
rect 26326 14560 26332 14572
rect 26384 14560 26390 14612
rect 26510 14560 26516 14612
rect 26568 14600 26574 14612
rect 30006 14600 30012 14612
rect 26568 14572 30012 14600
rect 26568 14560 26574 14572
rect 30006 14560 30012 14572
rect 30064 14560 30070 14612
rect 30469 14603 30527 14609
rect 30469 14569 30481 14603
rect 30515 14600 30527 14603
rect 33778 14600 33784 14612
rect 30515 14572 33784 14600
rect 30515 14569 30527 14572
rect 30469 14563 30527 14569
rect 33778 14560 33784 14572
rect 33836 14560 33842 14612
rect 36630 14560 36636 14612
rect 36688 14560 36694 14612
rect 37090 14560 37096 14612
rect 37148 14560 37154 14612
rect 38562 14560 38568 14612
rect 38620 14600 38626 14612
rect 38620 14572 38976 14600
rect 38620 14560 38626 14572
rect 25424 14504 25728 14532
rect 27430 14492 27436 14544
rect 27488 14532 27494 14544
rect 27488 14504 30696 14532
rect 27488 14492 27494 14504
rect 15378 14424 15384 14476
rect 15436 14464 15442 14476
rect 16945 14467 17003 14473
rect 16945 14464 16957 14467
rect 15436 14436 16957 14464
rect 15436 14424 15442 14436
rect 16945 14433 16957 14436
rect 16991 14433 17003 14467
rect 16945 14427 17003 14433
rect 17402 14424 17408 14476
rect 17460 14464 17466 14476
rect 17497 14467 17555 14473
rect 17497 14464 17509 14467
rect 17460 14436 17509 14464
rect 17460 14424 17466 14436
rect 17497 14433 17509 14436
rect 17543 14464 17555 14467
rect 18693 14467 18751 14473
rect 18693 14464 18705 14467
rect 17543 14436 18705 14464
rect 17543 14433 17555 14436
rect 17497 14427 17555 14433
rect 18693 14433 18705 14436
rect 18739 14433 18751 14467
rect 18693 14427 18751 14433
rect 19334 14424 19340 14476
rect 19392 14464 19398 14476
rect 20073 14467 20131 14473
rect 20073 14464 20085 14467
rect 19392 14436 20085 14464
rect 19392 14424 19398 14436
rect 20073 14433 20085 14436
rect 20119 14433 20131 14467
rect 20073 14427 20131 14433
rect 21085 14467 21143 14473
rect 21085 14433 21097 14467
rect 21131 14464 21143 14467
rect 21358 14464 21364 14476
rect 21131 14436 21364 14464
rect 21131 14433 21143 14436
rect 21085 14427 21143 14433
rect 21358 14424 21364 14436
rect 21416 14424 21422 14476
rect 21726 14424 21732 14476
rect 21784 14464 21790 14476
rect 21784 14436 27844 14464
rect 21784 14424 21790 14436
rect 16853 14399 16911 14405
rect 16853 14396 16865 14399
rect 15304 14368 16865 14396
rect 14921 14359 14979 14365
rect 16853 14365 16865 14368
rect 16899 14396 16911 14399
rect 17218 14396 17224 14408
rect 16899 14368 17224 14396
rect 16899 14365 16911 14368
rect 16853 14359 16911 14365
rect 17218 14356 17224 14368
rect 17276 14356 17282 14408
rect 17678 14356 17684 14408
rect 17736 14396 17742 14408
rect 18598 14396 18604 14408
rect 17736 14368 18604 14396
rect 17736 14356 17742 14368
rect 18598 14356 18604 14368
rect 18656 14356 18662 14408
rect 19886 14356 19892 14408
rect 19944 14396 19950 14408
rect 20438 14396 20444 14408
rect 19944 14368 20444 14396
rect 19944 14356 19950 14368
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 22646 14396 22652 14408
rect 22494 14368 22652 14396
rect 22646 14356 22652 14368
rect 22704 14396 22710 14408
rect 23014 14396 23020 14408
rect 22704 14368 23020 14396
rect 22704 14356 22710 14368
rect 23014 14356 23020 14368
rect 23072 14396 23078 14408
rect 23201 14399 23259 14405
rect 23201 14396 23213 14399
rect 23072 14368 23213 14396
rect 23072 14356 23078 14368
rect 23201 14365 23213 14368
rect 23247 14396 23259 14399
rect 23477 14399 23535 14405
rect 23477 14396 23489 14399
rect 23247 14368 23489 14396
rect 23247 14365 23259 14368
rect 23201 14359 23259 14365
rect 23477 14365 23489 14368
rect 23523 14365 23535 14399
rect 23477 14359 23535 14365
rect 27338 14356 27344 14408
rect 27396 14356 27402 14408
rect 27816 14396 27844 14436
rect 27890 14424 27896 14476
rect 27948 14424 27954 14476
rect 29362 14464 29368 14476
rect 28092 14436 29368 14464
rect 28092 14396 28120 14436
rect 29362 14424 29368 14436
rect 29420 14424 29426 14476
rect 29730 14424 29736 14476
rect 29788 14464 29794 14476
rect 29825 14467 29883 14473
rect 29825 14464 29837 14467
rect 29788 14436 29837 14464
rect 29788 14424 29794 14436
rect 29825 14433 29837 14436
rect 29871 14433 29883 14467
rect 29825 14427 29883 14433
rect 30006 14424 30012 14476
rect 30064 14424 30070 14476
rect 27816 14368 28120 14396
rect 28169 14399 28227 14405
rect 28169 14365 28181 14399
rect 28215 14396 28227 14399
rect 28626 14396 28632 14408
rect 28215 14368 28632 14396
rect 28215 14365 28227 14368
rect 28169 14359 28227 14365
rect 28626 14356 28632 14368
rect 28684 14356 28690 14408
rect 30668 14396 30696 14504
rect 31662 14492 31668 14544
rect 31720 14492 31726 14544
rect 32490 14492 32496 14544
rect 32548 14532 32554 14544
rect 34057 14535 34115 14541
rect 32548 14504 33640 14532
rect 32548 14492 32554 14504
rect 30742 14424 30748 14476
rect 30800 14464 30806 14476
rect 31021 14467 31079 14473
rect 31021 14464 31033 14467
rect 30800 14436 31033 14464
rect 30800 14424 30806 14436
rect 31021 14433 31033 14436
rect 31067 14433 31079 14467
rect 31021 14427 31079 14433
rect 31570 14424 31576 14476
rect 31628 14464 31634 14476
rect 33612 14473 33640 14504
rect 34057 14501 34069 14535
rect 34103 14532 34115 14535
rect 34103 14504 35020 14532
rect 34103 14501 34115 14504
rect 34057 14495 34115 14501
rect 32217 14467 32275 14473
rect 32217 14464 32229 14467
rect 31628 14436 32229 14464
rect 31628 14424 31634 14436
rect 32217 14433 32229 14436
rect 32263 14433 32275 14467
rect 33413 14467 33471 14473
rect 33413 14464 33425 14467
rect 32217 14427 32275 14433
rect 32324 14436 33425 14464
rect 30668 14368 31340 14396
rect 10008 14300 10640 14328
rect 10008 14288 10014 14300
rect 11238 14288 11244 14340
rect 11296 14288 11302 14340
rect 12161 14331 12219 14337
rect 12161 14297 12173 14331
rect 12207 14328 12219 14331
rect 12802 14328 12808 14340
rect 12207 14300 12808 14328
rect 12207 14297 12219 14300
rect 12161 14291 12219 14297
rect 12802 14288 12808 14300
rect 12860 14288 12866 14340
rect 13357 14331 13415 14337
rect 13357 14297 13369 14331
rect 13403 14328 13415 14331
rect 15933 14331 15991 14337
rect 13403 14300 15056 14328
rect 13403 14297 13415 14300
rect 13357 14291 13415 14297
rect 10502 14220 10508 14272
rect 10560 14260 10566 14272
rect 11149 14263 11207 14269
rect 11149 14260 11161 14263
rect 10560 14232 11161 14260
rect 10560 14220 10566 14232
rect 11149 14229 11161 14232
rect 11195 14229 11207 14263
rect 11149 14223 11207 14229
rect 12253 14263 12311 14269
rect 12253 14229 12265 14263
rect 12299 14260 12311 14263
rect 12710 14260 12716 14272
rect 12299 14232 12716 14260
rect 12299 14229 12311 14232
rect 12253 14223 12311 14229
rect 12710 14220 12716 14232
rect 12768 14220 12774 14272
rect 13449 14263 13507 14269
rect 13449 14229 13461 14263
rect 13495 14260 13507 14263
rect 13998 14260 14004 14272
rect 13495 14232 14004 14260
rect 13495 14229 13507 14232
rect 13449 14223 13507 14229
rect 13998 14220 14004 14232
rect 14056 14220 14062 14272
rect 14182 14220 14188 14272
rect 14240 14260 14246 14272
rect 14829 14263 14887 14269
rect 14829 14260 14841 14263
rect 14240 14232 14841 14260
rect 14240 14220 14246 14232
rect 14829 14229 14841 14232
rect 14875 14229 14887 14263
rect 15028 14260 15056 14300
rect 15933 14297 15945 14331
rect 15979 14328 15991 14331
rect 16761 14331 16819 14337
rect 16761 14328 16773 14331
rect 15979 14300 16773 14328
rect 15979 14297 15991 14300
rect 15933 14291 15991 14297
rect 16761 14297 16773 14300
rect 16807 14297 16819 14331
rect 16761 14291 16819 14297
rect 16942 14288 16948 14340
rect 17000 14328 17006 14340
rect 17310 14328 17316 14340
rect 17000 14300 17316 14328
rect 17000 14288 17006 14300
rect 17310 14288 17316 14300
rect 17368 14288 17374 14340
rect 17865 14331 17923 14337
rect 17865 14297 17877 14331
rect 17911 14328 17923 14331
rect 19426 14328 19432 14340
rect 17911 14300 19432 14328
rect 17911 14297 17923 14300
rect 17865 14291 17923 14297
rect 19426 14288 19432 14300
rect 19484 14288 19490 14340
rect 19996 14300 21220 14328
rect 16393 14263 16451 14269
rect 16393 14260 16405 14263
rect 15028 14232 16405 14260
rect 14829 14223 14887 14229
rect 16393 14229 16405 14232
rect 16439 14229 16451 14263
rect 16393 14223 16451 14229
rect 17494 14220 17500 14272
rect 17552 14260 17558 14272
rect 17954 14260 17960 14272
rect 17552 14232 17960 14260
rect 17552 14220 17558 14232
rect 17954 14220 17960 14232
rect 18012 14220 18018 14272
rect 18046 14220 18052 14272
rect 18104 14260 18110 14272
rect 18414 14260 18420 14272
rect 18104 14232 18420 14260
rect 18104 14220 18110 14232
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 18509 14263 18567 14269
rect 18509 14229 18521 14263
rect 18555 14260 18567 14263
rect 18966 14260 18972 14272
rect 18555 14232 18972 14260
rect 18555 14229 18567 14232
rect 18509 14223 18567 14229
rect 18966 14220 18972 14232
rect 19024 14220 19030 14272
rect 19518 14220 19524 14272
rect 19576 14220 19582 14272
rect 19794 14220 19800 14272
rect 19852 14260 19858 14272
rect 19996 14269 20024 14300
rect 19981 14263 20039 14269
rect 19981 14260 19993 14263
rect 19852 14232 19993 14260
rect 19852 14220 19858 14232
rect 19981 14229 19993 14232
rect 20027 14229 20039 14263
rect 19981 14223 20039 14229
rect 20530 14220 20536 14272
rect 20588 14220 20594 14272
rect 21192 14260 21220 14300
rect 21266 14288 21272 14340
rect 21324 14328 21330 14340
rect 21361 14331 21419 14337
rect 21361 14328 21373 14331
rect 21324 14300 21373 14328
rect 21324 14288 21330 14300
rect 21361 14297 21373 14300
rect 21407 14297 21419 14331
rect 21361 14291 21419 14297
rect 24486 14288 24492 14340
rect 24544 14328 24550 14340
rect 24544 14300 25268 14328
rect 24544 14288 24550 14300
rect 21726 14260 21732 14272
rect 21192 14232 21732 14260
rect 21726 14220 21732 14232
rect 21784 14220 21790 14272
rect 23842 14220 23848 14272
rect 23900 14220 23906 14272
rect 24394 14220 24400 14272
rect 24452 14220 24458 14272
rect 25130 14220 25136 14272
rect 25188 14220 25194 14272
rect 25240 14260 25268 14300
rect 25774 14288 25780 14340
rect 25832 14328 25838 14340
rect 25832 14300 25898 14328
rect 25832 14288 25838 14300
rect 27062 14288 27068 14340
rect 27120 14288 27126 14340
rect 31205 14331 31263 14337
rect 31205 14328 31217 14331
rect 28552 14300 31217 14328
rect 27706 14260 27712 14272
rect 25240 14232 27712 14260
rect 27706 14220 27712 14232
rect 27764 14260 27770 14272
rect 28077 14263 28135 14269
rect 28077 14260 28089 14263
rect 27764 14232 28089 14260
rect 27764 14220 27770 14232
rect 28077 14229 28089 14232
rect 28123 14260 28135 14263
rect 28442 14260 28448 14272
rect 28123 14232 28448 14260
rect 28123 14229 28135 14232
rect 28077 14223 28135 14229
rect 28442 14220 28448 14232
rect 28500 14220 28506 14272
rect 28552 14269 28580 14300
rect 31205 14297 31217 14300
rect 31251 14297 31263 14331
rect 31312 14328 31340 14368
rect 31846 14356 31852 14408
rect 31904 14396 31910 14408
rect 32324 14396 32352 14436
rect 33413 14433 33425 14436
rect 33459 14433 33471 14467
rect 33413 14427 33471 14433
rect 33597 14467 33655 14473
rect 33597 14433 33609 14467
rect 33643 14433 33655 14467
rect 33597 14427 33655 14433
rect 34790 14424 34796 14476
rect 34848 14464 34854 14476
rect 34885 14467 34943 14473
rect 34885 14464 34897 14467
rect 34848 14436 34897 14464
rect 34848 14424 34854 14436
rect 34885 14433 34897 14436
rect 34931 14433 34943 14467
rect 34992 14464 35020 14504
rect 36354 14492 36360 14544
rect 36412 14532 36418 14544
rect 37108 14532 37136 14560
rect 36412 14504 37136 14532
rect 36412 14492 36418 14504
rect 37090 14464 37096 14476
rect 34992 14436 37096 14464
rect 34885 14427 34943 14433
rect 37090 14424 37096 14436
rect 37148 14424 37154 14476
rect 37366 14424 37372 14476
rect 37424 14464 37430 14476
rect 38841 14467 38899 14473
rect 38841 14464 38853 14467
rect 37424 14436 38853 14464
rect 37424 14424 37430 14436
rect 38841 14433 38853 14436
rect 38887 14433 38899 14467
rect 38841 14427 38899 14433
rect 31904 14368 32352 14396
rect 31904 14356 31910 14368
rect 32950 14356 32956 14408
rect 33008 14396 33014 14408
rect 33689 14399 33747 14405
rect 33689 14396 33701 14399
rect 33008 14368 33701 14396
rect 33008 14356 33014 14368
rect 33689 14365 33701 14368
rect 33735 14365 33747 14399
rect 38948 14396 38976 14572
rect 39942 14560 39948 14612
rect 40000 14600 40006 14612
rect 40037 14603 40095 14609
rect 40037 14600 40049 14603
rect 40000 14572 40049 14600
rect 40000 14560 40006 14572
rect 40037 14569 40049 14572
rect 40083 14569 40095 14603
rect 40037 14563 40095 14569
rect 39301 14399 39359 14405
rect 39301 14396 39313 14399
rect 38948 14368 39313 14396
rect 33689 14359 33747 14365
rect 39301 14365 39313 14368
rect 39347 14365 39359 14399
rect 39301 14359 39359 14365
rect 49050 14356 49056 14408
rect 49108 14356 49114 14408
rect 49234 14356 49240 14408
rect 49292 14356 49298 14408
rect 32401 14331 32459 14337
rect 32401 14328 32413 14331
rect 31312 14300 32413 14328
rect 31205 14291 31263 14297
rect 32401 14297 32413 14300
rect 32447 14297 32459 14331
rect 32401 14291 32459 14297
rect 32493 14331 32551 14337
rect 32493 14297 32505 14331
rect 32539 14328 32551 14331
rect 33502 14328 33508 14340
rect 32539 14300 33508 14328
rect 32539 14297 32551 14300
rect 32493 14291 32551 14297
rect 33502 14288 33508 14300
rect 33560 14288 33566 14340
rect 34606 14288 34612 14340
rect 34664 14328 34670 14340
rect 35158 14328 35164 14340
rect 34664 14300 35164 14328
rect 34664 14288 34670 14300
rect 35158 14288 35164 14300
rect 35216 14288 35222 14340
rect 35618 14288 35624 14340
rect 35676 14288 35682 14340
rect 36814 14288 36820 14340
rect 36872 14328 36878 14340
rect 38565 14331 38623 14337
rect 36872 14300 37398 14328
rect 36872 14288 36878 14300
rect 38565 14297 38577 14331
rect 38611 14297 38623 14331
rect 38565 14291 38623 14297
rect 48593 14331 48651 14337
rect 48593 14297 48605 14331
rect 48639 14328 48651 14331
rect 49252 14328 49280 14356
rect 48639 14300 49280 14328
rect 48639 14297 48651 14300
rect 48593 14291 48651 14297
rect 28537 14263 28595 14269
rect 28537 14229 28549 14263
rect 28583 14229 28595 14263
rect 28537 14223 28595 14229
rect 28994 14220 29000 14272
rect 29052 14220 29058 14272
rect 29638 14220 29644 14272
rect 29696 14260 29702 14272
rect 30006 14260 30012 14272
rect 29696 14232 30012 14260
rect 29696 14220 29702 14232
rect 30006 14220 30012 14232
rect 30064 14220 30070 14272
rect 30101 14263 30159 14269
rect 30101 14229 30113 14263
rect 30147 14260 30159 14263
rect 30282 14260 30288 14272
rect 30147 14232 30288 14260
rect 30147 14229 30159 14232
rect 30101 14223 30159 14229
rect 30282 14220 30288 14232
rect 30340 14220 30346 14272
rect 31018 14220 31024 14272
rect 31076 14260 31082 14272
rect 31297 14263 31355 14269
rect 31297 14260 31309 14263
rect 31076 14232 31309 14260
rect 31076 14220 31082 14232
rect 31297 14229 31309 14232
rect 31343 14229 31355 14263
rect 31297 14223 31355 14229
rect 32766 14220 32772 14272
rect 32824 14260 32830 14272
rect 32861 14263 32919 14269
rect 32861 14260 32873 14263
rect 32824 14232 32873 14260
rect 32824 14220 32830 14232
rect 32861 14229 32873 14232
rect 32907 14229 32919 14263
rect 32861 14223 32919 14229
rect 33410 14220 33416 14272
rect 33468 14260 33474 14272
rect 34333 14263 34391 14269
rect 34333 14260 34345 14263
rect 33468 14232 34345 14260
rect 33468 14220 33474 14232
rect 34333 14229 34345 14232
rect 34379 14229 34391 14263
rect 34333 14223 34391 14229
rect 34882 14220 34888 14272
rect 34940 14260 34946 14272
rect 37550 14260 37556 14272
rect 34940 14232 37556 14260
rect 34940 14220 34946 14232
rect 37550 14220 37556 14232
rect 37608 14220 37614 14272
rect 37642 14220 37648 14272
rect 37700 14260 37706 14272
rect 38580 14260 38608 14291
rect 37700 14232 38608 14260
rect 37700 14220 37706 14232
rect 39482 14220 39488 14272
rect 39540 14220 39546 14272
rect 48314 14220 48320 14272
rect 48372 14260 48378 14272
rect 48685 14263 48743 14269
rect 48685 14260 48697 14263
rect 48372 14232 48697 14260
rect 48372 14220 48378 14232
rect 48685 14229 48697 14232
rect 48731 14229 48743 14263
rect 48685 14223 48743 14229
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 3605 14059 3663 14065
rect 3605 14025 3617 14059
rect 3651 14056 3663 14059
rect 9858 14056 9864 14068
rect 3651 14028 9864 14056
rect 3651 14025 3663 14028
rect 3605 14019 3663 14025
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 9950 14016 9956 14068
rect 10008 14016 10014 14068
rect 10410 14016 10416 14068
rect 10468 14016 10474 14068
rect 11882 14016 11888 14068
rect 11940 14056 11946 14068
rect 11977 14059 12035 14065
rect 11977 14056 11989 14059
rect 11940 14028 11989 14056
rect 11940 14016 11946 14028
rect 11977 14025 11989 14028
rect 12023 14025 12035 14059
rect 11977 14019 12035 14025
rect 12894 14016 12900 14068
rect 12952 14056 12958 14068
rect 14182 14056 14188 14068
rect 12952 14028 14188 14056
rect 12952 14016 12958 14028
rect 14182 14016 14188 14028
rect 14240 14016 14246 14068
rect 14274 14016 14280 14068
rect 14332 14056 14338 14068
rect 15565 14059 15623 14065
rect 15565 14056 15577 14059
rect 14332 14028 15577 14056
rect 14332 14016 14338 14028
rect 15565 14025 15577 14028
rect 15611 14025 15623 14059
rect 15565 14019 15623 14025
rect 15930 14016 15936 14068
rect 15988 14016 15994 14068
rect 16574 14016 16580 14068
rect 16632 14056 16638 14068
rect 17129 14059 17187 14065
rect 17129 14056 17141 14059
rect 16632 14028 17141 14056
rect 16632 14016 16638 14028
rect 17129 14025 17141 14028
rect 17175 14025 17187 14059
rect 17129 14019 17187 14025
rect 17494 14016 17500 14068
rect 17552 14016 17558 14068
rect 17586 14016 17592 14068
rect 17644 14016 17650 14068
rect 18322 14016 18328 14068
rect 18380 14016 18386 14068
rect 18693 14059 18751 14065
rect 18693 14025 18705 14059
rect 18739 14056 18751 14059
rect 18782 14056 18788 14068
rect 18739 14028 18788 14056
rect 18739 14025 18751 14028
rect 18693 14019 18751 14025
rect 18782 14016 18788 14028
rect 18840 14016 18846 14068
rect 19429 14059 19487 14065
rect 19429 14025 19441 14059
rect 19475 14056 19487 14059
rect 19886 14056 19892 14068
rect 19475 14028 19892 14056
rect 19475 14025 19487 14028
rect 19429 14019 19487 14025
rect 19886 14016 19892 14028
rect 19944 14016 19950 14068
rect 21266 14016 21272 14068
rect 21324 14056 21330 14068
rect 21453 14059 21511 14065
rect 21453 14056 21465 14059
rect 21324 14028 21465 14056
rect 21324 14016 21330 14028
rect 21453 14025 21465 14028
rect 21499 14025 21511 14059
rect 21453 14019 21511 14025
rect 21542 14016 21548 14068
rect 21600 14056 21606 14068
rect 24486 14056 24492 14068
rect 21600 14028 24492 14056
rect 21600 14016 21606 14028
rect 24486 14016 24492 14028
rect 24544 14016 24550 14068
rect 24857 14059 24915 14065
rect 24857 14025 24869 14059
rect 24903 14056 24915 14059
rect 25314 14056 25320 14068
rect 24903 14028 25320 14056
rect 24903 14025 24915 14028
rect 24857 14019 24915 14025
rect 25314 14016 25320 14028
rect 25372 14016 25378 14068
rect 25498 14016 25504 14068
rect 25556 14056 25562 14068
rect 25556 14028 26004 14056
rect 25556 14016 25562 14028
rect 1026 13948 1032 14000
rect 1084 13988 1090 14000
rect 1765 13991 1823 13997
rect 1765 13988 1777 13991
rect 1084 13960 1777 13988
rect 1084 13948 1090 13960
rect 1765 13957 1777 13960
rect 1811 13957 1823 13991
rect 10502 13988 10508 14000
rect 1765 13951 1823 13957
rect 2976 13960 10508 13988
rect 2976 13929 3004 13960
rect 10502 13948 10508 13960
rect 10560 13948 10566 14000
rect 10689 13991 10747 13997
rect 10689 13957 10701 13991
rect 10735 13988 10747 13991
rect 11238 13988 11244 14000
rect 10735 13960 11244 13988
rect 10735 13957 10747 13960
rect 10689 13951 10747 13957
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 13262 13948 13268 14000
rect 13320 13948 13326 14000
rect 13722 13948 13728 14000
rect 13780 13948 13786 14000
rect 15010 13988 15016 14000
rect 14660 13960 15016 13988
rect 2961 13923 3019 13929
rect 2961 13889 2973 13923
rect 3007 13889 3019 13923
rect 2961 13883 3019 13889
rect 3510 13880 3516 13932
rect 3568 13920 3574 13932
rect 3973 13923 4031 13929
rect 3973 13920 3985 13923
rect 3568 13892 3985 13920
rect 3568 13880 3574 13892
rect 3973 13889 3985 13892
rect 4019 13889 4031 13923
rect 3973 13883 4031 13889
rect 11149 13923 11207 13929
rect 11149 13889 11161 13923
rect 11195 13920 11207 13923
rect 12069 13923 12127 13929
rect 12069 13920 12081 13923
rect 11195 13892 12081 13920
rect 11195 13889 11207 13892
rect 11149 13883 11207 13889
rect 12069 13889 12081 13892
rect 12115 13889 12127 13923
rect 12069 13883 12127 13889
rect 11885 13855 11943 13861
rect 11885 13821 11897 13855
rect 11931 13852 11943 13855
rect 12250 13852 12256 13864
rect 11931 13824 12256 13852
rect 11931 13821 11943 13824
rect 11885 13815 11943 13821
rect 12250 13812 12256 13824
rect 12308 13812 12314 13864
rect 12989 13855 13047 13861
rect 12989 13821 13001 13855
rect 13035 13821 13047 13855
rect 12989 13815 13047 13821
rect 12342 13744 12348 13796
rect 12400 13784 12406 13796
rect 12437 13787 12495 13793
rect 12437 13784 12449 13787
rect 12400 13756 12449 13784
rect 12400 13744 12406 13756
rect 12437 13753 12449 13756
rect 12483 13753 12495 13787
rect 12437 13747 12495 13753
rect 10778 13676 10784 13728
rect 10836 13716 10842 13728
rect 13004 13716 13032 13815
rect 13722 13812 13728 13864
rect 13780 13852 13786 13864
rect 14458 13852 14464 13864
rect 13780 13824 14464 13852
rect 13780 13812 13786 13824
rect 14458 13812 14464 13824
rect 14516 13852 14522 13864
rect 14660 13852 14688 13960
rect 15010 13948 15016 13960
rect 15068 13948 15074 14000
rect 15286 13948 15292 14000
rect 15344 13948 15350 14000
rect 16025 13991 16083 13997
rect 16025 13957 16037 13991
rect 16071 13988 16083 13991
rect 19518 13988 19524 14000
rect 16071 13960 19524 13988
rect 16071 13957 16083 13960
rect 16025 13951 16083 13957
rect 19518 13948 19524 13960
rect 19576 13948 19582 14000
rect 20714 13948 20720 14000
rect 20772 13948 20778 14000
rect 23014 13948 23020 14000
rect 23072 13948 23078 14000
rect 25774 13948 25780 14000
rect 25832 13948 25838 14000
rect 25976 13988 26004 14028
rect 27614 14016 27620 14068
rect 27672 14016 27678 14068
rect 29365 14059 29423 14065
rect 29365 14025 29377 14059
rect 29411 14025 29423 14059
rect 29365 14019 29423 14025
rect 26329 13991 26387 13997
rect 26329 13988 26341 13991
rect 25976 13960 26341 13988
rect 26329 13957 26341 13960
rect 26375 13957 26387 13991
rect 26329 13951 26387 13957
rect 27062 13948 27068 14000
rect 27120 13988 27126 14000
rect 27522 13988 27528 14000
rect 27120 13960 27528 13988
rect 27120 13948 27126 13960
rect 27522 13948 27528 13960
rect 27580 13988 27586 14000
rect 29380 13988 29408 14019
rect 30006 14016 30012 14068
rect 30064 14056 30070 14068
rect 31110 14056 31116 14068
rect 30064 14028 31116 14056
rect 30064 14016 30070 14028
rect 31110 14016 31116 14028
rect 31168 14016 31174 14068
rect 31757 14059 31815 14065
rect 31757 14025 31769 14059
rect 31803 14056 31815 14059
rect 36081 14059 36139 14065
rect 36081 14056 36093 14059
rect 31803 14028 36093 14056
rect 31803 14025 31815 14028
rect 31757 14019 31815 14025
rect 36081 14025 36093 14028
rect 36127 14025 36139 14059
rect 36081 14019 36139 14025
rect 36449 14059 36507 14065
rect 36449 14025 36461 14059
rect 36495 14056 36507 14059
rect 37829 14059 37887 14065
rect 37829 14056 37841 14059
rect 36495 14028 37841 14056
rect 36495 14025 36507 14028
rect 36449 14019 36507 14025
rect 37829 14025 37841 14028
rect 37875 14025 37887 14059
rect 37829 14019 37887 14025
rect 38197 14059 38255 14065
rect 38197 14025 38209 14059
rect 38243 14056 38255 14059
rect 41322 14056 41328 14068
rect 38243 14028 41328 14056
rect 38243 14025 38255 14028
rect 38197 14019 38255 14025
rect 41322 14016 41328 14028
rect 41380 14016 41386 14068
rect 45833 14059 45891 14065
rect 45833 14025 45845 14059
rect 45879 14056 45891 14059
rect 47026 14056 47032 14068
rect 45879 14028 47032 14056
rect 45879 14025 45891 14028
rect 45833 14019 45891 14025
rect 47026 14016 47032 14028
rect 47084 14016 47090 14068
rect 48406 14016 48412 14068
rect 48464 14016 48470 14068
rect 49142 14016 49148 14068
rect 49200 14016 49206 14068
rect 27580 13960 29408 13988
rect 27580 13948 27586 13960
rect 31202 13948 31208 14000
rect 31260 13988 31266 14000
rect 31260 13960 32614 13988
rect 31260 13948 31266 13960
rect 33686 13948 33692 14000
rect 33744 13988 33750 14000
rect 34885 13991 34943 13997
rect 34885 13988 34897 13991
rect 33744 13960 34897 13988
rect 33744 13948 33750 13960
rect 34885 13957 34897 13960
rect 34931 13957 34943 13991
rect 34885 13951 34943 13957
rect 35158 13948 35164 14000
rect 35216 13988 35222 14000
rect 35216 13960 36216 13988
rect 35216 13948 35222 13960
rect 16482 13920 16488 13932
rect 14752 13892 16488 13920
rect 14752 13861 14780 13892
rect 16482 13880 16488 13892
rect 16540 13880 16546 13932
rect 16853 13923 16911 13929
rect 16853 13889 16865 13923
rect 16899 13920 16911 13923
rect 17034 13920 17040 13932
rect 16899 13892 17040 13920
rect 16899 13889 16911 13892
rect 16853 13883 16911 13889
rect 17034 13880 17040 13892
rect 17092 13920 17098 13932
rect 17586 13920 17592 13932
rect 17092 13892 17592 13920
rect 17092 13880 17098 13892
rect 17586 13880 17592 13892
rect 17644 13880 17650 13932
rect 18785 13923 18843 13929
rect 18785 13889 18797 13923
rect 18831 13920 18843 13923
rect 19426 13920 19432 13932
rect 18831 13892 19432 13920
rect 18831 13889 18843 13892
rect 18785 13883 18843 13889
rect 19426 13880 19432 13892
rect 19484 13880 19490 13932
rect 24302 13920 24308 13932
rect 23768 13892 24308 13920
rect 14516 13824 14688 13852
rect 14737 13855 14795 13861
rect 14516 13812 14522 13824
rect 14737 13821 14749 13855
rect 14783 13821 14795 13855
rect 14737 13815 14795 13821
rect 16206 13812 16212 13864
rect 16264 13812 16270 13864
rect 17773 13855 17831 13861
rect 17773 13821 17785 13855
rect 17819 13821 17831 13855
rect 17773 13815 17831 13821
rect 14936 13756 15148 13784
rect 13630 13716 13636 13728
rect 10836 13688 13636 13716
rect 10836 13676 10842 13688
rect 13630 13676 13636 13688
rect 13688 13676 13694 13728
rect 14642 13676 14648 13728
rect 14700 13716 14706 13728
rect 14936 13716 14964 13756
rect 14700 13688 14964 13716
rect 15120 13716 15148 13756
rect 15286 13744 15292 13796
rect 15344 13784 15350 13796
rect 17126 13784 17132 13796
rect 15344 13756 17132 13784
rect 15344 13744 15350 13756
rect 17126 13744 17132 13756
rect 17184 13744 17190 13796
rect 17788 13784 17816 13815
rect 18874 13812 18880 13864
rect 18932 13812 18938 13864
rect 18966 13812 18972 13864
rect 19024 13852 19030 13864
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 19024 13824 19717 13852
rect 19024 13812 19030 13824
rect 19705 13821 19717 13824
rect 19751 13821 19763 13855
rect 19705 13815 19763 13821
rect 20714 13812 20720 13864
rect 20772 13852 20778 13864
rect 22002 13852 22008 13864
rect 20772 13824 21128 13852
rect 20772 13812 20778 13824
rect 21100 13796 21128 13824
rect 21376 13824 22008 13852
rect 17954 13784 17960 13796
rect 17788 13756 17960 13784
rect 17954 13744 17960 13756
rect 18012 13744 18018 13796
rect 21082 13744 21088 13796
rect 21140 13744 21146 13796
rect 19794 13716 19800 13728
rect 15120 13688 19800 13716
rect 14700 13676 14706 13688
rect 19794 13676 19800 13688
rect 19852 13676 19858 13728
rect 19978 13725 19984 13728
rect 19968 13719 19984 13725
rect 19968 13685 19980 13719
rect 20036 13716 20042 13728
rect 21376 13716 21404 13824
rect 22002 13812 22008 13824
rect 22060 13812 22066 13864
rect 23768 13861 23796 13892
rect 24302 13880 24308 13892
rect 24360 13880 24366 13932
rect 28902 13880 28908 13932
rect 28960 13880 28966 13932
rect 29270 13880 29276 13932
rect 29328 13920 29334 13932
rect 29328 13892 29762 13920
rect 29328 13880 29334 13892
rect 31110 13880 31116 13932
rect 31168 13880 31174 13932
rect 31938 13880 31944 13932
rect 31996 13920 32002 13932
rect 32490 13920 32496 13932
rect 31996 13892 32496 13920
rect 31996 13880 32002 13892
rect 32490 13880 32496 13892
rect 32548 13880 32554 13932
rect 34146 13880 34152 13932
rect 34204 13920 34210 13932
rect 34793 13923 34851 13929
rect 34793 13920 34805 13923
rect 34204 13892 34805 13920
rect 34204 13880 34210 13892
rect 34793 13889 34805 13892
rect 34839 13889 34851 13923
rect 36078 13920 36084 13932
rect 34793 13883 34851 13889
rect 35268 13892 36084 13920
rect 23477 13855 23535 13861
rect 23477 13852 23489 13855
rect 22112 13824 23489 13852
rect 21910 13744 21916 13796
rect 21968 13784 21974 13796
rect 22112 13784 22140 13824
rect 23477 13821 23489 13824
rect 23523 13852 23535 13855
rect 23753 13855 23811 13861
rect 23523 13824 23704 13852
rect 23523 13821 23535 13824
rect 23477 13815 23535 13821
rect 21968 13756 22140 13784
rect 23676 13784 23704 13824
rect 23753 13821 23765 13855
rect 23799 13821 23811 13855
rect 23753 13815 23811 13821
rect 23934 13812 23940 13864
rect 23992 13852 23998 13864
rect 24213 13855 24271 13861
rect 24213 13852 24225 13855
rect 23992 13824 24225 13852
rect 23992 13812 23998 13824
rect 24213 13821 24225 13824
rect 24259 13821 24271 13855
rect 24213 13815 24271 13821
rect 26605 13855 26663 13861
rect 26605 13821 26617 13855
rect 26651 13852 26663 13855
rect 27338 13852 27344 13864
rect 26651 13824 27344 13852
rect 26651 13821 26663 13824
rect 26605 13815 26663 13821
rect 27338 13812 27344 13824
rect 27396 13812 27402 13864
rect 30282 13852 30288 13864
rect 29748 13824 30288 13852
rect 29748 13796 29776 13824
rect 30282 13812 30288 13824
rect 30340 13812 30346 13864
rect 30837 13855 30895 13861
rect 30837 13821 30849 13855
rect 30883 13852 30895 13855
rect 32306 13852 32312 13864
rect 30883 13824 31064 13852
rect 30883 13821 30895 13824
rect 30837 13815 30895 13821
rect 24578 13784 24584 13796
rect 23676 13756 24584 13784
rect 21968 13744 21974 13756
rect 24578 13744 24584 13756
rect 24636 13744 24642 13796
rect 29730 13744 29736 13796
rect 29788 13744 29794 13796
rect 31036 13784 31064 13824
rect 31726 13824 32312 13852
rect 31726 13784 31754 13824
rect 32306 13812 32312 13824
rect 32364 13812 32370 13864
rect 34054 13812 34060 13864
rect 34112 13812 34118 13864
rect 34609 13855 34667 13861
rect 34609 13821 34621 13855
rect 34655 13821 34667 13855
rect 34609 13815 34667 13821
rect 31036 13756 31754 13784
rect 34624 13784 34652 13815
rect 34698 13784 34704 13796
rect 34624 13756 34704 13784
rect 34698 13744 34704 13756
rect 34756 13744 34762 13796
rect 35268 13793 35296 13892
rect 36078 13880 36084 13892
rect 36136 13880 36142 13932
rect 36188 13920 36216 13960
rect 36722 13948 36728 14000
rect 36780 13988 36786 14000
rect 37737 13991 37795 13997
rect 37737 13988 37749 13991
rect 36780 13960 37749 13988
rect 36780 13948 36786 13960
rect 37737 13957 37749 13960
rect 37783 13957 37795 13991
rect 37737 13951 37795 13957
rect 38565 13991 38623 13997
rect 38565 13957 38577 13991
rect 38611 13988 38623 13991
rect 38654 13988 38660 14000
rect 38611 13960 38660 13988
rect 38611 13957 38623 13960
rect 38565 13951 38623 13957
rect 38654 13948 38660 13960
rect 38712 13988 38718 14000
rect 38933 13991 38991 13997
rect 38933 13988 38945 13991
rect 38712 13960 38945 13988
rect 38712 13948 38718 13960
rect 38933 13957 38945 13960
rect 38979 13957 38991 13991
rect 38933 13951 38991 13957
rect 39482 13948 39488 14000
rect 39540 13988 39546 14000
rect 45005 13991 45063 13997
rect 45005 13988 45017 13991
rect 39540 13960 45017 13988
rect 39540 13948 39546 13960
rect 45005 13957 45017 13960
rect 45051 13957 45063 13991
rect 45005 13951 45063 13957
rect 48133 13991 48191 13997
rect 48133 13957 48145 13991
rect 48179 13988 48191 13991
rect 49234 13988 49240 14000
rect 48179 13960 49240 13988
rect 48179 13957 48191 13960
rect 48133 13951 48191 13957
rect 49234 13948 49240 13960
rect 49292 13948 49298 14000
rect 36909 13923 36967 13929
rect 36909 13920 36921 13923
rect 36188 13892 36921 13920
rect 36909 13889 36921 13892
rect 36955 13889 36967 13923
rect 36909 13883 36967 13889
rect 45646 13880 45652 13932
rect 45704 13880 45710 13932
rect 48222 13880 48228 13932
rect 48280 13920 48286 13932
rect 48593 13923 48651 13929
rect 48593 13920 48605 13923
rect 48280 13892 48605 13920
rect 48280 13880 48286 13892
rect 48593 13889 48605 13892
rect 48639 13889 48651 13923
rect 48593 13883 48651 13889
rect 35897 13855 35955 13861
rect 35897 13821 35909 13855
rect 35943 13821 35955 13855
rect 35897 13815 35955 13821
rect 35253 13787 35311 13793
rect 35253 13753 35265 13787
rect 35299 13753 35311 13787
rect 35912 13784 35940 13815
rect 35986 13812 35992 13864
rect 36044 13812 36050 13864
rect 37645 13855 37703 13861
rect 37645 13821 37657 13855
rect 37691 13821 37703 13855
rect 37645 13815 37703 13821
rect 45189 13855 45247 13861
rect 45189 13821 45201 13855
rect 45235 13852 45247 13855
rect 46290 13852 46296 13864
rect 45235 13824 46296 13852
rect 45235 13821 45247 13824
rect 45189 13815 45247 13821
rect 36630 13784 36636 13796
rect 35912 13756 36636 13784
rect 35253 13747 35311 13753
rect 36630 13744 36636 13756
rect 36688 13744 36694 13796
rect 37660 13784 37688 13815
rect 46290 13812 46296 13824
rect 46348 13812 46354 13864
rect 38194 13784 38200 13796
rect 37660 13756 38200 13784
rect 38194 13744 38200 13756
rect 38252 13744 38258 13796
rect 20036 13688 21404 13716
rect 19968 13679 19984 13685
rect 19978 13676 19984 13679
rect 20036 13676 20042 13688
rect 22830 13676 22836 13728
rect 22888 13716 22894 13728
rect 26326 13716 26332 13728
rect 22888 13688 26332 13716
rect 22888 13676 22894 13688
rect 26326 13676 26332 13688
rect 26384 13676 26390 13728
rect 30834 13676 30840 13728
rect 30892 13716 30898 13728
rect 33799 13719 33857 13725
rect 33799 13716 33811 13719
rect 30892 13688 33811 13716
rect 30892 13676 30898 13688
rect 33799 13685 33811 13688
rect 33845 13716 33857 13719
rect 36354 13716 36360 13728
rect 33845 13688 36360 13716
rect 33845 13685 33857 13688
rect 33799 13679 33857 13685
rect 36354 13676 36360 13688
rect 36412 13676 36418 13728
rect 36722 13676 36728 13728
rect 36780 13676 36786 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 9646 13484 12112 13512
rect 9646 13444 9674 13484
rect 2976 13416 9674 13444
rect 1762 13336 1768 13388
rect 1820 13336 1826 13388
rect 2976 13317 3004 13416
rect 10502 13404 10508 13456
rect 10560 13444 10566 13456
rect 12084 13444 12112 13484
rect 12250 13472 12256 13524
rect 12308 13512 12314 13524
rect 12529 13515 12587 13521
rect 12529 13512 12541 13515
rect 12308 13484 12541 13512
rect 12308 13472 12314 13484
rect 12529 13481 12541 13484
rect 12575 13512 12587 13515
rect 12986 13512 12992 13524
rect 12575 13484 12992 13512
rect 12575 13481 12587 13484
rect 12529 13475 12587 13481
rect 12986 13472 12992 13484
rect 13044 13472 13050 13524
rect 13722 13472 13728 13524
rect 13780 13472 13786 13524
rect 14182 13472 14188 13524
rect 14240 13512 14246 13524
rect 14921 13515 14979 13521
rect 14240 13484 14412 13512
rect 14240 13472 14246 13484
rect 14277 13447 14335 13453
rect 14277 13444 14289 13447
rect 10560 13416 10916 13444
rect 12084 13416 14289 13444
rect 10560 13404 10566 13416
rect 10778 13336 10784 13388
rect 10836 13336 10842 13388
rect 10888 13376 10916 13416
rect 14277 13413 14289 13416
rect 14323 13413 14335 13447
rect 14384 13444 14412 13484
rect 14921 13481 14933 13515
rect 14967 13512 14979 13515
rect 15010 13512 15016 13524
rect 14967 13484 15016 13512
rect 14967 13481 14979 13484
rect 14921 13475 14979 13481
rect 15010 13472 15016 13484
rect 15068 13472 15074 13524
rect 17954 13512 17960 13524
rect 15396 13484 17960 13512
rect 15194 13444 15200 13456
rect 14384 13416 15200 13444
rect 14277 13407 14335 13413
rect 15194 13404 15200 13416
rect 15252 13404 15258 13456
rect 11146 13376 11152 13388
rect 10888 13348 11152 13376
rect 11146 13336 11152 13348
rect 11204 13336 11210 13388
rect 12894 13336 12900 13388
rect 12952 13376 12958 13388
rect 13081 13379 13139 13385
rect 13081 13376 13093 13379
rect 12952 13348 13093 13376
rect 12952 13336 12958 13348
rect 13081 13345 13093 13348
rect 13127 13345 13139 13379
rect 13081 13339 13139 13345
rect 13814 13336 13820 13388
rect 13872 13376 13878 13388
rect 13909 13379 13967 13385
rect 13909 13376 13921 13379
rect 13872 13348 13921 13376
rect 13872 13336 13878 13348
rect 13909 13345 13921 13348
rect 13955 13376 13967 13379
rect 14826 13376 14832 13388
rect 13955 13348 14832 13376
rect 13955 13345 13967 13348
rect 13909 13339 13967 13345
rect 14826 13336 14832 13348
rect 14884 13336 14890 13388
rect 15396 13385 15424 13484
rect 17954 13472 17960 13484
rect 18012 13512 18018 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 18012 13484 18153 13512
rect 18012 13472 18018 13484
rect 18141 13481 18153 13484
rect 18187 13512 18199 13515
rect 18414 13512 18420 13524
rect 18187 13484 18420 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 18414 13472 18420 13484
rect 18472 13472 18478 13524
rect 20254 13472 20260 13524
rect 20312 13512 20318 13524
rect 20441 13515 20499 13521
rect 20441 13512 20453 13515
rect 20312 13484 20453 13512
rect 20312 13472 20318 13484
rect 20441 13481 20453 13484
rect 20487 13481 20499 13515
rect 20441 13475 20499 13481
rect 20898 13472 20904 13524
rect 20956 13472 20962 13524
rect 22097 13515 22155 13521
rect 22097 13481 22109 13515
rect 22143 13512 22155 13515
rect 22186 13512 22192 13524
rect 22143 13484 22192 13512
rect 22143 13481 22155 13484
rect 22097 13475 22155 13481
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 22738 13512 22744 13524
rect 22664 13484 22744 13512
rect 17862 13404 17868 13456
rect 17920 13444 17926 13456
rect 22554 13444 22560 13456
rect 17920 13416 22560 13444
rect 17920 13404 17926 13416
rect 22554 13404 22560 13416
rect 22612 13404 22618 13456
rect 15381 13379 15439 13385
rect 15381 13345 15393 13379
rect 15427 13345 15439 13379
rect 15381 13339 15439 13345
rect 15470 13336 15476 13388
rect 15528 13336 15534 13388
rect 15746 13336 15752 13388
rect 15804 13376 15810 13388
rect 16393 13379 16451 13385
rect 16393 13376 16405 13379
rect 15804 13348 16405 13376
rect 15804 13336 15810 13348
rect 16393 13345 16405 13348
rect 16439 13376 16451 13379
rect 18966 13376 18972 13388
rect 16439 13348 18972 13376
rect 16439 13345 16451 13348
rect 16393 13339 16451 13345
rect 18966 13336 18972 13348
rect 19024 13336 19030 13388
rect 19889 13379 19947 13385
rect 19889 13345 19901 13379
rect 19935 13376 19947 13379
rect 19978 13376 19984 13388
rect 19935 13348 19984 13376
rect 19935 13345 19947 13348
rect 19889 13339 19947 13345
rect 19978 13336 19984 13348
rect 20036 13336 20042 13388
rect 21358 13336 21364 13388
rect 21416 13376 21422 13388
rect 21453 13379 21511 13385
rect 21453 13376 21465 13379
rect 21416 13348 21465 13376
rect 21416 13336 21422 13348
rect 21453 13345 21465 13348
rect 21499 13376 21511 13379
rect 22664 13376 22692 13484
rect 22738 13472 22744 13484
rect 22796 13472 22802 13524
rect 23658 13472 23664 13524
rect 23716 13512 23722 13524
rect 24029 13515 24087 13521
rect 24029 13512 24041 13515
rect 23716 13484 24041 13512
rect 23716 13472 23722 13484
rect 24029 13481 24041 13484
rect 24075 13481 24087 13515
rect 24029 13475 24087 13481
rect 25590 13472 25596 13524
rect 25648 13472 25654 13524
rect 25774 13472 25780 13524
rect 25832 13512 25838 13524
rect 26697 13515 26755 13521
rect 26697 13512 26709 13515
rect 25832 13484 26709 13512
rect 25832 13472 25838 13484
rect 26697 13481 26709 13484
rect 26743 13512 26755 13515
rect 27430 13512 27436 13524
rect 26743 13484 27436 13512
rect 26743 13481 26755 13484
rect 26697 13475 26755 13481
rect 27430 13472 27436 13484
rect 27488 13472 27494 13524
rect 27798 13472 27804 13524
rect 27856 13472 27862 13524
rect 28169 13515 28227 13521
rect 28169 13481 28181 13515
rect 28215 13512 28227 13515
rect 28350 13512 28356 13524
rect 28215 13484 28356 13512
rect 28215 13481 28227 13484
rect 28169 13475 28227 13481
rect 28350 13472 28356 13484
rect 28408 13512 28414 13524
rect 28902 13512 28908 13524
rect 28408 13484 28908 13512
rect 28408 13472 28414 13484
rect 28902 13472 28908 13484
rect 28960 13472 28966 13524
rect 29181 13515 29239 13521
rect 29181 13481 29193 13515
rect 29227 13512 29239 13515
rect 33778 13512 33784 13524
rect 29227 13484 33784 13512
rect 29227 13481 29239 13484
rect 29181 13475 29239 13481
rect 33778 13472 33784 13484
rect 33836 13472 33842 13524
rect 35621 13515 35679 13521
rect 35621 13481 35633 13515
rect 35667 13512 35679 13515
rect 35710 13512 35716 13524
rect 35667 13484 35716 13512
rect 35667 13481 35679 13484
rect 35621 13475 35679 13481
rect 35710 13472 35716 13484
rect 35768 13472 35774 13524
rect 38194 13472 38200 13524
rect 38252 13472 38258 13524
rect 38565 13515 38623 13521
rect 38565 13481 38577 13515
rect 38611 13512 38623 13515
rect 38654 13512 38660 13524
rect 38611 13484 38660 13512
rect 38611 13481 38623 13484
rect 38565 13475 38623 13481
rect 38654 13472 38660 13484
rect 38712 13512 38718 13524
rect 38838 13512 38844 13524
rect 38712 13484 38844 13512
rect 38712 13472 38718 13484
rect 38838 13472 38844 13484
rect 38896 13512 38902 13524
rect 39577 13515 39635 13521
rect 39577 13512 39589 13515
rect 38896 13484 39589 13512
rect 38896 13472 38902 13484
rect 39577 13481 39589 13484
rect 39623 13481 39635 13515
rect 39577 13475 39635 13481
rect 24486 13444 24492 13456
rect 22756 13416 24492 13444
rect 22756 13385 22784 13416
rect 24486 13404 24492 13416
rect 24544 13404 24550 13456
rect 29914 13444 29920 13456
rect 28644 13416 29920 13444
rect 21499 13348 22692 13376
rect 22741 13379 22799 13385
rect 21499 13345 21511 13348
rect 21453 13339 21511 13345
rect 22741 13345 22753 13379
rect 22787 13345 22799 13379
rect 22741 13339 22799 13345
rect 22830 13336 22836 13388
rect 22888 13376 22894 13388
rect 23477 13379 23535 13385
rect 23477 13376 23489 13379
rect 22888 13348 23489 13376
rect 22888 13336 22894 13348
rect 23477 13345 23489 13348
rect 23523 13345 23535 13379
rect 23477 13339 23535 13345
rect 23569 13379 23627 13385
rect 23569 13345 23581 13379
rect 23615 13376 23627 13379
rect 24394 13376 24400 13388
rect 23615 13348 24400 13376
rect 23615 13345 23627 13348
rect 23569 13339 23627 13345
rect 24394 13336 24400 13348
rect 24452 13336 24458 13388
rect 25041 13379 25099 13385
rect 25041 13345 25053 13379
rect 25087 13376 25099 13379
rect 27062 13376 27068 13388
rect 25087 13348 27068 13376
rect 25087 13345 25099 13348
rect 25041 13339 25099 13345
rect 27062 13336 27068 13348
rect 27120 13336 27126 13388
rect 28644 13385 28672 13416
rect 29914 13404 29920 13416
rect 29972 13404 29978 13456
rect 30374 13404 30380 13456
rect 30432 13444 30438 13456
rect 31113 13447 31171 13453
rect 31113 13444 31125 13447
rect 30432 13416 31125 13444
rect 30432 13404 30438 13416
rect 31113 13413 31125 13416
rect 31159 13413 31171 13447
rect 31113 13407 31171 13413
rect 33321 13447 33379 13453
rect 33321 13413 33333 13447
rect 33367 13413 33379 13447
rect 36081 13447 36139 13453
rect 36081 13444 36093 13447
rect 33321 13407 33379 13413
rect 34440 13416 36093 13444
rect 28629 13379 28687 13385
rect 28629 13345 28641 13379
rect 28675 13345 28687 13379
rect 28629 13339 28687 13345
rect 29822 13336 29828 13388
rect 29880 13336 29886 13388
rect 30009 13379 30067 13385
rect 30009 13345 30021 13379
rect 30055 13376 30067 13379
rect 30466 13376 30472 13388
rect 30055 13348 30472 13376
rect 30055 13345 30067 13348
rect 30009 13339 30067 13345
rect 30466 13336 30472 13348
rect 30524 13336 30530 13388
rect 31386 13336 31392 13388
rect 31444 13376 31450 13388
rect 33336 13376 33364 13407
rect 31444 13348 33364 13376
rect 31444 13336 31450 13348
rect 33870 13336 33876 13388
rect 33928 13376 33934 13388
rect 34333 13379 34391 13385
rect 34333 13376 34345 13379
rect 33928 13348 34345 13376
rect 33928 13336 33934 13348
rect 34333 13345 34345 13348
rect 34379 13345 34391 13379
rect 34333 13339 34391 13345
rect 2961 13311 3019 13317
rect 2961 13277 2973 13311
rect 3007 13277 3019 13311
rect 2961 13271 3019 13277
rect 14461 13311 14519 13317
rect 14461 13277 14473 13311
rect 14507 13308 14519 13311
rect 14550 13308 14556 13320
rect 14507 13280 14556 13308
rect 14507 13277 14519 13280
rect 14461 13271 14519 13277
rect 14550 13268 14556 13280
rect 14608 13268 14614 13320
rect 18322 13268 18328 13320
rect 18380 13308 18386 13320
rect 24489 13311 24547 13317
rect 24489 13308 24501 13311
rect 18380 13280 24501 13308
rect 18380 13268 18386 13280
rect 24489 13277 24501 13280
rect 24535 13277 24547 13311
rect 24489 13271 24547 13277
rect 9030 13200 9036 13252
rect 9088 13240 9094 13252
rect 11057 13243 11115 13249
rect 11057 13240 11069 13243
rect 9088 13212 11069 13240
rect 9088 13200 9094 13212
rect 11057 13209 11069 13212
rect 11103 13209 11115 13243
rect 11057 13203 11115 13209
rect 10962 13132 10968 13184
rect 11020 13172 11026 13184
rect 11072 13172 11100 13203
rect 11146 13200 11152 13252
rect 11204 13240 11210 13252
rect 11204 13212 11546 13240
rect 11204 13200 11210 13212
rect 12986 13200 12992 13252
rect 13044 13240 13050 13252
rect 14918 13240 14924 13252
rect 13044 13212 14924 13240
rect 13044 13200 13050 13212
rect 14918 13200 14924 13212
rect 14976 13200 14982 13252
rect 16206 13240 16212 13252
rect 15120 13212 16212 13240
rect 15120 13184 15148 13212
rect 16206 13200 16212 13212
rect 16264 13200 16270 13252
rect 16298 13200 16304 13252
rect 16356 13240 16362 13252
rect 16669 13243 16727 13249
rect 16669 13240 16681 13243
rect 16356 13212 16681 13240
rect 16356 13200 16362 13212
rect 16669 13209 16681 13212
rect 16715 13209 16727 13243
rect 16669 13203 16727 13209
rect 17126 13200 17132 13252
rect 17184 13200 17190 13252
rect 18877 13243 18935 13249
rect 18877 13209 18889 13243
rect 18923 13240 18935 13243
rect 20073 13243 20131 13249
rect 20073 13240 20085 13243
rect 18923 13212 20085 13240
rect 18923 13209 18935 13212
rect 18877 13203 18935 13209
rect 20073 13209 20085 13212
rect 20119 13209 20131 13243
rect 20073 13203 20131 13209
rect 21361 13243 21419 13249
rect 21361 13209 21373 13243
rect 21407 13240 21419 13243
rect 21450 13240 21456 13252
rect 21407 13212 21456 13240
rect 21407 13209 21419 13212
rect 21361 13203 21419 13209
rect 21450 13200 21456 13212
rect 21508 13240 21514 13252
rect 21634 13240 21640 13252
rect 21508 13212 21640 13240
rect 21508 13200 21514 13212
rect 21634 13200 21640 13212
rect 21692 13200 21698 13252
rect 22465 13243 22523 13249
rect 22465 13209 22477 13243
rect 22511 13240 22523 13243
rect 22830 13240 22836 13252
rect 22511 13212 22836 13240
rect 22511 13209 22523 13212
rect 22465 13203 22523 13209
rect 22830 13200 22836 13212
rect 22888 13200 22894 13252
rect 24026 13240 24032 13252
rect 23584 13212 24032 13240
rect 13814 13172 13820 13184
rect 11020 13144 13820 13172
rect 11020 13132 11026 13144
rect 13814 13132 13820 13144
rect 13872 13132 13878 13184
rect 14090 13132 14096 13184
rect 14148 13172 14154 13184
rect 15102 13172 15108 13184
rect 14148 13144 15108 13172
rect 14148 13132 14154 13144
rect 15102 13132 15108 13144
rect 15160 13132 15166 13184
rect 15562 13132 15568 13184
rect 15620 13132 15626 13184
rect 15930 13132 15936 13184
rect 15988 13132 15994 13184
rect 16758 13132 16764 13184
rect 16816 13172 16822 13184
rect 18506 13172 18512 13184
rect 16816 13144 18512 13172
rect 16816 13132 16822 13144
rect 18506 13132 18512 13144
rect 18564 13172 18570 13184
rect 19334 13172 19340 13184
rect 18564 13144 19340 13172
rect 18564 13132 18570 13144
rect 19334 13132 19340 13144
rect 19392 13132 19398 13184
rect 19978 13132 19984 13184
rect 20036 13132 20042 13184
rect 21269 13175 21327 13181
rect 21269 13141 21281 13175
rect 21315 13172 21327 13175
rect 21542 13172 21548 13184
rect 21315 13144 21548 13172
rect 21315 13141 21327 13144
rect 21269 13135 21327 13141
rect 21542 13132 21548 13144
rect 21600 13172 21606 13184
rect 21818 13172 21824 13184
rect 21600 13144 21824 13172
rect 21600 13132 21606 13144
rect 21818 13132 21824 13144
rect 21876 13132 21882 13184
rect 22557 13175 22615 13181
rect 22557 13141 22569 13175
rect 22603 13172 22615 13175
rect 23584 13172 23612 13212
rect 24026 13200 24032 13212
rect 24084 13200 24090 13252
rect 22603 13144 23612 13172
rect 22603 13141 22615 13144
rect 22557 13135 22615 13141
rect 23658 13132 23664 13184
rect 23716 13132 23722 13184
rect 23842 13132 23848 13184
rect 23900 13172 23906 13184
rect 24394 13172 24400 13184
rect 23900 13144 24400 13172
rect 23900 13132 23906 13144
rect 24394 13132 24400 13144
rect 24452 13132 24458 13184
rect 24504 13172 24532 13271
rect 25130 13268 25136 13320
rect 25188 13308 25194 13320
rect 25225 13311 25283 13317
rect 25225 13308 25237 13311
rect 25188 13280 25237 13308
rect 25188 13268 25194 13280
rect 25225 13277 25237 13280
rect 25271 13277 25283 13311
rect 25225 13271 25283 13277
rect 28813 13311 28871 13317
rect 28813 13277 28825 13311
rect 28859 13308 28871 13311
rect 28994 13308 29000 13320
rect 28859 13280 29000 13308
rect 28859 13277 28871 13280
rect 28813 13271 28871 13277
rect 28994 13268 29000 13280
rect 29052 13268 29058 13320
rect 30101 13311 30159 13317
rect 30101 13277 30113 13311
rect 30147 13308 30159 13311
rect 30190 13308 30196 13320
rect 30147 13280 30196 13308
rect 30147 13277 30159 13280
rect 30101 13271 30159 13277
rect 30190 13268 30196 13280
rect 30248 13268 30254 13320
rect 31202 13268 31208 13320
rect 31260 13308 31266 13320
rect 32861 13311 32919 13317
rect 31260 13280 31510 13308
rect 31260 13268 31266 13280
rect 32861 13277 32873 13311
rect 32907 13308 32919 13311
rect 34054 13308 34060 13320
rect 32907 13280 34060 13308
rect 32907 13277 32919 13280
rect 32861 13271 32919 13277
rect 34054 13268 34060 13280
rect 34112 13268 34118 13320
rect 24854 13200 24860 13252
rect 24912 13240 24918 13252
rect 25774 13240 25780 13252
rect 24912 13212 25780 13240
rect 24912 13200 24918 13212
rect 25774 13200 25780 13212
rect 25832 13200 25838 13252
rect 26050 13200 26056 13252
rect 26108 13200 26114 13252
rect 27709 13243 27767 13249
rect 27709 13209 27721 13243
rect 27755 13240 27767 13243
rect 28626 13240 28632 13252
rect 27755 13212 28632 13240
rect 27755 13209 27767 13212
rect 27709 13203 27767 13209
rect 28626 13200 28632 13212
rect 28684 13200 28690 13252
rect 32585 13243 32643 13249
rect 30484 13212 31340 13240
rect 25133 13175 25191 13181
rect 25133 13172 25145 13175
rect 24504 13144 25145 13172
rect 25133 13141 25145 13144
rect 25179 13172 25191 13175
rect 26510 13172 26516 13184
rect 25179 13144 26516 13172
rect 25179 13141 25191 13144
rect 25133 13135 25191 13141
rect 26510 13132 26516 13144
rect 26568 13132 26574 13184
rect 28718 13132 28724 13184
rect 28776 13132 28782 13184
rect 30484 13181 30512 13212
rect 30469 13175 30527 13181
rect 30469 13141 30481 13175
rect 30515 13141 30527 13175
rect 31312 13172 31340 13212
rect 32585 13209 32597 13243
rect 32631 13240 32643 13243
rect 33594 13240 33600 13252
rect 32631 13212 33600 13240
rect 32631 13209 32643 13212
rect 32585 13203 32643 13209
rect 33594 13200 33600 13212
rect 33652 13200 33658 13252
rect 33686 13200 33692 13252
rect 33744 13240 33750 13252
rect 34440 13240 34468 13416
rect 36081 13413 36093 13416
rect 36127 13413 36139 13447
rect 36081 13407 36139 13413
rect 35069 13379 35127 13385
rect 35069 13345 35081 13379
rect 35115 13376 35127 13379
rect 39206 13376 39212 13388
rect 35115 13348 39212 13376
rect 35115 13345 35127 13348
rect 35069 13339 35127 13345
rect 39206 13336 39212 13348
rect 39264 13336 39270 13388
rect 34882 13268 34888 13320
rect 34940 13308 34946 13320
rect 36449 13311 36507 13317
rect 36449 13308 36461 13311
rect 34940 13280 36461 13308
rect 34940 13268 34946 13280
rect 36449 13277 36461 13280
rect 36495 13277 36507 13311
rect 36449 13271 36507 13277
rect 33744 13212 34468 13240
rect 33744 13200 33750 13212
rect 35158 13200 35164 13252
rect 35216 13200 35222 13252
rect 35253 13243 35311 13249
rect 35253 13209 35265 13243
rect 35299 13240 35311 13243
rect 36354 13240 36360 13252
rect 35299 13212 36360 13240
rect 35299 13209 35311 13212
rect 35253 13203 35311 13209
rect 36354 13200 36360 13212
rect 36412 13200 36418 13252
rect 31662 13172 31668 13184
rect 31312 13144 31668 13172
rect 30469 13135 30527 13141
rect 31662 13132 31668 13144
rect 31720 13132 31726 13184
rect 33781 13175 33839 13181
rect 33781 13141 33793 13175
rect 33827 13172 33839 13175
rect 34422 13172 34428 13184
rect 33827 13144 34428 13172
rect 33827 13141 33839 13144
rect 33781 13135 33839 13141
rect 34422 13132 34428 13144
rect 34480 13132 34486 13184
rect 35618 13132 35624 13184
rect 35676 13172 35682 13184
rect 35897 13175 35955 13181
rect 35897 13172 35909 13175
rect 35676 13144 35909 13172
rect 35676 13132 35682 13144
rect 35897 13141 35909 13144
rect 35943 13141 35955 13175
rect 36464 13172 36492 13271
rect 41322 13268 41328 13320
rect 41380 13268 41386 13320
rect 46290 13268 46296 13320
rect 46348 13308 46354 13320
rect 47949 13311 48007 13317
rect 47949 13308 47961 13311
rect 46348 13280 47961 13308
rect 46348 13268 46354 13280
rect 47949 13277 47961 13280
rect 47995 13277 48007 13311
rect 47949 13271 48007 13277
rect 49142 13268 49148 13320
rect 49200 13268 49206 13320
rect 36630 13200 36636 13252
rect 36688 13240 36694 13252
rect 36725 13243 36783 13249
rect 36725 13240 36737 13243
rect 36688 13212 36737 13240
rect 36688 13200 36694 13212
rect 36725 13209 36737 13212
rect 36771 13209 36783 13243
rect 38838 13240 38844 13252
rect 37950 13212 38844 13240
rect 36725 13203 36783 13209
rect 38838 13200 38844 13212
rect 38896 13200 38902 13252
rect 37458 13172 37464 13184
rect 36464 13144 37464 13172
rect 35897 13135 35955 13141
rect 37458 13132 37464 13144
rect 37516 13132 37522 13184
rect 37642 13132 37648 13184
rect 37700 13172 37706 13184
rect 39574 13172 39580 13184
rect 37700 13144 39580 13172
rect 37700 13132 37706 13144
rect 39574 13132 39580 13144
rect 39632 13132 39638 13184
rect 41509 13175 41567 13181
rect 41509 13141 41521 13175
rect 41555 13172 41567 13175
rect 45922 13172 45928 13184
rect 41555 13144 45928 13172
rect 41555 13141 41567 13144
rect 41509 13135 41567 13141
rect 45922 13132 45928 13144
rect 45980 13132 45986 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 3053 12971 3111 12977
rect 3053 12937 3065 12971
rect 3099 12968 3111 12971
rect 5442 12968 5448 12980
rect 3099 12940 5448 12968
rect 3099 12937 3111 12940
rect 3053 12931 3111 12937
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 10962 12928 10968 12980
rect 11020 12928 11026 12980
rect 11146 12928 11152 12980
rect 11204 12928 11210 12980
rect 11330 12928 11336 12980
rect 11388 12968 11394 12980
rect 11977 12971 12035 12977
rect 11977 12968 11989 12971
rect 11388 12940 11989 12968
rect 11388 12928 11394 12940
rect 11977 12937 11989 12940
rect 12023 12937 12035 12971
rect 11977 12931 12035 12937
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12713 12971 12771 12977
rect 12713 12968 12725 12971
rect 12492 12940 12725 12968
rect 12492 12928 12498 12940
rect 12713 12937 12725 12940
rect 12759 12937 12771 12971
rect 12713 12931 12771 12937
rect 13081 12971 13139 12977
rect 13081 12937 13093 12971
rect 13127 12968 13139 12971
rect 13262 12968 13268 12980
rect 13127 12940 13268 12968
rect 13127 12937 13139 12940
rect 13081 12931 13139 12937
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 13630 12928 13636 12980
rect 13688 12968 13694 12980
rect 13688 12940 14872 12968
rect 13688 12928 13694 12940
rect 1302 12860 1308 12912
rect 1360 12900 1366 12912
rect 1673 12903 1731 12909
rect 1673 12900 1685 12903
rect 1360 12872 1685 12900
rect 1360 12860 1366 12872
rect 1673 12869 1685 12872
rect 1719 12900 1731 12903
rect 2133 12903 2191 12909
rect 2133 12900 2145 12903
rect 1719 12872 2145 12900
rect 1719 12869 1731 12872
rect 1673 12863 1731 12869
rect 2133 12869 2145 12872
rect 2179 12869 2191 12903
rect 14458 12900 14464 12912
rect 14122 12872 14464 12900
rect 2133 12863 2191 12869
rect 14458 12860 14464 12872
rect 14516 12860 14522 12912
rect 1210 12792 1216 12844
rect 1268 12832 1274 12844
rect 2869 12835 2927 12841
rect 2869 12832 2881 12835
rect 1268 12804 2881 12832
rect 1268 12792 1274 12804
rect 2869 12801 2881 12804
rect 2915 12832 2927 12835
rect 3329 12835 3387 12841
rect 3329 12832 3341 12835
rect 2915 12804 3341 12832
rect 2915 12801 2927 12804
rect 2869 12795 2927 12801
rect 3329 12801 3341 12804
rect 3375 12801 3387 12835
rect 3329 12795 3387 12801
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12832 12127 12835
rect 12115 12804 12434 12832
rect 12115 12801 12127 12804
rect 12069 12795 12127 12801
rect 1857 12767 1915 12773
rect 1857 12733 1869 12767
rect 1903 12764 1915 12767
rect 9490 12764 9496 12776
rect 1903 12736 9496 12764
rect 1903 12733 1915 12736
rect 1857 12727 1915 12733
rect 9490 12724 9496 12736
rect 9548 12724 9554 12776
rect 11790 12724 11796 12776
rect 11848 12724 11854 12776
rect 12406 12764 12434 12804
rect 13906 12764 13912 12776
rect 12406 12736 13912 12764
rect 13906 12724 13912 12736
rect 13964 12724 13970 12776
rect 14550 12724 14556 12776
rect 14608 12724 14614 12776
rect 14844 12773 14872 12940
rect 15286 12928 15292 12980
rect 15344 12928 15350 12980
rect 15841 12971 15899 12977
rect 15841 12937 15853 12971
rect 15887 12968 15899 12971
rect 18322 12968 18328 12980
rect 15887 12940 18328 12968
rect 15887 12937 15899 12940
rect 15841 12931 15899 12937
rect 15856 12832 15884 12931
rect 18322 12928 18328 12940
rect 18380 12928 18386 12980
rect 19058 12928 19064 12980
rect 19116 12968 19122 12980
rect 19245 12971 19303 12977
rect 19245 12968 19257 12971
rect 19116 12940 19257 12968
rect 19116 12928 19122 12940
rect 19245 12937 19257 12940
rect 19291 12937 19303 12971
rect 19245 12931 19303 12937
rect 22922 12928 22928 12980
rect 22980 12928 22986 12980
rect 23382 12928 23388 12980
rect 23440 12928 23446 12980
rect 24302 12928 24308 12980
rect 24360 12968 24366 12980
rect 24578 12968 24584 12980
rect 24360 12940 24584 12968
rect 24360 12928 24366 12940
rect 24578 12928 24584 12940
rect 24636 12968 24642 12980
rect 24636 12940 25636 12968
rect 24636 12928 24642 12940
rect 15933 12903 15991 12909
rect 15933 12869 15945 12903
rect 15979 12900 15991 12903
rect 16390 12900 16396 12912
rect 15979 12872 16396 12900
rect 15979 12869 15991 12872
rect 15933 12863 15991 12869
rect 16390 12860 16396 12872
rect 16448 12860 16454 12912
rect 18693 12903 18751 12909
rect 18693 12869 18705 12903
rect 18739 12900 18751 12903
rect 18966 12900 18972 12912
rect 18739 12872 18972 12900
rect 18739 12869 18751 12872
rect 18693 12863 18751 12869
rect 18966 12860 18972 12872
rect 19024 12860 19030 12912
rect 19886 12900 19892 12912
rect 19306 12872 19892 12900
rect 15672 12804 15884 12832
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12764 14887 12767
rect 15470 12764 15476 12776
rect 14875 12736 15476 12764
rect 14875 12733 14887 12736
rect 14829 12727 14887 12733
rect 15470 12724 15476 12736
rect 15528 12724 15534 12776
rect 15672 12696 15700 12804
rect 16298 12792 16304 12844
rect 16356 12792 16362 12844
rect 16850 12792 16856 12844
rect 16908 12832 16914 12844
rect 17770 12832 17776 12844
rect 16908 12804 17776 12832
rect 16908 12792 16914 12804
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 17865 12835 17923 12841
rect 17865 12801 17877 12835
rect 17911 12832 17923 12835
rect 18598 12832 18604 12844
rect 17911 12804 18604 12832
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 18598 12792 18604 12804
rect 18656 12832 18662 12844
rect 19058 12832 19064 12844
rect 18656 12804 19064 12832
rect 18656 12792 18662 12804
rect 19058 12792 19064 12804
rect 19116 12792 19122 12844
rect 15749 12767 15807 12773
rect 15749 12733 15761 12767
rect 15795 12764 15807 12767
rect 16316 12764 16344 12792
rect 15795 12736 16344 12764
rect 17405 12767 17463 12773
rect 15795 12733 15807 12736
rect 15749 12727 15807 12733
rect 17405 12733 17417 12767
rect 17451 12764 17463 12767
rect 19306 12764 19334 12872
rect 19886 12860 19892 12872
rect 19944 12860 19950 12912
rect 24854 12860 24860 12912
rect 24912 12860 24918 12912
rect 25314 12860 25320 12912
rect 25372 12860 25378 12912
rect 19518 12792 19524 12844
rect 19576 12832 19582 12844
rect 19613 12835 19671 12841
rect 19613 12832 19625 12835
rect 19576 12804 19625 12832
rect 19576 12792 19582 12804
rect 19613 12801 19625 12804
rect 19659 12801 19671 12835
rect 19613 12795 19671 12801
rect 21085 12835 21143 12841
rect 21085 12801 21097 12835
rect 21131 12832 21143 12835
rect 21910 12832 21916 12844
rect 21131 12804 21916 12832
rect 21131 12801 21143 12804
rect 21085 12795 21143 12801
rect 21910 12792 21916 12804
rect 21968 12792 21974 12844
rect 22186 12792 22192 12844
rect 22244 12832 22250 12844
rect 23014 12832 23020 12844
rect 22244 12804 23020 12832
rect 22244 12792 22250 12804
rect 23014 12792 23020 12804
rect 23072 12792 23078 12844
rect 25608 12841 25636 12940
rect 25774 12928 25780 12980
rect 25832 12968 25838 12980
rect 26053 12971 26111 12977
rect 26053 12968 26065 12971
rect 25832 12940 26065 12968
rect 25832 12928 25838 12940
rect 26053 12937 26065 12940
rect 26099 12937 26111 12971
rect 26053 12931 26111 12937
rect 26234 12928 26240 12980
rect 26292 12928 26298 12980
rect 26510 12928 26516 12980
rect 26568 12968 26574 12980
rect 26697 12971 26755 12977
rect 26697 12968 26709 12971
rect 26568 12940 26709 12968
rect 26568 12928 26574 12940
rect 26697 12937 26709 12940
rect 26743 12937 26755 12971
rect 26697 12931 26755 12937
rect 27890 12928 27896 12980
rect 27948 12968 27954 12980
rect 31757 12971 31815 12977
rect 27948 12940 31616 12968
rect 27948 12928 27954 12940
rect 27430 12860 27436 12912
rect 27488 12900 27494 12912
rect 27488 12872 27738 12900
rect 27488 12860 27494 12872
rect 29638 12860 29644 12912
rect 29696 12860 29702 12912
rect 30190 12860 30196 12912
rect 30248 12900 30254 12912
rect 30285 12903 30343 12909
rect 30285 12900 30297 12903
rect 30248 12872 30297 12900
rect 30248 12860 30254 12872
rect 30285 12869 30297 12872
rect 30331 12869 30343 12903
rect 30285 12863 30343 12869
rect 31294 12860 31300 12912
rect 31352 12860 31358 12912
rect 31588 12900 31616 12940
rect 31757 12937 31769 12971
rect 31803 12968 31815 12971
rect 31846 12968 31852 12980
rect 31803 12940 31852 12968
rect 31803 12937 31815 12940
rect 31757 12931 31815 12937
rect 31846 12928 31852 12940
rect 31904 12968 31910 12980
rect 32398 12968 32404 12980
rect 31904 12940 32404 12968
rect 31904 12928 31910 12940
rect 32398 12928 32404 12940
rect 32456 12928 32462 12980
rect 33413 12971 33471 12977
rect 33413 12937 33425 12971
rect 33459 12968 33471 12971
rect 33502 12968 33508 12980
rect 33459 12940 33508 12968
rect 33459 12937 33471 12940
rect 33413 12931 33471 12937
rect 33502 12928 33508 12940
rect 33560 12968 33566 12980
rect 33686 12968 33692 12980
rect 33560 12940 33692 12968
rect 33560 12928 33566 12940
rect 33686 12928 33692 12940
rect 33744 12928 33750 12980
rect 34054 12928 34060 12980
rect 34112 12968 34118 12980
rect 34112 12940 34836 12968
rect 34112 12928 34118 12940
rect 32677 12903 32735 12909
rect 32677 12900 32689 12903
rect 31588 12872 32689 12900
rect 32677 12869 32689 12872
rect 32723 12869 32735 12903
rect 33870 12900 33876 12912
rect 32677 12863 32735 12869
rect 32968 12872 33876 12900
rect 25593 12835 25651 12841
rect 25593 12801 25605 12835
rect 25639 12801 25651 12835
rect 25593 12795 25651 12801
rect 26418 12792 26424 12844
rect 26476 12832 26482 12844
rect 27154 12832 27160 12844
rect 26476 12804 27160 12832
rect 26476 12792 26482 12804
rect 27154 12792 27160 12804
rect 27212 12792 27218 12844
rect 29181 12835 29239 12841
rect 29181 12801 29193 12835
rect 29227 12832 29239 12835
rect 30006 12832 30012 12844
rect 29227 12804 30012 12832
rect 29227 12801 29239 12804
rect 29181 12795 29239 12801
rect 30006 12792 30012 12804
rect 30064 12792 30070 12844
rect 17451 12736 19334 12764
rect 17451 12733 17463 12736
rect 17405 12727 17463 12733
rect 19702 12724 19708 12776
rect 19760 12724 19766 12776
rect 19889 12767 19947 12773
rect 19889 12733 19901 12767
rect 19935 12764 19947 12767
rect 20254 12764 20260 12776
rect 19935 12736 20260 12764
rect 19935 12733 19947 12736
rect 19889 12727 19947 12733
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 21177 12767 21235 12773
rect 21177 12733 21189 12767
rect 21223 12733 21235 12767
rect 21177 12727 21235 12733
rect 11256 12668 13584 12696
rect 11256 12640 11284 12668
rect 11238 12588 11244 12640
rect 11296 12588 11302 12640
rect 12437 12631 12495 12637
rect 12437 12597 12449 12631
rect 12483 12628 12495 12631
rect 12526 12628 12532 12640
rect 12483 12600 12532 12628
rect 12483 12597 12495 12600
rect 12437 12591 12495 12597
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 13556 12628 13584 12668
rect 14752 12668 15700 12696
rect 16301 12699 16359 12705
rect 14752 12628 14780 12668
rect 16301 12665 16313 12699
rect 16347 12696 16359 12699
rect 17310 12696 17316 12708
rect 16347 12668 17316 12696
rect 16347 12665 16359 12668
rect 16301 12659 16359 12665
rect 17310 12656 17316 12668
rect 17368 12656 17374 12708
rect 17770 12656 17776 12708
rect 17828 12696 17834 12708
rect 20717 12699 20775 12705
rect 20717 12696 20729 12699
rect 17828 12668 20729 12696
rect 17828 12656 17834 12668
rect 20717 12665 20729 12668
rect 20763 12665 20775 12699
rect 21192 12696 21220 12727
rect 21266 12724 21272 12776
rect 21324 12724 21330 12776
rect 21726 12724 21732 12776
rect 21784 12764 21790 12776
rect 22005 12767 22063 12773
rect 22005 12764 22017 12767
rect 21784 12736 22017 12764
rect 21784 12724 21790 12736
rect 22005 12733 22017 12736
rect 22051 12733 22063 12767
rect 22005 12727 22063 12733
rect 22738 12724 22744 12776
rect 22796 12724 22802 12776
rect 23566 12724 23572 12776
rect 23624 12764 23630 12776
rect 23845 12767 23903 12773
rect 23845 12764 23857 12767
rect 23624 12736 23857 12764
rect 23624 12724 23630 12736
rect 23845 12733 23857 12736
rect 23891 12764 23903 12767
rect 24946 12764 24952 12776
rect 23891 12736 24952 12764
rect 23891 12733 23903 12736
rect 23845 12727 23903 12733
rect 24946 12724 24952 12736
rect 25004 12724 25010 12776
rect 28902 12724 28908 12776
rect 28960 12764 28966 12776
rect 32401 12767 32459 12773
rect 28960 12736 31340 12764
rect 28960 12724 28966 12736
rect 31312 12696 31340 12736
rect 32401 12733 32413 12767
rect 32447 12733 32459 12767
rect 32401 12727 32459 12733
rect 32585 12767 32643 12773
rect 32585 12733 32597 12767
rect 32631 12764 32643 12767
rect 32674 12764 32680 12776
rect 32631 12736 32680 12764
rect 32631 12733 32643 12736
rect 32585 12727 32643 12733
rect 32416 12696 32444 12727
rect 32674 12724 32680 12736
rect 32732 12724 32738 12776
rect 21192 12668 23980 12696
rect 31312 12668 32444 12696
rect 20717 12659 20775 12665
rect 13556 12600 14780 12628
rect 16758 12588 16764 12640
rect 16816 12588 16822 12640
rect 16850 12588 16856 12640
rect 16908 12628 16914 12640
rect 17126 12628 17132 12640
rect 16908 12600 17132 12628
rect 16908 12588 16914 12600
rect 17126 12588 17132 12600
rect 17184 12588 17190 12640
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 20441 12631 20499 12637
rect 20441 12628 20453 12631
rect 19392 12600 20453 12628
rect 19392 12588 19398 12600
rect 20441 12597 20453 12600
rect 20487 12628 20499 12631
rect 21174 12628 21180 12640
rect 20487 12600 21180 12628
rect 20487 12597 20499 12600
rect 20441 12591 20499 12597
rect 21174 12588 21180 12600
rect 21232 12628 21238 12640
rect 23842 12628 23848 12640
rect 21232 12600 23848 12628
rect 21232 12588 21238 12600
rect 23842 12588 23848 12600
rect 23900 12588 23906 12640
rect 23952 12628 23980 12668
rect 25682 12628 25688 12640
rect 23952 12600 25688 12628
rect 25682 12588 25688 12600
rect 25740 12588 25746 12640
rect 25958 12588 25964 12640
rect 26016 12588 26022 12640
rect 27798 12588 27804 12640
rect 27856 12628 27862 12640
rect 32968 12628 32996 12872
rect 33870 12860 33876 12872
rect 33928 12860 33934 12912
rect 34808 12909 34836 12940
rect 35158 12928 35164 12980
rect 35216 12968 35222 12980
rect 36449 12971 36507 12977
rect 36449 12968 36461 12971
rect 35216 12940 36461 12968
rect 35216 12928 35222 12940
rect 36449 12937 36461 12940
rect 36495 12968 36507 12971
rect 40310 12968 40316 12980
rect 36495 12940 40316 12968
rect 36495 12937 36507 12940
rect 36449 12931 36507 12937
rect 40310 12928 40316 12940
rect 40368 12928 40374 12980
rect 34793 12903 34851 12909
rect 34793 12869 34805 12903
rect 34839 12900 34851 12903
rect 34882 12900 34888 12912
rect 34839 12872 34888 12900
rect 34839 12869 34851 12872
rect 34793 12863 34851 12869
rect 34882 12860 34888 12872
rect 34940 12860 34946 12912
rect 35713 12903 35771 12909
rect 35713 12869 35725 12903
rect 35759 12900 35771 12903
rect 36998 12900 37004 12912
rect 35759 12872 37004 12900
rect 35759 12869 35771 12872
rect 35713 12863 35771 12869
rect 34054 12792 34060 12844
rect 34112 12792 34118 12844
rect 34330 12792 34336 12844
rect 34388 12832 34394 12844
rect 35728 12832 35756 12863
rect 36998 12860 37004 12872
rect 37056 12900 37062 12912
rect 37093 12903 37151 12909
rect 37093 12900 37105 12903
rect 37056 12872 37105 12900
rect 37056 12860 37062 12872
rect 37093 12869 37105 12872
rect 37139 12900 37151 12903
rect 37182 12900 37188 12912
rect 37139 12872 37188 12900
rect 37139 12869 37151 12872
rect 37093 12863 37151 12869
rect 37182 12860 37188 12872
rect 37240 12860 37246 12912
rect 37642 12900 37648 12912
rect 37292 12872 37648 12900
rect 34388 12804 35756 12832
rect 35805 12835 35863 12841
rect 34388 12792 34394 12804
rect 35805 12801 35817 12835
rect 35851 12832 35863 12835
rect 36725 12835 36783 12841
rect 36725 12832 36737 12835
rect 35851 12804 36737 12832
rect 35851 12801 35863 12804
rect 35805 12795 35863 12801
rect 36725 12801 36737 12804
rect 36771 12832 36783 12835
rect 37292 12832 37320 12872
rect 37642 12860 37648 12872
rect 37700 12860 37706 12912
rect 36771 12804 37320 12832
rect 36771 12801 36783 12804
rect 36725 12795 36783 12801
rect 33226 12724 33232 12776
rect 33284 12764 33290 12776
rect 33284 12736 34928 12764
rect 33284 12724 33290 12736
rect 33045 12699 33103 12705
rect 33045 12665 33057 12699
rect 33091 12696 33103 12699
rect 34790 12696 34796 12708
rect 33091 12668 34796 12696
rect 33091 12665 33103 12668
rect 33045 12659 33103 12665
rect 34790 12656 34796 12668
rect 34848 12656 34854 12708
rect 34900 12696 34928 12736
rect 35250 12724 35256 12776
rect 35308 12764 35314 12776
rect 35618 12764 35624 12776
rect 35308 12736 35624 12764
rect 35308 12724 35314 12736
rect 35618 12724 35624 12736
rect 35676 12724 35682 12776
rect 35820 12696 35848 12795
rect 37458 12792 37464 12844
rect 37516 12792 37522 12844
rect 38838 12792 38844 12844
rect 38896 12792 38902 12844
rect 40034 12792 40040 12844
rect 40092 12832 40098 12844
rect 40497 12835 40555 12841
rect 40497 12832 40509 12835
rect 40092 12804 40509 12832
rect 40092 12792 40098 12804
rect 40497 12801 40509 12804
rect 40543 12801 40555 12835
rect 40497 12795 40555 12801
rect 45922 12792 45928 12844
rect 45980 12792 45986 12844
rect 47026 12792 47032 12844
rect 47084 12832 47090 12844
rect 47949 12835 48007 12841
rect 47949 12832 47961 12835
rect 47084 12804 47961 12832
rect 47084 12792 47090 12804
rect 47949 12801 47961 12804
rect 47995 12801 48007 12835
rect 47949 12795 48007 12801
rect 49142 12792 49148 12844
rect 49200 12792 49206 12844
rect 37737 12767 37795 12773
rect 37737 12733 37749 12767
rect 37783 12764 37795 12767
rect 38286 12764 38292 12776
rect 37783 12736 38292 12764
rect 37783 12733 37795 12736
rect 37737 12727 37795 12733
rect 38286 12724 38292 12736
rect 38344 12724 38350 12776
rect 39298 12724 39304 12776
rect 39356 12764 39362 12776
rect 39485 12767 39543 12773
rect 39485 12764 39497 12767
rect 39356 12736 39497 12764
rect 39356 12724 39362 12736
rect 39485 12733 39497 12736
rect 39531 12733 39543 12767
rect 39485 12727 39543 12733
rect 34900 12668 35848 12696
rect 36173 12699 36231 12705
rect 36173 12665 36185 12699
rect 36219 12696 36231 12699
rect 37274 12696 37280 12708
rect 36219 12668 37280 12696
rect 36219 12665 36231 12668
rect 36173 12659 36231 12665
rect 37274 12656 37280 12668
rect 37332 12656 37338 12708
rect 40221 12699 40279 12705
rect 40221 12665 40233 12699
rect 40267 12696 40279 12699
rect 42702 12696 42708 12708
rect 40267 12668 42708 12696
rect 40267 12665 40279 12668
rect 40221 12659 40279 12665
rect 42702 12656 42708 12668
rect 42760 12656 42766 12708
rect 27856 12600 32996 12628
rect 27856 12588 27862 12600
rect 33318 12588 33324 12640
rect 33376 12628 33382 12640
rect 33505 12631 33563 12637
rect 33505 12628 33517 12631
rect 33376 12600 33517 12628
rect 33376 12588 33382 12600
rect 33505 12597 33517 12600
rect 33551 12628 33563 12631
rect 33689 12631 33747 12637
rect 33689 12628 33701 12631
rect 33551 12600 33701 12628
rect 33551 12597 33563 12600
rect 33505 12591 33563 12597
rect 33689 12597 33701 12600
rect 33735 12597 33747 12631
rect 33689 12591 33747 12597
rect 35618 12588 35624 12640
rect 35676 12628 35682 12640
rect 36909 12631 36967 12637
rect 36909 12628 36921 12631
rect 35676 12600 36921 12628
rect 35676 12588 35682 12600
rect 36909 12597 36921 12600
rect 36955 12628 36967 12631
rect 39298 12628 39304 12640
rect 36955 12600 39304 12628
rect 36955 12597 36967 12600
rect 36909 12591 36967 12597
rect 39298 12588 39304 12600
rect 39356 12588 39362 12640
rect 46109 12631 46167 12637
rect 46109 12597 46121 12631
rect 46155 12628 46167 12631
rect 47946 12628 47952 12640
rect 46155 12600 47952 12628
rect 46155 12597 46167 12600
rect 46109 12591 46167 12597
rect 47946 12588 47952 12600
rect 48004 12588 48010 12640
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 11241 12427 11299 12433
rect 11241 12393 11253 12427
rect 11287 12424 11299 12427
rect 11790 12424 11796 12436
rect 11287 12396 11796 12424
rect 11287 12393 11299 12396
rect 11241 12387 11299 12393
rect 11790 12384 11796 12396
rect 11848 12384 11854 12436
rect 14090 12384 14096 12436
rect 14148 12424 14154 12436
rect 14369 12427 14427 12433
rect 14369 12424 14381 12427
rect 14148 12396 14381 12424
rect 14148 12384 14154 12396
rect 14369 12393 14381 12396
rect 14415 12393 14427 12427
rect 14369 12387 14427 12393
rect 14550 12384 14556 12436
rect 14608 12384 14614 12436
rect 15286 12384 15292 12436
rect 15344 12424 15350 12436
rect 16022 12424 16028 12436
rect 15344 12396 16028 12424
rect 15344 12384 15350 12396
rect 16022 12384 16028 12396
rect 16080 12384 16086 12436
rect 16298 12384 16304 12436
rect 16356 12424 16362 12436
rect 16393 12427 16451 12433
rect 16393 12424 16405 12427
rect 16356 12396 16405 12424
rect 16356 12384 16362 12396
rect 16393 12393 16405 12396
rect 16439 12393 16451 12427
rect 21637 12427 21695 12433
rect 16393 12387 16451 12393
rect 17144 12396 21404 12424
rect 13814 12316 13820 12368
rect 13872 12356 13878 12368
rect 14568 12356 14596 12384
rect 13872 12328 14596 12356
rect 13872 12316 13878 12328
rect 14734 12316 14740 12368
rect 14792 12316 14798 12368
rect 1302 12248 1308 12300
rect 1360 12288 1366 12300
rect 2409 12291 2467 12297
rect 2409 12288 2421 12291
rect 1360 12260 2421 12288
rect 1360 12248 1366 12260
rect 2409 12257 2421 12260
rect 2455 12288 2467 12291
rect 2685 12291 2743 12297
rect 2685 12288 2697 12291
rect 2455 12260 2697 12288
rect 2455 12257 2467 12260
rect 2409 12251 2467 12257
rect 2685 12257 2697 12260
rect 2731 12257 2743 12291
rect 2685 12251 2743 12257
rect 9493 12291 9551 12297
rect 9493 12257 9505 12291
rect 9539 12288 9551 12291
rect 10778 12288 10784 12300
rect 9539 12260 10784 12288
rect 9539 12257 9551 12260
rect 9493 12251 9551 12257
rect 10778 12248 10784 12260
rect 10836 12288 10842 12300
rect 11701 12291 11759 12297
rect 11701 12288 11713 12291
rect 10836 12260 11713 12288
rect 10836 12248 10842 12260
rect 11701 12257 11713 12260
rect 11747 12257 11759 12291
rect 11701 12251 11759 12257
rect 13725 12291 13783 12297
rect 13725 12257 13737 12291
rect 13771 12288 13783 12291
rect 14752 12288 14780 12316
rect 13771 12260 14780 12288
rect 13771 12257 13783 12260
rect 13725 12251 13783 12257
rect 15470 12248 15476 12300
rect 15528 12288 15534 12300
rect 15746 12288 15752 12300
rect 15528 12260 15752 12288
rect 15528 12248 15534 12260
rect 15746 12248 15752 12260
rect 15804 12288 15810 12300
rect 16117 12291 16175 12297
rect 16117 12288 16129 12291
rect 15804 12260 16129 12288
rect 15804 12248 15810 12260
rect 16117 12257 16129 12260
rect 16163 12257 16175 12291
rect 16117 12251 16175 12257
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 5902 12220 5908 12232
rect 2179 12192 5908 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 5902 12180 5908 12192
rect 5960 12180 5966 12232
rect 16408 12220 16436 12387
rect 17144 12229 17172 12396
rect 21376 12356 21404 12396
rect 21637 12393 21649 12427
rect 21683 12424 21695 12427
rect 21683 12396 22508 12424
rect 21683 12393 21695 12396
rect 21637 12387 21695 12393
rect 22094 12356 22100 12368
rect 21008 12328 21312 12356
rect 21376 12328 22100 12356
rect 17402 12248 17408 12300
rect 17460 12248 17466 12300
rect 19886 12248 19892 12300
rect 19944 12288 19950 12300
rect 21008 12297 21036 12328
rect 19981 12291 20039 12297
rect 19981 12288 19993 12291
rect 19944 12260 19993 12288
rect 19944 12248 19950 12260
rect 19981 12257 19993 12260
rect 20027 12257 20039 12291
rect 19981 12251 20039 12257
rect 20625 12291 20683 12297
rect 20625 12257 20637 12291
rect 20671 12288 20683 12291
rect 20993 12291 21051 12297
rect 20993 12288 21005 12291
rect 20671 12260 21005 12288
rect 20671 12257 20683 12260
rect 20625 12251 20683 12257
rect 20993 12257 21005 12260
rect 21039 12257 21051 12291
rect 20993 12251 21051 12257
rect 21174 12248 21180 12300
rect 21232 12248 21238 12300
rect 21284 12288 21312 12328
rect 22094 12316 22100 12328
rect 22152 12316 22158 12368
rect 22480 12356 22508 12396
rect 22554 12384 22560 12436
rect 22612 12424 22618 12436
rect 23293 12427 23351 12433
rect 23293 12424 23305 12427
rect 22612 12396 23305 12424
rect 22612 12384 22618 12396
rect 23293 12393 23305 12396
rect 23339 12393 23351 12427
rect 26694 12424 26700 12436
rect 23293 12387 23351 12393
rect 23860 12396 26700 12424
rect 23474 12356 23480 12368
rect 22480 12328 23480 12356
rect 23474 12316 23480 12328
rect 23532 12316 23538 12368
rect 21284 12260 22232 12288
rect 17129 12223 17187 12229
rect 17129 12220 17141 12223
rect 16408 12192 17141 12220
rect 17129 12189 17141 12192
rect 17175 12189 17187 12223
rect 17129 12183 17187 12189
rect 18064 12192 19012 12220
rect 9766 12112 9772 12164
rect 9824 12112 9830 12164
rect 10502 12112 10508 12164
rect 10560 12112 10566 12164
rect 11054 12112 11060 12164
rect 11112 12152 11118 12164
rect 11977 12155 12035 12161
rect 11977 12152 11989 12155
rect 11112 12124 11989 12152
rect 11112 12112 11118 12124
rect 11977 12121 11989 12124
rect 12023 12121 12035 12155
rect 13630 12152 13636 12164
rect 13202 12124 13636 12152
rect 11977 12115 12035 12121
rect 13630 12112 13636 12124
rect 13688 12152 13694 12164
rect 14458 12152 14464 12164
rect 13688 12124 14464 12152
rect 13688 12112 13694 12124
rect 14458 12112 14464 12124
rect 14516 12152 14522 12164
rect 14516 12124 14674 12152
rect 14516 12112 14522 12124
rect 15838 12112 15844 12164
rect 15896 12112 15902 12164
rect 16316 12124 17356 12152
rect 9784 12084 9812 12112
rect 12250 12084 12256 12096
rect 9784 12056 12256 12084
rect 12250 12044 12256 12056
rect 12308 12044 12314 12096
rect 13446 12044 13452 12096
rect 13504 12084 13510 12096
rect 16316 12084 16344 12124
rect 13504 12056 16344 12084
rect 13504 12044 13510 12056
rect 16758 12044 16764 12096
rect 16816 12044 16822 12096
rect 17218 12044 17224 12096
rect 17276 12044 17282 12096
rect 17328 12084 17356 12124
rect 17586 12112 17592 12164
rect 17644 12152 17650 12164
rect 18064 12152 18092 12192
rect 17644 12124 18092 12152
rect 18141 12155 18199 12161
rect 17644 12112 17650 12124
rect 18141 12121 18153 12155
rect 18187 12152 18199 12155
rect 18782 12152 18788 12164
rect 18187 12124 18788 12152
rect 18187 12121 18199 12124
rect 18141 12115 18199 12121
rect 18782 12112 18788 12124
rect 18840 12112 18846 12164
rect 18874 12112 18880 12164
rect 18932 12112 18938 12164
rect 18984 12152 19012 12192
rect 19794 12180 19800 12232
rect 19852 12180 19858 12232
rect 20530 12220 20536 12232
rect 20088 12192 20536 12220
rect 20088 12152 20116 12192
rect 20530 12180 20536 12192
rect 20588 12220 20594 12232
rect 20898 12220 20904 12232
rect 20588 12192 20904 12220
rect 20588 12180 20594 12192
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 21269 12223 21327 12229
rect 21269 12189 21281 12223
rect 21315 12220 21327 12223
rect 21450 12220 21456 12232
rect 21315 12192 21456 12220
rect 21315 12189 21327 12192
rect 21269 12183 21327 12189
rect 21450 12180 21456 12192
rect 21508 12180 21514 12232
rect 22204 12220 22232 12260
rect 22278 12248 22284 12300
rect 22336 12248 22342 12300
rect 23753 12291 23811 12297
rect 23753 12257 23765 12291
rect 23799 12288 23811 12291
rect 23860 12288 23888 12396
rect 26694 12384 26700 12396
rect 26752 12384 26758 12436
rect 27709 12427 27767 12433
rect 27709 12393 27721 12427
rect 27755 12424 27767 12427
rect 27890 12424 27896 12436
rect 27755 12396 27896 12424
rect 27755 12393 27767 12396
rect 27709 12387 27767 12393
rect 27890 12384 27896 12396
rect 27948 12384 27954 12436
rect 32030 12384 32036 12436
rect 32088 12424 32094 12436
rect 34606 12424 34612 12436
rect 32088 12396 34612 12424
rect 32088 12384 32094 12396
rect 34606 12384 34612 12396
rect 34664 12384 34670 12436
rect 35148 12427 35206 12433
rect 35148 12424 35160 12427
rect 34716 12396 35160 12424
rect 26326 12316 26332 12368
rect 26384 12356 26390 12368
rect 26878 12356 26884 12368
rect 26384 12328 26884 12356
rect 26384 12316 26390 12328
rect 26878 12316 26884 12328
rect 26936 12316 26942 12368
rect 29454 12356 29460 12368
rect 27172 12328 29460 12356
rect 27172 12300 27200 12328
rect 29454 12316 29460 12328
rect 29512 12316 29518 12368
rect 34514 12316 34520 12368
rect 34572 12356 34578 12368
rect 34716 12356 34744 12396
rect 35148 12393 35160 12396
rect 35194 12424 35206 12427
rect 35618 12424 35624 12436
rect 35194 12396 35624 12424
rect 35194 12393 35206 12396
rect 35148 12387 35206 12393
rect 35618 12384 35624 12396
rect 35676 12384 35682 12436
rect 36630 12384 36636 12436
rect 36688 12424 36694 12436
rect 39206 12424 39212 12436
rect 36688 12396 39212 12424
rect 36688 12384 36694 12396
rect 39206 12384 39212 12396
rect 39264 12384 39270 12436
rect 39298 12384 39304 12436
rect 39356 12384 39362 12436
rect 34572 12328 34744 12356
rect 39025 12359 39083 12365
rect 34572 12316 34578 12328
rect 39025 12325 39037 12359
rect 39071 12325 39083 12359
rect 39025 12319 39083 12325
rect 40313 12359 40371 12365
rect 40313 12325 40325 12359
rect 40359 12356 40371 12359
rect 47118 12356 47124 12368
rect 40359 12328 47124 12356
rect 40359 12325 40371 12328
rect 40313 12319 40371 12325
rect 23799 12260 23888 12288
rect 23937 12291 23995 12297
rect 23799 12257 23811 12260
rect 23753 12251 23811 12257
rect 23937 12257 23949 12291
rect 23983 12288 23995 12291
rect 24394 12288 24400 12300
rect 23983 12260 24400 12288
rect 23983 12257 23995 12260
rect 23937 12251 23995 12257
rect 24394 12248 24400 12260
rect 24452 12248 24458 12300
rect 24857 12291 24915 12297
rect 24857 12257 24869 12291
rect 24903 12288 24915 12291
rect 24946 12288 24952 12300
rect 24903 12260 24952 12288
rect 24903 12257 24915 12260
rect 24857 12251 24915 12257
rect 24946 12248 24952 12260
rect 25004 12248 25010 12300
rect 27154 12248 27160 12300
rect 27212 12248 27218 12300
rect 27338 12248 27344 12300
rect 27396 12288 27402 12300
rect 28353 12291 28411 12297
rect 28353 12288 28365 12291
rect 27396 12260 28365 12288
rect 27396 12248 27402 12260
rect 28353 12257 28365 12260
rect 28399 12288 28411 12291
rect 29733 12291 29791 12297
rect 29733 12288 29745 12291
rect 28399 12260 29745 12288
rect 28399 12257 28411 12260
rect 28353 12251 28411 12257
rect 29733 12257 29745 12260
rect 29779 12288 29791 12291
rect 30006 12288 30012 12300
rect 29779 12260 30012 12288
rect 29779 12257 29791 12260
rect 29733 12251 29791 12257
rect 30006 12248 30012 12260
rect 30064 12248 30070 12300
rect 31294 12248 31300 12300
rect 31352 12288 31358 12300
rect 31754 12288 31760 12300
rect 31352 12260 31760 12288
rect 31352 12248 31358 12260
rect 31754 12248 31760 12260
rect 31812 12248 31818 12300
rect 33594 12248 33600 12300
rect 33652 12288 33658 12300
rect 33873 12291 33931 12297
rect 33873 12288 33885 12291
rect 33652 12260 33885 12288
rect 33652 12248 33658 12260
rect 33873 12257 33885 12260
rect 33919 12288 33931 12291
rect 37185 12291 37243 12297
rect 37185 12288 37197 12291
rect 33919 12260 37197 12288
rect 33919 12257 33931 12260
rect 33873 12251 33931 12257
rect 37185 12257 37197 12260
rect 37231 12257 37243 12291
rect 37185 12251 37243 12257
rect 38378 12248 38384 12300
rect 38436 12248 38442 12300
rect 38565 12291 38623 12297
rect 38565 12257 38577 12291
rect 38611 12288 38623 12291
rect 38746 12288 38752 12300
rect 38611 12260 38752 12288
rect 38611 12257 38623 12260
rect 38565 12251 38623 12257
rect 38746 12248 38752 12260
rect 38804 12248 38810 12300
rect 39040 12288 39068 12319
rect 47118 12316 47124 12328
rect 47176 12316 47182 12368
rect 39040 12260 41460 12288
rect 22738 12220 22744 12232
rect 22204 12192 22744 12220
rect 22738 12180 22744 12192
rect 22796 12180 22802 12232
rect 24578 12180 24584 12232
rect 24636 12180 24642 12232
rect 26510 12180 26516 12232
rect 26568 12220 26574 12232
rect 27249 12223 27307 12229
rect 27249 12220 27261 12223
rect 26568 12192 27261 12220
rect 26568 12180 26574 12192
rect 27249 12189 27261 12192
rect 27295 12220 27307 12223
rect 27522 12220 27528 12232
rect 27295 12192 27528 12220
rect 27295 12189 27307 12192
rect 27249 12183 27307 12189
rect 27522 12180 27528 12192
rect 27580 12180 27586 12232
rect 27614 12180 27620 12232
rect 27672 12220 27678 12232
rect 28810 12220 28816 12232
rect 27672 12192 28816 12220
rect 27672 12180 27678 12192
rect 28810 12180 28816 12192
rect 28868 12220 28874 12232
rect 29181 12223 29239 12229
rect 29181 12220 29193 12223
rect 28868 12192 29193 12220
rect 28868 12180 28874 12192
rect 29181 12189 29193 12192
rect 29227 12189 29239 12223
rect 31312 12220 31340 12248
rect 31142 12192 31340 12220
rect 29181 12183 29239 12189
rect 31478 12180 31484 12232
rect 31536 12180 31542 12232
rect 32122 12180 32128 12232
rect 32180 12180 32186 12232
rect 34882 12180 34888 12232
rect 34940 12180 34946 12232
rect 37090 12180 37096 12232
rect 37148 12220 37154 12232
rect 41432 12229 41460 12260
rect 49142 12248 49148 12300
rect 49200 12248 49206 12300
rect 37369 12223 37427 12229
rect 37369 12220 37381 12223
rect 37148 12192 37381 12220
rect 37148 12180 37154 12192
rect 37369 12189 37381 12192
rect 37415 12189 37427 12223
rect 40773 12223 40831 12229
rect 40773 12220 40785 12223
rect 37369 12183 37427 12189
rect 37844 12192 40785 12220
rect 18984 12124 20116 12152
rect 20162 12112 20168 12164
rect 20220 12152 20226 12164
rect 22465 12155 22523 12161
rect 22465 12152 22477 12155
rect 20220 12124 22477 12152
rect 20220 12112 20226 12124
rect 22465 12121 22477 12124
rect 22511 12121 22523 12155
rect 23661 12155 23719 12161
rect 23661 12152 23673 12155
rect 22465 12115 22523 12121
rect 22848 12124 23673 12152
rect 19429 12087 19487 12093
rect 19429 12084 19441 12087
rect 17328 12056 19441 12084
rect 19429 12053 19441 12056
rect 19475 12053 19487 12087
rect 19429 12047 19487 12053
rect 19794 12044 19800 12096
rect 19852 12084 19858 12096
rect 19889 12087 19947 12093
rect 19889 12084 19901 12087
rect 19852 12056 19901 12084
rect 19852 12044 19858 12056
rect 19889 12053 19901 12056
rect 19935 12053 19947 12087
rect 19889 12047 19947 12053
rect 20070 12044 20076 12096
rect 20128 12084 20134 12096
rect 22186 12084 22192 12096
rect 20128 12056 22192 12084
rect 20128 12044 20134 12056
rect 22186 12044 22192 12056
rect 22244 12044 22250 12096
rect 22373 12087 22431 12093
rect 22373 12053 22385 12087
rect 22419 12084 22431 12087
rect 22554 12084 22560 12096
rect 22419 12056 22560 12084
rect 22419 12053 22431 12056
rect 22373 12047 22431 12053
rect 22554 12044 22560 12056
rect 22612 12044 22618 12096
rect 22848 12093 22876 12124
rect 23661 12121 23673 12124
rect 23707 12121 23719 12155
rect 26697 12155 26755 12161
rect 26697 12152 26709 12155
rect 26082 12124 26709 12152
rect 23661 12115 23719 12121
rect 22833 12087 22891 12093
rect 22833 12053 22845 12087
rect 22879 12053 22891 12087
rect 22833 12047 22891 12053
rect 25498 12044 25504 12096
rect 25556 12084 25562 12096
rect 26160 12084 26188 12124
rect 26697 12121 26709 12124
rect 26743 12152 26755 12155
rect 27430 12152 27436 12164
rect 26743 12124 27436 12152
rect 26743 12121 26755 12124
rect 26697 12115 26755 12121
rect 27430 12112 27436 12124
rect 27488 12112 27494 12164
rect 29914 12112 29920 12164
rect 29972 12152 29978 12164
rect 30009 12155 30067 12161
rect 30009 12152 30021 12155
rect 29972 12124 30021 12152
rect 29972 12112 29978 12124
rect 30009 12121 30021 12124
rect 30055 12121 30067 12155
rect 31496 12152 31524 12180
rect 32306 12152 32312 12164
rect 31496 12124 32312 12152
rect 30009 12115 30067 12121
rect 32306 12112 32312 12124
rect 32364 12112 32370 12164
rect 32398 12112 32404 12164
rect 32456 12112 32462 12164
rect 32784 12124 32890 12152
rect 34256 12124 35650 12152
rect 25556 12056 26188 12084
rect 25556 12044 25562 12056
rect 27338 12044 27344 12096
rect 27396 12044 27402 12096
rect 27448 12084 27476 12112
rect 27614 12084 27620 12096
rect 27448 12056 27620 12084
rect 27614 12044 27620 12056
rect 27672 12044 27678 12096
rect 31386 12044 31392 12096
rect 31444 12084 31450 12096
rect 31481 12087 31539 12093
rect 31481 12084 31493 12087
rect 31444 12056 31493 12084
rect 31444 12044 31450 12056
rect 31481 12053 31493 12056
rect 31527 12053 31539 12087
rect 31481 12047 31539 12053
rect 31754 12044 31760 12096
rect 31812 12084 31818 12096
rect 32784 12084 32812 12124
rect 34256 12096 34284 12124
rect 33318 12084 33324 12096
rect 31812 12056 33324 12084
rect 31812 12044 31818 12056
rect 33318 12044 33324 12056
rect 33376 12084 33382 12096
rect 34149 12087 34207 12093
rect 34149 12084 34161 12087
rect 33376 12056 34161 12084
rect 33376 12044 33382 12056
rect 34149 12053 34161 12056
rect 34195 12084 34207 12087
rect 34238 12084 34244 12096
rect 34195 12056 34244 12084
rect 34195 12053 34207 12056
rect 34149 12047 34207 12053
rect 34238 12044 34244 12056
rect 34296 12044 34302 12096
rect 34330 12044 34336 12096
rect 34388 12044 34394 12096
rect 35434 12044 35440 12096
rect 35492 12084 35498 12096
rect 36170 12084 36176 12096
rect 35492 12056 36176 12084
rect 35492 12044 35498 12056
rect 36170 12044 36176 12056
rect 36228 12084 36234 12096
rect 36630 12084 36636 12096
rect 36228 12056 36636 12084
rect 36228 12044 36234 12056
rect 36630 12044 36636 12056
rect 36688 12044 36694 12096
rect 37366 12044 37372 12096
rect 37424 12084 37430 12096
rect 37844 12093 37872 12192
rect 40773 12189 40785 12192
rect 40819 12189 40831 12223
rect 40773 12183 40831 12189
rect 41417 12223 41475 12229
rect 41417 12189 41429 12223
rect 41463 12189 41475 12223
rect 45925 12223 45983 12229
rect 45925 12220 45937 12223
rect 41417 12183 41475 12189
rect 45526 12192 45937 12220
rect 38838 12112 38844 12164
rect 38896 12152 38902 12164
rect 39485 12155 39543 12161
rect 39485 12152 39497 12155
rect 38896 12124 39497 12152
rect 38896 12112 38902 12124
rect 39485 12121 39497 12124
rect 39531 12121 39543 12155
rect 39485 12115 39543 12121
rect 40126 12112 40132 12164
rect 40184 12112 40190 12164
rect 37461 12087 37519 12093
rect 37461 12084 37473 12087
rect 37424 12056 37473 12084
rect 37424 12044 37430 12056
rect 37461 12053 37473 12056
rect 37507 12053 37519 12087
rect 37461 12047 37519 12053
rect 37829 12087 37887 12093
rect 37829 12053 37841 12087
rect 37875 12053 37887 12087
rect 37829 12047 37887 12053
rect 38654 12044 38660 12096
rect 38712 12044 38718 12096
rect 40954 12044 40960 12096
rect 41012 12044 41018 12096
rect 41601 12087 41659 12093
rect 41601 12053 41613 12087
rect 41647 12084 41659 12087
rect 45526 12084 45554 12192
rect 45925 12189 45937 12192
rect 45971 12189 45983 12223
rect 45925 12183 45983 12189
rect 47946 12180 47952 12232
rect 48004 12180 48010 12232
rect 41647 12056 45554 12084
rect 41647 12053 41659 12056
rect 41601 12047 41659 12053
rect 46106 12044 46112 12096
rect 46164 12044 46170 12096
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 10502 11840 10508 11892
rect 10560 11880 10566 11892
rect 11330 11880 11336 11892
rect 10560 11852 11336 11880
rect 10560 11840 10566 11852
rect 11330 11840 11336 11852
rect 11388 11880 11394 11892
rect 11517 11883 11575 11889
rect 11517 11880 11529 11883
rect 11388 11852 11529 11880
rect 11388 11840 11394 11852
rect 11517 11849 11529 11852
rect 11563 11880 11575 11883
rect 11977 11883 12035 11889
rect 11977 11880 11989 11883
rect 11563 11852 11989 11880
rect 11563 11849 11575 11852
rect 11517 11843 11575 11849
rect 11977 11849 11989 11852
rect 12023 11849 12035 11883
rect 11977 11843 12035 11849
rect 13538 11840 13544 11892
rect 13596 11880 13602 11892
rect 14185 11883 14243 11889
rect 14185 11880 14197 11883
rect 13596 11852 14197 11880
rect 13596 11840 13602 11852
rect 14185 11849 14197 11852
rect 14231 11849 14243 11883
rect 14185 11843 14243 11849
rect 14274 11840 14280 11892
rect 14332 11840 14338 11892
rect 19245 11883 19303 11889
rect 14660 11852 15792 11880
rect 2498 11772 2504 11824
rect 2556 11812 2562 11824
rect 14660 11812 14688 11852
rect 2556 11784 14688 11812
rect 2556 11772 2562 11784
rect 14734 11772 14740 11824
rect 14792 11812 14798 11824
rect 15764 11812 15792 11852
rect 19245 11849 19257 11883
rect 19291 11880 19303 11883
rect 19334 11880 19340 11892
rect 19291 11852 19340 11880
rect 19291 11849 19303 11852
rect 19245 11843 19303 11849
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 19978 11840 19984 11892
rect 20036 11880 20042 11892
rect 20257 11883 20315 11889
rect 20257 11880 20269 11883
rect 20036 11852 20269 11880
rect 20036 11840 20042 11852
rect 20257 11849 20269 11852
rect 20303 11849 20315 11883
rect 20257 11843 20315 11849
rect 20714 11840 20720 11892
rect 20772 11840 20778 11892
rect 21174 11840 21180 11892
rect 21232 11840 21238 11892
rect 21634 11840 21640 11892
rect 21692 11880 21698 11892
rect 21821 11883 21879 11889
rect 21821 11880 21833 11883
rect 21692 11852 21833 11880
rect 21692 11840 21698 11852
rect 21821 11849 21833 11852
rect 21867 11849 21879 11883
rect 21821 11843 21879 11849
rect 22097 11883 22155 11889
rect 22097 11849 22109 11883
rect 22143 11880 22155 11883
rect 22554 11880 22560 11892
rect 22143 11852 22560 11880
rect 22143 11849 22155 11852
rect 22097 11843 22155 11849
rect 22554 11840 22560 11852
rect 22612 11840 22618 11892
rect 26605 11883 26663 11889
rect 22664 11852 25544 11880
rect 17034 11812 17040 11824
rect 14792 11784 15608 11812
rect 15764 11784 17040 11812
rect 14792 11772 14798 11784
rect 1210 11704 1216 11756
rect 1268 11744 1274 11756
rect 1581 11747 1639 11753
rect 1581 11744 1593 11747
rect 1268 11716 1593 11744
rect 1268 11704 1274 11716
rect 1581 11713 1593 11716
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11713 2375 11747
rect 2317 11707 2375 11713
rect 1302 11636 1308 11688
rect 1360 11676 1366 11688
rect 2332 11676 2360 11707
rect 12342 11704 12348 11756
rect 12400 11744 12406 11756
rect 12713 11747 12771 11753
rect 12713 11744 12725 11747
rect 12400 11716 12725 11744
rect 12400 11704 12406 11716
rect 12713 11713 12725 11716
rect 12759 11713 12771 11747
rect 12713 11707 12771 11713
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11744 12863 11747
rect 14366 11744 14372 11756
rect 12851 11716 14372 11744
rect 12851 11713 12863 11716
rect 12805 11707 12863 11713
rect 14366 11704 14372 11716
rect 14424 11704 14430 11756
rect 14642 11704 14648 11756
rect 14700 11744 14706 11756
rect 15102 11744 15108 11756
rect 14700 11716 15108 11744
rect 14700 11704 14706 11716
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 15286 11704 15292 11756
rect 15344 11744 15350 11756
rect 15473 11747 15531 11753
rect 15473 11744 15485 11747
rect 15344 11716 15485 11744
rect 15344 11704 15350 11716
rect 15473 11713 15485 11716
rect 15519 11713 15531 11747
rect 15580 11744 15608 11784
rect 17034 11772 17040 11784
rect 17092 11772 17098 11824
rect 19061 11815 19119 11821
rect 15580 11716 15700 11744
rect 15473 11707 15531 11713
rect 2777 11679 2835 11685
rect 2777 11676 2789 11679
rect 1360 11648 2789 11676
rect 1360 11636 1366 11648
rect 2777 11645 2789 11648
rect 2823 11645 2835 11679
rect 2777 11639 2835 11645
rect 11790 11636 11796 11688
rect 11848 11676 11854 11688
rect 12897 11679 12955 11685
rect 11848 11648 12434 11676
rect 11848 11636 11854 11648
rect 1765 11611 1823 11617
rect 1765 11577 1777 11611
rect 1811 11608 1823 11611
rect 11514 11608 11520 11620
rect 1811 11580 11520 11608
rect 1811 11577 1823 11580
rect 1765 11571 1823 11577
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 12406 11608 12434 11648
rect 12897 11645 12909 11679
rect 12943 11645 12955 11679
rect 12897 11639 12955 11645
rect 12912 11608 12940 11639
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 13630 11676 13636 11688
rect 13504 11648 13636 11676
rect 13504 11636 13510 11648
rect 13630 11636 13636 11648
rect 13688 11636 13694 11688
rect 13906 11636 13912 11688
rect 13964 11676 13970 11688
rect 14001 11679 14059 11685
rect 14001 11676 14013 11679
rect 13964 11648 14013 11676
rect 13964 11636 13970 11648
rect 14001 11645 14013 11648
rect 14047 11645 14059 11679
rect 14001 11639 14059 11645
rect 14568 11648 15516 11676
rect 12406 11580 12940 11608
rect 13262 11568 13268 11620
rect 13320 11608 13326 11620
rect 13538 11608 13544 11620
rect 13320 11580 13544 11608
rect 13320 11568 13326 11580
rect 13538 11568 13544 11580
rect 13596 11568 13602 11620
rect 13814 11568 13820 11620
rect 13872 11608 13878 11620
rect 14568 11608 14596 11648
rect 13872 11580 14596 11608
rect 14645 11611 14703 11617
rect 13872 11568 13878 11580
rect 14645 11577 14657 11611
rect 14691 11608 14703 11611
rect 15488 11608 15516 11648
rect 15562 11636 15568 11688
rect 15620 11636 15626 11688
rect 15672 11685 15700 11716
rect 16022 11704 16028 11756
rect 16080 11744 16086 11756
rect 16393 11747 16451 11753
rect 16393 11744 16405 11747
rect 16080 11716 16405 11744
rect 16080 11704 16086 11716
rect 16393 11713 16405 11716
rect 16439 11744 16451 11747
rect 16850 11744 16856 11756
rect 16439 11716 16856 11744
rect 16439 11713 16451 11716
rect 16393 11707 16451 11713
rect 16850 11704 16856 11716
rect 16908 11744 16914 11756
rect 17144 11744 17172 11798
rect 19061 11781 19073 11815
rect 19107 11812 19119 11815
rect 19797 11815 19855 11821
rect 19797 11812 19809 11815
rect 19107 11784 19809 11812
rect 19107 11781 19119 11784
rect 19061 11775 19119 11781
rect 19797 11781 19809 11784
rect 19843 11812 19855 11815
rect 20070 11812 20076 11824
rect 19843 11784 20076 11812
rect 19843 11781 19855 11784
rect 19797 11775 19855 11781
rect 20070 11772 20076 11784
rect 20128 11772 20134 11824
rect 21085 11815 21143 11821
rect 21085 11781 21097 11815
rect 21131 11812 21143 11815
rect 21726 11812 21732 11824
rect 21131 11784 21732 11812
rect 21131 11781 21143 11784
rect 21085 11775 21143 11781
rect 21726 11772 21732 11784
rect 21784 11772 21790 11824
rect 22664 11812 22692 11852
rect 24486 11812 24492 11824
rect 21836 11784 22692 11812
rect 23952 11784 24492 11812
rect 16908 11716 17172 11744
rect 16908 11704 16914 11716
rect 19518 11704 19524 11756
rect 19576 11744 19582 11756
rect 19889 11747 19947 11753
rect 19889 11744 19901 11747
rect 19576 11716 19901 11744
rect 19576 11704 19582 11716
rect 19889 11713 19901 11716
rect 19935 11744 19947 11747
rect 20622 11744 20628 11756
rect 19935 11716 20628 11744
rect 19935 11713 19947 11716
rect 19889 11707 19947 11713
rect 20622 11704 20628 11716
rect 20680 11704 20686 11756
rect 20898 11704 20904 11756
rect 20956 11744 20962 11756
rect 21836 11744 21864 11784
rect 20956 11716 21864 11744
rect 20956 11704 20962 11716
rect 22462 11704 22468 11756
rect 22520 11744 22526 11756
rect 23952 11753 23980 11784
rect 24486 11772 24492 11784
rect 24544 11772 24550 11824
rect 25516 11812 25544 11852
rect 26605 11849 26617 11883
rect 26651 11880 26663 11883
rect 27338 11880 27344 11892
rect 26651 11852 27344 11880
rect 26651 11849 26663 11852
rect 26605 11843 26663 11849
rect 27338 11840 27344 11852
rect 27396 11840 27402 11892
rect 27430 11840 27436 11892
rect 27488 11880 27494 11892
rect 27525 11883 27583 11889
rect 27525 11880 27537 11883
rect 27488 11852 27537 11880
rect 27488 11840 27494 11852
rect 27525 11849 27537 11852
rect 27571 11849 27583 11883
rect 27525 11843 27583 11849
rect 27893 11883 27951 11889
rect 27893 11849 27905 11883
rect 27939 11880 27951 11883
rect 28718 11880 28724 11892
rect 27939 11852 28724 11880
rect 27939 11849 27951 11852
rect 27893 11843 27951 11849
rect 28718 11840 28724 11852
rect 28776 11840 28782 11892
rect 31481 11883 31539 11889
rect 31481 11849 31493 11883
rect 31527 11880 31539 11883
rect 31846 11880 31852 11892
rect 31527 11852 31852 11880
rect 31527 11849 31539 11852
rect 31481 11843 31539 11849
rect 31846 11840 31852 11852
rect 31904 11840 31910 11892
rect 32214 11840 32220 11892
rect 32272 11880 32278 11892
rect 32585 11883 32643 11889
rect 32585 11880 32597 11883
rect 32272 11852 32597 11880
rect 32272 11840 32278 11852
rect 32585 11849 32597 11852
rect 32631 11849 32643 11883
rect 32585 11843 32643 11849
rect 32677 11883 32735 11889
rect 32677 11849 32689 11883
rect 32723 11880 32735 11883
rect 32766 11880 32772 11892
rect 32723 11852 32772 11880
rect 32723 11849 32735 11852
rect 32677 11843 32735 11849
rect 32766 11840 32772 11852
rect 32824 11840 32830 11892
rect 33778 11840 33784 11892
rect 33836 11880 33842 11892
rect 33873 11883 33931 11889
rect 33873 11880 33885 11883
rect 33836 11852 33885 11880
rect 33836 11840 33842 11852
rect 33873 11849 33885 11852
rect 33919 11849 33931 11883
rect 33873 11843 33931 11849
rect 34238 11840 34244 11892
rect 34296 11880 34302 11892
rect 34701 11883 34759 11889
rect 34701 11880 34713 11883
rect 34296 11852 34713 11880
rect 34296 11840 34302 11852
rect 34701 11849 34713 11852
rect 34747 11849 34759 11883
rect 34701 11843 34759 11849
rect 25516 11784 27476 11812
rect 22557 11747 22615 11753
rect 22557 11744 22569 11747
rect 22520 11716 22569 11744
rect 22520 11704 22526 11716
rect 22557 11713 22569 11716
rect 22603 11713 22615 11747
rect 22557 11707 22615 11713
rect 23385 11747 23443 11753
rect 23385 11713 23397 11747
rect 23431 11744 23443 11747
rect 23937 11747 23995 11753
rect 23937 11744 23949 11747
rect 23431 11716 23949 11744
rect 23431 11713 23443 11716
rect 23385 11707 23443 11713
rect 23937 11713 23949 11716
rect 23983 11713 23995 11747
rect 25498 11744 25504 11756
rect 25346 11716 25504 11744
rect 23937 11707 23995 11713
rect 25498 11704 25504 11716
rect 25556 11704 25562 11756
rect 25774 11704 25780 11756
rect 25832 11744 25838 11756
rect 26145 11747 26203 11753
rect 26145 11744 26157 11747
rect 25832 11716 26157 11744
rect 25832 11704 25838 11716
rect 26145 11713 26157 11716
rect 26191 11744 26203 11747
rect 27062 11744 27068 11756
rect 26191 11716 27068 11744
rect 26191 11713 26203 11716
rect 26145 11707 26203 11713
rect 27062 11704 27068 11716
rect 27120 11744 27126 11756
rect 27338 11744 27344 11756
rect 27120 11716 27344 11744
rect 27120 11704 27126 11716
rect 27338 11704 27344 11716
rect 27396 11704 27402 11756
rect 15657 11679 15715 11685
rect 15657 11645 15669 11679
rect 15703 11645 15715 11679
rect 15657 11639 15715 11645
rect 16114 11636 16120 11688
rect 16172 11676 16178 11688
rect 17586 11676 17592 11688
rect 16172 11648 17592 11676
rect 16172 11636 16178 11648
rect 17586 11636 17592 11648
rect 17644 11636 17650 11688
rect 18325 11679 18383 11685
rect 18325 11645 18337 11679
rect 18371 11676 18383 11679
rect 18601 11679 18659 11685
rect 18371 11648 18552 11676
rect 18371 11645 18383 11648
rect 18325 11639 18383 11645
rect 16853 11611 16911 11617
rect 16853 11608 16865 11611
rect 14691 11580 15424 11608
rect 15488 11580 16865 11608
rect 14691 11577 14703 11580
rect 14645 11571 14703 11577
rect 2501 11543 2559 11549
rect 2501 11509 2513 11543
rect 2547 11540 2559 11543
rect 4154 11540 4160 11552
rect 2547 11512 4160 11540
rect 2547 11509 2559 11512
rect 2501 11503 2559 11509
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 12342 11500 12348 11552
rect 12400 11500 12406 11552
rect 13354 11500 13360 11552
rect 13412 11500 13418 11552
rect 14826 11500 14832 11552
rect 14884 11540 14890 11552
rect 15105 11543 15163 11549
rect 15105 11540 15117 11543
rect 14884 11512 15117 11540
rect 14884 11500 14890 11512
rect 15105 11509 15117 11512
rect 15151 11509 15163 11543
rect 15396 11540 15424 11580
rect 16853 11577 16865 11580
rect 16899 11577 16911 11611
rect 16853 11571 16911 11577
rect 15470 11540 15476 11552
rect 15396 11512 15476 11540
rect 15105 11503 15163 11509
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 16206 11500 16212 11552
rect 16264 11540 16270 11552
rect 16301 11543 16359 11549
rect 16301 11540 16313 11543
rect 16264 11512 16313 11540
rect 16264 11500 16270 11512
rect 16301 11509 16313 11512
rect 16347 11540 16359 11543
rect 16482 11540 16488 11552
rect 16347 11512 16488 11540
rect 16347 11509 16359 11512
rect 16301 11503 16359 11509
rect 16482 11500 16488 11512
rect 16540 11500 16546 11552
rect 18524 11540 18552 11648
rect 18601 11645 18613 11679
rect 18647 11676 18659 11679
rect 18782 11676 18788 11688
rect 18647 11648 18788 11676
rect 18647 11645 18659 11648
rect 18601 11639 18659 11645
rect 18782 11636 18788 11648
rect 18840 11636 18846 11688
rect 19613 11679 19671 11685
rect 19613 11645 19625 11679
rect 19659 11645 19671 11679
rect 19613 11639 19671 11645
rect 19628 11608 19656 11639
rect 20070 11636 20076 11688
rect 20128 11676 20134 11688
rect 20128 11648 21128 11676
rect 20128 11636 20134 11648
rect 20990 11608 20996 11620
rect 19628 11580 20996 11608
rect 20990 11568 20996 11580
rect 21048 11568 21054 11620
rect 21100 11608 21128 11648
rect 21358 11636 21364 11688
rect 21416 11636 21422 11688
rect 22278 11636 22284 11688
rect 22336 11676 22342 11688
rect 24213 11679 24271 11685
rect 24213 11676 24225 11679
rect 22336 11648 24225 11676
rect 22336 11636 22342 11648
rect 24213 11645 24225 11648
rect 24259 11676 24271 11679
rect 26326 11676 26332 11688
rect 24259 11648 26332 11676
rect 24259 11645 24271 11648
rect 24213 11639 24271 11645
rect 26326 11636 26332 11648
rect 26384 11636 26390 11688
rect 27246 11636 27252 11688
rect 27304 11636 27310 11688
rect 27448 11685 27476 11784
rect 27614 11772 27620 11824
rect 27672 11812 27678 11824
rect 30009 11815 30067 11821
rect 27672 11784 28842 11812
rect 27672 11772 27678 11784
rect 30009 11781 30021 11815
rect 30055 11812 30067 11815
rect 31386 11812 31392 11824
rect 30055 11784 31392 11812
rect 30055 11781 30067 11784
rect 30009 11775 30067 11781
rect 31386 11772 31392 11784
rect 31444 11812 31450 11824
rect 31444 11784 31524 11812
rect 31444 11772 31450 11784
rect 31110 11704 31116 11756
rect 31168 11704 31174 11756
rect 31496 11744 31524 11784
rect 31570 11772 31576 11824
rect 31628 11812 31634 11824
rect 31754 11812 31760 11824
rect 31628 11784 31760 11812
rect 31628 11772 31634 11784
rect 31754 11772 31760 11784
rect 31812 11772 31818 11824
rect 32306 11772 32312 11824
rect 32364 11812 32370 11824
rect 34716 11812 34744 11843
rect 34790 11840 34796 11892
rect 34848 11880 34854 11892
rect 34974 11880 34980 11892
rect 34848 11852 34980 11880
rect 34848 11840 34854 11852
rect 34974 11840 34980 11852
rect 35032 11840 35038 11892
rect 36078 11840 36084 11892
rect 36136 11880 36142 11892
rect 37737 11883 37795 11889
rect 37737 11880 37749 11883
rect 36136 11852 37749 11880
rect 36136 11840 36142 11852
rect 37737 11849 37749 11852
rect 37783 11849 37795 11883
rect 37737 11843 37795 11849
rect 38654 11840 38660 11892
rect 38712 11840 38718 11892
rect 40126 11840 40132 11892
rect 40184 11880 40190 11892
rect 40405 11883 40463 11889
rect 40405 11880 40417 11883
rect 40184 11852 40417 11880
rect 40184 11840 40190 11852
rect 40405 11849 40417 11852
rect 40451 11849 40463 11883
rect 40405 11843 40463 11849
rect 35894 11812 35900 11824
rect 32364 11784 33824 11812
rect 34716 11784 35900 11812
rect 32364 11772 32370 11784
rect 33796 11753 33824 11784
rect 35894 11772 35900 11784
rect 35952 11772 35958 11824
rect 37274 11772 37280 11824
rect 37332 11812 37338 11824
rect 39117 11815 39175 11821
rect 39117 11812 39129 11815
rect 37332 11784 39129 11812
rect 37332 11772 37338 11784
rect 39117 11781 39129 11784
rect 39163 11781 39175 11815
rect 39117 11775 39175 11781
rect 40954 11772 40960 11824
rect 41012 11812 41018 11824
rect 45097 11815 45155 11821
rect 45097 11812 45109 11815
rect 41012 11784 45109 11812
rect 41012 11772 41018 11784
rect 45097 11781 45109 11784
rect 45143 11781 45155 11815
rect 45097 11775 45155 11781
rect 49142 11772 49148 11824
rect 49200 11772 49206 11824
rect 33781 11747 33839 11753
rect 31496 11716 33640 11744
rect 27433 11679 27491 11685
rect 27433 11645 27445 11679
rect 27479 11676 27491 11679
rect 27706 11676 27712 11688
rect 27479 11648 27712 11676
rect 27479 11645 27491 11648
rect 27433 11639 27491 11645
rect 27706 11636 27712 11648
rect 27764 11636 27770 11688
rect 28537 11679 28595 11685
rect 28537 11645 28549 11679
rect 28583 11676 28595 11679
rect 29546 11676 29552 11688
rect 28583 11648 29552 11676
rect 28583 11645 28595 11648
rect 28537 11639 28595 11645
rect 21100 11580 24072 11608
rect 24044 11552 24072 11580
rect 27338 11568 27344 11620
rect 27396 11608 27402 11620
rect 28552 11608 28580 11639
rect 29546 11636 29552 11648
rect 29604 11636 29610 11688
rect 29638 11636 29644 11688
rect 29696 11676 29702 11688
rect 30285 11679 30343 11685
rect 30285 11676 30297 11679
rect 29696 11648 30297 11676
rect 29696 11636 29702 11648
rect 30285 11645 30297 11648
rect 30331 11645 30343 11679
rect 30285 11639 30343 11645
rect 30834 11636 30840 11688
rect 30892 11636 30898 11688
rect 31021 11679 31079 11685
rect 31021 11645 31033 11679
rect 31067 11676 31079 11679
rect 31846 11676 31852 11688
rect 31067 11648 31852 11676
rect 31067 11645 31079 11648
rect 31021 11639 31079 11645
rect 31846 11636 31852 11648
rect 31904 11636 31910 11688
rect 32493 11679 32551 11685
rect 32493 11645 32505 11679
rect 32539 11676 32551 11679
rect 32582 11676 32588 11688
rect 32539 11648 32588 11676
rect 32539 11645 32551 11648
rect 32493 11639 32551 11645
rect 32582 11636 32588 11648
rect 32640 11636 32646 11688
rect 33502 11676 33508 11688
rect 32968 11648 33508 11676
rect 27396 11580 28580 11608
rect 27396 11568 27402 11580
rect 30466 11568 30472 11620
rect 30524 11608 30530 11620
rect 32968 11608 32996 11648
rect 33502 11636 33508 11648
rect 33560 11636 33566 11688
rect 33612 11685 33640 11716
rect 33781 11713 33793 11747
rect 33827 11713 33839 11747
rect 33781 11707 33839 11713
rect 36814 11704 36820 11756
rect 36872 11744 36878 11756
rect 37829 11747 37887 11753
rect 37829 11744 37841 11747
rect 36872 11716 37841 11744
rect 36872 11704 36878 11716
rect 37829 11713 37841 11716
rect 37875 11713 37887 11747
rect 38378 11744 38384 11756
rect 37829 11707 37887 11713
rect 37936 11716 38384 11744
rect 33597 11679 33655 11685
rect 33597 11645 33609 11679
rect 33643 11645 33655 11679
rect 33597 11639 33655 11645
rect 34882 11636 34888 11688
rect 34940 11676 34946 11688
rect 35161 11679 35219 11685
rect 35161 11676 35173 11679
rect 34940 11648 35173 11676
rect 34940 11636 34946 11648
rect 35161 11645 35173 11648
rect 35207 11645 35219 11679
rect 35161 11639 35219 11645
rect 30524 11580 32996 11608
rect 33045 11611 33103 11617
rect 30524 11568 30530 11580
rect 33045 11577 33057 11611
rect 33091 11608 33103 11611
rect 33870 11608 33876 11620
rect 33091 11580 33876 11608
rect 33091 11577 33103 11580
rect 33045 11571 33103 11577
rect 33870 11568 33876 11580
rect 33928 11568 33934 11620
rect 34241 11611 34299 11617
rect 34241 11577 34253 11611
rect 34287 11608 34299 11611
rect 35066 11608 35072 11620
rect 34287 11580 35072 11608
rect 34287 11577 34299 11580
rect 34241 11571 34299 11577
rect 35066 11568 35072 11580
rect 35124 11568 35130 11620
rect 21266 11540 21272 11552
rect 18524 11512 21272 11540
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 22281 11543 22339 11549
rect 22281 11509 22293 11543
rect 22327 11540 22339 11543
rect 22462 11540 22468 11552
rect 22327 11512 22468 11540
rect 22327 11509 22339 11512
rect 22281 11503 22339 11509
rect 22462 11500 22468 11512
rect 22520 11500 22526 11552
rect 24026 11500 24032 11552
rect 24084 11500 24090 11552
rect 24394 11500 24400 11552
rect 24452 11540 24458 11552
rect 25685 11543 25743 11549
rect 25685 11540 25697 11543
rect 24452 11512 25697 11540
rect 24452 11500 24458 11512
rect 25685 11509 25697 11512
rect 25731 11509 25743 11543
rect 25685 11503 25743 11509
rect 34606 11500 34612 11552
rect 34664 11500 34670 11552
rect 35176 11540 35204 11639
rect 35434 11636 35440 11688
rect 35492 11636 35498 11688
rect 36630 11636 36636 11688
rect 36688 11676 36694 11688
rect 37553 11679 37611 11685
rect 37553 11676 37565 11679
rect 36688 11648 37565 11676
rect 36688 11636 36694 11648
rect 37553 11645 37565 11648
rect 37599 11645 37611 11679
rect 37553 11639 37611 11645
rect 36909 11611 36967 11617
rect 36909 11577 36921 11611
rect 36955 11608 36967 11611
rect 37936 11608 37964 11716
rect 38378 11704 38384 11716
rect 38436 11704 38442 11756
rect 39022 11704 39028 11756
rect 39080 11704 39086 11756
rect 39945 11747 40003 11753
rect 39945 11713 39957 11747
rect 39991 11744 40003 11747
rect 40589 11747 40647 11753
rect 40589 11744 40601 11747
rect 39991 11716 40601 11744
rect 39991 11713 40003 11716
rect 39945 11707 40003 11713
rect 40589 11713 40601 11716
rect 40635 11713 40647 11747
rect 40589 11707 40647 11713
rect 39206 11636 39212 11688
rect 39264 11636 39270 11688
rect 36955 11580 37964 11608
rect 36955 11577 36967 11580
rect 36909 11571 36967 11577
rect 38010 11568 38016 11620
rect 38068 11608 38074 11620
rect 39960 11608 39988 11707
rect 46106 11704 46112 11756
rect 46164 11744 46170 11756
rect 47949 11747 48007 11753
rect 47949 11744 47961 11747
rect 46164 11716 47961 11744
rect 46164 11704 46170 11716
rect 47949 11713 47961 11716
rect 47995 11713 48007 11747
rect 47949 11707 48007 11713
rect 38068 11580 39988 11608
rect 40129 11611 40187 11617
rect 38068 11568 38074 11580
rect 40129 11577 40141 11611
rect 40175 11608 40187 11611
rect 45281 11611 45339 11617
rect 40175 11580 42840 11608
rect 40175 11577 40187 11580
rect 40129 11571 40187 11577
rect 35618 11540 35624 11552
rect 35176 11512 35624 11540
rect 35618 11500 35624 11512
rect 35676 11500 35682 11552
rect 38197 11543 38255 11549
rect 38197 11509 38209 11543
rect 38243 11540 38255 11543
rect 40218 11540 40224 11552
rect 38243 11512 40224 11540
rect 38243 11509 38255 11512
rect 38197 11503 38255 11509
rect 40218 11500 40224 11512
rect 40276 11500 40282 11552
rect 42812 11540 42840 11580
rect 45281 11577 45293 11611
rect 45327 11608 45339 11611
rect 46750 11608 46756 11620
rect 45327 11580 46756 11608
rect 45327 11577 45339 11580
rect 45281 11571 45339 11577
rect 46750 11568 46756 11580
rect 46808 11568 46814 11620
rect 47762 11540 47768 11552
rect 42812 11512 47768 11540
rect 47762 11500 47768 11512
rect 47820 11500 47826 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 1210 11296 1216 11348
rect 1268 11336 1274 11348
rect 2133 11339 2191 11345
rect 2133 11336 2145 11339
rect 1268 11308 2145 11336
rect 1268 11296 1274 11308
rect 2133 11305 2145 11308
rect 2179 11305 2191 11339
rect 2133 11299 2191 11305
rect 6886 11308 13400 11336
rect 1765 11271 1823 11277
rect 1765 11237 1777 11271
rect 1811 11268 1823 11271
rect 6886 11268 6914 11308
rect 1811 11240 6914 11268
rect 13372 11268 13400 11308
rect 13998 11296 14004 11348
rect 14056 11336 14062 11348
rect 14369 11339 14427 11345
rect 14369 11336 14381 11339
rect 14056 11308 14381 11336
rect 14056 11296 14062 11308
rect 14369 11305 14381 11308
rect 14415 11305 14427 11339
rect 15562 11336 15568 11348
rect 14369 11299 14427 11305
rect 14752 11308 15568 11336
rect 14458 11268 14464 11280
rect 13372 11240 14464 11268
rect 1811 11237 1823 11240
rect 1765 11231 1823 11237
rect 14458 11228 14464 11240
rect 14516 11228 14522 11280
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11200 11023 11203
rect 11054 11200 11060 11212
rect 11011 11172 11060 11200
rect 11011 11169 11023 11172
rect 10965 11163 11023 11169
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 11790 11160 11796 11212
rect 11848 11200 11854 11212
rect 12437 11203 12495 11209
rect 12437 11200 12449 11203
rect 11848 11172 12449 11200
rect 11848 11160 11854 11172
rect 12437 11169 12449 11172
rect 12483 11169 12495 11203
rect 12437 11163 12495 11169
rect 12894 11160 12900 11212
rect 12952 11200 12958 11212
rect 14752 11200 14780 11308
rect 15562 11296 15568 11308
rect 15620 11296 15626 11348
rect 16666 11296 16672 11348
rect 16724 11336 16730 11348
rect 16761 11339 16819 11345
rect 16761 11336 16773 11339
rect 16724 11308 16773 11336
rect 16724 11296 16730 11308
rect 16761 11305 16773 11308
rect 16807 11305 16819 11339
rect 17957 11339 18015 11345
rect 17957 11336 17969 11339
rect 16761 11299 16819 11305
rect 16868 11308 17969 11336
rect 15102 11228 15108 11280
rect 15160 11268 15166 11280
rect 16868 11268 16896 11308
rect 17957 11305 17969 11308
rect 18003 11305 18015 11339
rect 17957 11299 18015 11305
rect 18874 11296 18880 11348
rect 18932 11336 18938 11348
rect 19061 11339 19119 11345
rect 19061 11336 19073 11339
rect 18932 11308 19073 11336
rect 18932 11296 18938 11308
rect 19061 11305 19073 11308
rect 19107 11336 19119 11339
rect 19337 11339 19395 11345
rect 19337 11336 19349 11339
rect 19107 11308 19349 11336
rect 19107 11305 19119 11308
rect 19061 11299 19119 11305
rect 19337 11305 19349 11308
rect 19383 11336 19395 11339
rect 22462 11336 22468 11348
rect 19383 11308 22468 11336
rect 19383 11305 19395 11308
rect 19337 11299 19395 11305
rect 22462 11296 22468 11308
rect 22520 11296 22526 11348
rect 23290 11296 23296 11348
rect 23348 11296 23354 11348
rect 25222 11336 25228 11348
rect 24320 11308 25228 11336
rect 15160 11240 16896 11268
rect 15160 11228 15166 11240
rect 17586 11228 17592 11280
rect 17644 11268 17650 11280
rect 17644 11240 18644 11268
rect 17644 11228 17650 11240
rect 18616 11212 18644 11240
rect 19518 11228 19524 11280
rect 19576 11228 19582 11280
rect 20070 11268 20076 11280
rect 19904 11240 20076 11268
rect 12952 11172 14780 11200
rect 12952 11160 12958 11172
rect 14826 11160 14832 11212
rect 14884 11160 14890 11212
rect 15013 11203 15071 11209
rect 15013 11169 15025 11203
rect 15059 11200 15071 11203
rect 15378 11200 15384 11212
rect 15059 11172 15384 11200
rect 15059 11169 15071 11172
rect 15013 11163 15071 11169
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11169 15807 11203
rect 15749 11163 15807 11169
rect 15841 11203 15899 11209
rect 15841 11169 15853 11203
rect 15887 11200 15899 11203
rect 15930 11200 15936 11212
rect 15887 11172 15936 11200
rect 15887 11169 15899 11172
rect 15841 11163 15899 11169
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 2317 11135 2375 11141
rect 2317 11132 2329 11135
rect 1636 11104 2329 11132
rect 1636 11092 1642 11104
rect 2317 11101 2329 11104
rect 2363 11101 2375 11135
rect 2317 11095 2375 11101
rect 11330 11092 11336 11144
rect 11388 11092 11394 11144
rect 12713 11135 12771 11141
rect 12713 11101 12725 11135
rect 12759 11132 12771 11135
rect 13630 11132 13636 11144
rect 12759 11104 13636 11132
rect 12759 11101 12771 11104
rect 12713 11095 12771 11101
rect 13630 11092 13636 11104
rect 13688 11092 13694 11144
rect 15764 11132 15792 11163
rect 15930 11160 15936 11172
rect 15988 11160 15994 11212
rect 17405 11203 17463 11209
rect 17405 11169 17417 11203
rect 17451 11200 17463 11203
rect 17451 11172 18460 11200
rect 17451 11169 17463 11172
rect 17405 11163 17463 11169
rect 16390 11132 16396 11144
rect 15764 11104 16396 11132
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 16482 11092 16488 11144
rect 16540 11132 16546 11144
rect 17221 11135 17279 11141
rect 16540 11104 17080 11132
rect 16540 11092 16546 11104
rect 12894 11024 12900 11076
rect 12952 11064 12958 11076
rect 12989 11067 13047 11073
rect 12989 11064 13001 11067
rect 12952 11036 13001 11064
rect 12952 11024 12958 11036
rect 12989 11033 13001 11036
rect 13035 11033 13047 11067
rect 12989 11027 13047 11033
rect 13265 11067 13323 11073
rect 13265 11033 13277 11067
rect 13311 11064 13323 11067
rect 13446 11064 13452 11076
rect 13311 11036 13452 11064
rect 13311 11033 13323 11036
rect 13265 11027 13323 11033
rect 13446 11024 13452 11036
rect 13504 11024 13510 11076
rect 13725 11067 13783 11073
rect 13725 11033 13737 11067
rect 13771 11064 13783 11067
rect 15838 11064 15844 11076
rect 13771 11036 15844 11064
rect 13771 11033 13783 11036
rect 13725 11027 13783 11033
rect 15838 11024 15844 11036
rect 15896 11024 15902 11076
rect 15933 11067 15991 11073
rect 15933 11033 15945 11067
rect 15979 11064 15991 11067
rect 16574 11064 16580 11076
rect 15979 11036 16580 11064
rect 15979 11033 15991 11036
rect 15933 11027 15991 11033
rect 16574 11024 16580 11036
rect 16632 11024 16638 11076
rect 14734 10956 14740 11008
rect 14792 10956 14798 11008
rect 16298 10956 16304 11008
rect 16356 10956 16362 11008
rect 17052 10996 17080 11104
rect 17221 11101 17233 11135
rect 17267 11132 17279 11135
rect 18322 11132 18328 11144
rect 17267 11104 18328 11132
rect 17267 11101 17279 11104
rect 17221 11095 17279 11101
rect 18322 11092 18328 11104
rect 18380 11092 18386 11144
rect 18432 11132 18460 11172
rect 18598 11160 18604 11212
rect 18656 11160 18662 11212
rect 18690 11160 18696 11212
rect 18748 11200 18754 11212
rect 19904 11200 19932 11240
rect 20070 11228 20076 11240
rect 20128 11228 20134 11280
rect 18748 11172 19932 11200
rect 19981 11203 20039 11209
rect 18748 11160 18754 11172
rect 19981 11169 19993 11203
rect 20027 11200 20039 11203
rect 20162 11200 20168 11212
rect 20027 11172 20168 11200
rect 20027 11169 20039 11172
rect 19981 11163 20039 11169
rect 20162 11160 20168 11172
rect 20220 11160 20226 11212
rect 20441 11203 20499 11209
rect 20441 11169 20453 11203
rect 20487 11200 20499 11203
rect 21266 11200 21272 11212
rect 20487 11172 21272 11200
rect 20487 11169 20499 11172
rect 20441 11163 20499 11169
rect 21266 11160 21272 11172
rect 21324 11160 21330 11212
rect 21913 11203 21971 11209
rect 21913 11169 21925 11203
rect 21959 11200 21971 11203
rect 23750 11200 23756 11212
rect 21959 11172 23756 11200
rect 21959 11169 21971 11172
rect 21913 11163 21971 11169
rect 23750 11160 23756 11172
rect 23808 11160 23814 11212
rect 23937 11203 23995 11209
rect 23937 11169 23949 11203
rect 23983 11200 23995 11203
rect 24320 11200 24348 11308
rect 25222 11296 25228 11308
rect 25280 11296 25286 11348
rect 26329 11339 26387 11345
rect 26329 11305 26341 11339
rect 26375 11336 26387 11339
rect 26602 11336 26608 11348
rect 26375 11308 26608 11336
rect 26375 11305 26387 11308
rect 26329 11299 26387 11305
rect 26602 11296 26608 11308
rect 26660 11296 26666 11348
rect 28810 11296 28816 11348
rect 28868 11336 28874 11348
rect 28997 11339 29055 11345
rect 28997 11336 29009 11339
rect 28868 11308 29009 11336
rect 28868 11296 28874 11308
rect 28997 11305 29009 11308
rect 29043 11336 29055 11339
rect 34054 11336 34060 11348
rect 29043 11308 34060 11336
rect 29043 11305 29055 11308
rect 28997 11299 29055 11305
rect 28629 11271 28687 11277
rect 28629 11237 28641 11271
rect 28675 11268 28687 11271
rect 28902 11268 28908 11280
rect 28675 11240 28908 11268
rect 28675 11237 28687 11240
rect 28629 11231 28687 11237
rect 28902 11228 28908 11240
rect 28960 11228 28966 11280
rect 30466 11228 30472 11280
rect 30524 11228 30530 11280
rect 23983 11172 24348 11200
rect 23983 11169 23995 11172
rect 23937 11163 23995 11169
rect 24394 11160 24400 11212
rect 24452 11200 24458 11212
rect 24857 11203 24915 11209
rect 24857 11200 24869 11203
rect 24452 11172 24869 11200
rect 24452 11160 24458 11172
rect 24857 11169 24869 11172
rect 24903 11169 24915 11203
rect 24857 11163 24915 11169
rect 27154 11160 27160 11212
rect 27212 11160 27218 11212
rect 29917 11203 29975 11209
rect 29917 11169 29929 11203
rect 29963 11200 29975 11203
rect 32030 11200 32036 11212
rect 29963 11172 32036 11200
rect 29963 11169 29975 11172
rect 29917 11163 29975 11169
rect 32030 11160 32036 11172
rect 32088 11160 32094 11212
rect 32582 11160 32588 11212
rect 32640 11200 32646 11212
rect 32861 11203 32919 11209
rect 32861 11200 32873 11203
rect 32640 11172 32873 11200
rect 32640 11160 32646 11172
rect 32861 11169 32873 11172
rect 32907 11169 32919 11203
rect 32861 11163 32919 11169
rect 19518 11132 19524 11144
rect 18432 11104 19524 11132
rect 19518 11092 19524 11104
rect 19576 11092 19582 11144
rect 22189 11135 22247 11141
rect 22189 11101 22201 11135
rect 22235 11132 22247 11135
rect 24578 11132 24584 11144
rect 22235 11104 24584 11132
rect 22235 11101 22247 11104
rect 22189 11095 22247 11101
rect 24578 11092 24584 11104
rect 24636 11092 24642 11144
rect 26878 11092 26884 11144
rect 26936 11092 26942 11144
rect 29638 11092 29644 11144
rect 29696 11132 29702 11144
rect 33336 11141 33364 11308
rect 34054 11296 34060 11308
rect 34112 11336 34118 11348
rect 34606 11336 34612 11348
rect 34112 11308 34612 11336
rect 34112 11296 34118 11308
rect 34606 11296 34612 11308
rect 34664 11336 34670 11348
rect 34701 11339 34759 11345
rect 34701 11336 34713 11339
rect 34664 11308 34713 11336
rect 34664 11296 34670 11308
rect 34701 11305 34713 11308
rect 34747 11305 34759 11339
rect 34701 11299 34759 11305
rect 35066 11296 35072 11348
rect 35124 11336 35130 11348
rect 38749 11339 38807 11345
rect 35124 11308 38240 11336
rect 35124 11296 35130 11308
rect 33502 11228 33508 11280
rect 33560 11268 33566 11280
rect 35986 11268 35992 11280
rect 33560 11240 35992 11268
rect 33560 11228 33566 11240
rect 35986 11228 35992 11240
rect 36044 11228 36050 11280
rect 35894 11160 35900 11212
rect 35952 11200 35958 11212
rect 36906 11200 36912 11212
rect 35952 11172 36912 11200
rect 35952 11160 35958 11172
rect 31113 11135 31171 11141
rect 31113 11132 31125 11135
rect 29696 11104 31125 11132
rect 29696 11092 29702 11104
rect 31113 11101 31125 11104
rect 31159 11101 31171 11135
rect 31113 11095 31171 11101
rect 33321 11135 33379 11141
rect 33321 11101 33333 11135
rect 33367 11101 33379 11135
rect 33321 11095 33379 11101
rect 33962 11092 33968 11144
rect 34020 11132 34026 11144
rect 34020 11104 35756 11132
rect 36372 11118 36400 11172
rect 36906 11160 36912 11172
rect 36964 11160 36970 11212
rect 37458 11160 37464 11212
rect 37516 11200 37522 11212
rect 37737 11203 37795 11209
rect 37737 11200 37749 11203
rect 37516 11172 37749 11200
rect 37516 11160 37522 11172
rect 37737 11169 37749 11172
rect 37783 11169 37795 11203
rect 37737 11163 37795 11169
rect 38212 11141 38240 11308
rect 38749 11305 38761 11339
rect 38795 11336 38807 11339
rect 38838 11336 38844 11348
rect 38795 11308 38844 11336
rect 38795 11305 38807 11308
rect 38749 11299 38807 11305
rect 38838 11296 38844 11308
rect 38896 11296 38902 11348
rect 39574 11296 39580 11348
rect 39632 11296 39638 11348
rect 44082 11336 44088 11348
rect 39868 11308 44088 11336
rect 38381 11271 38439 11277
rect 38381 11237 38393 11271
rect 38427 11268 38439 11271
rect 39868 11268 39896 11308
rect 44082 11296 44088 11308
rect 44140 11296 44146 11348
rect 38427 11240 39896 11268
rect 40957 11271 41015 11277
rect 38427 11237 38439 11240
rect 38381 11231 38439 11237
rect 40957 11237 40969 11271
rect 41003 11268 41015 11271
rect 41003 11240 41414 11268
rect 41003 11237 41015 11240
rect 40957 11231 41015 11237
rect 38197 11135 38255 11141
rect 34020 11092 34026 11104
rect 17126 11024 17132 11076
rect 17184 11024 17190 11076
rect 20530 11064 20536 11076
rect 17236 11036 20536 11064
rect 17236 10996 17264 11036
rect 18340 11005 18368 11036
rect 20530 11024 20536 11036
rect 20588 11024 20594 11076
rect 21174 11024 21180 11076
rect 21232 11024 21238 11076
rect 23661 11067 23719 11073
rect 23661 11033 23673 11067
rect 23707 11064 23719 11067
rect 23934 11064 23940 11076
rect 23707 11036 23940 11064
rect 23707 11033 23719 11036
rect 23661 11027 23719 11033
rect 23934 11024 23940 11036
rect 23992 11024 23998 11076
rect 25498 11024 25504 11076
rect 25556 11024 25562 11076
rect 27614 11024 27620 11076
rect 27672 11024 27678 11076
rect 29012 11036 30144 11064
rect 17052 10968 17264 10996
rect 18325 10999 18383 11005
rect 18325 10965 18337 10999
rect 18371 10965 18383 10999
rect 18325 10959 18383 10965
rect 18417 10999 18475 11005
rect 18417 10965 18429 10999
rect 18463 10996 18475 10999
rect 18782 10996 18788 11008
rect 18463 10968 18788 10996
rect 18463 10965 18475 10968
rect 18417 10959 18475 10965
rect 18782 10956 18788 10968
rect 18840 10956 18846 11008
rect 19978 10956 19984 11008
rect 20036 10996 20042 11008
rect 22370 10996 22376 11008
rect 20036 10968 22376 10996
rect 20036 10956 20042 10968
rect 22370 10956 22376 10968
rect 22428 10956 22434 11008
rect 22646 10956 22652 11008
rect 22704 10956 22710 11008
rect 23753 10999 23811 11005
rect 23753 10965 23765 10999
rect 23799 10996 23811 10999
rect 24026 10996 24032 11008
rect 23799 10968 24032 10996
rect 23799 10965 23811 10968
rect 23753 10959 23811 10965
rect 24026 10956 24032 10968
rect 24084 10956 24090 11008
rect 24670 10956 24676 11008
rect 24728 10996 24734 11008
rect 29012 10996 29040 11036
rect 24728 10968 29040 10996
rect 24728 10956 24734 10968
rect 29178 10956 29184 11008
rect 29236 10996 29242 11008
rect 29273 10999 29331 11005
rect 29273 10996 29285 10999
rect 29236 10968 29285 10996
rect 29236 10956 29242 10968
rect 29273 10965 29285 10968
rect 29319 10965 29331 10999
rect 29273 10959 29331 10965
rect 29362 10956 29368 11008
rect 29420 10996 29426 11008
rect 30006 10996 30012 11008
rect 29420 10968 30012 10996
rect 29420 10956 29426 10968
rect 30006 10956 30012 10968
rect 30064 10956 30070 11008
rect 30116 11005 30144 11036
rect 31386 11024 31392 11076
rect 31444 11024 31450 11076
rect 31478 11024 31484 11076
rect 31536 11064 31542 11076
rect 35728 11073 35756 11104
rect 38197 11101 38209 11135
rect 38243 11101 38255 11135
rect 38197 11095 38255 11101
rect 39574 11092 39580 11144
rect 39632 11132 39638 11144
rect 40129 11135 40187 11141
rect 40129 11132 40141 11135
rect 39632 11104 40141 11132
rect 39632 11092 39638 11104
rect 40129 11101 40141 11104
rect 40175 11101 40187 11135
rect 40129 11095 40187 11101
rect 40218 11092 40224 11144
rect 40276 11132 40282 11144
rect 40773 11135 40831 11141
rect 40773 11132 40785 11135
rect 40276 11104 40785 11132
rect 40276 11092 40282 11104
rect 40773 11101 40785 11104
rect 40819 11101 40831 11135
rect 41386 11132 41414 11240
rect 42702 11160 42708 11212
rect 42760 11200 42766 11212
rect 42760 11172 47992 11200
rect 42760 11160 42766 11172
rect 47964 11141 47992 11172
rect 49142 11160 49148 11212
rect 49200 11160 49206 11212
rect 45649 11135 45707 11141
rect 45649 11132 45661 11135
rect 41386 11104 45661 11132
rect 40773 11095 40831 11101
rect 45649 11101 45661 11104
rect 45695 11101 45707 11135
rect 45649 11095 45707 11101
rect 47949 11135 48007 11141
rect 47949 11101 47961 11135
rect 47995 11101 48007 11135
rect 47949 11095 48007 11101
rect 34057 11067 34115 11073
rect 34057 11064 34069 11067
rect 31536 11036 31878 11064
rect 32784 11036 34069 11064
rect 31536 11024 31542 11036
rect 30101 10999 30159 11005
rect 30101 10965 30113 10999
rect 30147 10996 30159 10999
rect 30742 10996 30748 11008
rect 30147 10968 30748 10996
rect 30147 10965 30159 10968
rect 30101 10959 30159 10965
rect 30742 10956 30748 10968
rect 30800 10956 30806 11008
rect 30834 10956 30840 11008
rect 30892 10996 30898 11008
rect 32030 10996 32036 11008
rect 30892 10968 32036 10996
rect 30892 10956 30898 10968
rect 32030 10956 32036 10968
rect 32088 10956 32094 11008
rect 32122 10956 32128 11008
rect 32180 10996 32186 11008
rect 32784 10996 32812 11036
rect 34057 11033 34069 11036
rect 34103 11033 34115 11067
rect 34057 11027 34115 11033
rect 35713 11067 35771 11073
rect 35713 11033 35725 11067
rect 35759 11064 35771 11067
rect 35894 11064 35900 11076
rect 35759 11036 35900 11064
rect 35759 11033 35771 11036
rect 35713 11027 35771 11033
rect 35894 11024 35900 11036
rect 35952 11024 35958 11076
rect 37461 11067 37519 11073
rect 37461 11033 37473 11067
rect 37507 11064 37519 11067
rect 38378 11064 38384 11076
rect 37507 11036 38384 11064
rect 37507 11033 37519 11036
rect 37461 11027 37519 11033
rect 38378 11024 38384 11036
rect 38436 11024 38442 11076
rect 40313 11067 40371 11073
rect 40313 11033 40325 11067
rect 40359 11064 40371 11067
rect 45738 11064 45744 11076
rect 40359 11036 45744 11064
rect 40359 11033 40371 11036
rect 40313 11027 40371 11033
rect 45738 11024 45744 11036
rect 45796 11024 45802 11076
rect 45833 11067 45891 11073
rect 45833 11033 45845 11067
rect 45879 11064 45891 11067
rect 46934 11064 46940 11076
rect 45879 11036 46940 11064
rect 45879 11033 45891 11036
rect 45833 11027 45891 11033
rect 46934 11024 46940 11036
rect 46992 11024 46998 11076
rect 32180 10968 32812 10996
rect 32180 10956 32186 10968
rect 32950 10956 32956 11008
rect 33008 10996 33014 11008
rect 38930 10996 38936 11008
rect 33008 10968 38936 10996
rect 33008 10956 33014 10968
rect 38930 10956 38936 10968
rect 38988 10956 38994 11008
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 2498 10752 2504 10804
rect 2556 10752 2562 10804
rect 11330 10752 11336 10804
rect 11388 10792 11394 10804
rect 12437 10795 12495 10801
rect 12437 10792 12449 10795
rect 11388 10764 12449 10792
rect 11388 10752 11394 10764
rect 12437 10761 12449 10764
rect 12483 10761 12495 10795
rect 12437 10755 12495 10761
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 13173 10795 13231 10801
rect 13173 10792 13185 10795
rect 12860 10764 13185 10792
rect 12860 10752 12866 10764
rect 13173 10761 13185 10764
rect 13219 10761 13231 10795
rect 13173 10755 13231 10761
rect 14366 10752 14372 10804
rect 14424 10752 14430 10804
rect 15562 10752 15568 10804
rect 15620 10752 15626 10804
rect 15933 10795 15991 10801
rect 15933 10761 15945 10795
rect 15979 10792 15991 10795
rect 17129 10795 17187 10801
rect 17129 10792 17141 10795
rect 15979 10764 17141 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 17129 10761 17141 10764
rect 17175 10761 17187 10795
rect 17129 10755 17187 10761
rect 19521 10795 19579 10801
rect 19521 10761 19533 10795
rect 19567 10792 19579 10795
rect 19702 10792 19708 10804
rect 19567 10764 19708 10792
rect 19567 10761 19579 10764
rect 19521 10755 19579 10761
rect 19702 10752 19708 10764
rect 19760 10752 19766 10804
rect 21085 10795 21143 10801
rect 21085 10761 21097 10795
rect 21131 10792 21143 10795
rect 22646 10792 22652 10804
rect 21131 10764 22652 10792
rect 21131 10761 21143 10764
rect 21085 10755 21143 10761
rect 22646 10752 22652 10764
rect 22704 10752 22710 10804
rect 22922 10752 22928 10804
rect 22980 10792 22986 10804
rect 24213 10795 24271 10801
rect 24213 10792 24225 10795
rect 22980 10764 24225 10792
rect 22980 10752 22986 10764
rect 24213 10761 24225 10764
rect 24259 10761 24271 10795
rect 24213 10755 24271 10761
rect 25498 10752 25504 10804
rect 25556 10792 25562 10804
rect 25869 10795 25927 10801
rect 25869 10792 25881 10795
rect 25556 10764 25881 10792
rect 25556 10752 25562 10764
rect 25869 10761 25881 10764
rect 25915 10792 25927 10795
rect 26421 10795 26479 10801
rect 26421 10792 26433 10795
rect 25915 10764 26433 10792
rect 25915 10761 25927 10764
rect 25869 10755 25927 10761
rect 26421 10761 26433 10764
rect 26467 10792 26479 10795
rect 26694 10792 26700 10804
rect 26467 10764 26700 10792
rect 26467 10761 26479 10764
rect 26421 10755 26479 10761
rect 26694 10752 26700 10764
rect 26752 10752 26758 10804
rect 26789 10795 26847 10801
rect 26789 10761 26801 10795
rect 26835 10792 26847 10795
rect 27706 10792 27712 10804
rect 26835 10764 27712 10792
rect 26835 10761 26847 10764
rect 26789 10755 26847 10761
rect 27706 10752 27712 10764
rect 27764 10752 27770 10804
rect 28537 10795 28595 10801
rect 28537 10761 28549 10795
rect 28583 10792 28595 10795
rect 28583 10764 28948 10792
rect 28583 10761 28595 10764
rect 28537 10755 28595 10761
rect 1210 10684 1216 10736
rect 1268 10724 1274 10736
rect 14550 10724 14556 10736
rect 1268 10696 2360 10724
rect 1268 10684 1274 10696
rect 1302 10616 1308 10668
rect 1360 10656 1366 10668
rect 2332 10665 2360 10696
rect 6886 10696 14556 10724
rect 1581 10659 1639 10665
rect 1581 10656 1593 10659
rect 1360 10628 1593 10656
rect 1360 10616 1366 10628
rect 1581 10625 1593 10628
rect 1627 10625 1639 10659
rect 1581 10619 1639 10625
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 2363 10628 2881 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 2869 10625 2881 10628
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 1596 10588 1624 10619
rect 3053 10591 3111 10597
rect 3053 10588 3065 10591
rect 1596 10560 3065 10588
rect 3053 10557 3065 10560
rect 3099 10557 3111 10591
rect 3053 10551 3111 10557
rect 1765 10523 1823 10529
rect 1765 10489 1777 10523
rect 1811 10520 1823 10523
rect 6886 10520 6914 10696
rect 14550 10684 14556 10696
rect 14608 10684 14614 10736
rect 15746 10724 15752 10736
rect 14752 10696 15752 10724
rect 12250 10616 12256 10668
rect 12308 10656 12314 10668
rect 14752 10665 14780 10696
rect 15746 10684 15752 10696
rect 15804 10684 15810 10736
rect 15838 10684 15844 10736
rect 15896 10724 15902 10736
rect 17497 10727 17555 10733
rect 17497 10724 17509 10727
rect 15896 10696 17509 10724
rect 15896 10684 15902 10696
rect 17497 10693 17509 10696
rect 17543 10693 17555 10727
rect 19981 10727 20039 10733
rect 19981 10724 19993 10727
rect 17497 10687 17555 10693
rect 18616 10696 19993 10724
rect 13541 10659 13599 10665
rect 13541 10656 13553 10659
rect 12308 10628 13553 10656
rect 12308 10616 12314 10628
rect 13541 10625 13553 10628
rect 13587 10625 13599 10659
rect 14737 10659 14795 10665
rect 14737 10656 14749 10659
rect 13541 10619 13599 10625
rect 13740 10628 14749 10656
rect 12713 10591 12771 10597
rect 12713 10557 12725 10591
rect 12759 10588 12771 10591
rect 13446 10588 13452 10600
rect 12759 10560 13452 10588
rect 12759 10557 12771 10560
rect 12713 10551 12771 10557
rect 13446 10548 13452 10560
rect 13504 10588 13510 10600
rect 13633 10591 13691 10597
rect 13633 10588 13645 10591
rect 13504 10560 13645 10588
rect 13504 10548 13510 10560
rect 13633 10557 13645 10560
rect 13679 10557 13691 10591
rect 13633 10551 13691 10557
rect 13740 10520 13768 10628
rect 14737 10625 14749 10628
rect 14783 10625 14795 10659
rect 14737 10619 14795 10625
rect 14829 10659 14887 10665
rect 14829 10625 14841 10659
rect 14875 10656 14887 10659
rect 16758 10656 16764 10668
rect 14875 10628 16764 10656
rect 14875 10625 14887 10628
rect 14829 10619 14887 10625
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10656 16911 10659
rect 18616 10656 18644 10696
rect 19981 10693 19993 10696
rect 20027 10724 20039 10727
rect 20346 10724 20352 10736
rect 20027 10696 20352 10724
rect 20027 10693 20039 10696
rect 19981 10687 20039 10693
rect 20346 10684 20352 10696
rect 20404 10684 20410 10736
rect 21177 10727 21235 10733
rect 21177 10693 21189 10727
rect 21223 10724 21235 10727
rect 22278 10724 22284 10736
rect 21223 10696 22284 10724
rect 21223 10693 21235 10696
rect 21177 10687 21235 10693
rect 22278 10684 22284 10696
rect 22336 10684 22342 10736
rect 23934 10724 23940 10736
rect 23506 10696 23940 10724
rect 23934 10684 23940 10696
rect 23992 10724 23998 10736
rect 25516 10724 25544 10752
rect 27433 10727 27491 10733
rect 27433 10724 27445 10727
rect 23992 10696 25544 10724
rect 26068 10696 27445 10724
rect 23992 10684 23998 10696
rect 26068 10668 26096 10696
rect 27433 10693 27445 10696
rect 27479 10724 27491 10727
rect 27614 10724 27620 10736
rect 27479 10696 27620 10724
rect 27479 10693 27491 10696
rect 27433 10687 27491 10693
rect 27614 10684 27620 10696
rect 27672 10684 27678 10736
rect 16899 10628 18644 10656
rect 16899 10625 16911 10628
rect 16853 10619 16911 10625
rect 18690 10616 18696 10668
rect 18748 10616 18754 10668
rect 19889 10659 19947 10665
rect 18800 10628 19840 10656
rect 13814 10548 13820 10600
rect 13872 10548 13878 10600
rect 14918 10548 14924 10600
rect 14976 10548 14982 10600
rect 16022 10548 16028 10600
rect 16080 10548 16086 10600
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10557 16175 10591
rect 16117 10551 16175 10557
rect 1811 10492 6914 10520
rect 12820 10492 13768 10520
rect 1811 10489 1823 10492
rect 1765 10483 1823 10489
rect 12250 10412 12256 10464
rect 12308 10412 12314 10464
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 12820 10461 12848 10492
rect 13906 10480 13912 10532
rect 13964 10520 13970 10532
rect 16132 10520 16160 10551
rect 16666 10548 16672 10600
rect 16724 10588 16730 10600
rect 17589 10591 17647 10597
rect 17589 10588 17601 10591
rect 16724 10560 17601 10588
rect 16724 10548 16730 10560
rect 17589 10557 17601 10560
rect 17635 10557 17647 10591
rect 17589 10551 17647 10557
rect 17678 10548 17684 10600
rect 17736 10548 17742 10600
rect 18046 10548 18052 10600
rect 18104 10588 18110 10600
rect 18800 10597 18828 10628
rect 18785 10591 18843 10597
rect 18785 10588 18797 10591
rect 18104 10560 18797 10588
rect 18104 10548 18110 10560
rect 18785 10557 18797 10560
rect 18831 10557 18843 10591
rect 18785 10551 18843 10557
rect 18877 10591 18935 10597
rect 18877 10557 18889 10591
rect 18923 10557 18935 10591
rect 18877 10551 18935 10557
rect 13964 10492 16160 10520
rect 13964 10480 13970 10492
rect 16206 10480 16212 10532
rect 16264 10520 16270 10532
rect 16264 10492 18460 10520
rect 16264 10480 16270 10492
rect 12805 10455 12863 10461
rect 12805 10452 12817 10455
rect 12768 10424 12817 10452
rect 12768 10412 12774 10424
rect 12805 10421 12817 10424
rect 12851 10421 12863 10455
rect 12805 10415 12863 10421
rect 14734 10412 14740 10464
rect 14792 10452 14798 10464
rect 16574 10452 16580 10464
rect 14792 10424 16580 10452
rect 14792 10412 14798 10424
rect 16574 10412 16580 10424
rect 16632 10412 16638 10464
rect 17034 10412 17040 10464
rect 17092 10452 17098 10464
rect 18325 10455 18383 10461
rect 18325 10452 18337 10455
rect 17092 10424 18337 10452
rect 17092 10412 17098 10424
rect 18325 10421 18337 10424
rect 18371 10421 18383 10455
rect 18432 10452 18460 10492
rect 18506 10480 18512 10532
rect 18564 10520 18570 10532
rect 18892 10520 18920 10551
rect 18564 10492 18920 10520
rect 19812 10520 19840 10628
rect 19889 10625 19901 10659
rect 19935 10625 19947 10659
rect 19889 10619 19947 10625
rect 19904 10588 19932 10619
rect 20438 10616 20444 10668
rect 20496 10656 20502 10668
rect 24581 10659 24639 10665
rect 20496 10628 21496 10656
rect 20496 10616 20502 10628
rect 19978 10588 19984 10600
rect 19904 10560 19984 10588
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 20165 10591 20223 10597
rect 20165 10557 20177 10591
rect 20211 10588 20223 10591
rect 21082 10588 21088 10600
rect 20211 10560 21088 10588
rect 20211 10557 20223 10560
rect 20165 10551 20223 10557
rect 21082 10548 21088 10560
rect 21140 10548 21146 10600
rect 21361 10591 21419 10597
rect 21361 10557 21373 10591
rect 21407 10557 21419 10591
rect 21361 10551 21419 10557
rect 21266 10520 21272 10532
rect 19812 10492 21272 10520
rect 18564 10480 18570 10492
rect 21266 10480 21272 10492
rect 21324 10480 21330 10532
rect 20717 10455 20775 10461
rect 20717 10452 20729 10455
rect 18432 10424 20729 10452
rect 18325 10415 18383 10421
rect 20717 10421 20729 10424
rect 20763 10421 20775 10455
rect 21376 10452 21404 10551
rect 21468 10520 21496 10628
rect 24581 10625 24593 10659
rect 24627 10656 24639 10659
rect 25409 10659 25467 10665
rect 25409 10656 25421 10659
rect 24627 10628 25421 10656
rect 24627 10625 24639 10628
rect 24581 10619 24639 10625
rect 25409 10625 25421 10628
rect 25455 10625 25467 10659
rect 25409 10619 25467 10625
rect 26050 10616 26056 10668
rect 26108 10616 26114 10668
rect 27246 10616 27252 10668
rect 27304 10656 27310 10668
rect 27525 10659 27583 10665
rect 27525 10656 27537 10659
rect 27304 10628 27537 10656
rect 27304 10616 27310 10628
rect 27525 10625 27537 10628
rect 27571 10625 27583 10659
rect 27724 10656 27752 10752
rect 28810 10684 28816 10736
rect 28868 10724 28874 10736
rect 28920 10724 28948 10764
rect 31110 10752 31116 10804
rect 31168 10792 31174 10804
rect 31389 10795 31447 10801
rect 31389 10792 31401 10795
rect 31168 10764 31401 10792
rect 31168 10752 31174 10764
rect 31389 10761 31401 10764
rect 31435 10761 31447 10795
rect 32950 10792 32956 10804
rect 31389 10755 31447 10761
rect 31726 10764 32956 10792
rect 31726 10724 31754 10764
rect 32950 10752 32956 10764
rect 33008 10752 33014 10804
rect 33045 10795 33103 10801
rect 33045 10761 33057 10795
rect 33091 10792 33103 10795
rect 33091 10764 36768 10792
rect 33091 10761 33103 10764
rect 33045 10755 33103 10761
rect 28868 10696 28948 10724
rect 29012 10696 31754 10724
rect 28868 10684 28874 10696
rect 29012 10656 29040 10696
rect 32030 10684 32036 10736
rect 32088 10724 32094 10736
rect 32766 10724 32772 10736
rect 32088 10696 32772 10724
rect 32088 10684 32094 10696
rect 32766 10684 32772 10696
rect 32824 10724 32830 10736
rect 35345 10727 35403 10733
rect 32824 10696 33916 10724
rect 32824 10684 32830 10696
rect 27724 10628 29040 10656
rect 27525 10619 27583 10625
rect 29914 10616 29920 10668
rect 29972 10656 29978 10668
rect 30561 10659 30619 10665
rect 30561 10656 30573 10659
rect 29972 10628 30573 10656
rect 29972 10616 29978 10628
rect 30561 10625 30573 10628
rect 30607 10625 30619 10659
rect 32677 10659 32735 10665
rect 32677 10656 32689 10659
rect 30561 10619 30619 10625
rect 31864 10628 32689 10656
rect 22002 10548 22008 10600
rect 22060 10548 22066 10600
rect 22281 10591 22339 10597
rect 22281 10588 22293 10591
rect 22112 10560 22293 10588
rect 22112 10520 22140 10560
rect 22281 10557 22293 10560
rect 22327 10557 22339 10591
rect 22281 10551 22339 10557
rect 24118 10548 24124 10600
rect 24176 10588 24182 10600
rect 24670 10588 24676 10600
rect 24176 10560 24676 10588
rect 24176 10548 24182 10560
rect 24670 10548 24676 10560
rect 24728 10548 24734 10600
rect 24857 10591 24915 10597
rect 24857 10557 24869 10591
rect 24903 10588 24915 10591
rect 26602 10588 26608 10600
rect 24903 10560 26608 10588
rect 24903 10557 24915 10560
rect 24857 10551 24915 10557
rect 26602 10548 26608 10560
rect 26660 10548 26666 10600
rect 27341 10591 27399 10597
rect 27341 10557 27353 10591
rect 27387 10557 27399 10591
rect 27341 10551 27399 10557
rect 21468 10492 22140 10520
rect 23750 10480 23756 10532
rect 23808 10520 23814 10532
rect 24762 10520 24768 10532
rect 23808 10492 24768 10520
rect 23808 10480 23814 10492
rect 24762 10480 24768 10492
rect 24820 10480 24826 10532
rect 25774 10520 25780 10532
rect 24872 10492 25780 10520
rect 22094 10452 22100 10464
rect 21376 10424 22100 10452
rect 20717 10415 20775 10421
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 22370 10412 22376 10464
rect 22428 10452 22434 10464
rect 24872 10452 24900 10492
rect 25774 10480 25780 10492
rect 25832 10480 25838 10532
rect 26234 10480 26240 10532
rect 26292 10480 26298 10532
rect 22428 10424 24900 10452
rect 27356 10452 27384 10551
rect 29270 10548 29276 10600
rect 29328 10588 29334 10600
rect 29549 10591 29607 10597
rect 29549 10588 29561 10591
rect 29328 10560 29561 10588
rect 29328 10548 29334 10560
rect 29549 10557 29561 10560
rect 29595 10588 29607 10591
rect 29638 10588 29644 10600
rect 29595 10560 29644 10588
rect 29595 10557 29607 10560
rect 29549 10551 29607 10557
rect 29638 10548 29644 10560
rect 29696 10548 29702 10600
rect 29822 10548 29828 10600
rect 29880 10588 29886 10600
rect 30377 10591 30435 10597
rect 30377 10588 30389 10591
rect 29880 10560 30389 10588
rect 29880 10548 29886 10560
rect 30377 10557 30389 10560
rect 30423 10557 30435 10591
rect 30377 10551 30435 10557
rect 30466 10548 30472 10600
rect 30524 10548 30530 10600
rect 30650 10548 30656 10600
rect 30708 10588 30714 10600
rect 31864 10588 31892 10628
rect 32677 10625 32689 10628
rect 32723 10625 32735 10659
rect 32677 10619 32735 10625
rect 33318 10616 33324 10668
rect 33376 10616 33382 10668
rect 30708 10560 31892 10588
rect 30708 10548 30714 10560
rect 32398 10548 32404 10600
rect 32456 10548 32462 10600
rect 33888 10597 33916 10696
rect 35345 10693 35357 10727
rect 35391 10724 35403 10727
rect 36630 10724 36636 10736
rect 35391 10696 36636 10724
rect 35391 10693 35403 10696
rect 35345 10687 35403 10693
rect 36630 10684 36636 10696
rect 36688 10684 36694 10736
rect 36740 10724 36768 10764
rect 36814 10752 36820 10804
rect 36872 10752 36878 10804
rect 36906 10752 36912 10804
rect 36964 10792 36970 10804
rect 37277 10795 37335 10801
rect 37277 10792 37289 10795
rect 36964 10764 37289 10792
rect 36964 10752 36970 10764
rect 37277 10761 37289 10764
rect 37323 10792 37335 10795
rect 37461 10795 37519 10801
rect 37461 10792 37473 10795
rect 37323 10764 37473 10792
rect 37323 10761 37335 10764
rect 37277 10755 37335 10761
rect 37461 10761 37473 10764
rect 37507 10792 37519 10795
rect 38838 10792 38844 10804
rect 37507 10764 38844 10792
rect 37507 10761 37519 10764
rect 37461 10755 37519 10761
rect 38838 10752 38844 10764
rect 38896 10752 38902 10804
rect 37366 10724 37372 10736
rect 36740 10696 37372 10724
rect 37366 10684 37372 10696
rect 37424 10684 37430 10736
rect 49145 10727 49203 10733
rect 49145 10693 49157 10727
rect 49191 10724 49203 10727
rect 49234 10724 49240 10736
rect 49191 10696 49240 10724
rect 49191 10693 49203 10696
rect 49145 10687 49203 10693
rect 49234 10684 49240 10696
rect 49292 10684 49298 10736
rect 34238 10616 34244 10668
rect 34296 10616 34302 10668
rect 35618 10616 35624 10668
rect 35676 10616 35682 10668
rect 36446 10616 36452 10668
rect 36504 10616 36510 10668
rect 39761 10659 39819 10665
rect 39761 10625 39773 10659
rect 39807 10656 39819 10659
rect 40221 10659 40279 10665
rect 40221 10656 40233 10659
rect 39807 10628 40233 10656
rect 39807 10625 39819 10628
rect 39761 10619 39819 10625
rect 40221 10625 40233 10628
rect 40267 10625 40279 10659
rect 40221 10619 40279 10625
rect 32585 10591 32643 10597
rect 32585 10557 32597 10591
rect 32631 10557 32643 10591
rect 32585 10551 32643 10557
rect 33873 10591 33931 10597
rect 33873 10557 33885 10591
rect 33919 10557 33931 10591
rect 33873 10551 33931 10557
rect 27893 10523 27951 10529
rect 27893 10489 27905 10523
rect 27939 10520 27951 10523
rect 27939 10492 32168 10520
rect 27939 10489 27951 10492
rect 27893 10483 27951 10489
rect 30190 10452 30196 10464
rect 27356 10424 30196 10452
rect 22428 10412 22434 10424
rect 30190 10412 30196 10424
rect 30248 10452 30254 10464
rect 30834 10452 30840 10464
rect 30248 10424 30840 10452
rect 30248 10412 30254 10424
rect 30834 10412 30840 10424
rect 30892 10412 30898 10464
rect 30929 10455 30987 10461
rect 30929 10421 30941 10455
rect 30975 10452 30987 10455
rect 31754 10452 31760 10464
rect 30975 10424 31760 10452
rect 30975 10421 30987 10424
rect 30929 10415 30987 10421
rect 31754 10412 31760 10424
rect 31812 10412 31818 10464
rect 31846 10412 31852 10464
rect 31904 10452 31910 10464
rect 31941 10455 31999 10461
rect 31941 10452 31953 10455
rect 31904 10424 31953 10452
rect 31904 10412 31910 10424
rect 31941 10421 31953 10424
rect 31987 10452 31999 10455
rect 32030 10452 32036 10464
rect 31987 10424 32036 10452
rect 31987 10421 31999 10424
rect 31941 10415 31999 10421
rect 32030 10412 32036 10424
rect 32088 10412 32094 10464
rect 32140 10452 32168 10492
rect 32600 10452 32628 10551
rect 34698 10548 34704 10600
rect 34756 10588 34762 10600
rect 36173 10591 36231 10597
rect 36173 10588 36185 10591
rect 34756 10560 36185 10588
rect 34756 10548 34762 10560
rect 36173 10557 36185 10560
rect 36219 10557 36231 10591
rect 36173 10551 36231 10557
rect 36354 10548 36360 10600
rect 36412 10548 36418 10600
rect 39776 10588 39804 10619
rect 46934 10616 46940 10668
rect 46992 10656 46998 10668
rect 47949 10659 48007 10665
rect 47949 10656 47961 10659
rect 46992 10628 47961 10656
rect 46992 10616 46998 10628
rect 47949 10625 47961 10628
rect 47995 10625 48007 10659
rect 47949 10619 48007 10625
rect 36464 10560 39804 10588
rect 35618 10480 35624 10532
rect 35676 10520 35682 10532
rect 36464 10520 36492 10560
rect 35676 10492 36492 10520
rect 39945 10523 40003 10529
rect 35676 10480 35682 10492
rect 39945 10489 39957 10523
rect 39991 10520 40003 10523
rect 46934 10520 46940 10532
rect 39991 10492 46940 10520
rect 39991 10489 40003 10492
rect 39945 10483 40003 10489
rect 46934 10480 46940 10492
rect 46992 10480 46998 10532
rect 32140 10424 32628 10452
rect 33870 10412 33876 10464
rect 33928 10452 33934 10464
rect 34790 10452 34796 10464
rect 33928 10424 34796 10452
rect 33928 10412 33934 10424
rect 34790 10412 34796 10424
rect 34848 10412 34854 10464
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 13449 10251 13507 10257
rect 13449 10217 13461 10251
rect 13495 10248 13507 10251
rect 16022 10248 16028 10260
rect 13495 10220 16028 10248
rect 13495 10217 13507 10220
rect 13449 10211 13507 10217
rect 16022 10208 16028 10220
rect 16080 10208 16086 10260
rect 18046 10248 18052 10260
rect 16408 10220 18052 10248
rect 13909 10183 13967 10189
rect 13909 10149 13921 10183
rect 13955 10180 13967 10183
rect 14734 10180 14740 10192
rect 13955 10152 14740 10180
rect 13955 10149 13967 10152
rect 13909 10143 13967 10149
rect 14734 10140 14740 10152
rect 14792 10140 14798 10192
rect 2130 10072 2136 10124
rect 2188 10072 2194 10124
rect 12897 10115 12955 10121
rect 12897 10081 12909 10115
rect 12943 10081 12955 10115
rect 12897 10075 12955 10081
rect 12989 10115 13047 10121
rect 12989 10081 13001 10115
rect 13035 10112 13047 10115
rect 15102 10112 15108 10124
rect 13035 10084 15108 10112
rect 13035 10081 13047 10084
rect 12989 10075 13047 10081
rect 2406 10004 2412 10056
rect 2464 10004 2470 10056
rect 12912 10044 12940 10075
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 15194 10072 15200 10124
rect 15252 10112 15258 10124
rect 16408 10121 16436 10220
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 18141 10251 18199 10257
rect 18141 10217 18153 10251
rect 18187 10248 18199 10251
rect 18322 10248 18328 10260
rect 18187 10220 18328 10248
rect 18187 10217 18199 10220
rect 18141 10211 18199 10217
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 20257 10251 20315 10257
rect 20257 10217 20269 10251
rect 20303 10248 20315 10251
rect 20438 10248 20444 10260
rect 20303 10220 20444 10248
rect 20303 10217 20315 10220
rect 20257 10211 20315 10217
rect 20438 10208 20444 10220
rect 20496 10208 20502 10260
rect 21634 10248 21640 10260
rect 20548 10220 21640 10248
rect 16574 10140 16580 10192
rect 16632 10180 16638 10192
rect 17494 10180 17500 10192
rect 16632 10152 17500 10180
rect 16632 10140 16638 10152
rect 17494 10140 17500 10152
rect 17552 10140 17558 10192
rect 17862 10180 17868 10192
rect 17604 10152 17868 10180
rect 16393 10115 16451 10121
rect 16393 10112 16405 10115
rect 15252 10084 16405 10112
rect 15252 10072 15258 10084
rect 16393 10081 16405 10084
rect 16439 10081 16451 10115
rect 16393 10075 16451 10081
rect 17310 10072 17316 10124
rect 17368 10112 17374 10124
rect 17604 10121 17632 10152
rect 17862 10140 17868 10152
rect 17920 10180 17926 10192
rect 18506 10180 18512 10192
rect 17920 10152 18512 10180
rect 17920 10140 17926 10152
rect 18506 10140 18512 10152
rect 18564 10140 18570 10192
rect 19150 10180 19156 10192
rect 18616 10152 19156 10180
rect 17405 10115 17463 10121
rect 17405 10112 17417 10115
rect 17368 10084 17417 10112
rect 17368 10072 17374 10084
rect 17405 10081 17417 10084
rect 17451 10081 17463 10115
rect 17405 10075 17463 10081
rect 17589 10115 17647 10121
rect 17589 10081 17601 10115
rect 17635 10081 17647 10115
rect 17589 10075 17647 10081
rect 18414 10072 18420 10124
rect 18472 10112 18478 10124
rect 18616 10121 18644 10152
rect 19150 10140 19156 10152
rect 19208 10140 19214 10192
rect 18601 10115 18659 10121
rect 18601 10112 18613 10115
rect 18472 10084 18613 10112
rect 18472 10072 18478 10084
rect 18601 10081 18613 10084
rect 18647 10081 18659 10115
rect 18601 10075 18659 10081
rect 18785 10115 18843 10121
rect 18785 10081 18797 10115
rect 18831 10112 18843 10115
rect 19426 10112 19432 10124
rect 18831 10084 19432 10112
rect 18831 10081 18843 10084
rect 18785 10075 18843 10081
rect 19426 10072 19432 10084
rect 19484 10072 19490 10124
rect 19610 10072 19616 10124
rect 19668 10112 19674 10124
rect 19705 10115 19763 10121
rect 19705 10112 19717 10115
rect 19668 10084 19717 10112
rect 19668 10072 19674 10084
rect 19705 10081 19717 10084
rect 19751 10081 19763 10115
rect 19705 10075 19763 10081
rect 14458 10044 14464 10056
rect 12912 10016 14464 10044
rect 14458 10004 14464 10016
rect 14516 10004 14522 10056
rect 14642 10004 14648 10056
rect 14700 10004 14706 10056
rect 16022 10004 16028 10056
rect 16080 10004 16086 10056
rect 16666 10004 16672 10056
rect 16724 10044 16730 10056
rect 20548 10044 20576 10220
rect 21634 10208 21640 10220
rect 21692 10248 21698 10260
rect 22186 10248 22192 10260
rect 21692 10220 22192 10248
rect 21692 10208 21698 10220
rect 22186 10208 22192 10220
rect 22244 10208 22250 10260
rect 23753 10251 23811 10257
rect 23753 10217 23765 10251
rect 23799 10248 23811 10251
rect 24026 10248 24032 10260
rect 23799 10220 24032 10248
rect 23799 10217 23811 10220
rect 23753 10211 23811 10217
rect 24026 10208 24032 10220
rect 24084 10208 24090 10260
rect 24302 10208 24308 10260
rect 24360 10248 24366 10260
rect 24581 10251 24639 10257
rect 24581 10248 24593 10251
rect 24360 10220 24593 10248
rect 24360 10208 24366 10220
rect 24581 10217 24593 10220
rect 24627 10217 24639 10251
rect 24581 10211 24639 10217
rect 26694 10208 26700 10260
rect 26752 10208 26758 10260
rect 27614 10208 27620 10260
rect 27672 10248 27678 10260
rect 28721 10251 28779 10257
rect 27672 10220 28672 10248
rect 27672 10208 27678 10220
rect 23474 10140 23480 10192
rect 23532 10180 23538 10192
rect 23934 10180 23940 10192
rect 23532 10152 23940 10180
rect 23532 10140 23538 10152
rect 23934 10140 23940 10152
rect 23992 10140 23998 10192
rect 26602 10180 26608 10192
rect 26252 10152 26608 10180
rect 21082 10072 21088 10124
rect 21140 10112 21146 10124
rect 21729 10115 21787 10121
rect 21729 10112 21741 10115
rect 21140 10084 21741 10112
rect 21140 10072 21146 10084
rect 21729 10081 21741 10084
rect 21775 10081 21787 10115
rect 21729 10075 21787 10081
rect 26053 10115 26111 10121
rect 26053 10081 26065 10115
rect 26099 10112 26111 10115
rect 26252 10112 26280 10152
rect 26602 10140 26608 10152
rect 26660 10140 26666 10192
rect 28644 10180 28672 10220
rect 28721 10217 28733 10251
rect 28767 10248 28779 10251
rect 29086 10248 29092 10260
rect 28767 10220 29092 10248
rect 28767 10217 28779 10220
rect 28721 10211 28779 10217
rect 29086 10208 29092 10220
rect 29144 10248 29150 10260
rect 29822 10248 29828 10260
rect 29144 10220 29828 10248
rect 29144 10208 29150 10220
rect 29822 10208 29828 10220
rect 29880 10208 29886 10260
rect 30377 10251 30435 10257
rect 30377 10217 30389 10251
rect 30423 10248 30435 10251
rect 31386 10248 31392 10260
rect 30423 10220 31392 10248
rect 30423 10217 30435 10220
rect 30377 10211 30435 10217
rect 31386 10208 31392 10220
rect 31444 10208 31450 10260
rect 32858 10248 32864 10260
rect 32048 10220 32864 10248
rect 28644 10152 30788 10180
rect 26099 10084 26280 10112
rect 26329 10115 26387 10121
rect 26099 10081 26111 10084
rect 26053 10075 26111 10081
rect 26329 10081 26341 10115
rect 26375 10112 26387 10115
rect 26878 10112 26884 10124
rect 26375 10084 26884 10112
rect 26375 10081 26387 10084
rect 26329 10075 26387 10081
rect 26878 10072 26884 10084
rect 26936 10112 26942 10124
rect 26973 10115 27031 10121
rect 26973 10112 26985 10115
rect 26936 10084 26985 10112
rect 26936 10072 26942 10084
rect 26973 10081 26985 10084
rect 27019 10112 27031 10115
rect 29270 10112 29276 10124
rect 27019 10084 29276 10112
rect 27019 10081 27031 10084
rect 26973 10075 27031 10081
rect 29270 10072 29276 10084
rect 29328 10072 29334 10124
rect 29362 10072 29368 10124
rect 29420 10072 29426 10124
rect 29917 10115 29975 10121
rect 29917 10081 29929 10115
rect 29963 10112 29975 10115
rect 30650 10112 30656 10124
rect 29963 10084 30656 10112
rect 29963 10081 29975 10084
rect 29917 10075 29975 10081
rect 30650 10072 30656 10084
rect 30708 10072 30714 10124
rect 30760 10112 30788 10152
rect 32048 10112 32076 10220
rect 32858 10208 32864 10220
rect 32916 10248 32922 10260
rect 32916 10220 36400 10248
rect 32916 10208 32922 10220
rect 34422 10180 34428 10192
rect 32324 10152 34428 10180
rect 30760 10084 32076 10112
rect 32122 10072 32128 10124
rect 32180 10072 32186 10124
rect 16724 10016 20576 10044
rect 16724 10004 16730 10016
rect 20622 10004 20628 10056
rect 20680 10004 20686 10056
rect 22005 10047 22063 10053
rect 22005 10013 22017 10047
rect 22051 10044 22063 10047
rect 23293 10047 23351 10053
rect 23293 10044 23305 10047
rect 22051 10016 23305 10044
rect 22051 10013 22063 10016
rect 22005 10007 22063 10013
rect 15749 9979 15807 9985
rect 13096 9948 14504 9976
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 13096 9917 13124 9948
rect 13081 9911 13139 9917
rect 13081 9908 13093 9911
rect 12492 9880 13093 9908
rect 12492 9868 12498 9880
rect 13081 9877 13093 9880
rect 13127 9877 13139 9911
rect 13081 9871 13139 9877
rect 13906 9868 13912 9920
rect 13964 9908 13970 9920
rect 14277 9911 14335 9917
rect 14277 9908 14289 9911
rect 13964 9880 14289 9908
rect 13964 9868 13970 9880
rect 14277 9877 14289 9880
rect 14323 9877 14335 9911
rect 14476 9908 14504 9948
rect 15749 9945 15761 9979
rect 15795 9976 15807 9979
rect 17678 9976 17684 9988
rect 15795 9948 17684 9976
rect 15795 9945 15807 9948
rect 15749 9939 15807 9945
rect 15010 9908 15016 9920
rect 14476 9880 15016 9908
rect 14277 9871 14335 9877
rect 15010 9868 15016 9880
rect 15068 9868 15074 9920
rect 15102 9868 15108 9920
rect 15160 9908 15166 9920
rect 15764 9908 15792 9939
rect 17678 9936 17684 9948
rect 17736 9936 17742 9988
rect 19978 9976 19984 9988
rect 18432 9948 19984 9976
rect 15160 9880 15792 9908
rect 15160 9868 15166 9880
rect 16942 9868 16948 9920
rect 17000 9868 17006 9920
rect 17310 9868 17316 9920
rect 17368 9868 17374 9920
rect 17494 9868 17500 9920
rect 17552 9908 17558 9920
rect 18432 9908 18460 9948
rect 19978 9936 19984 9948
rect 20036 9936 20042 9988
rect 17552 9880 18460 9908
rect 17552 9868 17558 9880
rect 18506 9868 18512 9920
rect 18564 9908 18570 9920
rect 21358 9908 21364 9920
rect 18564 9880 21364 9908
rect 18564 9868 18570 9880
rect 21358 9868 21364 9880
rect 21416 9868 21422 9920
rect 21450 9868 21456 9920
rect 21508 9908 21514 9920
rect 22002 9908 22008 9920
rect 21508 9880 22008 9908
rect 21508 9868 21514 9880
rect 22002 9868 22008 9880
rect 22060 9908 22066 9920
rect 22112 9908 22140 10016
rect 23293 10013 23305 10016
rect 23339 10044 23351 10047
rect 24026 10044 24032 10056
rect 23339 10016 24032 10044
rect 23339 10013 23351 10016
rect 23293 10007 23351 10013
rect 24026 10004 24032 10016
rect 24084 10004 24090 10056
rect 22462 9936 22468 9988
rect 22520 9936 22526 9988
rect 25498 9936 25504 9988
rect 25556 9936 25562 9988
rect 27249 9979 27307 9985
rect 27249 9945 27261 9979
rect 27295 9976 27307 9979
rect 27338 9976 27344 9988
rect 27295 9948 27344 9976
rect 27295 9945 27307 9948
rect 27249 9939 27307 9945
rect 27338 9936 27344 9948
rect 27396 9936 27402 9988
rect 27706 9976 27712 9988
rect 27448 9948 27712 9976
rect 22060 9880 22140 9908
rect 22060 9868 22066 9880
rect 24118 9868 24124 9920
rect 24176 9868 24182 9920
rect 26694 9868 26700 9920
rect 26752 9908 26758 9920
rect 27448 9908 27476 9948
rect 27706 9936 27712 9948
rect 27764 9936 27770 9988
rect 29089 9979 29147 9985
rect 29089 9945 29101 9979
rect 29135 9976 29147 9979
rect 29178 9976 29184 9988
rect 29135 9948 29184 9976
rect 29135 9945 29147 9948
rect 29089 9939 29147 9945
rect 29178 9936 29184 9948
rect 29236 9976 29242 9988
rect 30374 9976 30380 9988
rect 29236 9948 30380 9976
rect 29236 9936 29242 9948
rect 30374 9936 30380 9948
rect 30432 9976 30438 9988
rect 30432 9948 30682 9976
rect 30432 9936 30438 9948
rect 31846 9936 31852 9988
rect 31904 9936 31910 9988
rect 26752 9880 27476 9908
rect 26752 9868 26758 9880
rect 29730 9868 29736 9920
rect 29788 9908 29794 9920
rect 32324 9908 32352 10152
rect 34422 10140 34428 10152
rect 34480 10140 34486 10192
rect 32766 10072 32772 10124
rect 32824 10072 32830 10124
rect 34698 10072 34704 10124
rect 34756 10112 34762 10124
rect 35158 10112 35164 10124
rect 34756 10084 35164 10112
rect 34756 10072 34762 10084
rect 35158 10072 35164 10084
rect 35216 10072 35222 10124
rect 32490 10004 32496 10056
rect 32548 10044 32554 10056
rect 32861 10047 32919 10053
rect 32861 10044 32873 10047
rect 32548 10016 32873 10044
rect 32548 10004 32554 10016
rect 32861 10013 32873 10016
rect 32907 10013 32919 10047
rect 32861 10007 32919 10013
rect 34882 10004 34888 10056
rect 34940 10004 34946 10056
rect 36372 10044 36400 10220
rect 36630 10208 36636 10260
rect 36688 10208 36694 10260
rect 36906 10208 36912 10260
rect 36964 10208 36970 10260
rect 38473 10115 38531 10121
rect 38473 10081 38485 10115
rect 38519 10112 38531 10115
rect 47026 10112 47032 10124
rect 38519 10084 47032 10112
rect 38519 10081 38531 10084
rect 38473 10075 38531 10081
rect 47026 10072 47032 10084
rect 47084 10072 47090 10124
rect 49142 10072 49148 10124
rect 49200 10072 49206 10124
rect 38289 10047 38347 10053
rect 38289 10044 38301 10047
rect 36372 10016 38301 10044
rect 38289 10013 38301 10016
rect 38335 10044 38347 10047
rect 38749 10047 38807 10053
rect 38749 10044 38761 10047
rect 38335 10016 38761 10044
rect 38335 10013 38347 10016
rect 38289 10007 38347 10013
rect 38749 10013 38761 10016
rect 38795 10013 38807 10047
rect 38749 10007 38807 10013
rect 38930 10004 38936 10056
rect 38988 10044 38994 10056
rect 40129 10047 40187 10053
rect 40129 10044 40141 10047
rect 38988 10016 40141 10044
rect 38988 10004 38994 10016
rect 40129 10013 40141 10016
rect 40175 10044 40187 10047
rect 40589 10047 40647 10053
rect 40589 10044 40601 10047
rect 40175 10016 40601 10044
rect 40175 10013 40187 10016
rect 40129 10007 40187 10013
rect 40589 10013 40601 10016
rect 40635 10013 40647 10047
rect 40589 10007 40647 10013
rect 44082 10004 44088 10056
rect 44140 10044 44146 10056
rect 44361 10047 44419 10053
rect 44361 10044 44373 10047
rect 44140 10016 44373 10044
rect 44140 10004 44146 10016
rect 44361 10013 44373 10016
rect 44407 10013 44419 10047
rect 44361 10007 44419 10013
rect 45738 10004 45744 10056
rect 45796 10044 45802 10056
rect 46109 10047 46167 10053
rect 46109 10044 46121 10047
rect 45796 10016 46121 10044
rect 45796 10004 45802 10016
rect 46109 10013 46121 10016
rect 46155 10013 46167 10047
rect 46109 10007 46167 10013
rect 46750 10004 46756 10056
rect 46808 10044 46814 10056
rect 47949 10047 48007 10053
rect 47949 10044 47961 10047
rect 46808 10016 47961 10044
rect 46808 10004 46814 10016
rect 47949 10013 47961 10016
rect 47995 10013 48007 10047
rect 47949 10007 48007 10013
rect 32674 9936 32680 9988
rect 32732 9976 32738 9988
rect 33781 9979 33839 9985
rect 33781 9976 33793 9979
rect 32732 9948 33793 9976
rect 32732 9936 32738 9948
rect 33781 9945 33793 9948
rect 33827 9945 33839 9979
rect 33781 9939 33839 9945
rect 34238 9936 34244 9988
rect 34296 9976 34302 9988
rect 35434 9976 35440 9988
rect 34296 9948 35440 9976
rect 34296 9936 34302 9948
rect 35434 9936 35440 9948
rect 35492 9936 35498 9988
rect 36906 9976 36912 9988
rect 36386 9948 36912 9976
rect 29788 9880 32352 9908
rect 29788 9868 29794 9880
rect 32398 9868 32404 9920
rect 32456 9908 32462 9920
rect 32953 9911 33011 9917
rect 32953 9908 32965 9911
rect 32456 9880 32965 9908
rect 32456 9868 32462 9880
rect 32953 9877 32965 9880
rect 32999 9877 33011 9911
rect 32953 9871 33011 9877
rect 33321 9911 33379 9917
rect 33321 9877 33333 9911
rect 33367 9908 33379 9911
rect 35802 9908 35808 9920
rect 33367 9880 35808 9908
rect 33367 9877 33379 9880
rect 33321 9871 33379 9877
rect 35802 9868 35808 9880
rect 35860 9868 35866 9920
rect 36078 9868 36084 9920
rect 36136 9908 36142 9920
rect 36464 9908 36492 9948
rect 36906 9936 36912 9948
rect 36964 9936 36970 9988
rect 40313 9979 40371 9985
rect 40313 9945 40325 9979
rect 40359 9976 40371 9979
rect 42702 9976 42708 9988
rect 40359 9948 42708 9976
rect 40359 9945 40371 9948
rect 40313 9939 40371 9945
rect 42702 9936 42708 9948
rect 42760 9936 42766 9988
rect 44545 9979 44603 9985
rect 44545 9945 44557 9979
rect 44591 9976 44603 9979
rect 46198 9976 46204 9988
rect 44591 9948 46204 9976
rect 44591 9945 44603 9948
rect 44545 9939 44603 9945
rect 46198 9936 46204 9948
rect 46256 9936 46262 9988
rect 47302 9936 47308 9988
rect 47360 9936 47366 9988
rect 36136 9880 36492 9908
rect 36136 9868 36142 9880
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 1302 9664 1308 9716
rect 1360 9704 1366 9716
rect 2133 9707 2191 9713
rect 2133 9704 2145 9707
rect 1360 9676 2145 9704
rect 1360 9664 1366 9676
rect 2133 9673 2145 9676
rect 2179 9704 2191 9707
rect 2406 9704 2412 9716
rect 2179 9676 2412 9704
rect 2179 9673 2191 9676
rect 2133 9667 2191 9673
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 14458 9664 14464 9716
rect 14516 9704 14522 9716
rect 15102 9704 15108 9716
rect 14516 9676 15108 9704
rect 14516 9664 14522 9676
rect 15102 9664 15108 9676
rect 15160 9664 15166 9716
rect 15746 9664 15752 9716
rect 15804 9704 15810 9716
rect 16482 9704 16488 9716
rect 15804 9676 16488 9704
rect 15804 9664 15810 9676
rect 13357 9639 13415 9645
rect 13357 9605 13369 9639
rect 13403 9636 13415 9639
rect 13722 9636 13728 9648
rect 13403 9608 13728 9636
rect 13403 9605 13415 9608
rect 13357 9599 13415 9605
rect 13722 9596 13728 9608
rect 13780 9596 13786 9648
rect 14642 9596 14648 9648
rect 14700 9636 14706 9648
rect 14826 9636 14832 9648
rect 14700 9608 14832 9636
rect 14700 9596 14706 9608
rect 14826 9596 14832 9608
rect 14884 9596 14890 9648
rect 15378 9596 15384 9648
rect 15436 9636 15442 9648
rect 16040 9645 16068 9676
rect 16482 9664 16488 9676
rect 16540 9664 16546 9716
rect 17218 9664 17224 9716
rect 17276 9704 17282 9716
rect 17276 9676 21036 9704
rect 17276 9664 17282 9676
rect 15841 9639 15899 9645
rect 15841 9636 15853 9639
rect 15436 9608 15853 9636
rect 15436 9596 15442 9608
rect 15841 9605 15853 9608
rect 15887 9605 15899 9639
rect 15841 9599 15899 9605
rect 16025 9639 16083 9645
rect 16025 9605 16037 9639
rect 16071 9605 16083 9639
rect 16025 9599 16083 9605
rect 16301 9639 16359 9645
rect 16301 9605 16313 9639
rect 16347 9636 16359 9639
rect 16666 9636 16672 9648
rect 16347 9608 16672 9636
rect 16347 9605 16359 9608
rect 16301 9599 16359 9605
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 18322 9636 18328 9648
rect 18170 9608 18328 9636
rect 18322 9596 18328 9608
rect 18380 9596 18386 9648
rect 19518 9596 19524 9648
rect 19576 9636 19582 9648
rect 19613 9639 19671 9645
rect 19613 9636 19625 9639
rect 19576 9608 19625 9636
rect 19576 9596 19582 9608
rect 19613 9605 19625 9608
rect 19659 9605 19671 9639
rect 21008 9636 21036 9676
rect 21082 9664 21088 9716
rect 21140 9664 21146 9716
rect 21192 9676 22232 9704
rect 21192 9636 21220 9676
rect 21008 9608 21220 9636
rect 19613 9599 19671 9605
rect 21266 9596 21272 9648
rect 21324 9636 21330 9648
rect 21361 9639 21419 9645
rect 21361 9636 21373 9639
rect 21324 9608 21373 9636
rect 21324 9596 21330 9608
rect 21361 9605 21373 9608
rect 21407 9605 21419 9639
rect 22204 9636 22232 9676
rect 22278 9664 22284 9716
rect 22336 9664 22342 9716
rect 26050 9704 26056 9716
rect 22388 9676 26056 9704
rect 22388 9636 22416 9676
rect 26050 9664 26056 9676
rect 26108 9664 26114 9716
rect 31754 9664 31760 9716
rect 31812 9704 31818 9716
rect 32953 9707 33011 9713
rect 32953 9704 32965 9707
rect 31812 9676 32965 9704
rect 31812 9664 31818 9676
rect 32953 9673 32965 9676
rect 32999 9673 33011 9707
rect 34882 9704 34888 9716
rect 32953 9667 33011 9673
rect 34532 9676 34888 9704
rect 22204 9608 22416 9636
rect 21361 9599 21419 9605
rect 1302 9528 1308 9580
rect 1360 9568 1366 9580
rect 1581 9571 1639 9577
rect 1581 9568 1593 9571
rect 1360 9540 1593 9568
rect 1360 9528 1366 9540
rect 1581 9537 1593 9540
rect 1627 9568 1639 9571
rect 2317 9571 2375 9577
rect 2317 9568 2329 9571
rect 1627 9540 2329 9568
rect 1627 9537 1639 9540
rect 1581 9531 1639 9537
rect 2317 9537 2329 9540
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 12342 9528 12348 9580
rect 12400 9568 12406 9580
rect 12529 9571 12587 9577
rect 12529 9568 12541 9571
rect 12400 9540 12541 9568
rect 12400 9528 12406 9540
rect 12529 9537 12541 9540
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 20622 9528 20628 9580
rect 20680 9568 20686 9580
rect 20680 9554 20746 9568
rect 20680 9540 20760 9554
rect 20680 9528 20686 9540
rect 11054 9460 11060 9512
rect 11112 9500 11118 9512
rect 12253 9503 12311 9509
rect 12253 9500 12265 9503
rect 11112 9472 12265 9500
rect 11112 9460 11118 9472
rect 12253 9469 12265 9472
rect 12299 9469 12311 9503
rect 12253 9463 12311 9469
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 1762 9392 1768 9444
rect 1820 9392 1826 9444
rect 12452 9432 12480 9463
rect 15102 9460 15108 9512
rect 15160 9460 15166 9512
rect 15381 9503 15439 9509
rect 15381 9469 15393 9503
rect 15427 9500 15439 9503
rect 16022 9500 16028 9512
rect 15427 9472 16028 9500
rect 15427 9469 15439 9472
rect 15381 9463 15439 9469
rect 12526 9432 12532 9444
rect 12452 9404 12532 9432
rect 12526 9392 12532 9404
rect 12584 9392 12590 9444
rect 12897 9435 12955 9441
rect 12897 9401 12909 9435
rect 12943 9432 12955 9435
rect 14090 9432 14096 9444
rect 12943 9404 14096 9432
rect 12943 9401 12955 9404
rect 12897 9395 12955 9401
rect 14090 9392 14096 9404
rect 14148 9392 14154 9444
rect 13630 9324 13636 9376
rect 13688 9364 13694 9376
rect 15396 9364 15424 9463
rect 16022 9460 16028 9472
rect 16080 9460 16086 9512
rect 16853 9503 16911 9509
rect 16853 9469 16865 9503
rect 16899 9500 16911 9503
rect 17586 9500 17592 9512
rect 16899 9472 17592 9500
rect 16899 9469 16911 9472
rect 16853 9463 16911 9469
rect 17586 9460 17592 9472
rect 17644 9460 17650 9512
rect 18598 9460 18604 9512
rect 18656 9460 18662 9512
rect 18874 9460 18880 9512
rect 18932 9500 18938 9512
rect 19337 9503 19395 9509
rect 19337 9500 19349 9503
rect 18932 9472 19349 9500
rect 18932 9460 18938 9472
rect 19337 9469 19349 9472
rect 19383 9469 19395 9503
rect 19337 9463 19395 9469
rect 17310 9432 17316 9444
rect 15672 9404 17316 9432
rect 15672 9376 15700 9404
rect 17310 9392 17316 9404
rect 17368 9392 17374 9444
rect 20732 9432 20760 9540
rect 21376 9500 21404 9599
rect 23474 9596 23480 9648
rect 23532 9636 23538 9648
rect 23532 9608 23782 9636
rect 23532 9596 23538 9608
rect 24670 9596 24676 9648
rect 24728 9636 24734 9648
rect 27338 9636 27344 9648
rect 24728 9608 25268 9636
rect 24728 9596 24734 9608
rect 22646 9528 22652 9580
rect 22704 9528 22710 9580
rect 25240 9577 25268 9608
rect 25884 9608 27344 9636
rect 22741 9571 22799 9577
rect 22741 9537 22753 9571
rect 22787 9568 22799 9571
rect 25225 9571 25283 9577
rect 22787 9540 23612 9568
rect 22787 9537 22799 9540
rect 22741 9531 22799 9537
rect 22756 9500 22784 9531
rect 21376 9472 22784 9500
rect 22925 9503 22983 9509
rect 22925 9469 22937 9503
rect 22971 9500 22983 9503
rect 22971 9472 23520 9500
rect 22971 9469 22983 9472
rect 22925 9463 22983 9469
rect 21637 9435 21695 9441
rect 21637 9432 21649 9435
rect 20732 9404 21649 9432
rect 21637 9401 21649 9404
rect 21683 9432 21695 9435
rect 22002 9432 22008 9444
rect 21683 9404 22008 9432
rect 21683 9401 21695 9404
rect 21637 9395 21695 9401
rect 22002 9392 22008 9404
rect 22060 9392 22066 9444
rect 13688 9336 15424 9364
rect 13688 9324 13694 9336
rect 15654 9324 15660 9376
rect 15712 9324 15718 9376
rect 16206 9324 16212 9376
rect 16264 9364 16270 9376
rect 16393 9367 16451 9373
rect 16393 9364 16405 9367
rect 16264 9336 16405 9364
rect 16264 9324 16270 9336
rect 16393 9333 16405 9336
rect 16439 9333 16451 9367
rect 16393 9327 16451 9333
rect 16482 9324 16488 9376
rect 16540 9364 16546 9376
rect 18506 9364 18512 9376
rect 16540 9336 18512 9364
rect 16540 9324 16546 9336
rect 18506 9324 18512 9336
rect 18564 9324 18570 9376
rect 21542 9324 21548 9376
rect 21600 9364 21606 9376
rect 21818 9364 21824 9376
rect 21600 9336 21824 9364
rect 21600 9324 21606 9336
rect 21818 9324 21824 9336
rect 21876 9324 21882 9376
rect 23492 9373 23520 9472
rect 23584 9432 23612 9540
rect 25225 9537 25237 9571
rect 25271 9537 25283 9571
rect 25225 9531 25283 9537
rect 24302 9460 24308 9512
rect 24360 9500 24366 9512
rect 25884 9509 25912 9608
rect 27338 9596 27344 9608
rect 27396 9596 27402 9648
rect 27706 9596 27712 9648
rect 27764 9636 27770 9648
rect 28997 9639 29055 9645
rect 27764 9608 27830 9636
rect 27764 9596 27770 9608
rect 28997 9605 29009 9639
rect 29043 9636 29055 9639
rect 30098 9636 30104 9648
rect 29043 9608 30104 9636
rect 29043 9605 29055 9608
rect 28997 9599 29055 9605
rect 30098 9596 30104 9608
rect 30156 9596 30162 9648
rect 30650 9596 30656 9648
rect 30708 9596 30714 9648
rect 31849 9639 31907 9645
rect 31849 9605 31861 9639
rect 31895 9636 31907 9639
rect 31938 9636 31944 9648
rect 31895 9608 31944 9636
rect 31895 9605 31907 9608
rect 31849 9599 31907 9605
rect 31938 9596 31944 9608
rect 31996 9596 32002 9648
rect 32122 9596 32128 9648
rect 32180 9636 32186 9648
rect 32490 9636 32496 9648
rect 32180 9608 32496 9636
rect 32180 9596 32186 9608
rect 32490 9596 32496 9608
rect 32548 9636 32554 9648
rect 34532 9636 34560 9676
rect 34882 9664 34888 9676
rect 34940 9664 34946 9716
rect 35158 9664 35164 9716
rect 35216 9704 35222 9716
rect 35621 9707 35679 9713
rect 35621 9704 35633 9707
rect 35216 9676 35633 9704
rect 35216 9664 35222 9676
rect 35621 9673 35633 9676
rect 35667 9673 35679 9707
rect 35621 9667 35679 9673
rect 36078 9664 36084 9716
rect 36136 9704 36142 9716
rect 36136 9676 36216 9704
rect 36136 9664 36142 9676
rect 35986 9636 35992 9648
rect 32548 9608 34560 9636
rect 35374 9608 35992 9636
rect 32548 9596 32554 9608
rect 26053 9571 26111 9577
rect 26053 9537 26065 9571
rect 26099 9537 26111 9571
rect 26053 9531 26111 9537
rect 24949 9503 25007 9509
rect 24949 9500 24961 9503
rect 24360 9472 24961 9500
rect 24360 9460 24366 9472
rect 24949 9469 24961 9472
rect 24995 9469 25007 9503
rect 24949 9463 25007 9469
rect 25869 9503 25927 9509
rect 25869 9469 25881 9503
rect 25915 9469 25927 9503
rect 25869 9463 25927 9469
rect 25958 9460 25964 9512
rect 26016 9460 26022 9512
rect 23584 9404 23888 9432
rect 23477 9367 23535 9373
rect 23477 9333 23489 9367
rect 23523 9364 23535 9367
rect 23750 9364 23756 9376
rect 23523 9336 23756 9364
rect 23523 9333 23535 9336
rect 23477 9327 23535 9333
rect 23750 9324 23756 9336
rect 23808 9324 23814 9376
rect 23860 9364 23888 9404
rect 25682 9392 25688 9444
rect 25740 9432 25746 9444
rect 26068 9432 26096 9531
rect 31662 9528 31668 9580
rect 31720 9568 31726 9580
rect 33888 9577 33916 9608
rect 35986 9596 35992 9608
rect 36044 9636 36050 9648
rect 36188 9636 36216 9676
rect 36044 9608 36216 9636
rect 49145 9639 49203 9645
rect 36044 9596 36050 9608
rect 49145 9605 49157 9639
rect 49191 9636 49203 9639
rect 49234 9636 49240 9648
rect 49191 9608 49240 9636
rect 49191 9605 49203 9608
rect 49145 9599 49203 9605
rect 49234 9596 49240 9608
rect 49292 9596 49298 9648
rect 32861 9571 32919 9577
rect 32861 9568 32873 9571
rect 31720 9540 32873 9568
rect 31720 9528 31726 9540
rect 32861 9537 32873 9540
rect 32907 9537 32919 9571
rect 32861 9531 32919 9537
rect 33873 9571 33931 9577
rect 33873 9537 33885 9571
rect 33919 9537 33931 9571
rect 33873 9531 33931 9537
rect 47118 9528 47124 9580
rect 47176 9568 47182 9580
rect 47949 9571 48007 9577
rect 47949 9568 47961 9571
rect 47176 9540 47961 9568
rect 47176 9528 47182 9540
rect 47949 9537 47961 9540
rect 47995 9537 48007 9571
rect 47949 9531 48007 9537
rect 26436 9472 29224 9500
rect 26436 9441 26464 9472
rect 25740 9404 26096 9432
rect 26421 9435 26479 9441
rect 25740 9392 25746 9404
rect 26421 9401 26433 9435
rect 26467 9401 26479 9435
rect 26421 9395 26479 9401
rect 27154 9392 27160 9444
rect 27212 9432 27218 9444
rect 27525 9435 27583 9441
rect 27525 9432 27537 9435
rect 27212 9404 27537 9432
rect 27212 9392 27218 9404
rect 27525 9401 27537 9404
rect 27571 9401 27583 9435
rect 29196 9432 29224 9472
rect 29270 9460 29276 9512
rect 29328 9500 29334 9512
rect 29733 9503 29791 9509
rect 29733 9500 29745 9503
rect 29328 9472 29745 9500
rect 29328 9460 29334 9472
rect 29733 9469 29745 9472
rect 29779 9469 29791 9503
rect 29733 9463 29791 9469
rect 30006 9460 30012 9512
rect 30064 9460 30070 9512
rect 30098 9460 30104 9512
rect 30156 9500 30162 9512
rect 31481 9503 31539 9509
rect 31481 9500 31493 9503
rect 30156 9472 31493 9500
rect 30156 9460 30162 9472
rect 31481 9469 31493 9472
rect 31527 9469 31539 9503
rect 31481 9463 31539 9469
rect 31496 9432 31524 9463
rect 31570 9460 31576 9512
rect 31628 9500 31634 9512
rect 31754 9500 31760 9512
rect 31628 9472 31760 9500
rect 31628 9460 31634 9472
rect 31754 9460 31760 9472
rect 31812 9460 31818 9512
rect 31938 9460 31944 9512
rect 31996 9500 32002 9512
rect 32677 9503 32735 9509
rect 32677 9500 32689 9503
rect 31996 9472 32689 9500
rect 31996 9460 32002 9472
rect 32677 9469 32689 9472
rect 32723 9469 32735 9503
rect 32677 9463 32735 9469
rect 34146 9460 34152 9512
rect 34204 9500 34210 9512
rect 35894 9500 35900 9512
rect 34204 9472 35900 9500
rect 34204 9460 34210 9472
rect 35894 9460 35900 9472
rect 35952 9460 35958 9512
rect 32766 9432 32772 9444
rect 29196 9404 29500 9432
rect 31496 9404 32772 9432
rect 27525 9395 27583 9401
rect 25406 9364 25412 9376
rect 23860 9336 25412 9364
rect 25406 9324 25412 9336
rect 25464 9324 25470 9376
rect 29472 9364 29500 9404
rect 32766 9392 32772 9404
rect 32824 9392 32830 9444
rect 30466 9364 30472 9376
rect 29472 9336 30472 9364
rect 30466 9324 30472 9336
rect 30524 9324 30530 9376
rect 30650 9324 30656 9376
rect 30708 9364 30714 9376
rect 31570 9364 31576 9376
rect 30708 9336 31576 9364
rect 30708 9324 30714 9336
rect 31570 9324 31576 9336
rect 31628 9324 31634 9376
rect 31754 9324 31760 9376
rect 31812 9364 31818 9376
rect 32217 9367 32275 9373
rect 32217 9364 32229 9367
rect 31812 9336 32229 9364
rect 31812 9324 31818 9336
rect 32217 9333 32229 9336
rect 32263 9364 32275 9367
rect 32858 9364 32864 9376
rect 32263 9336 32864 9364
rect 32263 9333 32275 9336
rect 32217 9327 32275 9333
rect 32858 9324 32864 9336
rect 32916 9324 32922 9376
rect 33321 9367 33379 9373
rect 33321 9333 33333 9367
rect 33367 9364 33379 9367
rect 35526 9364 35532 9376
rect 33367 9336 35532 9364
rect 33367 9333 33379 9336
rect 33321 9327 33379 9333
rect 35526 9324 35532 9336
rect 35584 9324 35590 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 17218 9160 17224 9172
rect 6886 9132 17224 9160
rect 1857 9095 1915 9101
rect 1857 9061 1869 9095
rect 1903 9092 1915 9095
rect 6886 9092 6914 9132
rect 17218 9120 17224 9132
rect 17276 9120 17282 9172
rect 17862 9120 17868 9172
rect 17920 9169 17926 9172
rect 17920 9163 17935 9169
rect 17923 9129 17935 9163
rect 17920 9123 17935 9129
rect 19429 9163 19487 9169
rect 19429 9129 19441 9163
rect 19475 9160 19487 9163
rect 19518 9160 19524 9172
rect 19475 9132 19524 9160
rect 19475 9129 19487 9132
rect 19429 9123 19487 9129
rect 17920 9120 17926 9123
rect 19518 9120 19524 9132
rect 19576 9120 19582 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 22281 9163 22339 9169
rect 22281 9160 22293 9163
rect 22152 9132 22293 9160
rect 22152 9120 22158 9132
rect 22281 9129 22293 9132
rect 22327 9129 22339 9163
rect 22281 9123 22339 9129
rect 22462 9120 22468 9172
rect 22520 9160 22526 9172
rect 24397 9163 24455 9169
rect 24397 9160 24409 9163
rect 22520 9132 24409 9160
rect 22520 9120 22526 9132
rect 24397 9129 24409 9132
rect 24443 9129 24455 9163
rect 24397 9123 24455 9129
rect 28905 9163 28963 9169
rect 28905 9129 28917 9163
rect 28951 9160 28963 9163
rect 32398 9160 32404 9172
rect 28951 9132 32404 9160
rect 28951 9129 28963 9132
rect 28905 9123 28963 9129
rect 32398 9120 32404 9132
rect 32456 9120 32462 9172
rect 34057 9163 34115 9169
rect 34057 9129 34069 9163
rect 34103 9160 34115 9163
rect 36354 9160 36360 9172
rect 34103 9132 36360 9160
rect 34103 9129 34115 9132
rect 34057 9123 34115 9129
rect 36354 9120 36360 9132
rect 36412 9120 36418 9172
rect 36725 9163 36783 9169
rect 36725 9129 36737 9163
rect 36771 9160 36783 9163
rect 43714 9160 43720 9172
rect 36771 9132 43720 9160
rect 36771 9129 36783 9132
rect 36725 9123 36783 9129
rect 43714 9120 43720 9132
rect 43772 9120 43778 9172
rect 1903 9064 6914 9092
rect 14461 9095 14519 9101
rect 1903 9061 1915 9064
rect 1857 9055 1915 9061
rect 14461 9061 14473 9095
rect 14507 9092 14519 9095
rect 16850 9092 16856 9104
rect 14507 9064 16856 9092
rect 14507 9061 14519 9064
rect 14461 9055 14519 9061
rect 16850 9052 16856 9064
rect 16908 9052 16914 9104
rect 30006 9092 30012 9104
rect 28368 9064 30012 9092
rect 2869 9027 2927 9033
rect 2869 9024 2881 9027
rect 2332 8996 2881 9024
rect 1210 8916 1216 8968
rect 1268 8956 1274 8968
rect 2332 8965 2360 8996
rect 2869 8993 2881 8996
rect 2915 8993 2927 9027
rect 2869 8987 2927 8993
rect 15102 8984 15108 9036
rect 15160 9024 15166 9036
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 15160 8996 15301 9024
rect 15160 8984 15166 8996
rect 15289 8993 15301 8996
rect 15335 8993 15347 9027
rect 15289 8987 15347 8993
rect 15470 8984 15476 9036
rect 15528 8984 15534 9036
rect 16022 8984 16028 9036
rect 16080 9024 16086 9036
rect 18141 9027 18199 9033
rect 18141 9024 18153 9027
rect 16080 8996 18153 9024
rect 16080 8984 16086 8996
rect 18141 8993 18153 8996
rect 18187 9024 18199 9027
rect 18874 9024 18880 9036
rect 18187 8996 18880 9024
rect 18187 8993 18199 8996
rect 18141 8987 18199 8993
rect 18874 8984 18880 8996
rect 18932 8984 18938 9036
rect 19426 8984 19432 9036
rect 19484 9024 19490 9036
rect 20901 9027 20959 9033
rect 20901 9024 20913 9027
rect 19484 8996 20913 9024
rect 19484 8984 19490 8996
rect 20901 8993 20913 8996
rect 20947 8993 20959 9027
rect 23382 9024 23388 9036
rect 20901 8987 20959 8993
rect 22664 8996 23388 9024
rect 2317 8959 2375 8965
rect 2317 8956 2329 8959
rect 1268 8928 2329 8956
rect 1268 8916 1274 8928
rect 2317 8925 2329 8928
rect 2363 8925 2375 8959
rect 3053 8959 3111 8965
rect 3053 8956 3065 8959
rect 2317 8919 2375 8925
rect 2424 8928 3065 8956
rect 1302 8848 1308 8900
rect 1360 8888 1366 8900
rect 1673 8891 1731 8897
rect 1673 8888 1685 8891
rect 1360 8860 1685 8888
rect 1360 8848 1366 8860
rect 1673 8857 1685 8860
rect 1719 8888 1731 8891
rect 2424 8888 2452 8928
rect 3053 8925 3065 8928
rect 3099 8925 3111 8959
rect 3053 8919 3111 8925
rect 11974 8916 11980 8968
rect 12032 8956 12038 8968
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 12032 8928 14289 8956
rect 12032 8916 12038 8928
rect 14277 8925 14289 8928
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 15562 8916 15568 8968
rect 15620 8916 15626 8968
rect 18690 8916 18696 8968
rect 18748 8916 18754 8968
rect 21177 8959 21235 8965
rect 21177 8925 21189 8959
rect 21223 8956 21235 8959
rect 21450 8956 21456 8968
rect 21223 8928 21456 8956
rect 21223 8925 21235 8928
rect 21177 8919 21235 8925
rect 21450 8916 21456 8928
rect 21508 8916 21514 8968
rect 22002 8916 22008 8968
rect 22060 8956 22066 8968
rect 22664 8956 22692 8996
rect 23382 8984 23388 8996
rect 23440 8984 23446 9036
rect 23750 8984 23756 9036
rect 23808 8984 23814 9036
rect 28368 9033 28396 9064
rect 30006 9052 30012 9064
rect 30064 9092 30070 9104
rect 30745 9095 30803 9101
rect 30745 9092 30757 9095
rect 30064 9064 30757 9092
rect 30064 9052 30070 9064
rect 30745 9061 30757 9064
rect 30791 9061 30803 9095
rect 33870 9092 33876 9104
rect 30745 9055 30803 9061
rect 32416 9064 33876 9092
rect 28353 9027 28411 9033
rect 28353 8993 28365 9027
rect 28399 8993 28411 9027
rect 28353 8987 28411 8993
rect 28442 8984 28448 9036
rect 28500 9024 28506 9036
rect 31754 9024 31760 9036
rect 28500 8996 31760 9024
rect 28500 8984 28506 8996
rect 31754 8984 31760 8996
rect 31812 8984 31818 9036
rect 32217 9027 32275 9033
rect 32217 8993 32229 9027
rect 32263 9024 32275 9027
rect 32416 9024 32444 9064
rect 33870 9052 33876 9064
rect 33928 9052 33934 9104
rect 34238 9052 34244 9104
rect 34296 9092 34302 9104
rect 34333 9095 34391 9101
rect 34333 9092 34345 9095
rect 34296 9064 34345 9092
rect 34296 9052 34302 9064
rect 34333 9061 34345 9064
rect 34379 9061 34391 9095
rect 34333 9055 34391 9061
rect 36262 9052 36268 9104
rect 36320 9092 36326 9104
rect 37829 9095 37887 9101
rect 36320 9064 37780 9092
rect 36320 9052 36326 9064
rect 32263 8996 32444 9024
rect 32263 8993 32275 8996
rect 32217 8987 32275 8993
rect 32490 8984 32496 9036
rect 32548 8984 32554 9036
rect 33042 8984 33048 9036
rect 33100 9024 33106 9036
rect 33413 9027 33471 9033
rect 33413 9024 33425 9027
rect 33100 8996 33425 9024
rect 33100 8984 33106 8996
rect 33413 8993 33425 8996
rect 33459 9024 33471 9027
rect 34146 9024 34152 9036
rect 33459 8996 34152 9024
rect 33459 8993 33471 8996
rect 33413 8987 33471 8993
rect 34146 8984 34152 8996
rect 34204 8984 34210 9036
rect 34974 8984 34980 9036
rect 35032 8984 35038 9036
rect 35066 8984 35072 9036
rect 35124 9024 35130 9036
rect 35124 8996 35296 9024
rect 35124 8984 35130 8996
rect 22060 8942 22692 8956
rect 22060 8928 22678 8942
rect 22060 8916 22066 8928
rect 24026 8916 24032 8968
rect 24084 8916 24090 8968
rect 25593 8959 25651 8965
rect 25593 8925 25605 8959
rect 25639 8956 25651 8959
rect 25958 8956 25964 8968
rect 25639 8928 25964 8956
rect 25639 8925 25651 8928
rect 25593 8919 25651 8925
rect 16114 8888 16120 8900
rect 1719 8860 2452 8888
rect 2516 8860 16120 8888
rect 1719 8857 1731 8860
rect 1673 8851 1731 8857
rect 2516 8829 2544 8860
rect 16114 8848 16120 8860
rect 16172 8848 16178 8900
rect 16206 8848 16212 8900
rect 16264 8888 16270 8900
rect 16264 8860 16620 8888
rect 16264 8848 16270 8860
rect 2501 8823 2559 8829
rect 2501 8789 2513 8823
rect 2547 8789 2559 8823
rect 2501 8783 2559 8789
rect 14918 8780 14924 8832
rect 14976 8780 14982 8832
rect 15930 8780 15936 8832
rect 15988 8780 15994 8832
rect 16390 8780 16396 8832
rect 16448 8780 16454 8832
rect 16592 8820 16620 8860
rect 17402 8848 17408 8900
rect 17460 8888 17466 8900
rect 18322 8888 18328 8900
rect 17460 8860 18328 8888
rect 17460 8848 17466 8860
rect 18322 8848 18328 8860
rect 18380 8848 18386 8900
rect 20438 8848 20444 8900
rect 20496 8848 20502 8900
rect 25608 8888 25636 8919
rect 25958 8916 25964 8928
rect 26016 8956 26022 8968
rect 30834 8956 30840 8968
rect 26016 8928 30840 8956
rect 26016 8916 26022 8928
rect 30834 8916 30840 8928
rect 30892 8916 30898 8968
rect 34790 8916 34796 8968
rect 34848 8956 34854 8968
rect 35161 8959 35219 8965
rect 35161 8956 35173 8959
rect 34848 8928 35173 8956
rect 34848 8916 34854 8928
rect 35161 8925 35173 8928
rect 35207 8925 35219 8959
rect 35268 8956 35296 8996
rect 35526 8984 35532 9036
rect 35584 9024 35590 9036
rect 35584 8996 37688 9024
rect 35584 8984 35590 8996
rect 37660 8965 37688 8996
rect 36541 8959 36599 8965
rect 36541 8956 36553 8959
rect 35268 8928 36553 8956
rect 35161 8919 35219 8925
rect 36541 8925 36553 8928
rect 36587 8925 36599 8959
rect 36541 8919 36599 8925
rect 37645 8959 37703 8965
rect 37645 8925 37657 8959
rect 37691 8925 37703 8959
rect 37752 8956 37780 9064
rect 37829 9061 37841 9095
rect 37875 9092 37887 9095
rect 37875 9064 41414 9092
rect 37875 9061 37887 9064
rect 37829 9055 37887 9061
rect 39853 9027 39911 9033
rect 39853 9024 39865 9027
rect 39316 8996 39865 9024
rect 39316 8965 39344 8996
rect 39853 8993 39865 8996
rect 39899 8993 39911 9027
rect 41386 9024 41414 9064
rect 44174 9024 44180 9036
rect 41386 8996 44180 9024
rect 39853 8987 39911 8993
rect 44174 8984 44180 8996
rect 44232 8984 44238 9036
rect 49145 9027 49203 9033
rect 49145 8993 49157 9027
rect 49191 9024 49203 9027
rect 49326 9024 49332 9036
rect 49191 8996 49332 9024
rect 49191 8993 49203 8996
rect 49145 8987 49203 8993
rect 49326 8984 49332 8996
rect 49384 8984 49390 9036
rect 39301 8959 39359 8965
rect 39301 8956 39313 8959
rect 37752 8928 39313 8956
rect 37645 8919 37703 8925
rect 39301 8925 39313 8928
rect 39347 8925 39359 8959
rect 39301 8919 39359 8925
rect 39485 8959 39543 8965
rect 39485 8925 39497 8959
rect 39531 8956 39543 8959
rect 47670 8956 47676 8968
rect 39531 8928 47676 8956
rect 39531 8925 39543 8928
rect 39485 8919 39543 8925
rect 47670 8916 47676 8928
rect 47728 8916 47734 8968
rect 47762 8916 47768 8968
rect 47820 8956 47826 8968
rect 47949 8959 48007 8965
rect 47949 8956 47961 8959
rect 47820 8928 47961 8956
rect 47820 8916 47826 8928
rect 47949 8925 47961 8928
rect 47995 8925 48007 8959
rect 47949 8919 48007 8925
rect 20548 8860 22508 8888
rect 18782 8820 18788 8832
rect 16592 8792 18788 8820
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 18874 8780 18880 8832
rect 18932 8820 18938 8832
rect 20548 8820 20576 8860
rect 18932 8792 20576 8820
rect 21821 8823 21879 8829
rect 18932 8780 18938 8792
rect 21821 8789 21833 8823
rect 21867 8820 21879 8823
rect 22186 8820 22192 8832
rect 21867 8792 22192 8820
rect 21867 8789 21879 8792
rect 21821 8783 21879 8789
rect 22186 8780 22192 8792
rect 22244 8780 22250 8832
rect 22480 8820 22508 8860
rect 23400 8860 25636 8888
rect 28537 8891 28595 8897
rect 23400 8820 23428 8860
rect 28537 8857 28549 8891
rect 28583 8888 28595 8891
rect 29733 8891 29791 8897
rect 29733 8888 29745 8891
rect 28583 8860 29745 8888
rect 28583 8857 28595 8860
rect 28537 8851 28595 8857
rect 29733 8857 29745 8860
rect 29779 8857 29791 8891
rect 29733 8851 29791 8857
rect 30926 8848 30932 8900
rect 30984 8888 30990 8900
rect 30984 8860 31050 8888
rect 30984 8848 30990 8860
rect 32766 8848 32772 8900
rect 32824 8888 32830 8900
rect 36446 8888 36452 8900
rect 32824 8860 36452 8888
rect 32824 8848 32830 8860
rect 36446 8848 36452 8860
rect 36504 8848 36510 8900
rect 22480 8792 23428 8820
rect 23474 8780 23480 8832
rect 23532 8820 23538 8832
rect 24581 8823 24639 8829
rect 24581 8820 24593 8823
rect 23532 8792 24593 8820
rect 23532 8780 23538 8792
rect 24581 8789 24593 8792
rect 24627 8820 24639 8823
rect 24765 8823 24823 8829
rect 24765 8820 24777 8823
rect 24627 8792 24777 8820
rect 24627 8789 24639 8792
rect 24581 8783 24639 8789
rect 24765 8789 24777 8792
rect 24811 8820 24823 8823
rect 25317 8823 25375 8829
rect 25317 8820 25329 8823
rect 24811 8792 25329 8820
rect 24811 8789 24823 8792
rect 24765 8783 24823 8789
rect 25317 8789 25329 8792
rect 25363 8789 25375 8823
rect 25317 8783 25375 8789
rect 25682 8780 25688 8832
rect 25740 8780 25746 8832
rect 27798 8780 27804 8832
rect 27856 8820 27862 8832
rect 28442 8820 28448 8832
rect 27856 8792 28448 8820
rect 27856 8780 27862 8792
rect 28442 8780 28448 8792
rect 28500 8780 28506 8832
rect 30285 8823 30343 8829
rect 30285 8789 30297 8823
rect 30331 8820 30343 8823
rect 30374 8820 30380 8832
rect 30331 8792 30380 8820
rect 30331 8789 30343 8792
rect 30285 8783 30343 8789
rect 30374 8780 30380 8792
rect 30432 8820 30438 8832
rect 30650 8820 30656 8832
rect 30432 8792 30656 8820
rect 30432 8780 30438 8792
rect 30650 8780 30656 8792
rect 30708 8780 30714 8832
rect 32858 8780 32864 8832
rect 32916 8820 32922 8832
rect 33045 8823 33103 8829
rect 33045 8820 33057 8823
rect 32916 8792 33057 8820
rect 32916 8780 32922 8792
rect 33045 8789 33057 8792
rect 33091 8820 33103 8823
rect 33134 8820 33140 8832
rect 33091 8792 33140 8820
rect 33091 8789 33103 8792
rect 33045 8783 33103 8789
rect 33134 8780 33140 8792
rect 33192 8780 33198 8832
rect 33594 8780 33600 8832
rect 33652 8780 33658 8832
rect 33689 8823 33747 8829
rect 33689 8789 33701 8823
rect 33735 8820 33747 8823
rect 34238 8820 34244 8832
rect 33735 8792 34244 8820
rect 33735 8789 33747 8792
rect 33689 8783 33747 8789
rect 34238 8780 34244 8792
rect 34296 8780 34302 8832
rect 35250 8780 35256 8832
rect 35308 8780 35314 8832
rect 35618 8780 35624 8832
rect 35676 8780 35682 8832
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 13538 8576 13544 8628
rect 13596 8616 13602 8628
rect 13722 8616 13728 8628
rect 13596 8588 13728 8616
rect 13596 8576 13602 8588
rect 13722 8576 13728 8588
rect 13780 8616 13786 8628
rect 13780 8588 15240 8616
rect 13780 8576 13786 8588
rect 13906 8508 13912 8560
rect 13964 8508 13970 8560
rect 15212 8548 15240 8588
rect 15488 8588 18460 8616
rect 15488 8548 15516 8588
rect 15212 8520 15516 8548
rect 16390 8508 16396 8560
rect 16448 8548 16454 8560
rect 16758 8548 16764 8560
rect 16448 8520 16764 8548
rect 16448 8508 16454 8520
rect 16758 8508 16764 8520
rect 16816 8548 16822 8560
rect 17129 8551 17187 8557
rect 17129 8548 17141 8551
rect 16816 8520 17141 8548
rect 16816 8508 16822 8520
rect 17129 8517 17141 8520
rect 17175 8517 17187 8551
rect 18432 8548 18460 8588
rect 18598 8576 18604 8628
rect 18656 8576 18662 8628
rect 19705 8619 19763 8625
rect 19705 8585 19717 8619
rect 19751 8616 19763 8619
rect 19886 8616 19892 8628
rect 19751 8588 19892 8616
rect 19751 8585 19763 8588
rect 19705 8579 19763 8585
rect 19886 8576 19892 8588
rect 19944 8576 19950 8628
rect 22005 8619 22063 8625
rect 22005 8616 22017 8619
rect 21192 8588 22017 8616
rect 18874 8548 18880 8560
rect 18432 8520 18880 8548
rect 17129 8511 17187 8517
rect 18874 8508 18880 8520
rect 18932 8508 18938 8560
rect 20438 8508 20444 8560
rect 20496 8508 20502 8560
rect 21192 8557 21220 8588
rect 21177 8551 21235 8557
rect 21177 8517 21189 8551
rect 21223 8517 21235 8551
rect 21177 8511 21235 8517
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 2682 8480 2688 8492
rect 2179 8452 2688 8480
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 2682 8440 2688 8452
rect 2740 8440 2746 8492
rect 14918 8440 14924 8492
rect 14976 8480 14982 8492
rect 14976 8466 15042 8480
rect 14976 8452 15056 8466
rect 14976 8440 14982 8452
rect 2406 8372 2412 8424
rect 2464 8372 2470 8424
rect 13630 8372 13636 8424
rect 13688 8372 13694 8424
rect 15028 8344 15056 8452
rect 16022 8440 16028 8492
rect 16080 8480 16086 8492
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16080 8452 16865 8480
rect 16080 8440 16086 8452
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 18230 8440 18236 8492
rect 18288 8480 18294 8492
rect 18506 8480 18512 8492
rect 18288 8452 18512 8480
rect 18288 8440 18294 8452
rect 18506 8440 18512 8452
rect 18564 8440 18570 8492
rect 15102 8372 15108 8424
rect 15160 8412 15166 8424
rect 15381 8415 15439 8421
rect 15381 8412 15393 8415
rect 15160 8384 15393 8412
rect 15160 8372 15166 8384
rect 15381 8381 15393 8384
rect 15427 8381 15439 8415
rect 15381 8375 15439 8381
rect 17126 8372 17132 8424
rect 17184 8412 17190 8424
rect 19061 8415 19119 8421
rect 19061 8412 19073 8415
rect 17184 8384 19073 8412
rect 17184 8372 17190 8384
rect 19061 8381 19073 8384
rect 19107 8381 19119 8415
rect 19061 8375 19119 8381
rect 21450 8372 21456 8424
rect 21508 8372 21514 8424
rect 15749 8347 15807 8353
rect 15749 8344 15761 8347
rect 15028 8316 15761 8344
rect 15749 8313 15761 8316
rect 15795 8344 15807 8347
rect 16209 8347 16267 8353
rect 16209 8344 16221 8347
rect 15795 8316 16221 8344
rect 15795 8313 15807 8316
rect 15749 8307 15807 8313
rect 16209 8313 16221 8316
rect 16255 8344 16267 8347
rect 21928 8344 21956 8588
rect 22005 8585 22017 8588
rect 22051 8585 22063 8619
rect 22005 8579 22063 8585
rect 23474 8576 23480 8628
rect 23532 8616 23538 8628
rect 24029 8619 24087 8625
rect 24029 8616 24041 8619
rect 23532 8588 24041 8616
rect 23532 8576 23538 8588
rect 24029 8585 24041 8588
rect 24075 8585 24087 8619
rect 24029 8579 24087 8585
rect 31757 8619 31815 8625
rect 31757 8585 31769 8619
rect 31803 8616 31815 8619
rect 32766 8616 32772 8628
rect 31803 8588 32772 8616
rect 31803 8585 31815 8588
rect 31757 8579 31815 8585
rect 32766 8576 32772 8588
rect 32824 8576 32830 8628
rect 33870 8576 33876 8628
rect 33928 8616 33934 8628
rect 34057 8619 34115 8625
rect 34057 8616 34069 8619
rect 33928 8588 34069 8616
rect 33928 8576 33934 8588
rect 34057 8585 34069 8588
rect 34103 8616 34115 8619
rect 34974 8616 34980 8628
rect 34103 8588 34980 8616
rect 34103 8585 34115 8588
rect 34057 8579 34115 8585
rect 34974 8576 34980 8588
rect 35032 8576 35038 8628
rect 35986 8616 35992 8628
rect 35544 8588 35992 8616
rect 29086 8508 29092 8560
rect 29144 8508 29150 8560
rect 30466 8508 30472 8560
rect 30524 8548 30530 8560
rect 31297 8551 31355 8557
rect 31297 8548 31309 8551
rect 30524 8520 31309 8548
rect 30524 8508 30530 8520
rect 31297 8517 31309 8520
rect 31343 8517 31355 8551
rect 32030 8548 32036 8560
rect 31297 8511 31355 8517
rect 31772 8520 32036 8548
rect 31772 8492 31800 8520
rect 32030 8508 32036 8520
rect 32088 8548 32094 8560
rect 32858 8548 32864 8560
rect 32088 8520 32864 8548
rect 32088 8508 32094 8520
rect 32858 8508 32864 8520
rect 32916 8508 32922 8560
rect 33134 8508 33140 8560
rect 33192 8508 33198 8560
rect 34793 8551 34851 8557
rect 34793 8517 34805 8551
rect 34839 8548 34851 8551
rect 35544 8548 35572 8588
rect 35986 8576 35992 8588
rect 36044 8576 36050 8628
rect 37645 8619 37703 8625
rect 37645 8585 37657 8619
rect 37691 8616 37703 8619
rect 40034 8616 40040 8628
rect 37691 8588 40040 8616
rect 37691 8585 37703 8588
rect 37645 8579 37703 8585
rect 40034 8576 40040 8588
rect 40092 8576 40098 8628
rect 42702 8576 42708 8628
rect 42760 8616 42766 8628
rect 42760 8588 45416 8616
rect 42760 8576 42766 8588
rect 34839 8520 35572 8548
rect 34839 8517 34851 8520
rect 34793 8511 34851 8517
rect 35618 8508 35624 8560
rect 35676 8548 35682 8560
rect 35676 8520 38976 8548
rect 35676 8508 35682 8520
rect 22002 8440 22008 8492
rect 22060 8480 22066 8492
rect 23753 8483 23811 8489
rect 22060 8452 22402 8480
rect 22060 8440 22066 8452
rect 23753 8449 23765 8483
rect 23799 8480 23811 8483
rect 24026 8480 24032 8492
rect 23799 8452 24032 8480
rect 23799 8449 23811 8452
rect 23753 8443 23811 8449
rect 24026 8440 24032 8452
rect 24084 8440 24090 8492
rect 30650 8480 30656 8492
rect 30222 8452 30656 8480
rect 30650 8440 30656 8452
rect 30708 8480 30714 8492
rect 30926 8480 30932 8492
rect 30708 8452 30932 8480
rect 30708 8440 30714 8452
rect 30926 8440 30932 8452
rect 30984 8440 30990 8492
rect 31110 8440 31116 8492
rect 31168 8480 31174 8492
rect 31389 8483 31447 8489
rect 31389 8480 31401 8483
rect 31168 8452 31401 8480
rect 31168 8440 31174 8452
rect 31389 8449 31401 8452
rect 31435 8449 31447 8483
rect 31389 8443 31447 8449
rect 31754 8440 31760 8492
rect 31812 8440 31818 8492
rect 32306 8440 32312 8492
rect 32364 8440 32370 8492
rect 35802 8440 35808 8492
rect 35860 8480 35866 8492
rect 38948 8489 38976 8520
rect 40310 8508 40316 8560
rect 40368 8548 40374 8560
rect 40773 8551 40831 8557
rect 40773 8548 40785 8551
rect 40368 8520 40785 8548
rect 40368 8508 40374 8520
rect 40773 8517 40785 8520
rect 40819 8517 40831 8551
rect 40773 8511 40831 8517
rect 44174 8508 44180 8560
rect 44232 8508 44238 8560
rect 45388 8548 45416 8588
rect 45462 8576 45468 8628
rect 45520 8616 45526 8628
rect 47578 8616 47584 8628
rect 45520 8588 47584 8616
rect 45520 8576 45526 8588
rect 47578 8576 47584 8588
rect 47636 8576 47642 8628
rect 45388 8520 45876 8548
rect 37461 8483 37519 8489
rect 37461 8480 37473 8483
rect 35860 8452 37473 8480
rect 35860 8440 35866 8452
rect 37461 8449 37473 8452
rect 37507 8449 37519 8483
rect 37461 8443 37519 8449
rect 38933 8483 38991 8489
rect 38933 8449 38945 8483
rect 38979 8449 38991 8483
rect 38933 8443 38991 8449
rect 40497 8483 40555 8489
rect 40497 8449 40509 8483
rect 40543 8480 40555 8483
rect 45462 8480 45468 8492
rect 40543 8452 45468 8480
rect 40543 8449 40555 8452
rect 40497 8443 40555 8449
rect 45462 8440 45468 8452
rect 45520 8440 45526 8492
rect 45848 8489 45876 8520
rect 49142 8508 49148 8560
rect 49200 8508 49206 8560
rect 45833 8483 45891 8489
rect 45833 8449 45845 8483
rect 45879 8449 45891 8483
rect 45833 8443 45891 8449
rect 46198 8440 46204 8492
rect 46256 8480 46262 8492
rect 47949 8483 48007 8489
rect 47949 8480 47961 8483
rect 46256 8452 47961 8480
rect 46256 8440 46262 8452
rect 47949 8449 47961 8452
rect 47995 8449 48007 8483
rect 47949 8443 48007 8449
rect 22094 8372 22100 8424
rect 22152 8412 22158 8424
rect 23477 8415 23535 8421
rect 23477 8412 23489 8415
rect 22152 8384 23489 8412
rect 22152 8372 22158 8384
rect 23477 8381 23489 8384
rect 23523 8381 23535 8415
rect 23477 8375 23535 8381
rect 28810 8372 28816 8424
rect 28868 8412 28874 8424
rect 29178 8412 29184 8424
rect 28868 8384 29184 8412
rect 28868 8372 28874 8384
rect 29178 8372 29184 8384
rect 29236 8372 29242 8424
rect 31205 8415 31263 8421
rect 31205 8381 31217 8415
rect 31251 8412 31263 8415
rect 31938 8412 31944 8424
rect 31251 8384 31944 8412
rect 31251 8381 31263 8384
rect 31205 8375 31263 8381
rect 31938 8372 31944 8384
rect 31996 8372 32002 8424
rect 32214 8372 32220 8424
rect 32272 8412 32278 8424
rect 32582 8412 32588 8424
rect 32272 8384 32588 8412
rect 32272 8372 32278 8384
rect 32582 8372 32588 8384
rect 32640 8372 32646 8424
rect 32950 8372 32956 8424
rect 33008 8412 33014 8424
rect 38746 8412 38752 8424
rect 33008 8384 38752 8412
rect 33008 8372 33014 8384
rect 38746 8372 38752 8384
rect 38804 8372 38810 8424
rect 40218 8412 40224 8424
rect 38856 8384 40224 8412
rect 22462 8344 22468 8356
rect 16255 8316 16988 8344
rect 21928 8316 22468 8344
rect 16255 8313 16267 8316
rect 16209 8307 16267 8313
rect 16960 8276 16988 8316
rect 22462 8304 22468 8316
rect 22520 8304 22526 8356
rect 30561 8347 30619 8353
rect 30561 8313 30573 8347
rect 30607 8344 30619 8347
rect 31846 8344 31852 8356
rect 30607 8316 31852 8344
rect 30607 8313 30619 8316
rect 30561 8307 30619 8313
rect 31846 8304 31852 8316
rect 31904 8304 31910 8356
rect 34333 8347 34391 8353
rect 34333 8344 34345 8347
rect 33612 8316 34345 8344
rect 17310 8276 17316 8288
rect 16960 8248 17316 8276
rect 17310 8236 17316 8248
rect 17368 8236 17374 8288
rect 31938 8236 31944 8288
rect 31996 8276 32002 8288
rect 33042 8276 33048 8288
rect 31996 8248 33048 8276
rect 31996 8236 32002 8248
rect 33042 8236 33048 8248
rect 33100 8276 33106 8288
rect 33612 8276 33640 8316
rect 34333 8313 34345 8316
rect 34379 8313 34391 8347
rect 34609 8347 34667 8353
rect 34609 8344 34621 8347
rect 34333 8307 34391 8313
rect 34440 8316 34621 8344
rect 33100 8248 33640 8276
rect 33100 8236 33106 8248
rect 33686 8236 33692 8288
rect 33744 8276 33750 8288
rect 34440 8276 34468 8316
rect 34609 8313 34621 8316
rect 34655 8344 34667 8347
rect 38856 8344 38884 8384
rect 40218 8372 40224 8384
rect 40276 8372 40282 8424
rect 44361 8415 44419 8421
rect 44361 8381 44373 8415
rect 44407 8412 44419 8415
rect 44407 8384 45554 8412
rect 44407 8381 44419 8384
rect 44361 8375 44419 8381
rect 34655 8316 38884 8344
rect 39117 8347 39175 8353
rect 34655 8313 34667 8316
rect 34609 8307 34667 8313
rect 39117 8313 39129 8347
rect 39163 8344 39175 8347
rect 44910 8344 44916 8356
rect 39163 8316 44916 8344
rect 39163 8313 39175 8316
rect 39117 8307 39175 8313
rect 44910 8304 44916 8316
rect 44968 8304 44974 8356
rect 45526 8344 45554 8384
rect 46842 8372 46848 8424
rect 46900 8372 46906 8424
rect 47762 8344 47768 8356
rect 45526 8316 47768 8344
rect 47762 8304 47768 8316
rect 47820 8304 47826 8356
rect 33744 8248 34468 8276
rect 33744 8236 33750 8248
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 1302 8032 1308 8084
rect 1360 8072 1366 8084
rect 2133 8075 2191 8081
rect 2133 8072 2145 8075
rect 1360 8044 2145 8072
rect 1360 8032 1366 8044
rect 2133 8041 2145 8044
rect 2179 8072 2191 8075
rect 2406 8072 2412 8084
rect 2179 8044 2412 8072
rect 2179 8041 2191 8044
rect 2133 8035 2191 8041
rect 2406 8032 2412 8044
rect 2464 8032 2470 8084
rect 18414 8032 18420 8084
rect 18472 8072 18478 8084
rect 18969 8075 19027 8081
rect 18969 8072 18981 8075
rect 18472 8044 18981 8072
rect 18472 8032 18478 8044
rect 18969 8041 18981 8044
rect 19015 8041 19027 8075
rect 18969 8035 19027 8041
rect 19426 8032 19432 8084
rect 19484 8032 19490 8084
rect 21910 8032 21916 8084
rect 21968 8072 21974 8084
rect 22005 8075 22063 8081
rect 22005 8072 22017 8075
rect 21968 8044 22017 8072
rect 21968 8032 21974 8044
rect 22005 8041 22017 8044
rect 22051 8041 22063 8075
rect 22005 8035 22063 8041
rect 30377 8075 30435 8081
rect 30377 8041 30389 8075
rect 30423 8072 30435 8075
rect 30558 8072 30564 8084
rect 30423 8044 30564 8072
rect 30423 8041 30435 8044
rect 30377 8035 30435 8041
rect 30558 8032 30564 8044
rect 30616 8032 30622 8084
rect 31757 8075 31815 8081
rect 31757 8041 31769 8075
rect 31803 8072 31815 8075
rect 35250 8072 35256 8084
rect 31803 8044 35256 8072
rect 31803 8041 31815 8044
rect 31757 8035 31815 8041
rect 35250 8032 35256 8044
rect 35308 8032 35314 8084
rect 15749 8007 15807 8013
rect 15749 7973 15761 8007
rect 15795 8004 15807 8007
rect 18874 8004 18880 8016
rect 15795 7976 18880 8004
rect 15795 7973 15807 7976
rect 15749 7967 15807 7973
rect 18874 7964 18880 7976
rect 18932 7964 18938 8016
rect 21634 7964 21640 8016
rect 21692 8004 21698 8016
rect 22646 8004 22652 8016
rect 21692 7976 22652 8004
rect 21692 7964 21698 7976
rect 22646 7964 22652 7976
rect 22704 8004 22710 8016
rect 32582 8004 32588 8016
rect 22704 7976 32588 8004
rect 22704 7964 22710 7976
rect 32582 7964 32588 7976
rect 32640 7964 32646 8016
rect 33045 8007 33103 8013
rect 33045 7973 33057 8007
rect 33091 8004 33103 8007
rect 39022 8004 39028 8016
rect 33091 7976 39028 8004
rect 33091 7973 33103 7976
rect 33045 7967 33103 7973
rect 39022 7964 39028 7976
rect 39080 7964 39086 8016
rect 16758 7896 16764 7948
rect 16816 7896 16822 7948
rect 16942 7896 16948 7948
rect 17000 7896 17006 7948
rect 18049 7939 18107 7945
rect 18049 7905 18061 7939
rect 18095 7936 18107 7939
rect 18598 7936 18604 7948
rect 18095 7908 18604 7936
rect 18095 7905 18107 7908
rect 18049 7899 18107 7905
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 19886 7896 19892 7948
rect 19944 7936 19950 7948
rect 20901 7939 20959 7945
rect 20901 7936 20913 7939
rect 19944 7908 20913 7936
rect 19944 7896 19950 7908
rect 20901 7905 20913 7908
rect 20947 7905 20959 7939
rect 20901 7899 20959 7905
rect 22557 7939 22615 7945
rect 22557 7905 22569 7939
rect 22603 7936 22615 7939
rect 23658 7936 23664 7948
rect 22603 7908 23664 7936
rect 22603 7905 22615 7908
rect 22557 7899 22615 7905
rect 23658 7896 23664 7908
rect 23716 7896 23722 7948
rect 29914 7896 29920 7948
rect 29972 7896 29978 7948
rect 31205 7939 31263 7945
rect 31205 7905 31217 7939
rect 31251 7936 31263 7939
rect 32214 7936 32220 7948
rect 31251 7908 32220 7936
rect 31251 7905 31263 7908
rect 31205 7899 31263 7905
rect 32214 7896 32220 7908
rect 32272 7896 32278 7948
rect 32493 7939 32551 7945
rect 32493 7905 32505 7939
rect 32539 7936 32551 7939
rect 33413 7939 33471 7945
rect 33413 7936 33425 7939
rect 32539 7908 33425 7936
rect 32539 7905 32551 7908
rect 32493 7899 32551 7905
rect 33413 7905 33425 7908
rect 33459 7936 33471 7939
rect 34514 7936 34520 7948
rect 33459 7908 34520 7936
rect 33459 7905 33471 7908
rect 33413 7899 33471 7905
rect 34514 7896 34520 7908
rect 34572 7896 34578 7948
rect 49145 7939 49203 7945
rect 49145 7905 49157 7939
rect 49191 7936 49203 7939
rect 49234 7936 49240 7948
rect 49191 7908 49240 7936
rect 49191 7905 49203 7908
rect 49145 7899 49203 7905
rect 49234 7896 49240 7908
rect 49292 7896 49298 7948
rect 1302 7828 1308 7880
rect 1360 7868 1366 7880
rect 1581 7871 1639 7877
rect 1581 7868 1593 7871
rect 1360 7840 1593 7868
rect 1360 7828 1366 7840
rect 1581 7837 1593 7840
rect 1627 7868 1639 7871
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 1627 7840 2329 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 2317 7837 2329 7840
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 14090 7828 14096 7880
rect 14148 7868 14154 7880
rect 15565 7871 15623 7877
rect 15565 7868 15577 7871
rect 14148 7840 15577 7868
rect 14148 7828 14154 7840
rect 15565 7837 15577 7840
rect 15611 7837 15623 7871
rect 15565 7831 15623 7837
rect 17034 7828 17040 7880
rect 17092 7828 17098 7880
rect 18141 7871 18199 7877
rect 18141 7868 18153 7871
rect 17236 7840 18153 7868
rect 13722 7800 13728 7812
rect 1780 7772 13728 7800
rect 1780 7741 1808 7772
rect 13722 7760 13728 7772
rect 13780 7760 13786 7812
rect 16298 7760 16304 7812
rect 16356 7800 16362 7812
rect 17236 7800 17264 7840
rect 18141 7837 18153 7840
rect 18187 7837 18199 7871
rect 18141 7831 18199 7837
rect 21177 7871 21235 7877
rect 21177 7837 21189 7871
rect 21223 7868 21235 7871
rect 21450 7868 21456 7880
rect 21223 7840 21456 7868
rect 21223 7837 21235 7840
rect 21177 7831 21235 7837
rect 18233 7803 18291 7809
rect 18233 7800 18245 7803
rect 16356 7772 17264 7800
rect 17420 7772 18245 7800
rect 16356 7760 16362 7772
rect 17420 7741 17448 7772
rect 18233 7769 18245 7772
rect 18279 7769 18291 7803
rect 19610 7800 19616 7812
rect 18233 7763 18291 7769
rect 18616 7772 19616 7800
rect 18616 7741 18644 7772
rect 19610 7760 19616 7772
rect 19668 7760 19674 7812
rect 20438 7760 20444 7812
rect 20496 7800 20502 7812
rect 20496 7772 20576 7800
rect 20496 7760 20502 7772
rect 1765 7735 1823 7741
rect 1765 7701 1777 7735
rect 1811 7701 1823 7735
rect 1765 7695 1823 7701
rect 17405 7735 17463 7741
rect 17405 7701 17417 7735
rect 17451 7701 17463 7735
rect 17405 7695 17463 7701
rect 18601 7735 18659 7741
rect 18601 7701 18613 7735
rect 18647 7701 18659 7735
rect 20548 7732 20576 7772
rect 20990 7760 20996 7812
rect 21048 7800 21054 7812
rect 21192 7800 21220 7831
rect 21450 7828 21456 7840
rect 21508 7828 21514 7880
rect 22186 7828 22192 7880
rect 22244 7868 22250 7880
rect 22373 7871 22431 7877
rect 22373 7868 22385 7871
rect 22244 7840 22385 7868
rect 22244 7828 22250 7840
rect 22373 7837 22385 7840
rect 22419 7837 22431 7871
rect 22373 7831 22431 7837
rect 30558 7828 30564 7880
rect 30616 7868 30622 7880
rect 31297 7871 31355 7877
rect 31297 7868 31309 7871
rect 30616 7840 31309 7868
rect 30616 7828 30622 7840
rect 31297 7837 31309 7840
rect 31343 7837 31355 7871
rect 31297 7831 31355 7837
rect 32674 7828 32680 7880
rect 32732 7828 32738 7880
rect 38746 7828 38752 7880
rect 38804 7868 38810 7880
rect 39209 7871 39267 7877
rect 39209 7868 39221 7871
rect 38804 7840 39221 7868
rect 38804 7828 38810 7840
rect 39209 7837 39221 7840
rect 39255 7837 39267 7871
rect 39209 7831 39267 7837
rect 46934 7828 46940 7880
rect 46992 7868 46998 7880
rect 47949 7871 48007 7877
rect 47949 7868 47961 7871
rect 46992 7840 47961 7868
rect 46992 7828 46998 7840
rect 47949 7837 47961 7840
rect 47995 7837 48007 7871
rect 47949 7831 48007 7837
rect 30466 7800 30472 7812
rect 21048 7772 21220 7800
rect 22388 7772 30472 7800
rect 21048 7760 21054 7772
rect 22388 7744 22416 7772
rect 30466 7760 30472 7772
rect 30524 7760 30530 7812
rect 37553 7803 37611 7809
rect 37553 7800 37565 7803
rect 30576 7772 37565 7800
rect 21450 7732 21456 7744
rect 20548 7704 21456 7732
rect 18601 7695 18659 7701
rect 21450 7692 21456 7704
rect 21508 7692 21514 7744
rect 21634 7692 21640 7744
rect 21692 7692 21698 7744
rect 22370 7692 22376 7744
rect 22428 7692 22434 7744
rect 22462 7692 22468 7744
rect 22520 7732 22526 7744
rect 23017 7735 23075 7741
rect 23017 7732 23029 7735
rect 22520 7704 23029 7732
rect 22520 7692 22526 7704
rect 23017 7701 23029 7704
rect 23063 7732 23075 7735
rect 25682 7732 25688 7744
rect 23063 7704 25688 7732
rect 23063 7701 23075 7704
rect 23017 7695 23075 7701
rect 25682 7692 25688 7704
rect 25740 7692 25746 7744
rect 27522 7692 27528 7744
rect 27580 7732 27586 7744
rect 30576 7732 30604 7772
rect 37553 7769 37565 7772
rect 37599 7800 37611 7803
rect 38013 7803 38071 7809
rect 38013 7800 38025 7803
rect 37599 7772 38025 7800
rect 37599 7769 37611 7772
rect 37553 7763 37611 7769
rect 38013 7769 38025 7772
rect 38059 7769 38071 7803
rect 38013 7763 38071 7769
rect 38933 7803 38991 7809
rect 38933 7769 38945 7803
rect 38979 7800 38991 7803
rect 40126 7800 40132 7812
rect 38979 7772 40132 7800
rect 38979 7769 38991 7772
rect 38933 7763 38991 7769
rect 40126 7760 40132 7772
rect 40184 7760 40190 7812
rect 27580 7704 30604 7732
rect 27580 7692 27586 7704
rect 30650 7692 30656 7744
rect 30708 7692 30714 7744
rect 31386 7692 31392 7744
rect 31444 7692 31450 7744
rect 32582 7692 32588 7744
rect 32640 7692 32646 7744
rect 38105 7735 38163 7741
rect 38105 7701 38117 7735
rect 38151 7732 38163 7735
rect 38654 7732 38660 7744
rect 38151 7704 38660 7732
rect 38151 7701 38163 7704
rect 38105 7695 38163 7701
rect 38654 7692 38660 7704
rect 38712 7692 38718 7744
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 19794 7488 19800 7540
rect 19852 7528 19858 7540
rect 22005 7531 22063 7537
rect 22005 7528 22017 7531
rect 19852 7500 22017 7528
rect 19852 7488 19858 7500
rect 22005 7497 22017 7500
rect 22051 7497 22063 7531
rect 22005 7491 22063 7497
rect 22278 7488 22284 7540
rect 22336 7528 22342 7540
rect 22465 7531 22523 7537
rect 22465 7528 22477 7531
rect 22336 7500 22477 7528
rect 22336 7488 22342 7500
rect 22465 7497 22477 7500
rect 22511 7528 22523 7531
rect 23017 7531 23075 7537
rect 23017 7528 23029 7531
rect 22511 7500 23029 7528
rect 22511 7497 22523 7500
rect 22465 7491 22523 7497
rect 23017 7497 23029 7500
rect 23063 7497 23075 7531
rect 23017 7491 23075 7497
rect 31110 7488 31116 7540
rect 31168 7488 31174 7540
rect 31386 7488 31392 7540
rect 31444 7528 31450 7540
rect 32309 7531 32367 7537
rect 32309 7528 32321 7531
rect 31444 7500 32321 7528
rect 31444 7488 31450 7500
rect 32309 7497 32321 7500
rect 32355 7497 32367 7531
rect 39025 7531 39083 7537
rect 39025 7528 39037 7531
rect 32309 7491 32367 7497
rect 38580 7500 39037 7528
rect 17862 7420 17868 7472
rect 17920 7460 17926 7472
rect 18325 7463 18383 7469
rect 18325 7460 18337 7463
rect 17920 7432 18337 7460
rect 17920 7420 17926 7432
rect 18325 7429 18337 7432
rect 18371 7460 18383 7463
rect 18506 7460 18512 7472
rect 18371 7432 18512 7460
rect 18371 7429 18383 7432
rect 18325 7423 18383 7429
rect 18506 7420 18512 7432
rect 18564 7460 18570 7472
rect 18785 7463 18843 7469
rect 18785 7460 18797 7463
rect 18564 7432 18797 7460
rect 18564 7420 18570 7432
rect 18785 7429 18797 7432
rect 18831 7460 18843 7463
rect 19061 7463 19119 7469
rect 19061 7460 19073 7463
rect 18831 7432 19073 7460
rect 18831 7429 18843 7432
rect 18785 7423 18843 7429
rect 19061 7429 19073 7432
rect 19107 7460 19119 7463
rect 20438 7460 20444 7472
rect 19107 7432 20444 7460
rect 19107 7429 19119 7432
rect 19061 7423 19119 7429
rect 20438 7420 20444 7432
rect 20496 7420 20502 7472
rect 31938 7420 31944 7472
rect 31996 7420 32002 7472
rect 34422 7420 34428 7472
rect 34480 7460 34486 7472
rect 38580 7469 38608 7500
rect 39025 7497 39037 7500
rect 39071 7497 39083 7531
rect 39025 7491 39083 7497
rect 38565 7463 38623 7469
rect 38565 7460 38577 7463
rect 34480 7432 38577 7460
rect 34480 7420 34486 7432
rect 38565 7429 38577 7432
rect 38611 7429 38623 7463
rect 38565 7423 38623 7429
rect 38654 7420 38660 7472
rect 38712 7460 38718 7472
rect 47302 7460 47308 7472
rect 38712 7432 47308 7460
rect 38712 7420 38718 7432
rect 47302 7420 47308 7432
rect 47360 7420 47366 7472
rect 49145 7463 49203 7469
rect 49145 7429 49157 7463
rect 49191 7460 49203 7463
rect 49326 7460 49332 7472
rect 49191 7432 49332 7460
rect 49191 7429 49203 7432
rect 49145 7423 49203 7429
rect 49326 7420 49332 7432
rect 49384 7420 49390 7472
rect 1302 7352 1308 7404
rect 1360 7392 1366 7404
rect 1581 7395 1639 7401
rect 1581 7392 1593 7395
rect 1360 7364 1593 7392
rect 1360 7352 1366 7364
rect 1581 7361 1593 7364
rect 1627 7392 1639 7395
rect 2133 7395 2191 7401
rect 2133 7392 2145 7395
rect 1627 7364 2145 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 2133 7361 2145 7364
rect 2179 7361 2191 7395
rect 2133 7355 2191 7361
rect 22370 7352 22376 7404
rect 22428 7352 22434 7404
rect 37829 7395 37887 7401
rect 37829 7392 37841 7395
rect 37384 7364 37841 7392
rect 22554 7284 22560 7336
rect 22612 7284 22618 7336
rect 1765 7259 1823 7265
rect 1765 7225 1777 7259
rect 1811 7256 1823 7259
rect 19242 7256 19248 7268
rect 1811 7228 19248 7256
rect 1811 7225 1823 7228
rect 1765 7219 1823 7225
rect 19242 7216 19248 7228
rect 19300 7216 19306 7268
rect 28626 7216 28632 7268
rect 28684 7256 28690 7268
rect 37384 7265 37412 7364
rect 37829 7361 37841 7364
rect 37875 7361 37887 7395
rect 37829 7355 37887 7361
rect 44910 7352 44916 7404
rect 44968 7352 44974 7404
rect 47026 7352 47032 7404
rect 47084 7392 47090 7404
rect 47949 7395 48007 7401
rect 47949 7392 47961 7395
rect 47084 7364 47961 7392
rect 47084 7352 47090 7364
rect 47949 7361 47961 7364
rect 47995 7361 48007 7395
rect 47949 7355 48007 7361
rect 37369 7259 37427 7265
rect 37369 7256 37381 7259
rect 28684 7228 37381 7256
rect 28684 7216 28690 7228
rect 37369 7225 37381 7228
rect 37415 7225 37427 7259
rect 37369 7219 37427 7225
rect 38749 7259 38807 7265
rect 38749 7225 38761 7259
rect 38795 7256 38807 7259
rect 45097 7259 45155 7265
rect 38795 7228 42104 7256
rect 38795 7225 38807 7228
rect 38749 7219 38807 7225
rect 21177 7191 21235 7197
rect 21177 7157 21189 7191
rect 21223 7188 21235 7191
rect 21361 7191 21419 7197
rect 21361 7188 21373 7191
rect 21223 7160 21373 7188
rect 21223 7157 21235 7160
rect 21177 7151 21235 7157
rect 21361 7157 21373 7160
rect 21407 7188 21419 7191
rect 21450 7188 21456 7200
rect 21407 7160 21456 7188
rect 21407 7157 21419 7160
rect 21361 7151 21419 7157
rect 21450 7148 21456 7160
rect 21508 7188 21514 7200
rect 21637 7191 21695 7197
rect 21637 7188 21649 7191
rect 21508 7160 21649 7188
rect 21508 7148 21514 7160
rect 21637 7157 21649 7160
rect 21683 7188 21695 7191
rect 22002 7188 22008 7200
rect 21683 7160 22008 7188
rect 21683 7157 21695 7160
rect 21637 7151 21695 7157
rect 22002 7148 22008 7160
rect 22060 7148 22066 7200
rect 32582 7148 32588 7200
rect 32640 7188 32646 7200
rect 32861 7191 32919 7197
rect 32861 7188 32873 7191
rect 32640 7160 32873 7188
rect 32640 7148 32646 7160
rect 32861 7157 32873 7160
rect 32907 7188 32919 7191
rect 37274 7188 37280 7200
rect 32907 7160 37280 7188
rect 32907 7157 32919 7160
rect 32861 7151 32919 7157
rect 37274 7148 37280 7160
rect 37332 7148 37338 7200
rect 37918 7148 37924 7200
rect 37976 7148 37982 7200
rect 42076 7188 42104 7228
rect 45097 7225 45109 7259
rect 45143 7256 45155 7259
rect 47854 7256 47860 7268
rect 45143 7228 47860 7256
rect 45143 7225 45155 7228
rect 45097 7219 45155 7225
rect 47854 7216 47860 7228
rect 47912 7216 47918 7268
rect 45830 7188 45836 7200
rect 42076 7160 45836 7188
rect 45830 7148 45836 7160
rect 45888 7148 45894 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 30466 6944 30472 6996
rect 30524 6984 30530 6996
rect 38470 6984 38476 6996
rect 30524 6956 38476 6984
rect 30524 6944 30530 6956
rect 38470 6944 38476 6956
rect 38528 6944 38534 6996
rect 37918 6876 37924 6928
rect 37976 6916 37982 6928
rect 46934 6916 46940 6928
rect 37976 6888 46940 6916
rect 37976 6876 37982 6888
rect 46934 6876 46940 6888
rect 46992 6876 46998 6928
rect 15654 6808 15660 6860
rect 15712 6848 15718 6860
rect 21821 6851 21879 6857
rect 21821 6848 21833 6851
rect 15712 6820 21833 6848
rect 15712 6808 15718 6820
rect 21821 6817 21833 6820
rect 21867 6848 21879 6851
rect 22370 6848 22376 6860
rect 21867 6820 22376 6848
rect 21867 6817 21879 6820
rect 21821 6811 21879 6817
rect 22370 6808 22376 6820
rect 22428 6808 22434 6860
rect 49142 6808 49148 6860
rect 49200 6808 49206 6860
rect 1302 6740 1308 6792
rect 1360 6780 1366 6792
rect 2317 6783 2375 6789
rect 2317 6780 2329 6783
rect 1360 6752 2329 6780
rect 1360 6740 1366 6752
rect 2317 6749 2329 6752
rect 2363 6780 2375 6783
rect 2777 6783 2835 6789
rect 2777 6780 2789 6783
rect 2363 6752 2789 6780
rect 2363 6749 2375 6752
rect 2317 6743 2375 6749
rect 2777 6749 2789 6752
rect 2823 6749 2835 6783
rect 2777 6743 2835 6749
rect 15930 6740 15936 6792
rect 15988 6780 15994 6792
rect 17681 6783 17739 6789
rect 17681 6780 17693 6783
rect 15988 6752 17693 6780
rect 15988 6740 15994 6752
rect 17681 6749 17693 6752
rect 17727 6749 17739 6783
rect 17681 6743 17739 6749
rect 19610 6740 19616 6792
rect 19668 6740 19674 6792
rect 40126 6740 40132 6792
rect 40184 6780 40190 6792
rect 46109 6783 46167 6789
rect 46109 6780 46121 6783
rect 40184 6752 46121 6780
rect 40184 6740 40190 6752
rect 46109 6749 46121 6752
rect 46155 6749 46167 6783
rect 46109 6743 46167 6749
rect 47762 6740 47768 6792
rect 47820 6780 47826 6792
rect 47949 6783 48007 6789
rect 47949 6780 47961 6783
rect 47820 6752 47961 6780
rect 47820 6740 47826 6752
rect 47949 6749 47961 6752
rect 47995 6749 48007 6783
rect 47949 6743 48007 6749
rect 1210 6672 1216 6724
rect 1268 6712 1274 6724
rect 1673 6715 1731 6721
rect 1673 6712 1685 6715
rect 1268 6684 1685 6712
rect 1268 6672 1274 6684
rect 1673 6681 1685 6684
rect 1719 6681 1731 6715
rect 10594 6712 10600 6724
rect 1673 6675 1731 6681
rect 2516 6684 10600 6712
rect 1762 6604 1768 6656
rect 1820 6604 1826 6656
rect 2516 6653 2544 6684
rect 10594 6672 10600 6684
rect 10652 6672 10658 6724
rect 47305 6715 47363 6721
rect 47305 6681 47317 6715
rect 47351 6712 47363 6715
rect 48682 6712 48688 6724
rect 47351 6684 48688 6712
rect 47351 6681 47363 6684
rect 47305 6675 47363 6681
rect 48682 6672 48688 6684
rect 48740 6672 48746 6724
rect 2501 6647 2559 6653
rect 2501 6613 2513 6647
rect 2547 6613 2559 6647
rect 2501 6607 2559 6613
rect 17865 6647 17923 6653
rect 17865 6613 17877 6647
rect 17911 6644 17923 6647
rect 19242 6644 19248 6656
rect 17911 6616 19248 6644
rect 17911 6613 17923 6616
rect 17865 6607 17923 6613
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 19797 6647 19855 6653
rect 19797 6613 19809 6647
rect 19843 6644 19855 6647
rect 21726 6644 21732 6656
rect 19843 6616 21732 6644
rect 19843 6613 19855 6616
rect 19797 6607 19855 6613
rect 21726 6604 21732 6616
rect 21784 6604 21790 6656
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 1210 6400 1216 6452
rect 1268 6440 1274 6452
rect 2133 6443 2191 6449
rect 2133 6440 2145 6443
rect 1268 6412 2145 6440
rect 1268 6400 1274 6412
rect 2133 6409 2145 6412
rect 2179 6409 2191 6443
rect 2133 6403 2191 6409
rect 1762 6332 1768 6384
rect 1820 6372 1826 6384
rect 27798 6372 27804 6384
rect 1820 6344 27804 6372
rect 1820 6332 1826 6344
rect 27798 6332 27804 6344
rect 27856 6332 27862 6384
rect 30742 6332 30748 6384
rect 30800 6372 30806 6384
rect 37553 6375 37611 6381
rect 37553 6372 37565 6375
rect 30800 6344 37565 6372
rect 30800 6332 30806 6344
rect 37553 6341 37565 6344
rect 37599 6372 37611 6375
rect 38013 6375 38071 6381
rect 38013 6372 38025 6375
rect 37599 6344 38025 6372
rect 37599 6341 37611 6344
rect 37553 6335 37611 6341
rect 38013 6341 38025 6344
rect 38059 6341 38071 6375
rect 38013 6335 38071 6341
rect 40034 6332 40040 6384
rect 40092 6372 40098 6384
rect 43993 6375 44051 6381
rect 43993 6372 44005 6375
rect 40092 6344 44005 6372
rect 40092 6332 40098 6344
rect 43993 6341 44005 6344
rect 44039 6341 44051 6375
rect 43993 6335 44051 6341
rect 49145 6375 49203 6381
rect 49145 6341 49157 6375
rect 49191 6372 49203 6375
rect 49326 6372 49332 6384
rect 49191 6344 49332 6372
rect 49191 6341 49203 6344
rect 49145 6335 49203 6341
rect 49326 6332 49332 6344
rect 49384 6332 49390 6384
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 1581 6307 1639 6313
rect 1581 6304 1593 6307
rect 1360 6276 1593 6304
rect 1360 6264 1366 6276
rect 1581 6273 1593 6276
rect 1627 6304 1639 6307
rect 2317 6307 2375 6313
rect 2317 6304 2329 6307
rect 1627 6276 2329 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 2317 6273 2329 6276
rect 2363 6273 2375 6307
rect 2317 6267 2375 6273
rect 16850 6264 16856 6316
rect 16908 6304 16914 6316
rect 18049 6307 18107 6313
rect 18049 6304 18061 6307
rect 16908 6276 18061 6304
rect 16908 6264 16914 6276
rect 18049 6273 18061 6276
rect 18095 6273 18107 6307
rect 18049 6267 18107 6273
rect 47670 6264 47676 6316
rect 47728 6304 47734 6316
rect 47949 6307 48007 6313
rect 47949 6304 47961 6307
rect 47728 6276 47961 6304
rect 47728 6264 47734 6276
rect 47949 6273 47961 6276
rect 47995 6273 48007 6307
rect 47949 6267 48007 6273
rect 18233 6239 18291 6245
rect 18233 6205 18245 6239
rect 18279 6236 18291 6239
rect 18322 6236 18328 6248
rect 18279 6208 18328 6236
rect 18279 6205 18291 6208
rect 18233 6199 18291 6205
rect 18322 6196 18328 6208
rect 18380 6196 18386 6248
rect 1765 6171 1823 6177
rect 1765 6137 1777 6171
rect 1811 6168 1823 6171
rect 11238 6168 11244 6180
rect 1811 6140 11244 6168
rect 1811 6137 1823 6140
rect 1765 6131 1823 6137
rect 11238 6128 11244 6140
rect 11296 6128 11302 6180
rect 44177 6171 44235 6177
rect 44177 6137 44189 6171
rect 44223 6168 44235 6171
rect 47026 6168 47032 6180
rect 44223 6140 47032 6168
rect 44223 6137 44235 6140
rect 44177 6131 44235 6137
rect 47026 6128 47032 6140
rect 47084 6128 47090 6180
rect 18693 6103 18751 6109
rect 18693 6069 18705 6103
rect 18739 6100 18751 6103
rect 19426 6100 19432 6112
rect 18739 6072 19432 6100
rect 18739 6069 18751 6072
rect 18693 6063 18751 6069
rect 19426 6060 19432 6072
rect 19484 6060 19490 6112
rect 37642 6060 37648 6112
rect 37700 6060 37706 6112
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 37642 5856 37648 5908
rect 37700 5896 37706 5908
rect 47210 5896 47216 5908
rect 37700 5868 47216 5896
rect 37700 5856 37706 5868
rect 47210 5856 47216 5868
rect 47268 5856 47274 5908
rect 2501 5831 2559 5837
rect 2501 5797 2513 5831
rect 2547 5828 2559 5831
rect 13354 5828 13360 5840
rect 2547 5800 13360 5828
rect 2547 5797 2559 5800
rect 2501 5791 2559 5797
rect 13354 5788 13360 5800
rect 13412 5788 13418 5840
rect 3053 5763 3111 5769
rect 3053 5760 3065 5763
rect 1596 5732 3065 5760
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 1596 5701 1624 5732
rect 3053 5729 3065 5732
rect 3099 5729 3111 5763
rect 3053 5723 3111 5729
rect 49145 5763 49203 5769
rect 49145 5729 49157 5763
rect 49191 5760 49203 5763
rect 49234 5760 49240 5772
rect 49191 5732 49240 5760
rect 49191 5729 49203 5732
rect 49145 5723 49203 5729
rect 49234 5720 49240 5732
rect 49292 5720 49298 5772
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1360 5664 1593 5692
rect 1360 5652 1366 5664
rect 1581 5661 1593 5664
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5692 2375 5695
rect 2774 5692 2780 5704
rect 2363 5664 2780 5692
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 2774 5652 2780 5664
rect 2832 5692 2838 5704
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 2832 5664 2881 5692
rect 2832 5652 2838 5664
rect 2869 5661 2881 5664
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 43714 5652 43720 5704
rect 43772 5652 43778 5704
rect 47578 5652 47584 5704
rect 47636 5692 47642 5704
rect 47949 5695 48007 5701
rect 47949 5692 47961 5695
rect 47636 5664 47961 5692
rect 47636 5652 47642 5664
rect 47949 5661 47961 5664
rect 47995 5661 48007 5695
rect 47949 5655 48007 5661
rect 16206 5624 16212 5636
rect 1780 5596 16212 5624
rect 1780 5565 1808 5596
rect 16206 5584 16212 5596
rect 16264 5584 16270 5636
rect 43901 5627 43959 5633
rect 43901 5593 43913 5627
rect 43947 5624 43959 5627
rect 45738 5624 45744 5636
rect 43947 5596 45744 5624
rect 43947 5593 43959 5596
rect 43901 5587 43959 5593
rect 45738 5584 45744 5596
rect 45796 5584 45802 5636
rect 1765 5559 1823 5565
rect 1765 5525 1777 5559
rect 1811 5525 1823 5559
rect 1765 5519 1823 5525
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 37274 5244 37280 5296
rect 37332 5284 37338 5296
rect 37369 5287 37427 5293
rect 37369 5284 37381 5287
rect 37332 5256 37381 5284
rect 37332 5244 37338 5256
rect 37369 5253 37381 5256
rect 37415 5284 37427 5287
rect 37737 5287 37795 5293
rect 37737 5284 37749 5287
rect 37415 5256 37749 5284
rect 37415 5253 37427 5256
rect 37369 5247 37427 5253
rect 37737 5253 37749 5256
rect 37783 5253 37795 5287
rect 37737 5247 37795 5253
rect 38470 5244 38476 5296
rect 38528 5284 38534 5296
rect 38933 5287 38991 5293
rect 38933 5284 38945 5287
rect 38528 5256 38945 5284
rect 38528 5244 38534 5256
rect 38933 5253 38945 5256
rect 38979 5253 38991 5287
rect 38933 5247 38991 5253
rect 49142 5244 49148 5296
rect 49200 5244 49206 5296
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 12802 5216 12808 5228
rect 2179 5188 12808 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 12802 5176 12808 5188
rect 12860 5176 12866 5228
rect 18874 5176 18880 5228
rect 18932 5176 18938 5228
rect 45830 5176 45836 5228
rect 45888 5176 45894 5228
rect 47854 5176 47860 5228
rect 47912 5216 47918 5228
rect 47949 5219 48007 5225
rect 47949 5216 47961 5219
rect 47912 5188 47961 5216
rect 47912 5176 47918 5188
rect 47949 5185 47961 5188
rect 47995 5185 48007 5219
rect 47949 5179 48007 5185
rect 1302 5108 1308 5160
rect 1360 5148 1366 5160
rect 2409 5151 2467 5157
rect 2409 5148 2421 5151
rect 1360 5120 2421 5148
rect 1360 5108 1366 5120
rect 2409 5117 2421 5120
rect 2455 5117 2467 5151
rect 2409 5111 2467 5117
rect 19058 5108 19064 5160
rect 19116 5108 19122 5160
rect 46845 5151 46903 5157
rect 46845 5117 46857 5151
rect 46891 5148 46903 5151
rect 48314 5148 48320 5160
rect 46891 5120 48320 5148
rect 46891 5117 46903 5120
rect 46845 5111 46903 5117
rect 48314 5108 48320 5120
rect 48372 5108 48378 5160
rect 38657 5083 38715 5089
rect 38657 5049 38669 5083
rect 38703 5080 38715 5083
rect 40034 5080 40040 5092
rect 38703 5052 40040 5080
rect 38703 5049 38715 5052
rect 38657 5043 38715 5049
rect 40034 5040 40040 5052
rect 40092 5040 40098 5092
rect 19521 5015 19579 5021
rect 19521 4981 19533 5015
rect 19567 5012 19579 5015
rect 20622 5012 20628 5024
rect 19567 4984 20628 5012
rect 19567 4981 19579 4984
rect 19521 4975 19579 4981
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 37826 4972 37832 5024
rect 37884 4972 37890 5024
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 1302 4768 1308 4820
rect 1360 4808 1366 4820
rect 2133 4811 2191 4817
rect 2133 4808 2145 4811
rect 1360 4780 2145 4808
rect 1360 4768 1366 4780
rect 2133 4777 2145 4780
rect 2179 4777 2191 4811
rect 24118 4808 24124 4820
rect 2133 4771 2191 4777
rect 22066 4780 24124 4808
rect 1765 4743 1823 4749
rect 1765 4709 1777 4743
rect 1811 4740 1823 4743
rect 22066 4740 22094 4780
rect 24118 4768 24124 4780
rect 24176 4768 24182 4820
rect 37826 4768 37832 4820
rect 37884 4808 37890 4820
rect 47118 4808 47124 4820
rect 37884 4780 47124 4808
rect 37884 4768 37890 4780
rect 47118 4768 47124 4780
rect 47176 4768 47182 4820
rect 1811 4712 22094 4740
rect 22557 4743 22615 4749
rect 1811 4709 1823 4712
rect 1765 4703 1823 4709
rect 22557 4709 22569 4743
rect 22603 4740 22615 4743
rect 26142 4740 26148 4752
rect 22603 4712 26148 4740
rect 22603 4709 22615 4712
rect 22557 4703 22615 4709
rect 26142 4700 26148 4712
rect 26200 4700 26206 4752
rect 36998 4700 37004 4752
rect 37056 4740 37062 4752
rect 37056 4712 37412 4740
rect 37056 4700 37062 4712
rect 19242 4632 19248 4684
rect 19300 4672 19306 4684
rect 20441 4675 20499 4681
rect 20441 4672 20453 4675
rect 19300 4644 20453 4672
rect 19300 4632 19306 4644
rect 20441 4641 20453 4644
rect 20487 4641 20499 4675
rect 20441 4635 20499 4641
rect 21726 4632 21732 4684
rect 21784 4672 21790 4684
rect 21913 4675 21971 4681
rect 21913 4672 21925 4675
rect 21784 4644 21925 4672
rect 21784 4632 21790 4644
rect 21913 4641 21925 4644
rect 21959 4641 21971 4675
rect 22922 4672 22928 4684
rect 21913 4635 21971 4641
rect 22020 4644 22928 4672
rect 1302 4564 1308 4616
rect 1360 4604 1366 4616
rect 1581 4607 1639 4613
rect 1581 4604 1593 4607
rect 1360 4576 1593 4604
rect 1360 4564 1366 4576
rect 1581 4573 1593 4576
rect 1627 4604 1639 4607
rect 2317 4607 2375 4613
rect 2317 4604 2329 4607
rect 1627 4576 2329 4604
rect 1627 4573 1639 4576
rect 1581 4567 1639 4573
rect 2317 4573 2329 4576
rect 2363 4573 2375 4607
rect 2317 4567 2375 4573
rect 19978 4564 19984 4616
rect 20036 4604 20042 4616
rect 20625 4607 20683 4613
rect 20625 4604 20637 4607
rect 20036 4576 20637 4604
rect 20036 4564 20042 4576
rect 20625 4573 20637 4576
rect 20671 4604 20683 4607
rect 22020 4604 22048 4644
rect 22922 4632 22928 4644
rect 22980 4632 22986 4684
rect 23198 4632 23204 4684
rect 23256 4672 23262 4684
rect 26789 4675 26847 4681
rect 26789 4672 26801 4675
rect 23256 4644 26801 4672
rect 23256 4632 23262 4644
rect 26789 4641 26801 4644
rect 26835 4641 26847 4675
rect 26789 4635 26847 4641
rect 27246 4632 27252 4684
rect 27304 4672 27310 4684
rect 36817 4675 36875 4681
rect 36817 4672 36829 4675
rect 27304 4644 36829 4672
rect 27304 4632 27310 4644
rect 36817 4641 36829 4644
rect 36863 4672 36875 4675
rect 37384 4672 37412 4712
rect 40218 4700 40224 4752
rect 40276 4740 40282 4752
rect 46477 4743 46535 4749
rect 46477 4740 46489 4743
rect 40276 4712 46489 4740
rect 40276 4700 40282 4712
rect 46477 4709 46489 4712
rect 46523 4709 46535 4743
rect 46477 4703 46535 4709
rect 47213 4675 47271 4681
rect 47213 4672 47225 4675
rect 36863 4644 37320 4672
rect 37384 4644 47225 4672
rect 36863 4641 36875 4644
rect 36817 4635 36875 4641
rect 20671 4576 22048 4604
rect 20671 4573 20683 4576
rect 20625 4567 20683 4573
rect 22094 4564 22100 4616
rect 22152 4564 22158 4616
rect 23084 4607 23142 4613
rect 23084 4604 23096 4607
rect 22388 4576 23096 4604
rect 19058 4496 19064 4548
rect 19116 4536 19122 4548
rect 22388 4536 22416 4576
rect 23084 4573 23096 4576
rect 23130 4604 23142 4607
rect 23566 4604 23572 4616
rect 23130 4576 23572 4604
rect 23130 4573 23142 4576
rect 23084 4567 23142 4573
rect 23566 4564 23572 4576
rect 23624 4564 23630 4616
rect 26973 4607 27031 4613
rect 26973 4573 26985 4607
rect 27019 4604 27031 4607
rect 32766 4604 32772 4616
rect 27019 4576 32772 4604
rect 27019 4573 27031 4576
rect 26973 4567 27031 4573
rect 32766 4564 32772 4576
rect 32824 4564 32830 4616
rect 37292 4613 37320 4644
rect 47213 4641 47225 4644
rect 47259 4641 47271 4675
rect 47213 4635 47271 4641
rect 49145 4675 49203 4681
rect 49145 4641 49157 4675
rect 49191 4672 49203 4675
rect 49418 4672 49424 4684
rect 49191 4644 49424 4672
rect 49191 4641 49203 4644
rect 49145 4635 49203 4641
rect 49418 4632 49424 4644
rect 49476 4632 49482 4684
rect 37277 4607 37335 4613
rect 37277 4573 37289 4607
rect 37323 4573 37335 4607
rect 37277 4567 37335 4573
rect 47302 4564 47308 4616
rect 47360 4604 47366 4616
rect 47949 4607 48007 4613
rect 47949 4604 47961 4607
rect 47360 4576 47961 4604
rect 47360 4564 47366 4576
rect 47949 4573 47961 4576
rect 47995 4573 48007 4607
rect 47949 4567 48007 4573
rect 25133 4539 25191 4545
rect 25133 4536 25145 4539
rect 19116 4508 22416 4536
rect 22480 4508 25145 4536
rect 19116 4496 19122 4508
rect 21085 4471 21143 4477
rect 21085 4437 21097 4471
rect 21131 4468 21143 4471
rect 21266 4468 21272 4480
rect 21131 4440 21272 4468
rect 21131 4437 21143 4440
rect 21085 4431 21143 4437
rect 21266 4428 21272 4440
rect 21324 4428 21330 4480
rect 21450 4428 21456 4480
rect 21508 4468 21514 4480
rect 21818 4468 21824 4480
rect 21508 4440 21824 4468
rect 21508 4428 21514 4440
rect 21818 4428 21824 4440
rect 21876 4468 21882 4480
rect 22480 4468 22508 4508
rect 25133 4505 25145 4508
rect 25179 4505 25191 4539
rect 25133 4499 25191 4505
rect 27062 4496 27068 4548
rect 27120 4536 27126 4548
rect 38013 4539 38071 4545
rect 38013 4536 38025 4539
rect 27120 4508 38025 4536
rect 27120 4496 27126 4508
rect 38013 4505 38025 4508
rect 38059 4536 38071 4539
rect 38473 4539 38531 4545
rect 38473 4536 38485 4539
rect 38059 4508 38485 4536
rect 38059 4505 38071 4508
rect 38013 4499 38071 4505
rect 38473 4505 38485 4508
rect 38519 4505 38531 4539
rect 38473 4499 38531 4505
rect 46661 4539 46719 4545
rect 46661 4505 46673 4539
rect 46707 4505 46719 4539
rect 46661 4499 46719 4505
rect 47397 4539 47455 4545
rect 47397 4505 47409 4539
rect 47443 4536 47455 4539
rect 47670 4536 47676 4548
rect 47443 4508 47676 4536
rect 47443 4505 47455 4508
rect 47397 4499 47455 4505
rect 21876 4440 22508 4468
rect 23155 4471 23213 4477
rect 21876 4428 21882 4440
rect 23155 4437 23167 4471
rect 23201 4468 23213 4471
rect 25866 4468 25872 4480
rect 23201 4440 25872 4468
rect 23201 4437 23213 4440
rect 23155 4431 23213 4437
rect 25866 4428 25872 4440
rect 25924 4428 25930 4480
rect 37366 4428 37372 4480
rect 37424 4428 37430 4480
rect 38105 4471 38163 4477
rect 38105 4437 38117 4471
rect 38151 4468 38163 4471
rect 39758 4468 39764 4480
rect 38151 4440 39764 4468
rect 38151 4437 38163 4440
rect 38105 4431 38163 4437
rect 39758 4428 39764 4440
rect 39816 4428 39822 4480
rect 46201 4471 46259 4477
rect 46201 4437 46213 4471
rect 46247 4468 46259 4471
rect 46676 4468 46704 4499
rect 47670 4496 47676 4508
rect 47728 4496 47734 4548
rect 49786 4468 49792 4480
rect 46247 4440 49792 4468
rect 46247 4437 46259 4440
rect 46201 4431 46259 4437
rect 49786 4428 49792 4440
rect 49844 4428 49850 4480
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 2501 4267 2559 4273
rect 2501 4233 2513 4267
rect 2547 4233 2559 4267
rect 2501 4227 2559 4233
rect 1394 4156 1400 4208
rect 1452 4196 1458 4208
rect 1673 4199 1731 4205
rect 1673 4196 1685 4199
rect 1452 4168 1685 4196
rect 1452 4156 1458 4168
rect 1673 4165 1685 4168
rect 1719 4196 1731 4199
rect 1719 4168 2452 4196
rect 1719 4165 1731 4168
rect 1673 4159 1731 4165
rect 2317 4131 2375 4137
rect 2317 4128 2329 4131
rect 1780 4100 2329 4128
rect 1302 3952 1308 4004
rect 1360 3992 1366 4004
rect 1780 3992 1808 4100
rect 2317 4097 2329 4100
rect 2363 4097 2375 4131
rect 2317 4091 2375 4097
rect 2424 4060 2452 4168
rect 2516 4128 2544 4227
rect 37366 4224 37372 4276
rect 37424 4264 37430 4276
rect 45646 4264 45652 4276
rect 37424 4236 45652 4264
rect 37424 4224 37430 4236
rect 45646 4224 45652 4236
rect 45704 4224 45710 4276
rect 22094 4156 22100 4208
rect 22152 4196 22158 4208
rect 22152 4168 23647 4196
rect 22152 4156 22158 4168
rect 15654 4128 15660 4140
rect 2516 4100 15660 4128
rect 15654 4088 15660 4100
rect 15712 4088 15718 4140
rect 22348 4130 22406 4136
rect 22348 4096 22360 4130
rect 22394 4127 22406 4130
rect 22394 4099 22462 4127
rect 22394 4096 22406 4099
rect 22348 4090 22406 4096
rect 3053 4063 3111 4069
rect 3053 4060 3065 4063
rect 2424 4032 3065 4060
rect 3053 4029 3065 4032
rect 3099 4029 3111 4063
rect 3053 4023 3111 4029
rect 1360 3964 1808 3992
rect 1360 3952 1366 3964
rect 1780 3924 1808 3964
rect 1857 3995 1915 4001
rect 1857 3961 1869 3995
rect 1903 3992 1915 3995
rect 1903 3964 6914 3992
rect 1903 3961 1915 3964
rect 1857 3955 1915 3961
rect 2869 3927 2927 3933
rect 2869 3924 2881 3927
rect 1780 3896 2881 3924
rect 2869 3893 2881 3896
rect 2915 3893 2927 3927
rect 6886 3924 6914 3964
rect 17954 3952 17960 4004
rect 18012 3992 18018 4004
rect 18322 3992 18328 4004
rect 18012 3964 18328 3992
rect 18012 3952 18018 3964
rect 18322 3952 18328 3964
rect 18380 3992 18386 4004
rect 22434 3992 22462 4099
rect 22922 4088 22928 4140
rect 22980 4137 22986 4140
rect 22980 4131 23018 4137
rect 23006 4097 23018 4131
rect 22980 4091 23018 4097
rect 23063 4131 23121 4137
rect 23063 4097 23075 4131
rect 23109 4128 23121 4131
rect 23198 4128 23204 4140
rect 23109 4100 23204 4128
rect 23109 4097 23121 4100
rect 23063 4091 23121 4097
rect 22980 4088 23003 4091
rect 23198 4088 23204 4100
rect 23256 4088 23262 4140
rect 23619 4137 23647 4168
rect 25866 4156 25872 4208
rect 25924 4156 25930 4208
rect 23604 4131 23662 4137
rect 23604 4097 23616 4131
rect 23650 4097 23662 4131
rect 23604 4091 23662 4097
rect 26053 4131 26111 4137
rect 26053 4097 26065 4131
rect 26099 4128 26111 4131
rect 27614 4128 27620 4140
rect 26099 4100 27620 4128
rect 26099 4097 26111 4100
rect 26053 4091 26111 4097
rect 27614 4088 27620 4100
rect 27672 4088 27678 4140
rect 45830 4088 45836 4140
rect 45888 4088 45894 4140
rect 46934 4088 46940 4140
rect 46992 4128 46998 4140
rect 47949 4131 48007 4137
rect 47949 4128 47961 4131
rect 46992 4100 47961 4128
rect 46992 4088 46998 4100
rect 47949 4097 47961 4100
rect 47995 4097 48007 4131
rect 47949 4091 48007 4097
rect 49145 4131 49203 4137
rect 49145 4097 49157 4131
rect 49191 4128 49203 4131
rect 49326 4128 49332 4140
rect 49191 4100 49332 4128
rect 49191 4097 49203 4100
rect 49145 4091 49203 4097
rect 49326 4088 49332 4100
rect 49384 4088 49390 4140
rect 22975 4060 23003 4088
rect 23290 4060 23296 4072
rect 22975 4032 23296 4060
rect 23290 4020 23296 4032
rect 23348 4020 23354 4072
rect 24854 4020 24860 4072
rect 24912 4020 24918 4072
rect 25774 4020 25780 4072
rect 25832 4060 25838 4072
rect 27157 4063 27215 4069
rect 27157 4060 27169 4063
rect 25832 4032 27169 4060
rect 25832 4020 25838 4032
rect 27157 4029 27169 4032
rect 27203 4029 27215 4063
rect 27157 4023 27215 4029
rect 28813 4063 28871 4069
rect 28813 4029 28825 4063
rect 28859 4029 28871 4063
rect 28813 4023 28871 4029
rect 28997 4063 29055 4069
rect 28997 4029 29009 4063
rect 29043 4060 29055 4063
rect 32858 4060 32864 4072
rect 29043 4032 32864 4060
rect 29043 4029 29055 4032
rect 28997 4023 29055 4029
rect 23707 3995 23765 4001
rect 18380 3964 22968 3992
rect 18380 3952 18386 3964
rect 21634 3924 21640 3936
rect 6886 3896 21640 3924
rect 2869 3887 2927 3893
rect 21634 3884 21640 3896
rect 21692 3884 21698 3936
rect 22419 3927 22477 3933
rect 22419 3893 22431 3927
rect 22465 3924 22477 3927
rect 22830 3924 22836 3936
rect 22465 3896 22836 3924
rect 22465 3893 22477 3896
rect 22419 3887 22477 3893
rect 22830 3884 22836 3896
rect 22888 3884 22894 3936
rect 22940 3924 22968 3964
rect 23707 3961 23719 3995
rect 23753 3992 23765 3995
rect 28828 3992 28856 4023
rect 32858 4020 32864 4032
rect 32916 4020 32922 4072
rect 46658 4020 46664 4072
rect 46716 4020 46722 4072
rect 23753 3964 28856 3992
rect 23753 3961 23765 3964
rect 23707 3955 23765 3961
rect 27522 3924 27528 3936
rect 22940 3896 27528 3924
rect 27522 3884 27528 3896
rect 27580 3884 27586 3936
rect 47670 3884 47676 3936
rect 47728 3884 47734 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 7524 3692 16620 3720
rect 7524 3680 7530 3692
rect 3326 3612 3332 3664
rect 3384 3652 3390 3664
rect 3384 3624 13860 3652
rect 3384 3612 3390 3624
rect 2133 3587 2191 3593
rect 2133 3553 2145 3587
rect 2179 3584 2191 3587
rect 12434 3584 12440 3596
rect 2179 3556 12440 3584
rect 2179 3553 2191 3556
rect 2133 3547 2191 3553
rect 12434 3544 12440 3556
rect 12492 3544 12498 3596
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 2409 3519 2467 3525
rect 2409 3516 2421 3519
rect 1360 3488 2421 3516
rect 1360 3476 1366 3488
rect 2409 3485 2421 3488
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 13832 3380 13860 3624
rect 16592 3584 16620 3692
rect 22002 3680 22008 3732
rect 22060 3720 22066 3732
rect 23017 3723 23075 3729
rect 23017 3720 23029 3723
rect 22060 3692 23029 3720
rect 22060 3680 22066 3692
rect 23017 3689 23029 3692
rect 23063 3689 23075 3723
rect 23017 3683 23075 3689
rect 23032 3652 23060 3683
rect 23566 3680 23572 3732
rect 23624 3680 23630 3732
rect 23937 3723 23995 3729
rect 23937 3689 23949 3723
rect 23983 3720 23995 3723
rect 25958 3720 25964 3732
rect 23983 3692 25964 3720
rect 23983 3689 23995 3692
rect 23937 3683 23995 3689
rect 25958 3680 25964 3692
rect 26016 3680 26022 3732
rect 24946 3652 24952 3664
rect 23032 3624 24952 3652
rect 24946 3612 24952 3624
rect 25004 3652 25010 3664
rect 26326 3652 26332 3664
rect 25004 3624 26332 3652
rect 25004 3612 25010 3624
rect 26326 3612 26332 3624
rect 26384 3652 26390 3664
rect 29638 3652 29644 3664
rect 26384 3624 29644 3652
rect 26384 3612 26390 3624
rect 29638 3612 29644 3624
rect 29696 3612 29702 3664
rect 33410 3612 33416 3664
rect 33468 3652 33474 3664
rect 45373 3655 45431 3661
rect 45373 3652 45385 3655
rect 33468 3624 45385 3652
rect 33468 3612 33474 3624
rect 45373 3621 45385 3624
rect 45419 3621 45431 3655
rect 45373 3615 45431 3621
rect 16592 3556 22784 3584
rect 16577 3519 16635 3525
rect 16577 3485 16589 3519
rect 16623 3516 16635 3519
rect 17954 3516 17960 3528
rect 16623 3488 17960 3516
rect 16623 3485 16635 3488
rect 16577 3479 16635 3485
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 20990 3476 20996 3528
rect 21048 3476 21054 3528
rect 13906 3408 13912 3460
rect 13964 3448 13970 3460
rect 16393 3451 16451 3457
rect 16393 3448 16405 3451
rect 13964 3420 16405 3448
rect 13964 3408 13970 3420
rect 16393 3417 16405 3420
rect 16439 3417 16451 3451
rect 16393 3411 16451 3417
rect 19334 3408 19340 3460
rect 19392 3448 19398 3460
rect 21269 3451 21327 3457
rect 21269 3448 21281 3451
rect 19392 3420 21281 3448
rect 19392 3408 19398 3420
rect 21269 3417 21281 3420
rect 21315 3448 21327 3451
rect 21358 3448 21364 3460
rect 21315 3420 21364 3448
rect 21315 3417 21327 3420
rect 21269 3411 21327 3417
rect 21358 3408 21364 3420
rect 21416 3408 21422 3460
rect 22002 3408 22008 3460
rect 22060 3408 22066 3460
rect 22756 3448 22784 3556
rect 22830 3544 22836 3596
rect 22888 3584 22894 3596
rect 26237 3587 26295 3593
rect 26237 3584 26249 3587
rect 22888 3556 26249 3584
rect 22888 3544 22894 3556
rect 26237 3553 26249 3556
rect 26283 3553 26295 3587
rect 26237 3547 26295 3553
rect 26421 3587 26479 3593
rect 26421 3553 26433 3587
rect 26467 3584 26479 3587
rect 28994 3584 29000 3596
rect 26467 3556 29000 3584
rect 26467 3553 26479 3556
rect 26421 3547 26479 3553
rect 28994 3544 29000 3556
rect 29052 3544 29058 3596
rect 40034 3544 40040 3596
rect 40092 3584 40098 3596
rect 40092 3556 46152 3584
rect 40092 3544 40098 3556
rect 23293 3519 23351 3525
rect 23293 3485 23305 3519
rect 23339 3516 23351 3519
rect 24026 3516 24032 3528
rect 23339 3488 24032 3516
rect 23339 3485 23351 3488
rect 23293 3479 23351 3485
rect 24026 3476 24032 3488
rect 24084 3476 24090 3528
rect 28350 3476 28356 3528
rect 28408 3516 28414 3528
rect 39206 3516 39212 3528
rect 28408 3488 39212 3516
rect 28408 3476 28414 3488
rect 39206 3476 39212 3488
rect 39264 3476 39270 3528
rect 45830 3516 45836 3528
rect 41386 3488 45836 3516
rect 23934 3448 23940 3460
rect 22756 3420 23940 3448
rect 23934 3408 23940 3420
rect 23992 3448 23998 3460
rect 24581 3451 24639 3457
rect 24581 3448 24593 3451
rect 23992 3420 24593 3448
rect 23992 3408 23998 3420
rect 24581 3417 24593 3420
rect 24627 3417 24639 3451
rect 36449 3451 36507 3457
rect 36449 3448 36461 3451
rect 24581 3411 24639 3417
rect 31726 3420 36461 3448
rect 21450 3380 21456 3392
rect 13832 3352 21456 3380
rect 21450 3340 21456 3352
rect 21508 3340 21514 3392
rect 22738 3340 22744 3392
rect 22796 3340 22802 3392
rect 23106 3340 23112 3392
rect 23164 3380 23170 3392
rect 31726 3380 31754 3420
rect 36449 3417 36461 3420
rect 36495 3417 36507 3451
rect 36449 3411 36507 3417
rect 36633 3451 36691 3457
rect 36633 3417 36645 3451
rect 36679 3448 36691 3451
rect 41386 3448 41414 3488
rect 45830 3476 45836 3488
rect 45888 3476 45894 3528
rect 46124 3525 46152 3556
rect 49142 3544 49148 3596
rect 49200 3544 49206 3596
rect 46109 3519 46167 3525
rect 46109 3485 46121 3519
rect 46155 3485 46167 3519
rect 46109 3479 46167 3485
rect 47026 3476 47032 3528
rect 47084 3516 47090 3528
rect 47949 3519 48007 3525
rect 47949 3516 47961 3519
rect 47084 3488 47961 3516
rect 47084 3476 47090 3488
rect 47949 3485 47961 3488
rect 47995 3485 48007 3519
rect 47949 3479 48007 3485
rect 36679 3420 41414 3448
rect 45097 3451 45155 3457
rect 36679 3417 36691 3420
rect 36633 3411 36691 3417
rect 45097 3417 45109 3451
rect 45143 3448 45155 3451
rect 45554 3448 45560 3460
rect 45143 3420 45560 3448
rect 45143 3417 45155 3420
rect 45097 3411 45155 3417
rect 23164 3352 31754 3380
rect 36464 3380 36492 3411
rect 45554 3408 45560 3420
rect 45612 3448 45618 3460
rect 47305 3451 47363 3457
rect 45612 3420 45657 3448
rect 45612 3408 45618 3420
rect 47305 3417 47317 3451
rect 47351 3448 47363 3451
rect 48682 3448 48688 3460
rect 47351 3420 48688 3448
rect 47351 3417 47363 3420
rect 47305 3411 47363 3417
rect 48682 3408 48688 3420
rect 48740 3408 48746 3460
rect 36909 3383 36967 3389
rect 36909 3380 36921 3383
rect 36464 3352 36921 3380
rect 23164 3340 23170 3352
rect 36909 3349 36921 3352
rect 36955 3349 36967 3383
rect 36909 3343 36967 3349
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 1302 3136 1308 3188
rect 1360 3176 1366 3188
rect 2133 3179 2191 3185
rect 2133 3176 2145 3179
rect 1360 3148 2145 3176
rect 1360 3136 1366 3148
rect 2133 3145 2145 3148
rect 2179 3145 2191 3179
rect 2133 3139 2191 3145
rect 9861 3179 9919 3185
rect 9861 3145 9873 3179
rect 9907 3145 9919 3179
rect 9861 3139 9919 3145
rect 16301 3179 16359 3185
rect 16301 3145 16313 3179
rect 16347 3176 16359 3179
rect 19334 3176 19340 3188
rect 16347 3148 19340 3176
rect 16347 3145 16359 3148
rect 16301 3139 16359 3145
rect 1302 3000 1308 3052
rect 1360 3040 1366 3052
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 1360 3012 1593 3040
rect 1360 3000 1366 3012
rect 1581 3009 1593 3012
rect 1627 3040 1639 3043
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 1627 3012 2513 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 9674 3000 9680 3052
rect 9732 3000 9738 3052
rect 9876 3040 9904 3139
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 19981 3179 20039 3185
rect 19981 3176 19993 3179
rect 19536 3148 19993 3176
rect 16761 3111 16819 3117
rect 16761 3108 16773 3111
rect 16054 3080 16773 3108
rect 16761 3077 16773 3080
rect 16807 3108 16819 3111
rect 17862 3108 17868 3120
rect 16807 3080 17868 3108
rect 16807 3077 16819 3080
rect 16761 3071 16819 3077
rect 17862 3068 17868 3080
rect 17920 3068 17926 3120
rect 12345 3043 12403 3049
rect 12345 3040 12357 3043
rect 9876 3012 12357 3040
rect 12345 3009 12357 3012
rect 12391 3009 12403 3043
rect 12345 3003 12403 3009
rect 13630 3000 13636 3052
rect 13688 3040 13694 3052
rect 14553 3043 14611 3049
rect 14553 3040 14565 3043
rect 13688 3012 14565 3040
rect 13688 3000 13694 3012
rect 14553 3009 14565 3012
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 17589 3043 17647 3049
rect 17589 3009 17601 3043
rect 17635 3040 17647 3043
rect 19058 3040 19064 3052
rect 17635 3012 19064 3040
rect 17635 3009 17647 3012
rect 17589 3003 17647 3009
rect 19058 3000 19064 3012
rect 19116 3000 19122 3052
rect 19536 3049 19564 3148
rect 19981 3145 19993 3148
rect 20027 3145 20039 3179
rect 19981 3139 20039 3145
rect 21450 3136 21456 3188
rect 21508 3136 21514 3188
rect 28353 3179 28411 3185
rect 28353 3176 28365 3179
rect 24688 3148 28365 3176
rect 24026 3108 24032 3120
rect 20180 3080 22232 3108
rect 20180 3049 20208 3080
rect 22204 3052 22232 3080
rect 23768 3080 24032 3108
rect 19521 3043 19579 3049
rect 19521 3009 19533 3043
rect 19567 3009 19579 3043
rect 19521 3003 19579 3009
rect 20165 3043 20223 3049
rect 20165 3009 20177 3043
rect 20211 3009 20223 3043
rect 20165 3003 20223 3009
rect 20622 3000 20628 3052
rect 20680 3000 20686 3052
rect 21266 3000 21272 3052
rect 21324 3000 21330 3052
rect 22186 3000 22192 3052
rect 22244 3000 22250 3052
rect 23768 3049 23796 3080
rect 24026 3068 24032 3080
rect 24084 3108 24090 3120
rect 24688 3108 24716 3148
rect 28353 3145 28365 3148
rect 28399 3176 28411 3179
rect 37734 3176 37740 3188
rect 28399 3148 37740 3176
rect 28399 3145 28411 3148
rect 28353 3139 28411 3145
rect 24084 3080 24716 3108
rect 24084 3068 24090 3080
rect 24946 3068 24952 3120
rect 25004 3068 25010 3120
rect 22649 3043 22707 3049
rect 22649 3009 22661 3043
rect 22695 3040 22707 3043
rect 23017 3043 23075 3049
rect 23017 3040 23029 3043
rect 22695 3012 23029 3040
rect 22695 3009 22707 3012
rect 22649 3003 22707 3009
rect 23017 3009 23029 3012
rect 23063 3040 23075 3043
rect 23753 3043 23811 3049
rect 23753 3040 23765 3043
rect 23063 3012 23765 3040
rect 23063 3009 23075 3012
rect 23017 3003 23075 3009
rect 23753 3009 23765 3012
rect 23799 3009 23811 3043
rect 23753 3003 23811 3009
rect 26142 3000 26148 3052
rect 26200 3040 26206 3052
rect 26421 3043 26479 3049
rect 26421 3040 26433 3043
rect 26200 3012 26433 3040
rect 26200 3000 26206 3012
rect 26421 3009 26433 3012
rect 26467 3009 26479 3043
rect 26421 3003 26479 3009
rect 27985 3043 28043 3049
rect 27985 3009 27997 3043
rect 28031 3040 28043 3043
rect 28368 3040 28396 3139
rect 37734 3136 37740 3148
rect 37792 3136 37798 3188
rect 29638 3068 29644 3120
rect 29696 3068 29702 3120
rect 49145 3111 49203 3117
rect 49145 3077 49157 3111
rect 49191 3108 49203 3111
rect 49234 3108 49240 3120
rect 49191 3080 49240 3108
rect 49191 3077 49203 3080
rect 49145 3071 49203 3077
rect 49234 3068 49240 3080
rect 49292 3068 49298 3120
rect 28031 3012 28396 3040
rect 28031 3009 28043 3012
rect 27985 3003 28043 3009
rect 28810 3000 28816 3052
rect 28868 3040 28874 3052
rect 28905 3043 28963 3049
rect 28905 3040 28917 3043
rect 28868 3012 28917 3040
rect 28868 3000 28874 3012
rect 28905 3009 28917 3012
rect 28951 3009 28963 3043
rect 28905 3003 28963 3009
rect 39758 3000 39764 3052
rect 39816 3040 39822 3052
rect 43993 3043 44051 3049
rect 43993 3040 44005 3043
rect 39816 3012 44005 3040
rect 39816 3000 39822 3012
rect 43993 3009 44005 3012
rect 44039 3009 44051 3043
rect 43993 3003 44051 3009
rect 45738 3000 45744 3052
rect 45796 3040 45802 3052
rect 45833 3043 45891 3049
rect 45833 3040 45845 3043
rect 45796 3012 45845 3040
rect 45796 3000 45802 3012
rect 45833 3009 45845 3012
rect 45879 3009 45891 3043
rect 45833 3003 45891 3009
rect 47210 3000 47216 3052
rect 47268 3040 47274 3052
rect 47949 3043 48007 3049
rect 47949 3040 47961 3043
rect 47268 3012 47961 3040
rect 47268 3000 47274 3012
rect 47949 3009 47961 3012
rect 47995 3009 48007 3043
rect 47949 3003 48007 3009
rect 12989 2975 13047 2981
rect 12989 2941 13001 2975
rect 13035 2972 13047 2975
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 13035 2944 14841 2972
rect 13035 2941 13047 2944
rect 12989 2935 13047 2941
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 18322 2932 18328 2984
rect 18380 2932 18386 2984
rect 20990 2932 20996 2984
rect 21048 2972 21054 2984
rect 24213 2975 24271 2981
rect 24213 2972 24225 2975
rect 21048 2944 24225 2972
rect 21048 2932 21054 2944
rect 24213 2941 24225 2944
rect 24259 2941 24271 2975
rect 24489 2975 24547 2981
rect 24489 2972 24501 2975
rect 24213 2935 24271 2941
rect 24320 2944 24501 2972
rect 1765 2907 1823 2913
rect 1765 2873 1777 2907
rect 1811 2904 1823 2907
rect 12710 2904 12716 2916
rect 1811 2876 12716 2904
rect 1811 2873 1823 2876
rect 1765 2867 1823 2873
rect 12710 2864 12716 2876
rect 12768 2864 12774 2916
rect 20809 2907 20867 2913
rect 20809 2873 20821 2907
rect 20855 2904 20867 2907
rect 22094 2904 22100 2916
rect 20855 2876 22100 2904
rect 20855 2873 20867 2876
rect 20809 2867 20867 2873
rect 22094 2864 22100 2876
rect 22152 2864 22158 2916
rect 22186 2864 22192 2916
rect 22244 2864 22250 2916
rect 22738 2864 22744 2916
rect 22796 2904 22802 2916
rect 24320 2904 24348 2944
rect 24489 2941 24501 2944
rect 24535 2941 24547 2975
rect 24489 2935 24547 2941
rect 25958 2932 25964 2984
rect 26016 2972 26022 2984
rect 29181 2975 29239 2981
rect 29181 2972 29193 2975
rect 26016 2944 29193 2972
rect 26016 2932 26022 2944
rect 29181 2941 29193 2944
rect 29227 2941 29239 2975
rect 29181 2935 29239 2941
rect 29638 2932 29644 2984
rect 29696 2972 29702 2984
rect 30650 2972 30656 2984
rect 29696 2944 30656 2972
rect 29696 2932 29702 2944
rect 30650 2932 30656 2944
rect 30708 2972 30714 2984
rect 31021 2975 31079 2981
rect 31021 2972 31033 2975
rect 30708 2944 31033 2972
rect 30708 2932 30714 2944
rect 31021 2941 31033 2944
rect 31067 2941 31079 2975
rect 31021 2935 31079 2941
rect 45189 2975 45247 2981
rect 45189 2941 45201 2975
rect 45235 2972 45247 2975
rect 46750 2972 46756 2984
rect 45235 2944 46756 2972
rect 45235 2941 45247 2944
rect 45189 2935 45247 2941
rect 46750 2932 46756 2944
rect 46808 2932 46814 2984
rect 46842 2932 46848 2984
rect 46900 2932 46906 2984
rect 22796 2876 24348 2904
rect 22796 2864 22802 2876
rect 2314 2796 2320 2848
rect 2372 2796 2378 2848
rect 2774 2796 2780 2848
rect 2832 2796 2838 2848
rect 17402 2796 17408 2848
rect 17460 2796 17466 2848
rect 21358 2796 21364 2848
rect 21416 2836 21422 2848
rect 22373 2839 22431 2845
rect 22373 2836 22385 2839
rect 21416 2808 22385 2836
rect 21416 2796 21422 2808
rect 22373 2805 22385 2808
rect 22419 2805 22431 2839
rect 22373 2799 22431 2805
rect 23290 2796 23296 2848
rect 23348 2796 23354 2848
rect 23492 2845 23520 2876
rect 27522 2864 27528 2916
rect 27580 2864 27586 2916
rect 38286 2904 38292 2916
rect 27908 2876 29040 2904
rect 23477 2839 23535 2845
rect 23477 2805 23489 2839
rect 23523 2805 23535 2839
rect 23477 2799 23535 2805
rect 26605 2839 26663 2845
rect 26605 2805 26617 2839
rect 26651 2836 26663 2839
rect 27154 2836 27160 2848
rect 26651 2808 27160 2836
rect 26651 2805 26663 2808
rect 26605 2799 26663 2805
rect 27154 2796 27160 2808
rect 27212 2796 27218 2848
rect 27908 2845 27936 2876
rect 27893 2839 27951 2845
rect 27893 2805 27905 2839
rect 27939 2805 27951 2839
rect 29012 2836 29040 2876
rect 30668 2876 38292 2904
rect 30668 2845 30696 2876
rect 38286 2864 38292 2876
rect 38344 2864 38350 2916
rect 30653 2839 30711 2845
rect 30653 2836 30665 2839
rect 29012 2808 30665 2836
rect 27893 2799 27951 2805
rect 30653 2805 30665 2808
rect 30699 2805 30711 2839
rect 30653 2799 30711 2805
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 2501 2635 2559 2641
rect 2501 2601 2513 2635
rect 2547 2632 2559 2635
rect 2547 2604 16574 2632
rect 2547 2601 2559 2604
rect 2501 2595 2559 2601
rect 1765 2567 1823 2573
rect 1765 2533 1777 2567
rect 1811 2533 1823 2567
rect 1765 2527 1823 2533
rect 3237 2567 3295 2573
rect 3237 2533 3249 2567
rect 3283 2564 3295 2567
rect 3283 2536 6914 2564
rect 3283 2533 3295 2536
rect 3237 2527 3295 2533
rect 1780 2496 1808 2527
rect 6886 2496 6914 2536
rect 9674 2524 9680 2576
rect 9732 2564 9738 2576
rect 10321 2567 10379 2573
rect 10321 2564 10333 2567
rect 9732 2536 10333 2564
rect 9732 2524 9738 2536
rect 10321 2533 10333 2536
rect 10367 2533 10379 2567
rect 16546 2564 16574 2604
rect 24026 2592 24032 2644
rect 24084 2592 24090 2644
rect 26326 2592 26332 2644
rect 26384 2592 26390 2644
rect 27614 2592 27620 2644
rect 27672 2592 27678 2644
rect 28994 2592 29000 2644
rect 29052 2592 29058 2644
rect 32858 2592 32864 2644
rect 32916 2632 32922 2644
rect 35069 2635 35127 2641
rect 35069 2632 35081 2635
rect 32916 2604 35081 2632
rect 32916 2592 32922 2604
rect 35069 2601 35081 2604
rect 35115 2601 35127 2635
rect 35069 2595 35127 2601
rect 22462 2564 22468 2576
rect 16546 2536 22468 2564
rect 10321 2527 10379 2533
rect 22462 2524 22468 2536
rect 22520 2524 22526 2576
rect 27632 2564 27660 2592
rect 30837 2567 30895 2573
rect 30837 2564 30849 2567
rect 27632 2536 30849 2564
rect 30837 2533 30849 2536
rect 30883 2533 30895 2567
rect 30837 2527 30895 2533
rect 32766 2524 32772 2576
rect 32824 2564 32830 2576
rect 32953 2567 33011 2573
rect 32953 2564 32965 2567
rect 32824 2536 32965 2564
rect 32824 2524 32830 2536
rect 32953 2533 32965 2536
rect 32999 2533 33011 2567
rect 32953 2527 33011 2533
rect 34422 2524 34428 2576
rect 34480 2564 34486 2576
rect 34480 2536 43852 2564
rect 34480 2524 34486 2536
rect 12250 2496 12256 2508
rect 1780 2468 4384 2496
rect 6886 2468 12256 2496
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 1360 2400 1593 2428
rect 1360 2388 1366 2400
rect 1581 2397 1593 2400
rect 1627 2428 1639 2431
rect 2774 2428 2780 2440
rect 1627 2400 2780 2428
rect 1627 2397 1639 2400
rect 1581 2391 1639 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 3053 2431 3111 2437
rect 3053 2428 3065 2431
rect 2884 2400 3065 2428
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 2314 2360 2320 2372
rect 1268 2332 2320 2360
rect 1268 2320 1274 2332
rect 2314 2320 2320 2332
rect 2372 2360 2378 2372
rect 2409 2363 2467 2369
rect 2409 2360 2421 2363
rect 2372 2332 2421 2360
rect 2372 2320 2378 2332
rect 2409 2329 2421 2332
rect 2455 2329 2467 2363
rect 2409 2323 2467 2329
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 2884 2292 2912 2400
rect 3053 2397 3065 2400
rect 3099 2428 3111 2431
rect 3513 2431 3571 2437
rect 3513 2428 3525 2431
rect 3099 2400 3525 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 3513 2397 3525 2400
rect 3559 2397 3571 2431
rect 3513 2391 3571 2397
rect 4356 2360 4384 2468
rect 12250 2456 12256 2468
rect 12308 2456 12314 2508
rect 19978 2496 19984 2508
rect 19306 2468 19984 2496
rect 9582 2388 9588 2440
rect 9640 2428 9646 2440
rect 9677 2431 9735 2437
rect 9677 2428 9689 2431
rect 9640 2400 9689 2428
rect 9640 2388 9646 2400
rect 9677 2397 9689 2400
rect 9723 2397 9735 2431
rect 9677 2391 9735 2397
rect 13173 2431 13231 2437
rect 13173 2397 13185 2431
rect 13219 2428 13231 2431
rect 13906 2428 13912 2440
rect 13219 2400 13912 2428
rect 13219 2397 13231 2400
rect 13173 2391 13231 2397
rect 13906 2388 13912 2400
rect 13964 2388 13970 2440
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2428 15715 2431
rect 17402 2428 17408 2440
rect 15703 2400 17408 2428
rect 15703 2397 15715 2400
rect 15657 2391 15715 2397
rect 17402 2388 17408 2400
rect 17460 2388 17466 2440
rect 18233 2431 18291 2437
rect 18233 2397 18245 2431
rect 18279 2428 18291 2431
rect 18877 2431 18935 2437
rect 18279 2400 18736 2428
rect 18279 2397 18291 2400
rect 18233 2391 18291 2397
rect 4356 2332 10824 2360
rect 1360 2264 2912 2292
rect 9401 2295 9459 2301
rect 1360 2252 1366 2264
rect 9401 2261 9413 2295
rect 9447 2292 9459 2295
rect 9582 2292 9588 2304
rect 9447 2264 9588 2292
rect 9447 2261 9459 2264
rect 9401 2255 9459 2261
rect 9582 2252 9588 2264
rect 9640 2252 9646 2304
rect 10796 2292 10824 2332
rect 11698 2320 11704 2372
rect 11756 2360 11762 2372
rect 11977 2363 12035 2369
rect 11977 2360 11989 2363
rect 11756 2332 11989 2360
rect 11756 2320 11762 2332
rect 11977 2329 11989 2332
rect 12023 2329 12035 2363
rect 11977 2323 12035 2329
rect 13814 2320 13820 2372
rect 13872 2360 13878 2372
rect 14461 2363 14519 2369
rect 14461 2360 14473 2363
rect 13872 2332 14473 2360
rect 13872 2320 13878 2332
rect 14461 2329 14473 2332
rect 14507 2329 14519 2363
rect 14461 2323 14519 2329
rect 15930 2320 15936 2372
rect 15988 2360 15994 2372
rect 17037 2363 17095 2369
rect 17037 2360 17049 2363
rect 15988 2332 17049 2360
rect 15988 2320 15994 2332
rect 17037 2329 17049 2332
rect 17083 2329 17095 2363
rect 17037 2323 17095 2329
rect 14734 2292 14740 2304
rect 10796 2264 14740 2292
rect 14734 2252 14740 2264
rect 14792 2252 14798 2304
rect 18708 2301 18736 2400
rect 18877 2397 18889 2431
rect 18923 2428 18935 2431
rect 19306 2428 19334 2468
rect 19978 2456 19984 2468
rect 20036 2456 20042 2508
rect 20162 2456 20168 2508
rect 20220 2496 20226 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20220 2468 20545 2496
rect 20220 2456 20226 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 22278 2456 22284 2508
rect 22336 2496 22342 2508
rect 22833 2499 22891 2505
rect 22833 2496 22845 2499
rect 22336 2468 22845 2496
rect 22336 2456 22342 2468
rect 22833 2465 22845 2468
rect 22879 2465 22891 2499
rect 22833 2459 22891 2465
rect 24394 2456 24400 2508
rect 24452 2496 24458 2508
rect 25041 2499 25099 2505
rect 25041 2496 25053 2499
rect 24452 2468 25053 2496
rect 24452 2456 24458 2468
rect 25041 2465 25053 2468
rect 25087 2465 25099 2499
rect 25041 2459 25099 2465
rect 26510 2456 26516 2508
rect 26568 2496 26574 2508
rect 27617 2499 27675 2505
rect 27617 2496 27629 2499
rect 26568 2468 27629 2496
rect 26568 2456 26574 2468
rect 27617 2465 27629 2468
rect 27663 2465 27675 2499
rect 27617 2459 27675 2465
rect 37734 2456 37740 2508
rect 37792 2456 37798 2508
rect 41322 2456 41328 2508
rect 41380 2496 41386 2508
rect 43824 2505 43852 2536
rect 41417 2499 41475 2505
rect 41417 2496 41429 2499
rect 41380 2468 41429 2496
rect 41380 2456 41386 2468
rect 41417 2465 41429 2468
rect 41463 2465 41475 2499
rect 41417 2459 41475 2465
rect 43809 2499 43867 2505
rect 43809 2465 43821 2499
rect 43855 2465 43867 2499
rect 43809 2459 43867 2465
rect 49142 2456 49148 2508
rect 49200 2456 49206 2508
rect 18923 2400 19334 2428
rect 18923 2397 18935 2400
rect 18877 2391 18935 2397
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 20073 2431 20131 2437
rect 20073 2428 20085 2431
rect 19628 2400 20085 2428
rect 19628 2301 19656 2400
rect 20073 2397 20085 2400
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 22094 2388 22100 2440
rect 22152 2428 22158 2440
rect 22373 2431 22431 2437
rect 22373 2428 22385 2431
rect 22152 2400 22385 2428
rect 22152 2388 22158 2400
rect 22373 2397 22385 2400
rect 22419 2397 22431 2431
rect 22373 2391 22431 2397
rect 24581 2431 24639 2437
rect 24581 2397 24593 2431
rect 24627 2397 24639 2431
rect 24581 2391 24639 2397
rect 21450 2320 21456 2372
rect 21508 2360 21514 2372
rect 24596 2360 24624 2391
rect 27154 2388 27160 2440
rect 27212 2388 27218 2440
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29181 2431 29239 2437
rect 29181 2428 29193 2431
rect 29052 2400 29193 2428
rect 29052 2388 29058 2400
rect 29181 2397 29193 2400
rect 29227 2428 29239 2431
rect 29549 2431 29607 2437
rect 29549 2428 29561 2431
rect 29227 2400 29561 2428
rect 29227 2397 29239 2400
rect 29181 2391 29239 2397
rect 29549 2397 29561 2400
rect 29595 2397 29607 2431
rect 29549 2391 29607 2397
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30800 2400 31033 2428
rect 30800 2388 30806 2400
rect 31021 2397 31033 2400
rect 31067 2428 31079 2431
rect 31297 2431 31355 2437
rect 31297 2428 31309 2431
rect 31067 2400 31309 2428
rect 31067 2397 31079 2400
rect 31021 2391 31079 2397
rect 31297 2397 31309 2400
rect 31343 2397 31355 2431
rect 31297 2391 31355 2397
rect 33134 2388 33140 2440
rect 33192 2428 33198 2440
rect 33413 2431 33471 2437
rect 33413 2428 33425 2431
rect 33192 2400 33425 2428
rect 33192 2388 33198 2400
rect 33413 2397 33425 2400
rect 33459 2397 33471 2431
rect 33413 2391 33471 2397
rect 34974 2388 34980 2440
rect 35032 2428 35038 2440
rect 35253 2431 35311 2437
rect 35253 2428 35265 2431
rect 35032 2400 35265 2428
rect 35032 2388 35038 2400
rect 35253 2397 35265 2400
rect 35299 2428 35311 2431
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 35299 2400 35541 2428
rect 35299 2397 35311 2400
rect 35253 2391 35311 2397
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 35529 2391 35587 2397
rect 37108 2400 37473 2428
rect 21508 2332 24624 2360
rect 21508 2320 21514 2332
rect 37108 2304 37136 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 38286 2388 38292 2440
rect 38344 2428 38350 2440
rect 40681 2431 40739 2437
rect 40681 2428 40693 2431
rect 38344 2400 40693 2428
rect 38344 2388 38350 2400
rect 40681 2397 40693 2400
rect 40727 2397 40739 2431
rect 43533 2431 43591 2437
rect 43533 2428 43545 2431
rect 40681 2391 40739 2397
rect 43456 2400 43545 2428
rect 43456 2304 43484 2400
rect 43533 2397 43545 2400
rect 43579 2397 43591 2431
rect 43533 2391 43591 2397
rect 45646 2388 45652 2440
rect 45704 2428 45710 2440
rect 45833 2431 45891 2437
rect 45833 2428 45845 2431
rect 45704 2400 45845 2428
rect 45704 2388 45710 2400
rect 45833 2397 45845 2400
rect 45879 2397 45891 2431
rect 45833 2391 45891 2397
rect 47118 2388 47124 2440
rect 47176 2428 47182 2440
rect 47949 2431 48007 2437
rect 47949 2428 47961 2431
rect 47176 2400 47961 2428
rect 47176 2388 47182 2400
rect 47949 2397 47961 2400
rect 47995 2397 48007 2431
rect 47949 2391 48007 2397
rect 47029 2363 47087 2369
rect 47029 2329 47041 2363
rect 47075 2360 47087 2363
rect 48498 2360 48504 2372
rect 47075 2332 48504 2360
rect 47075 2329 47087 2332
rect 47029 2323 47087 2329
rect 48498 2320 48504 2332
rect 48556 2320 48562 2372
rect 18693 2295 18751 2301
rect 18693 2261 18705 2295
rect 18739 2261 18751 2295
rect 18693 2255 18751 2261
rect 19613 2295 19671 2301
rect 19613 2261 19625 2295
rect 19659 2261 19671 2295
rect 19613 2255 19671 2261
rect 37090 2252 37096 2304
rect 37148 2252 37154 2304
rect 43257 2295 43315 2301
rect 43257 2261 43269 2295
rect 43303 2292 43315 2295
rect 43438 2292 43444 2304
rect 43303 2264 43444 2292
rect 43303 2261 43315 2264
rect 43257 2255 43315 2261
rect 43438 2252 43444 2264
rect 43496 2252 43502 2304
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
<< via1 >>
rect 30564 25236 30616 25288
rect 37924 25236 37976 25288
rect 3424 24828 3476 24880
rect 9772 24828 9824 24880
rect 3608 24760 3660 24812
rect 5908 24760 5960 24812
rect 17224 24760 17276 24812
rect 24032 24760 24084 24812
rect 24768 24760 24820 24812
rect 30380 24760 30432 24812
rect 18880 24692 18932 24744
rect 27252 24692 27304 24744
rect 29920 24692 29972 24744
rect 33324 24828 33376 24880
rect 39580 24828 39632 24880
rect 45284 24828 45336 24880
rect 38936 24760 38988 24812
rect 42064 24760 42116 24812
rect 22560 24624 22612 24676
rect 26332 24624 26384 24676
rect 26424 24624 26476 24676
rect 34612 24692 34664 24744
rect 34888 24692 34940 24744
rect 40316 24692 40368 24744
rect 33140 24624 33192 24676
rect 39948 24624 40000 24676
rect 40224 24624 40276 24676
rect 43996 24624 44048 24676
rect 20536 24556 20588 24608
rect 29736 24556 29788 24608
rect 29828 24556 29880 24608
rect 31576 24556 31628 24608
rect 31852 24556 31904 24608
rect 39488 24556 39540 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 3516 24216 3568 24268
rect 6736 24216 6788 24268
rect 3884 24148 3936 24200
rect 4620 24191 4672 24200
rect 4620 24157 4629 24191
rect 4629 24157 4663 24191
rect 4663 24157 4672 24191
rect 4620 24148 4672 24157
rect 9588 24352 9640 24404
rect 12348 24352 12400 24404
rect 17224 24352 17276 24404
rect 18604 24352 18656 24404
rect 8668 24216 8720 24268
rect 11888 24284 11940 24336
rect 15476 24284 15528 24336
rect 16028 24284 16080 24336
rect 7196 24148 7248 24200
rect 7932 24148 7984 24200
rect 13820 24216 13872 24268
rect 17684 24216 17736 24268
rect 10140 24080 10192 24132
rect 12624 24080 12676 24132
rect 14280 24148 14332 24200
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 19616 24284 19668 24336
rect 20260 24284 20312 24336
rect 14924 24080 14976 24132
rect 18880 24191 18932 24200
rect 18880 24157 18889 24191
rect 18889 24157 18923 24191
rect 18923 24157 18932 24191
rect 18880 24148 18932 24157
rect 20536 24148 20588 24200
rect 20628 24080 20680 24132
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 22376 24216 22428 24268
rect 26424 24395 26476 24404
rect 26424 24361 26433 24395
rect 26433 24361 26467 24395
rect 26467 24361 26476 24395
rect 26424 24352 26476 24361
rect 27252 24395 27304 24404
rect 27252 24361 27261 24395
rect 27261 24361 27295 24395
rect 27295 24361 27304 24395
rect 27252 24352 27304 24361
rect 29736 24395 29788 24404
rect 29736 24361 29745 24395
rect 29745 24361 29779 24395
rect 29779 24361 29788 24395
rect 29736 24352 29788 24361
rect 30380 24352 30432 24404
rect 25780 24327 25832 24336
rect 25780 24293 25789 24327
rect 25789 24293 25823 24327
rect 25823 24293 25832 24327
rect 25780 24284 25832 24293
rect 21456 24148 21508 24200
rect 28632 24284 28684 24336
rect 25412 24148 25464 24200
rect 27344 24216 27396 24268
rect 26240 24148 26292 24200
rect 25320 24080 25372 24132
rect 26608 24123 26660 24132
rect 5540 24012 5592 24064
rect 7472 24012 7524 24064
rect 9128 24055 9180 24064
rect 9128 24021 9137 24055
rect 9137 24021 9171 24055
rect 9171 24021 9180 24055
rect 9128 24012 9180 24021
rect 11152 24012 11204 24064
rect 11796 24012 11848 24064
rect 18420 24012 18472 24064
rect 19432 24055 19484 24064
rect 19432 24021 19441 24055
rect 19441 24021 19475 24055
rect 19475 24021 19484 24055
rect 19432 24012 19484 24021
rect 20260 24012 20312 24064
rect 23848 24012 23900 24064
rect 24676 24012 24728 24064
rect 26608 24089 26617 24123
rect 26617 24089 26651 24123
rect 26651 24089 26660 24123
rect 26608 24080 26660 24089
rect 27252 24080 27304 24132
rect 27344 24123 27396 24132
rect 27344 24089 27353 24123
rect 27353 24089 27387 24123
rect 27387 24089 27396 24123
rect 27344 24080 27396 24089
rect 30380 24191 30432 24200
rect 30380 24157 30389 24191
rect 30389 24157 30423 24191
rect 30423 24157 30432 24191
rect 30380 24148 30432 24157
rect 31116 24216 31168 24268
rect 33508 24284 33560 24336
rect 31576 24148 31628 24200
rect 33324 24148 33376 24200
rect 36728 24259 36780 24268
rect 36728 24225 36737 24259
rect 36737 24225 36771 24259
rect 36771 24225 36780 24259
rect 36728 24216 36780 24225
rect 37280 24216 37332 24268
rect 36360 24148 36412 24200
rect 37832 24216 37884 24268
rect 38660 24395 38712 24404
rect 38660 24361 38669 24395
rect 38669 24361 38703 24395
rect 38703 24361 38712 24395
rect 38660 24352 38712 24361
rect 39304 24395 39356 24404
rect 39304 24361 39313 24395
rect 39313 24361 39347 24395
rect 39347 24361 39356 24395
rect 39304 24352 39356 24361
rect 39856 24352 39908 24404
rect 42248 24352 42300 24404
rect 42616 24352 42668 24404
rect 43904 24352 43956 24404
rect 39764 24284 39816 24336
rect 42524 24284 42576 24336
rect 45376 24216 45428 24268
rect 47492 24216 47544 24268
rect 48228 24216 48280 24268
rect 37740 24148 37792 24200
rect 37924 24148 37976 24200
rect 26976 24012 27028 24064
rect 27804 24012 27856 24064
rect 28540 24012 28592 24064
rect 28724 24055 28776 24064
rect 28724 24021 28733 24055
rect 28733 24021 28767 24055
rect 28767 24021 28776 24055
rect 28724 24012 28776 24021
rect 30564 24055 30616 24064
rect 30564 24021 30573 24055
rect 30573 24021 30607 24055
rect 30607 24021 30616 24055
rect 30564 24012 30616 24021
rect 30932 24012 30984 24064
rect 32128 24012 32180 24064
rect 32312 24055 32364 24064
rect 32312 24021 32321 24055
rect 32321 24021 32355 24055
rect 32355 24021 32364 24055
rect 32312 24012 32364 24021
rect 34152 24080 34204 24132
rect 34612 24080 34664 24132
rect 35164 24123 35216 24132
rect 35164 24089 35173 24123
rect 35173 24089 35207 24123
rect 35207 24089 35216 24123
rect 35164 24080 35216 24089
rect 36820 24080 36872 24132
rect 38108 24080 38160 24132
rect 39488 24191 39540 24200
rect 39488 24157 39497 24191
rect 39497 24157 39531 24191
rect 39531 24157 39540 24191
rect 39488 24148 39540 24157
rect 40132 24148 40184 24200
rect 34060 24055 34112 24064
rect 34060 24021 34069 24055
rect 34069 24021 34103 24055
rect 34103 24021 34112 24055
rect 34060 24012 34112 24021
rect 34796 24012 34848 24064
rect 35256 24055 35308 24064
rect 35256 24021 35265 24055
rect 35265 24021 35299 24055
rect 35299 24021 35308 24055
rect 35256 24012 35308 24021
rect 35624 24055 35676 24064
rect 35624 24021 35633 24055
rect 35633 24021 35667 24055
rect 35667 24021 35676 24055
rect 35624 24012 35676 24021
rect 36084 24055 36136 24064
rect 36084 24021 36093 24055
rect 36093 24021 36127 24055
rect 36127 24021 36136 24055
rect 36084 24012 36136 24021
rect 37740 24055 37792 24064
rect 37740 24021 37749 24055
rect 37749 24021 37783 24055
rect 37783 24021 37792 24055
rect 37740 24012 37792 24021
rect 38660 24012 38712 24064
rect 39672 24080 39724 24132
rect 41144 24080 41196 24132
rect 42800 24148 42852 24200
rect 43812 24148 43864 24200
rect 43904 24191 43956 24200
rect 43904 24157 43913 24191
rect 43913 24157 43947 24191
rect 43947 24157 43956 24191
rect 43904 24148 43956 24157
rect 44456 24148 44508 24200
rect 45560 24148 45612 24200
rect 46204 24191 46256 24200
rect 46204 24157 46213 24191
rect 46213 24157 46247 24191
rect 46247 24157 46256 24191
rect 46204 24148 46256 24157
rect 46296 24148 46348 24200
rect 48044 24191 48096 24200
rect 48044 24157 48053 24191
rect 48053 24157 48087 24191
rect 48087 24157 48096 24191
rect 48044 24148 48096 24157
rect 48780 24191 48832 24200
rect 48780 24157 48789 24191
rect 48789 24157 48823 24191
rect 48823 24157 48832 24191
rect 48780 24148 48832 24157
rect 44272 24080 44324 24132
rect 44732 24080 44784 24132
rect 47400 24080 47452 24132
rect 39856 24012 39908 24064
rect 40040 24055 40092 24064
rect 40040 24021 40049 24055
rect 40049 24021 40083 24055
rect 40083 24021 40092 24055
rect 40040 24012 40092 24021
rect 40316 24012 40368 24064
rect 42616 24012 42668 24064
rect 42708 24012 42760 24064
rect 46020 24055 46072 24064
rect 46020 24021 46029 24055
rect 46029 24021 46063 24055
rect 46063 24021 46072 24055
rect 46020 24012 46072 24021
rect 46112 24012 46164 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 4620 23808 4672 23860
rect 10324 23808 10376 23860
rect 4068 23715 4120 23724
rect 4068 23681 4077 23715
rect 4077 23681 4111 23715
rect 4111 23681 4120 23715
rect 4068 23672 4120 23681
rect 4712 23715 4764 23724
rect 4712 23681 4721 23715
rect 4721 23681 4755 23715
rect 4755 23681 4764 23715
rect 4712 23672 4764 23681
rect 4160 23604 4212 23656
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 8484 23672 8536 23724
rect 11796 23740 11848 23792
rect 8392 23604 8444 23656
rect 9220 23604 9272 23656
rect 10600 23647 10652 23656
rect 10600 23613 10609 23647
rect 10609 23613 10643 23647
rect 10643 23613 10652 23647
rect 10600 23604 10652 23613
rect 12348 23715 12400 23724
rect 12348 23681 12357 23715
rect 12357 23681 12391 23715
rect 12391 23681 12400 23715
rect 12348 23672 12400 23681
rect 12716 23672 12768 23724
rect 14188 23740 14240 23792
rect 14372 23740 14424 23792
rect 19616 23808 19668 23860
rect 20260 23783 20312 23792
rect 20260 23749 20269 23783
rect 20269 23749 20303 23783
rect 20303 23749 20312 23783
rect 20260 23740 20312 23749
rect 21456 23851 21508 23860
rect 21456 23817 21465 23851
rect 21465 23817 21499 23851
rect 21499 23817 21508 23851
rect 21456 23808 21508 23817
rect 27896 23808 27948 23860
rect 28448 23851 28500 23860
rect 28448 23817 28457 23851
rect 28457 23817 28491 23851
rect 28491 23817 28500 23851
rect 28448 23808 28500 23817
rect 21640 23740 21692 23792
rect 25872 23740 25924 23792
rect 27712 23740 27764 23792
rect 28264 23740 28316 23792
rect 3424 23536 3476 23588
rect 5816 23536 5868 23588
rect 16396 23604 16448 23656
rect 18328 23604 18380 23656
rect 2780 23468 2832 23520
rect 5724 23468 5776 23520
rect 6000 23468 6052 23520
rect 18788 23511 18840 23520
rect 18788 23477 18797 23511
rect 18797 23477 18831 23511
rect 18831 23477 18840 23511
rect 18788 23468 18840 23477
rect 21272 23715 21324 23724
rect 21272 23681 21281 23715
rect 21281 23681 21315 23715
rect 21315 23681 21324 23715
rect 21272 23672 21324 23681
rect 23480 23672 23532 23724
rect 23664 23715 23716 23724
rect 23664 23681 23673 23715
rect 23673 23681 23707 23715
rect 23707 23681 23716 23715
rect 23664 23672 23716 23681
rect 21732 23604 21784 23656
rect 22560 23647 22612 23656
rect 22560 23613 22569 23647
rect 22569 23613 22603 23647
rect 22603 23613 22612 23647
rect 22560 23604 22612 23613
rect 23848 23647 23900 23656
rect 23848 23613 23857 23647
rect 23857 23613 23891 23647
rect 23891 23613 23900 23647
rect 23848 23604 23900 23613
rect 26608 23647 26660 23656
rect 26608 23613 26617 23647
rect 26617 23613 26651 23647
rect 26651 23613 26660 23647
rect 26608 23604 26660 23613
rect 23388 23536 23440 23588
rect 27804 23715 27856 23724
rect 27804 23681 27813 23715
rect 27813 23681 27847 23715
rect 27847 23681 27856 23715
rect 27804 23672 27856 23681
rect 40040 23808 40092 23860
rect 40132 23808 40184 23860
rect 42248 23851 42300 23860
rect 42248 23817 42257 23851
rect 42257 23817 42291 23851
rect 42291 23817 42300 23851
rect 42248 23808 42300 23817
rect 32404 23740 32456 23792
rect 28356 23604 28408 23656
rect 30380 23672 30432 23724
rect 32680 23715 32732 23724
rect 32680 23681 32689 23715
rect 32689 23681 32723 23715
rect 32723 23681 32732 23715
rect 32680 23672 32732 23681
rect 29368 23604 29420 23656
rect 20996 23468 21048 23520
rect 23480 23468 23532 23520
rect 24400 23511 24452 23520
rect 24400 23477 24409 23511
rect 24409 23477 24443 23511
rect 24443 23477 24452 23511
rect 24400 23468 24452 23477
rect 24860 23511 24912 23520
rect 24860 23477 24869 23511
rect 24869 23477 24903 23511
rect 24903 23477 24912 23511
rect 24860 23468 24912 23477
rect 29644 23536 29696 23588
rect 31760 23647 31812 23656
rect 31760 23613 31769 23647
rect 31769 23613 31803 23647
rect 31803 23613 31812 23647
rect 31760 23604 31812 23613
rect 33784 23740 33836 23792
rect 34980 23740 35032 23792
rect 32312 23536 32364 23588
rect 27804 23468 27856 23520
rect 29092 23468 29144 23520
rect 30288 23468 30340 23520
rect 34980 23604 35032 23656
rect 34520 23468 34572 23520
rect 35348 23647 35400 23656
rect 35348 23613 35357 23647
rect 35357 23613 35391 23647
rect 35391 23613 35400 23647
rect 35348 23604 35400 23613
rect 35624 23740 35676 23792
rect 39672 23740 39724 23792
rect 42708 23740 42760 23792
rect 35992 23672 36044 23724
rect 35440 23536 35492 23588
rect 35532 23468 35584 23520
rect 39212 23715 39264 23724
rect 39212 23681 39221 23715
rect 39221 23681 39255 23715
rect 39255 23681 39264 23715
rect 39212 23672 39264 23681
rect 39948 23672 40000 23724
rect 38568 23647 38620 23656
rect 38568 23613 38577 23647
rect 38577 23613 38611 23647
rect 38611 23613 38620 23647
rect 38568 23604 38620 23613
rect 39396 23604 39448 23656
rect 39488 23647 39540 23656
rect 39488 23613 39497 23647
rect 39497 23613 39531 23647
rect 39531 23613 39540 23647
rect 39488 23604 39540 23613
rect 40316 23672 40368 23724
rect 40592 23604 40644 23656
rect 40224 23536 40276 23588
rect 40776 23604 40828 23656
rect 42800 23672 42852 23724
rect 44824 23715 44876 23724
rect 44824 23681 44833 23715
rect 44833 23681 44867 23715
rect 44867 23681 44876 23715
rect 44824 23672 44876 23681
rect 45928 23715 45980 23724
rect 45928 23681 45937 23715
rect 45937 23681 45971 23715
rect 45971 23681 45980 23715
rect 45928 23672 45980 23681
rect 46204 23808 46256 23860
rect 47860 23808 47912 23860
rect 46940 23783 46992 23792
rect 46940 23749 46949 23783
rect 46949 23749 46983 23783
rect 46983 23749 46992 23783
rect 46940 23740 46992 23749
rect 47400 23715 47452 23724
rect 47400 23681 47409 23715
rect 47409 23681 47443 23715
rect 47443 23681 47452 23715
rect 47400 23672 47452 23681
rect 49240 23672 49292 23724
rect 47308 23604 47360 23656
rect 36912 23511 36964 23520
rect 36912 23477 36921 23511
rect 36921 23477 36955 23511
rect 36955 23477 36964 23511
rect 36912 23468 36964 23477
rect 37372 23468 37424 23520
rect 42708 23536 42760 23588
rect 45928 23536 45980 23588
rect 46940 23536 46992 23588
rect 47124 23536 47176 23588
rect 40684 23468 40736 23520
rect 43536 23468 43588 23520
rect 46204 23511 46256 23520
rect 46204 23477 46213 23511
rect 46213 23477 46247 23511
rect 46247 23477 46256 23511
rect 46204 23468 46256 23477
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 4712 23307 4764 23316
rect 4712 23273 4721 23307
rect 4721 23273 4755 23307
rect 4755 23273 4764 23307
rect 4712 23264 4764 23273
rect 5264 23196 5316 23248
rect 5632 23128 5684 23180
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 15844 23264 15896 23316
rect 14188 23239 14240 23248
rect 14188 23205 14197 23239
rect 14197 23205 14231 23239
rect 14231 23205 14240 23239
rect 14188 23196 14240 23205
rect 19616 23239 19668 23248
rect 19616 23205 19625 23239
rect 19625 23205 19659 23239
rect 19659 23205 19668 23239
rect 19616 23196 19668 23205
rect 19892 23264 19944 23316
rect 20260 23264 20312 23316
rect 22836 23264 22888 23316
rect 25136 23264 25188 23316
rect 25412 23264 25464 23316
rect 27896 23307 27948 23316
rect 27896 23273 27905 23307
rect 27905 23273 27939 23307
rect 27939 23273 27948 23307
rect 27896 23264 27948 23273
rect 28356 23264 28408 23316
rect 30380 23264 30432 23316
rect 31484 23264 31536 23316
rect 33324 23264 33376 23316
rect 35072 23264 35124 23316
rect 37372 23264 37424 23316
rect 37464 23264 37516 23316
rect 11244 23171 11296 23180
rect 11244 23137 11253 23171
rect 11253 23137 11287 23171
rect 11287 23137 11296 23171
rect 11244 23128 11296 23137
rect 13360 23128 13412 23180
rect 15752 23171 15804 23180
rect 15752 23137 15761 23171
rect 15761 23137 15795 23171
rect 15795 23137 15804 23171
rect 15752 23128 15804 23137
rect 4436 23060 4488 23112
rect 1768 23035 1820 23044
rect 1768 23001 1777 23035
rect 1777 23001 1811 23035
rect 1811 23001 1820 23035
rect 1768 22992 1820 23001
rect 4620 22924 4672 22976
rect 5356 23103 5408 23112
rect 5356 23069 5365 23103
rect 5365 23069 5399 23103
rect 5399 23069 5408 23103
rect 5356 23060 5408 23069
rect 5540 23060 5592 23112
rect 9128 23060 9180 23112
rect 11888 23103 11940 23112
rect 11888 23069 11897 23103
rect 11897 23069 11931 23103
rect 11931 23069 11940 23103
rect 11888 23060 11940 23069
rect 13820 23060 13872 23112
rect 19524 23128 19576 23180
rect 21732 23128 21784 23180
rect 19340 23060 19392 23112
rect 23388 23196 23440 23248
rect 28264 23196 28316 23248
rect 33784 23196 33836 23248
rect 34612 23196 34664 23248
rect 36360 23196 36412 23248
rect 37188 23196 37240 23248
rect 40040 23239 40092 23248
rect 40040 23205 40049 23239
rect 40049 23205 40083 23239
rect 40083 23205 40092 23239
rect 40040 23196 40092 23205
rect 24860 23128 24912 23180
rect 26056 23128 26108 23180
rect 29644 23128 29696 23180
rect 30196 23171 30248 23180
rect 30196 23137 30205 23171
rect 30205 23137 30239 23171
rect 30239 23137 30248 23171
rect 30196 23128 30248 23137
rect 30288 23171 30340 23180
rect 30288 23137 30297 23171
rect 30297 23137 30331 23171
rect 30331 23137 30340 23171
rect 30288 23128 30340 23137
rect 16580 22992 16632 23044
rect 17868 22992 17920 23044
rect 18604 23035 18656 23044
rect 18604 23001 18613 23035
rect 18613 23001 18647 23035
rect 18647 23001 18656 23035
rect 18604 22992 18656 23001
rect 19800 23035 19852 23044
rect 19800 23001 19809 23035
rect 19809 23001 19843 23035
rect 19843 23001 19852 23035
rect 19800 22992 19852 23001
rect 21732 22992 21784 23044
rect 21824 23035 21876 23044
rect 21824 23001 21833 23035
rect 21833 23001 21867 23035
rect 21867 23001 21876 23035
rect 21824 22992 21876 23001
rect 22560 23035 22612 23044
rect 22560 23001 22569 23035
rect 22569 23001 22603 23035
rect 22603 23001 22612 23035
rect 22560 22992 22612 23001
rect 24768 23035 24820 23044
rect 24768 23001 24777 23035
rect 24777 23001 24811 23035
rect 24811 23001 24820 23035
rect 24768 22992 24820 23001
rect 25688 23103 25740 23112
rect 25688 23069 25697 23103
rect 25697 23069 25731 23103
rect 25731 23069 25740 23103
rect 25688 23060 25740 23069
rect 30104 23060 30156 23112
rect 26240 22992 26292 23044
rect 27252 22992 27304 23044
rect 9220 22924 9272 22976
rect 14372 22967 14424 22976
rect 14372 22933 14381 22967
rect 14381 22933 14415 22967
rect 14415 22933 14424 22967
rect 14372 22924 14424 22933
rect 14648 22967 14700 22976
rect 14648 22933 14657 22967
rect 14657 22933 14691 22967
rect 14691 22933 14700 22967
rect 14648 22924 14700 22933
rect 17132 22967 17184 22976
rect 17132 22933 17141 22967
rect 17141 22933 17175 22967
rect 17175 22933 17184 22967
rect 17132 22924 17184 22933
rect 18880 22924 18932 22976
rect 20812 22924 20864 22976
rect 21548 22924 21600 22976
rect 23204 22924 23256 22976
rect 23296 22967 23348 22976
rect 23296 22933 23305 22967
rect 23305 22933 23339 22967
rect 23339 22933 23348 22967
rect 23296 22924 23348 22933
rect 23756 22967 23808 22976
rect 23756 22933 23765 22967
rect 23765 22933 23799 22967
rect 23799 22933 23808 22967
rect 23756 22924 23808 22933
rect 25320 22967 25372 22976
rect 25320 22933 25329 22967
rect 25329 22933 25363 22967
rect 25363 22933 25372 22967
rect 25320 22924 25372 22933
rect 25412 22924 25464 22976
rect 26056 22924 26108 22976
rect 26332 22924 26384 22976
rect 29920 22992 29972 23044
rect 31760 23128 31812 23180
rect 33508 23128 33560 23180
rect 34336 23128 34388 23180
rect 35348 23128 35400 23180
rect 35716 23128 35768 23180
rect 38384 23128 38436 23180
rect 38660 23128 38712 23180
rect 39488 23171 39540 23180
rect 39488 23137 39497 23171
rect 39497 23137 39531 23171
rect 39531 23137 39540 23171
rect 39488 23128 39540 23137
rect 42800 23264 42852 23316
rect 44824 23264 44876 23316
rect 46664 23307 46716 23316
rect 46664 23273 46673 23307
rect 46673 23273 46707 23307
rect 46707 23273 46716 23307
rect 46664 23264 46716 23273
rect 46940 23307 46992 23316
rect 46940 23273 46949 23307
rect 46949 23273 46983 23307
rect 46983 23273 46992 23307
rect 46940 23264 46992 23273
rect 43720 23196 43772 23248
rect 46112 23196 46164 23248
rect 31392 23103 31444 23112
rect 31392 23069 31401 23103
rect 31401 23069 31435 23103
rect 31435 23069 31444 23103
rect 31392 23060 31444 23069
rect 30104 22967 30156 22976
rect 30104 22933 30113 22967
rect 30113 22933 30147 22967
rect 30147 22933 30156 22967
rect 30104 22924 30156 22933
rect 32128 22992 32180 23044
rect 30380 22924 30432 22976
rect 31208 22924 31260 22976
rect 44088 23060 44140 23112
rect 45376 23103 45428 23112
rect 45376 23069 45385 23103
rect 45385 23069 45419 23103
rect 45419 23069 45428 23103
rect 45376 23060 45428 23069
rect 46664 23060 46716 23112
rect 47124 23103 47176 23112
rect 47124 23069 47133 23103
rect 47133 23069 47167 23103
rect 47167 23069 47176 23103
rect 47124 23060 47176 23069
rect 47308 23060 47360 23112
rect 48688 23060 48740 23112
rect 49424 23060 49476 23112
rect 33416 22992 33468 23044
rect 33784 22924 33836 22976
rect 34520 22992 34572 23044
rect 36912 22992 36964 23044
rect 35164 22924 35216 22976
rect 37096 22924 37148 22976
rect 40224 22992 40276 23044
rect 41512 23035 41564 23044
rect 41512 23001 41521 23035
rect 41521 23001 41555 23035
rect 41555 23001 41564 23035
rect 41512 22992 41564 23001
rect 42708 22992 42760 23044
rect 43536 22992 43588 23044
rect 43628 22992 43680 23044
rect 38660 22924 38712 22976
rect 39672 22924 39724 22976
rect 41236 22924 41288 22976
rect 46112 22967 46164 22976
rect 46112 22933 46121 22967
rect 46121 22933 46155 22967
rect 46155 22933 46164 22967
rect 46112 22924 46164 22933
rect 47032 22924 47084 22976
rect 47492 22924 47544 22976
rect 47676 22967 47728 22976
rect 47676 22933 47685 22967
rect 47685 22933 47719 22967
rect 47719 22933 47728 22967
rect 47676 22924 47728 22933
rect 48412 22967 48464 22976
rect 48412 22933 48421 22967
rect 48421 22933 48455 22967
rect 48455 22933 48464 22967
rect 48412 22924 48464 22933
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 1584 22720 1636 22772
rect 3424 22720 3476 22772
rect 3608 22720 3660 22772
rect 5356 22720 5408 22772
rect 7196 22763 7248 22772
rect 7196 22729 7205 22763
rect 7205 22729 7239 22763
rect 7239 22729 7248 22763
rect 7196 22720 7248 22729
rect 4804 22695 4856 22704
rect 4804 22661 4813 22695
rect 4813 22661 4847 22695
rect 4847 22661 4856 22695
rect 4804 22652 4856 22661
rect 7104 22652 7156 22704
rect 2780 22516 2832 22568
rect 6000 22627 6052 22636
rect 6000 22593 6009 22627
rect 6009 22593 6043 22627
rect 6043 22593 6052 22627
rect 6000 22584 6052 22593
rect 7196 22584 7248 22636
rect 15752 22720 15804 22772
rect 18604 22763 18656 22772
rect 18604 22729 18613 22763
rect 18613 22729 18647 22763
rect 18647 22729 18656 22763
rect 18604 22720 18656 22729
rect 19340 22720 19392 22772
rect 9956 22695 10008 22704
rect 9956 22661 9965 22695
rect 9965 22661 9999 22695
rect 9999 22661 10008 22695
rect 9956 22652 10008 22661
rect 7472 22627 7524 22636
rect 7472 22593 7481 22627
rect 7481 22593 7515 22627
rect 7515 22593 7524 22627
rect 7472 22584 7524 22593
rect 11152 22627 11204 22636
rect 11152 22593 11161 22627
rect 11161 22593 11195 22627
rect 11195 22593 11204 22627
rect 11152 22584 11204 22593
rect 12808 22695 12860 22704
rect 12808 22661 12817 22695
rect 12817 22661 12851 22695
rect 12851 22661 12860 22695
rect 12808 22652 12860 22661
rect 15108 22695 15160 22704
rect 15108 22661 15117 22695
rect 15117 22661 15151 22695
rect 15151 22661 15160 22695
rect 15108 22652 15160 22661
rect 15200 22652 15252 22704
rect 17868 22652 17920 22704
rect 13452 22584 13504 22636
rect 14648 22584 14700 22636
rect 7380 22516 7432 22568
rect 11796 22516 11848 22568
rect 5448 22448 5500 22500
rect 9128 22448 9180 22500
rect 11060 22448 11112 22500
rect 13912 22448 13964 22500
rect 3056 22380 3108 22432
rect 6000 22380 6052 22432
rect 12072 22380 12124 22432
rect 14372 22423 14424 22432
rect 14372 22389 14381 22423
rect 14381 22389 14415 22423
rect 14415 22389 14424 22423
rect 14372 22380 14424 22389
rect 18788 22584 18840 22636
rect 20812 22584 20864 22636
rect 21364 22720 21416 22772
rect 21824 22720 21876 22772
rect 23204 22720 23256 22772
rect 25504 22720 25556 22772
rect 24032 22652 24084 22704
rect 24860 22652 24912 22704
rect 25872 22652 25924 22704
rect 26332 22695 26384 22704
rect 26332 22661 26341 22695
rect 26341 22661 26375 22695
rect 26375 22661 26384 22695
rect 26332 22652 26384 22661
rect 26608 22720 26660 22772
rect 27252 22652 27304 22704
rect 27620 22652 27672 22704
rect 27896 22652 27948 22704
rect 28264 22652 28316 22704
rect 21916 22584 21968 22636
rect 24400 22627 24452 22636
rect 24400 22593 24409 22627
rect 24409 22593 24443 22627
rect 24443 22593 24452 22627
rect 24400 22584 24452 22593
rect 16764 22516 16816 22568
rect 17868 22516 17920 22568
rect 18880 22559 18932 22568
rect 18880 22525 18889 22559
rect 18889 22525 18923 22559
rect 18923 22525 18932 22559
rect 18880 22516 18932 22525
rect 19340 22448 19392 22500
rect 19708 22559 19760 22568
rect 19708 22525 19717 22559
rect 19717 22525 19751 22559
rect 19751 22525 19760 22559
rect 19708 22516 19760 22525
rect 23296 22516 23348 22568
rect 23572 22516 23624 22568
rect 26608 22627 26660 22636
rect 26608 22593 26617 22627
rect 26617 22593 26651 22627
rect 26651 22593 26660 22627
rect 26608 22584 26660 22593
rect 31392 22720 31444 22772
rect 30656 22695 30708 22704
rect 30656 22661 30665 22695
rect 30665 22661 30699 22695
rect 30699 22661 30708 22695
rect 30656 22652 30708 22661
rect 30748 22695 30800 22704
rect 30748 22661 30757 22695
rect 30757 22661 30791 22695
rect 30791 22661 30800 22695
rect 30748 22652 30800 22661
rect 30472 22584 30524 22636
rect 34244 22720 34296 22772
rect 34336 22720 34388 22772
rect 35532 22720 35584 22772
rect 37464 22763 37516 22772
rect 37464 22729 37473 22763
rect 37473 22729 37507 22763
rect 37507 22729 37516 22763
rect 37464 22720 37516 22729
rect 37648 22720 37700 22772
rect 38568 22720 38620 22772
rect 38752 22720 38804 22772
rect 33600 22652 33652 22704
rect 32772 22584 32824 22636
rect 33416 22627 33468 22636
rect 33416 22593 33425 22627
rect 33425 22593 33459 22627
rect 33459 22593 33468 22627
rect 33416 22584 33468 22593
rect 34612 22652 34664 22704
rect 35256 22584 35308 22636
rect 21824 22448 21876 22500
rect 20812 22380 20864 22432
rect 21640 22423 21692 22432
rect 21640 22389 21649 22423
rect 21649 22389 21683 22423
rect 21683 22389 21692 22423
rect 21640 22380 21692 22389
rect 24216 22448 24268 22500
rect 24952 22448 25004 22500
rect 24492 22423 24544 22432
rect 24492 22389 24501 22423
rect 24501 22389 24535 22423
rect 24535 22389 24544 22423
rect 24492 22380 24544 22389
rect 25780 22516 25832 22568
rect 27252 22516 27304 22568
rect 27620 22516 27672 22568
rect 27712 22516 27764 22568
rect 28080 22559 28132 22568
rect 28080 22525 28089 22559
rect 28089 22525 28123 22559
rect 28123 22525 28132 22559
rect 28080 22516 28132 22525
rect 28356 22516 28408 22568
rect 29184 22516 29236 22568
rect 27344 22491 27396 22500
rect 27344 22457 27353 22491
rect 27353 22457 27387 22491
rect 27387 22457 27396 22491
rect 27344 22448 27396 22457
rect 29920 22516 29972 22568
rect 31024 22448 31076 22500
rect 26332 22380 26384 22432
rect 26608 22380 26660 22432
rect 30380 22380 30432 22432
rect 31116 22380 31168 22432
rect 31484 22423 31536 22432
rect 31484 22389 31493 22423
rect 31493 22389 31527 22423
rect 31527 22389 31536 22423
rect 31484 22380 31536 22389
rect 33508 22516 33560 22568
rect 34060 22516 34112 22568
rect 38660 22652 38712 22704
rect 38844 22652 38896 22704
rect 39488 22627 39540 22636
rect 39488 22593 39497 22627
rect 39497 22593 39531 22627
rect 39531 22593 39540 22627
rect 39488 22584 39540 22593
rect 40592 22652 40644 22704
rect 48688 22720 48740 22772
rect 46112 22652 46164 22704
rect 46756 22652 46808 22704
rect 40684 22584 40736 22636
rect 41420 22627 41472 22636
rect 41420 22593 41429 22627
rect 41429 22593 41463 22627
rect 41463 22593 41472 22627
rect 41420 22584 41472 22593
rect 42064 22627 42116 22636
rect 42064 22593 42073 22627
rect 42073 22593 42107 22627
rect 42107 22593 42116 22627
rect 42064 22584 42116 22593
rect 43996 22584 44048 22636
rect 44732 22627 44784 22636
rect 44732 22593 44741 22627
rect 44741 22593 44775 22627
rect 44775 22593 44784 22627
rect 44732 22584 44784 22593
rect 45284 22584 45336 22636
rect 47768 22627 47820 22636
rect 47768 22593 47777 22627
rect 47777 22593 47811 22627
rect 47811 22593 47820 22627
rect 47768 22584 47820 22593
rect 49332 22627 49384 22636
rect 49332 22593 49341 22627
rect 49341 22593 49375 22627
rect 49375 22593 49384 22627
rect 49332 22584 49384 22593
rect 34152 22380 34204 22432
rect 36360 22448 36412 22500
rect 37096 22448 37148 22500
rect 42616 22559 42668 22568
rect 42616 22525 42625 22559
rect 42625 22525 42659 22559
rect 42659 22525 42668 22559
rect 42616 22516 42668 22525
rect 43444 22516 43496 22568
rect 41880 22491 41932 22500
rect 41880 22457 41889 22491
rect 41889 22457 41923 22491
rect 41923 22457 41932 22491
rect 41880 22448 41932 22457
rect 45192 22491 45244 22500
rect 45192 22457 45201 22491
rect 45201 22457 45235 22491
rect 45235 22457 45244 22491
rect 45192 22448 45244 22457
rect 35164 22380 35216 22432
rect 37556 22380 37608 22432
rect 38752 22380 38804 22432
rect 39120 22380 39172 22432
rect 40040 22423 40092 22432
rect 40040 22389 40049 22423
rect 40049 22389 40083 22423
rect 40083 22389 40092 22423
rect 40040 22380 40092 22389
rect 41236 22423 41288 22432
rect 41236 22389 41245 22423
rect 41245 22389 41279 22423
rect 41279 22389 41288 22423
rect 41236 22380 41288 22389
rect 43904 22423 43956 22432
rect 43904 22389 43913 22423
rect 43913 22389 43947 22423
rect 43947 22389 43956 22423
rect 43904 22380 43956 22389
rect 44548 22423 44600 22432
rect 44548 22389 44557 22423
rect 44557 22389 44591 22423
rect 44591 22389 44600 22423
rect 44548 22380 44600 22389
rect 45376 22380 45428 22432
rect 46940 22380 46992 22432
rect 47584 22448 47636 22500
rect 49240 22448 49292 22500
rect 48320 22380 48372 22432
rect 48688 22380 48740 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 2228 22176 2280 22228
rect 4252 22176 4304 22228
rect 11888 22176 11940 22228
rect 2872 22108 2924 22160
rect 7104 22108 7156 22160
rect 7840 22108 7892 22160
rect 10232 22108 10284 22160
rect 1032 21904 1084 21956
rect 3240 21904 3292 21956
rect 6736 21972 6788 22024
rect 7748 21972 7800 22024
rect 9680 22040 9732 22092
rect 9772 22083 9824 22092
rect 9772 22049 9781 22083
rect 9781 22049 9815 22083
rect 9815 22049 9824 22083
rect 9772 22040 9824 22049
rect 11888 22083 11940 22092
rect 11888 22049 11897 22083
rect 11897 22049 11931 22083
rect 11931 22049 11940 22083
rect 11888 22040 11940 22049
rect 5632 21904 5684 21956
rect 8392 21879 8444 21888
rect 8392 21845 8401 21879
rect 8401 21845 8435 21879
rect 8435 21845 8444 21879
rect 8392 21836 8444 21845
rect 8944 21836 8996 21888
rect 9128 22015 9180 22024
rect 9128 21981 9137 22015
rect 9137 21981 9171 22015
rect 9171 21981 9180 22015
rect 9128 21972 9180 21981
rect 12532 22015 12584 22024
rect 12532 21981 12541 22015
rect 12541 21981 12575 22015
rect 12575 21981 12584 22015
rect 12532 21972 12584 21981
rect 14188 22151 14240 22160
rect 14188 22117 14197 22151
rect 14197 22117 14231 22151
rect 14231 22117 14240 22151
rect 14188 22108 14240 22117
rect 14372 22108 14424 22160
rect 15108 22108 15160 22160
rect 19616 22176 19668 22228
rect 22192 22176 22244 22228
rect 24676 22176 24728 22228
rect 14280 22040 14332 22092
rect 15200 22083 15252 22092
rect 15200 22049 15209 22083
rect 15209 22049 15243 22083
rect 15243 22049 15252 22083
rect 15200 22040 15252 22049
rect 15660 22108 15712 22160
rect 17040 22108 17092 22160
rect 15384 22040 15436 22092
rect 20168 22108 20220 22160
rect 17132 21972 17184 22024
rect 18972 22040 19024 22092
rect 22744 22040 22796 22092
rect 23572 22040 23624 22092
rect 23664 22040 23716 22092
rect 24860 22108 24912 22160
rect 24952 22108 25004 22160
rect 14648 21947 14700 21956
rect 14648 21913 14657 21947
rect 14657 21913 14691 21947
rect 14691 21913 14700 21947
rect 14648 21904 14700 21913
rect 16120 21904 16172 21956
rect 16672 21947 16724 21956
rect 16672 21913 16681 21947
rect 16681 21913 16715 21947
rect 16715 21913 16724 21947
rect 16672 21904 16724 21913
rect 19248 21972 19300 22024
rect 19432 22015 19484 22024
rect 19432 21981 19441 22015
rect 19441 21981 19475 22015
rect 19475 21981 19484 22015
rect 19432 21972 19484 21981
rect 22560 21972 22612 22024
rect 24032 22015 24084 22024
rect 24032 21981 24041 22015
rect 24041 21981 24075 22015
rect 24075 21981 24084 22015
rect 24032 21972 24084 21981
rect 25412 22040 25464 22092
rect 25320 21972 25372 22024
rect 28264 22176 28316 22228
rect 26700 22108 26752 22160
rect 28724 22176 28776 22228
rect 30196 22176 30248 22228
rect 31852 22176 31904 22228
rect 32772 22176 32824 22228
rect 35440 22176 35492 22228
rect 35532 22176 35584 22228
rect 26332 22040 26384 22092
rect 27620 22083 27672 22092
rect 27620 22049 27629 22083
rect 27629 22049 27663 22083
rect 27663 22049 27672 22083
rect 27620 22040 27672 22049
rect 27712 22083 27764 22092
rect 27712 22049 27721 22083
rect 27721 22049 27755 22083
rect 27755 22049 27764 22083
rect 27712 22040 27764 22049
rect 28080 22040 28132 22092
rect 28908 22083 28960 22092
rect 28908 22049 28917 22083
rect 28917 22049 28951 22083
rect 28951 22049 28960 22083
rect 28908 22040 28960 22049
rect 29552 22040 29604 22092
rect 30564 22040 30616 22092
rect 31484 22040 31536 22092
rect 32312 22040 32364 22092
rect 33876 22040 33928 22092
rect 34796 22040 34848 22092
rect 34980 22083 35032 22092
rect 34980 22049 34989 22083
rect 34989 22049 35023 22083
rect 35023 22049 35032 22083
rect 34980 22040 35032 22049
rect 38660 22176 38712 22228
rect 38844 22176 38896 22228
rect 39488 22219 39540 22228
rect 39488 22185 39497 22219
rect 39497 22185 39531 22219
rect 39531 22185 39540 22219
rect 39488 22176 39540 22185
rect 40224 22219 40276 22228
rect 40224 22185 40233 22219
rect 40233 22185 40267 22219
rect 40267 22185 40276 22219
rect 40224 22176 40276 22185
rect 41052 22176 41104 22228
rect 42708 22176 42760 22228
rect 43536 22176 43588 22228
rect 44088 22176 44140 22228
rect 47032 22219 47084 22228
rect 47032 22185 47041 22219
rect 47041 22185 47075 22219
rect 47075 22185 47084 22219
rect 47032 22176 47084 22185
rect 49424 22176 49476 22228
rect 38844 22083 38896 22092
rect 38844 22049 38853 22083
rect 38853 22049 38887 22083
rect 38887 22049 38896 22083
rect 38844 22040 38896 22049
rect 26608 21972 26660 22024
rect 27804 21972 27856 22024
rect 29828 21972 29880 22024
rect 30656 21972 30708 22024
rect 30840 22015 30892 22024
rect 30840 21981 30849 22015
rect 30849 21981 30883 22015
rect 30883 21981 30892 22015
rect 30840 21972 30892 21981
rect 32128 21972 32180 22024
rect 39396 22040 39448 22092
rect 21548 21904 21600 21956
rect 22928 21904 22980 21956
rect 24584 21904 24636 21956
rect 24952 21947 25004 21956
rect 24952 21913 24961 21947
rect 24961 21913 24995 21947
rect 24995 21913 25004 21947
rect 24952 21904 25004 21913
rect 26056 21904 26108 21956
rect 26332 21947 26384 21956
rect 26332 21913 26341 21947
rect 26341 21913 26375 21947
rect 26375 21913 26384 21947
rect 26332 21904 26384 21913
rect 30472 21904 30524 21956
rect 31024 21904 31076 21956
rect 31392 21904 31444 21956
rect 21272 21836 21324 21888
rect 21456 21879 21508 21888
rect 21456 21845 21465 21879
rect 21465 21845 21499 21879
rect 21499 21845 21508 21879
rect 21456 21836 21508 21845
rect 21916 21879 21968 21888
rect 21916 21845 21925 21879
rect 21925 21845 21959 21879
rect 21959 21845 21968 21879
rect 21916 21836 21968 21845
rect 22652 21879 22704 21888
rect 22652 21845 22661 21879
rect 22661 21845 22695 21879
rect 22695 21845 22704 21879
rect 22652 21836 22704 21845
rect 23112 21879 23164 21888
rect 23112 21845 23121 21879
rect 23121 21845 23155 21879
rect 23155 21845 23164 21879
rect 23112 21836 23164 21845
rect 23756 21836 23808 21888
rect 25964 21879 26016 21888
rect 25964 21845 25973 21879
rect 25973 21845 26007 21879
rect 26007 21845 26016 21879
rect 25964 21836 26016 21845
rect 26148 21836 26200 21888
rect 29552 21836 29604 21888
rect 29736 21879 29788 21888
rect 29736 21845 29745 21879
rect 29745 21845 29779 21879
rect 29779 21845 29788 21879
rect 29736 21836 29788 21845
rect 30380 21879 30432 21888
rect 30380 21845 30389 21879
rect 30389 21845 30423 21879
rect 30423 21845 30432 21879
rect 30380 21836 30432 21845
rect 32128 21836 32180 21888
rect 32404 21836 32456 21888
rect 32680 21836 32732 21888
rect 33416 21879 33468 21888
rect 33416 21845 33425 21879
rect 33425 21845 33459 21879
rect 33459 21845 33468 21879
rect 33416 21836 33468 21845
rect 34336 21879 34388 21888
rect 34336 21845 34345 21879
rect 34345 21845 34379 21879
rect 34379 21845 34388 21879
rect 34336 21836 34388 21845
rect 34612 21836 34664 21888
rect 35808 21904 35860 21956
rect 39580 21972 39632 22024
rect 42432 21972 42484 22024
rect 43720 22108 43772 22160
rect 44272 22108 44324 22160
rect 42892 22040 42944 22092
rect 43812 22040 43864 22092
rect 44732 22040 44784 22092
rect 42800 22015 42852 22024
rect 42800 21981 42809 22015
rect 42809 21981 42843 22015
rect 42843 21981 42852 22015
rect 42800 21972 42852 21981
rect 43260 22015 43312 22024
rect 43260 21981 43269 22015
rect 43269 21981 43303 22015
rect 43303 21981 43312 22015
rect 43260 21972 43312 21981
rect 47584 21972 47636 22024
rect 48504 22015 48556 22024
rect 48504 21981 48513 22015
rect 48513 21981 48547 22015
rect 48547 21981 48556 22015
rect 48504 21972 48556 21981
rect 37188 21904 37240 21956
rect 37556 21904 37608 21956
rect 38384 21904 38436 21956
rect 35992 21836 36044 21888
rect 36268 21836 36320 21888
rect 36544 21836 36596 21888
rect 36820 21879 36872 21888
rect 36820 21845 36829 21879
rect 36829 21845 36863 21879
rect 36863 21845 36872 21879
rect 36820 21836 36872 21845
rect 37280 21836 37332 21888
rect 37464 21836 37516 21888
rect 40040 21904 40092 21956
rect 39672 21879 39724 21888
rect 39672 21845 39681 21879
rect 39681 21845 39715 21879
rect 39715 21845 39724 21879
rect 39672 21836 39724 21845
rect 39948 21836 40000 21888
rect 40868 21836 40920 21888
rect 40960 21836 41012 21888
rect 42708 21904 42760 21956
rect 49056 21947 49108 21956
rect 49056 21913 49065 21947
rect 49065 21913 49099 21947
rect 49099 21913 49108 21947
rect 49056 21904 49108 21913
rect 49240 21947 49292 21956
rect 49240 21913 49249 21947
rect 49249 21913 49283 21947
rect 49283 21913 49292 21947
rect 49240 21904 49292 21913
rect 41328 21836 41380 21888
rect 41788 21879 41840 21888
rect 41788 21845 41797 21879
rect 41797 21845 41831 21879
rect 41831 21845 41840 21879
rect 41788 21836 41840 21845
rect 41880 21836 41932 21888
rect 47860 21836 47912 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 9588 21632 9640 21684
rect 3332 21564 3384 21616
rect 6736 21564 6788 21616
rect 1768 21471 1820 21480
rect 1768 21437 1777 21471
rect 1777 21437 1811 21471
rect 1811 21437 1820 21471
rect 1768 21428 1820 21437
rect 4620 21539 4672 21548
rect 4620 21505 4629 21539
rect 4629 21505 4663 21539
rect 4663 21505 4672 21539
rect 4620 21496 4672 21505
rect 6552 21496 6604 21548
rect 6644 21539 6696 21548
rect 6644 21505 6653 21539
rect 6653 21505 6687 21539
rect 6687 21505 6696 21539
rect 6644 21496 6696 21505
rect 5632 21428 5684 21480
rect 5816 21428 5868 21480
rect 9036 21496 9088 21548
rect 9956 21496 10008 21548
rect 12440 21632 12492 21684
rect 10968 21564 11020 21616
rect 12624 21564 12676 21616
rect 13820 21632 13872 21684
rect 20996 21632 21048 21684
rect 21916 21632 21968 21684
rect 22560 21632 22612 21684
rect 22928 21632 22980 21684
rect 14280 21564 14332 21616
rect 3792 21292 3844 21344
rect 12072 21496 12124 21548
rect 12164 21496 12216 21548
rect 14004 21496 14056 21548
rect 14372 21496 14424 21548
rect 11428 21428 11480 21480
rect 11704 21471 11756 21480
rect 11704 21437 11713 21471
rect 11713 21437 11747 21471
rect 11747 21437 11756 21471
rect 11704 21428 11756 21437
rect 12624 21428 12676 21480
rect 12808 21471 12860 21480
rect 12808 21437 12817 21471
rect 12817 21437 12851 21471
rect 12851 21437 12860 21471
rect 12808 21428 12860 21437
rect 13912 21428 13964 21480
rect 13728 21360 13780 21412
rect 8944 21292 8996 21344
rect 10876 21292 10928 21344
rect 11796 21292 11848 21344
rect 12256 21335 12308 21344
rect 12256 21301 12265 21335
rect 12265 21301 12299 21335
rect 12299 21301 12308 21335
rect 12256 21292 12308 21301
rect 15200 21428 15252 21480
rect 16120 21564 16172 21616
rect 16948 21564 17000 21616
rect 18328 21496 18380 21548
rect 16672 21428 16724 21480
rect 17500 21428 17552 21480
rect 18788 21564 18840 21616
rect 19156 21564 19208 21616
rect 20628 21564 20680 21616
rect 16764 21403 16816 21412
rect 16764 21369 16773 21403
rect 16773 21369 16807 21403
rect 16807 21369 16816 21403
rect 16764 21360 16816 21369
rect 18880 21471 18932 21480
rect 18880 21437 18889 21471
rect 18889 21437 18923 21471
rect 18923 21437 18932 21471
rect 18880 21428 18932 21437
rect 19248 21428 19300 21480
rect 27068 21632 27120 21684
rect 16948 21335 17000 21344
rect 16948 21301 16957 21335
rect 16957 21301 16991 21335
rect 16991 21301 17000 21335
rect 16948 21292 17000 21301
rect 17868 21292 17920 21344
rect 21088 21360 21140 21412
rect 21548 21428 21600 21480
rect 22284 21496 22336 21548
rect 23848 21496 23900 21548
rect 22192 21428 22244 21480
rect 25044 21564 25096 21616
rect 27436 21632 27488 21684
rect 31760 21632 31812 21684
rect 33416 21632 33468 21684
rect 35900 21632 35952 21684
rect 37464 21632 37516 21684
rect 37556 21632 37608 21684
rect 39120 21632 39172 21684
rect 39212 21632 39264 21684
rect 39948 21632 40000 21684
rect 29368 21564 29420 21616
rect 33692 21564 33744 21616
rect 34888 21564 34940 21616
rect 37280 21564 37332 21616
rect 38292 21607 38344 21616
rect 38292 21573 38301 21607
rect 38301 21573 38335 21607
rect 38335 21573 38344 21607
rect 38292 21564 38344 21573
rect 39672 21564 39724 21616
rect 41052 21632 41104 21684
rect 42064 21632 42116 21684
rect 43536 21632 43588 21684
rect 43996 21632 44048 21684
rect 46204 21632 46256 21684
rect 47860 21632 47912 21684
rect 40868 21564 40920 21616
rect 42524 21607 42576 21616
rect 42524 21573 42533 21607
rect 42533 21573 42567 21607
rect 42567 21573 42576 21607
rect 42524 21564 42576 21573
rect 42708 21607 42760 21616
rect 42708 21573 42717 21607
rect 42717 21573 42751 21607
rect 42751 21573 42760 21607
rect 42708 21564 42760 21573
rect 42800 21564 42852 21616
rect 25872 21496 25924 21548
rect 26056 21539 26108 21548
rect 26056 21505 26065 21539
rect 26065 21505 26099 21539
rect 26099 21505 26108 21539
rect 26056 21496 26108 21505
rect 24492 21428 24544 21480
rect 25412 21471 25464 21480
rect 25412 21437 25421 21471
rect 25421 21437 25455 21471
rect 25455 21437 25464 21471
rect 25412 21428 25464 21437
rect 19340 21292 19392 21344
rect 19616 21292 19668 21344
rect 21640 21292 21692 21344
rect 22376 21292 22428 21344
rect 22560 21292 22612 21344
rect 24676 21292 24728 21344
rect 25136 21360 25188 21412
rect 27896 21496 27948 21548
rect 30748 21496 30800 21548
rect 31208 21539 31260 21548
rect 31208 21505 31217 21539
rect 31217 21505 31251 21539
rect 31251 21505 31260 21539
rect 31208 21496 31260 21505
rect 33508 21539 33560 21548
rect 33508 21505 33517 21539
rect 33517 21505 33551 21539
rect 33551 21505 33560 21539
rect 33508 21496 33560 21505
rect 28816 21471 28868 21480
rect 28816 21437 28825 21471
rect 28825 21437 28859 21471
rect 28859 21437 28868 21471
rect 28816 21428 28868 21437
rect 28908 21471 28960 21480
rect 28908 21437 28917 21471
rect 28917 21437 28951 21471
rect 28951 21437 28960 21471
rect 28908 21428 28960 21437
rect 29736 21428 29788 21480
rect 31576 21428 31628 21480
rect 33416 21471 33468 21480
rect 33416 21437 33425 21471
rect 33425 21437 33459 21471
rect 33459 21437 33468 21471
rect 33416 21428 33468 21437
rect 34244 21428 34296 21480
rect 30472 21360 30524 21412
rect 30564 21360 30616 21412
rect 31484 21360 31536 21412
rect 34704 21360 34756 21412
rect 25872 21335 25924 21344
rect 25872 21301 25881 21335
rect 25881 21301 25915 21335
rect 25915 21301 25924 21335
rect 25872 21292 25924 21301
rect 26240 21292 26292 21344
rect 29552 21335 29604 21344
rect 29552 21301 29561 21335
rect 29561 21301 29595 21335
rect 29595 21301 29604 21335
rect 29552 21292 29604 21301
rect 29644 21292 29696 21344
rect 29920 21292 29972 21344
rect 30748 21335 30800 21344
rect 30748 21301 30757 21335
rect 30757 21301 30791 21335
rect 30791 21301 30800 21335
rect 30748 21292 30800 21301
rect 31944 21292 31996 21344
rect 37740 21496 37792 21548
rect 40684 21496 40736 21548
rect 43260 21539 43312 21548
rect 43260 21505 43269 21539
rect 43269 21505 43303 21539
rect 43303 21505 43312 21539
rect 43260 21496 43312 21505
rect 46848 21496 46900 21548
rect 48596 21539 48648 21548
rect 48596 21505 48605 21539
rect 48605 21505 48639 21539
rect 48639 21505 48648 21539
rect 48596 21496 48648 21505
rect 49332 21539 49384 21548
rect 49332 21505 49341 21539
rect 49341 21505 49375 21539
rect 49375 21505 49384 21539
rect 49332 21496 49384 21505
rect 34888 21428 34940 21480
rect 36176 21471 36228 21480
rect 36176 21437 36185 21471
rect 36185 21437 36219 21471
rect 36219 21437 36228 21471
rect 36176 21428 36228 21437
rect 36912 21428 36964 21480
rect 37188 21428 37240 21480
rect 37556 21428 37608 21480
rect 40316 21428 40368 21480
rect 35164 21335 35216 21344
rect 35164 21301 35173 21335
rect 35173 21301 35207 21335
rect 35207 21301 35216 21335
rect 35164 21292 35216 21301
rect 35716 21335 35768 21344
rect 35716 21301 35725 21335
rect 35725 21301 35759 21335
rect 35759 21301 35768 21335
rect 35716 21292 35768 21301
rect 35808 21292 35860 21344
rect 37556 21335 37608 21344
rect 37556 21301 37565 21335
rect 37565 21301 37599 21335
rect 37599 21301 37608 21335
rect 37556 21292 37608 21301
rect 37740 21292 37792 21344
rect 38108 21292 38160 21344
rect 38844 21292 38896 21344
rect 39028 21292 39080 21344
rect 40868 21335 40920 21344
rect 40868 21301 40877 21335
rect 40877 21301 40911 21335
rect 40911 21301 40920 21335
rect 41512 21471 41564 21480
rect 41512 21437 41521 21471
rect 41521 21437 41555 21471
rect 41555 21437 41564 21471
rect 41512 21428 41564 21437
rect 41604 21428 41656 21480
rect 41788 21360 41840 21412
rect 40868 21292 40920 21301
rect 41328 21292 41380 21344
rect 43536 21292 43588 21344
rect 49148 21335 49200 21344
rect 49148 21301 49157 21335
rect 49157 21301 49191 21335
rect 49191 21301 49200 21335
rect 49148 21292 49200 21301
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 2872 20952 2924 21004
rect 9128 21088 9180 21140
rect 9220 21131 9272 21140
rect 9220 21097 9229 21131
rect 9229 21097 9263 21131
rect 9263 21097 9272 21131
rect 9220 21088 9272 21097
rect 12256 21088 12308 21140
rect 12808 21088 12860 21140
rect 14280 21131 14332 21140
rect 14280 21097 14289 21131
rect 14289 21097 14323 21131
rect 14323 21097 14332 21131
rect 14280 21088 14332 21097
rect 14372 21088 14424 21140
rect 15292 21088 15344 21140
rect 16304 21088 16356 21140
rect 19708 21088 19760 21140
rect 22560 21088 22612 21140
rect 24124 21088 24176 21140
rect 4160 20995 4212 21004
rect 4160 20961 4169 20995
rect 4169 20961 4203 20995
rect 4203 20961 4212 20995
rect 4160 20952 4212 20961
rect 6000 20995 6052 21004
rect 6000 20961 6009 20995
rect 6009 20961 6043 20995
rect 6043 20961 6052 20995
rect 6000 20952 6052 20961
rect 7748 20952 7800 21004
rect 7288 20748 7340 20800
rect 7564 20791 7616 20800
rect 7564 20757 7573 20791
rect 7573 20757 7607 20791
rect 7607 20757 7616 20791
rect 7564 20748 7616 20757
rect 8392 20927 8444 20936
rect 8392 20893 8401 20927
rect 8401 20893 8435 20927
rect 8435 20893 8444 20927
rect 8392 20884 8444 20893
rect 19248 21020 19300 21072
rect 19616 21020 19668 21072
rect 10232 20952 10284 21004
rect 12716 20995 12768 21004
rect 12716 20961 12725 20995
rect 12725 20961 12759 20995
rect 12759 20961 12768 20995
rect 12716 20952 12768 20961
rect 23296 21020 23348 21072
rect 23848 21020 23900 21072
rect 25504 21088 25556 21140
rect 27068 21088 27120 21140
rect 29460 21088 29512 21140
rect 11336 20923 11388 20936
rect 11336 20889 11345 20923
rect 11345 20889 11379 20923
rect 11379 20889 11388 20923
rect 11336 20884 11388 20889
rect 10600 20748 10652 20800
rect 10692 20791 10744 20800
rect 10692 20757 10701 20791
rect 10701 20757 10735 20791
rect 10735 20757 10744 20791
rect 10692 20748 10744 20757
rect 11060 20748 11112 20800
rect 12624 20884 12676 20936
rect 16764 20884 16816 20936
rect 19340 20884 19392 20936
rect 12072 20816 12124 20868
rect 12624 20748 12676 20800
rect 15200 20816 15252 20868
rect 16120 20816 16172 20868
rect 13544 20791 13596 20800
rect 13544 20757 13553 20791
rect 13553 20757 13587 20791
rect 13587 20757 13596 20791
rect 13544 20748 13596 20757
rect 17868 20816 17920 20868
rect 19432 20816 19484 20868
rect 18512 20748 18564 20800
rect 19340 20791 19392 20800
rect 19340 20757 19349 20791
rect 19349 20757 19383 20791
rect 19383 20757 19392 20791
rect 19340 20748 19392 20757
rect 19800 20884 19852 20936
rect 22652 20952 22704 21004
rect 25228 21063 25280 21072
rect 25228 21029 25237 21063
rect 25237 21029 25271 21063
rect 25271 21029 25280 21063
rect 25228 21020 25280 21029
rect 25780 21020 25832 21072
rect 26148 21020 26200 21072
rect 29552 21020 29604 21072
rect 29920 21088 29972 21140
rect 30012 21088 30064 21140
rect 26240 20952 26292 21004
rect 26332 20995 26384 21004
rect 26332 20961 26341 20995
rect 26341 20961 26375 20995
rect 26375 20961 26384 20995
rect 26332 20952 26384 20961
rect 27896 20995 27948 21004
rect 27896 20961 27905 20995
rect 27905 20961 27939 20995
rect 27939 20961 27948 20995
rect 27896 20952 27948 20961
rect 35716 21088 35768 21140
rect 36728 21088 36780 21140
rect 37648 21131 37700 21140
rect 37648 21097 37657 21131
rect 37657 21097 37691 21131
rect 37691 21097 37700 21131
rect 37648 21088 37700 21097
rect 31944 21063 31996 21072
rect 31944 21029 31953 21063
rect 31953 21029 31987 21063
rect 31987 21029 31996 21063
rect 31944 21020 31996 21029
rect 34888 21063 34940 21072
rect 34888 21029 34897 21063
rect 34897 21029 34931 21063
rect 34931 21029 34940 21063
rect 34888 21020 34940 21029
rect 38384 21088 38436 21140
rect 40132 21088 40184 21140
rect 40500 21088 40552 21140
rect 41328 21088 41380 21140
rect 41420 21088 41472 21140
rect 42616 21088 42668 21140
rect 46848 21088 46900 21140
rect 48596 21131 48648 21140
rect 48596 21097 48605 21131
rect 48605 21097 48639 21131
rect 48639 21097 48648 21131
rect 48596 21088 48648 21097
rect 40224 21020 40276 21072
rect 41052 21020 41104 21072
rect 49332 21020 49384 21072
rect 22928 20927 22980 20936
rect 22928 20893 22937 20927
rect 22937 20893 22971 20927
rect 22971 20893 22980 20927
rect 22928 20884 22980 20893
rect 24124 20884 24176 20936
rect 26976 20884 27028 20936
rect 29736 20884 29788 20936
rect 29920 20927 29972 20936
rect 29920 20893 29929 20927
rect 29929 20893 29963 20927
rect 29963 20893 29972 20927
rect 29920 20884 29972 20893
rect 32312 20952 32364 21004
rect 33140 20952 33192 21004
rect 33508 20952 33560 21004
rect 34336 20952 34388 21004
rect 32404 20884 32456 20936
rect 32496 20927 32548 20936
rect 32496 20893 32505 20927
rect 32505 20893 32539 20927
rect 32539 20893 32548 20927
rect 32496 20884 32548 20893
rect 19616 20791 19668 20800
rect 19616 20757 19625 20791
rect 19625 20757 19659 20791
rect 19659 20757 19668 20791
rect 19616 20748 19668 20757
rect 22376 20816 22428 20868
rect 22560 20816 22612 20868
rect 22744 20816 22796 20868
rect 23572 20859 23624 20868
rect 23572 20825 23581 20859
rect 23581 20825 23615 20859
rect 23615 20825 23624 20859
rect 23572 20816 23624 20825
rect 25964 20816 26016 20868
rect 26792 20816 26844 20868
rect 27436 20859 27488 20868
rect 27436 20825 27445 20859
rect 27445 20825 27479 20859
rect 27479 20825 27488 20859
rect 27436 20816 27488 20825
rect 28356 20816 28408 20868
rect 24124 20748 24176 20800
rect 26148 20791 26200 20800
rect 26148 20757 26157 20791
rect 26157 20757 26191 20791
rect 26191 20757 26200 20791
rect 26148 20748 26200 20757
rect 26884 20748 26936 20800
rect 27160 20748 27212 20800
rect 27620 20748 27672 20800
rect 28724 20791 28776 20800
rect 28724 20757 28733 20791
rect 28733 20757 28767 20791
rect 28767 20757 28776 20791
rect 28724 20748 28776 20757
rect 30104 20748 30156 20800
rect 32128 20816 32180 20868
rect 31208 20791 31260 20800
rect 31208 20757 31217 20791
rect 31217 20757 31251 20791
rect 31251 20757 31260 20791
rect 31208 20748 31260 20757
rect 31484 20748 31536 20800
rect 32956 20748 33008 20800
rect 35072 20816 35124 20868
rect 36360 20859 36412 20868
rect 36360 20825 36369 20859
rect 36369 20825 36403 20859
rect 36403 20825 36412 20859
rect 36360 20816 36412 20825
rect 34336 20748 34388 20800
rect 37004 20791 37056 20800
rect 37004 20757 37013 20791
rect 37013 20757 37047 20791
rect 37047 20757 37056 20791
rect 37004 20748 37056 20757
rect 37556 20816 37608 20868
rect 38660 20952 38712 21004
rect 39120 20952 39172 21004
rect 39580 20952 39632 21004
rect 39764 20952 39816 21004
rect 40684 20952 40736 21004
rect 42432 20952 42484 21004
rect 43352 20952 43404 21004
rect 38384 20816 38436 20868
rect 39028 20816 39080 20868
rect 41604 20927 41656 20936
rect 41604 20893 41613 20927
rect 41613 20893 41647 20927
rect 41647 20893 41656 20927
rect 41604 20884 41656 20893
rect 49332 20927 49384 20936
rect 49332 20893 49341 20927
rect 49341 20893 49375 20927
rect 49375 20893 49384 20927
rect 49332 20884 49384 20893
rect 38292 20748 38344 20800
rect 40684 20748 40736 20800
rect 49424 20816 49476 20868
rect 41328 20748 41380 20800
rect 46204 20748 46256 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 6644 20544 6696 20596
rect 9680 20587 9732 20596
rect 9680 20553 9689 20587
rect 9689 20553 9723 20587
rect 9723 20553 9732 20587
rect 9680 20544 9732 20553
rect 10324 20587 10376 20596
rect 10324 20553 10333 20587
rect 10333 20553 10367 20587
rect 10367 20553 10376 20587
rect 10324 20544 10376 20553
rect 1308 20476 1360 20528
rect 3976 20408 4028 20460
rect 4804 20451 4856 20460
rect 4804 20417 4813 20451
rect 4813 20417 4847 20451
rect 4847 20417 4856 20451
rect 4804 20408 4856 20417
rect 8300 20476 8352 20528
rect 5448 20408 5500 20460
rect 9680 20408 9732 20460
rect 10968 20476 11020 20528
rect 12348 20476 12400 20528
rect 12716 20544 12768 20596
rect 14096 20587 14148 20596
rect 14096 20553 14105 20587
rect 14105 20553 14139 20587
rect 14139 20553 14148 20587
rect 14096 20544 14148 20553
rect 14924 20587 14976 20596
rect 14924 20553 14933 20587
rect 14933 20553 14967 20587
rect 14967 20553 14976 20587
rect 14924 20544 14976 20553
rect 15476 20544 15528 20596
rect 15844 20544 15896 20596
rect 16028 20587 16080 20596
rect 16028 20553 16037 20587
rect 16037 20553 16071 20587
rect 16071 20553 16080 20587
rect 16028 20544 16080 20553
rect 13912 20476 13964 20528
rect 16396 20544 16448 20596
rect 17132 20544 17184 20596
rect 17960 20544 18012 20596
rect 18880 20544 18932 20596
rect 19432 20544 19484 20596
rect 19708 20587 19760 20596
rect 19708 20553 19717 20587
rect 19717 20553 19751 20587
rect 19751 20553 19760 20587
rect 19708 20544 19760 20553
rect 20168 20544 20220 20596
rect 21088 20544 21140 20596
rect 21732 20544 21784 20596
rect 22744 20544 22796 20596
rect 22928 20544 22980 20596
rect 5908 20340 5960 20392
rect 10876 20408 10928 20460
rect 11796 20408 11848 20460
rect 12348 20340 12400 20392
rect 12900 20408 12952 20460
rect 15016 20408 15068 20460
rect 14280 20383 14332 20392
rect 14280 20349 14289 20383
rect 14289 20349 14323 20383
rect 14323 20349 14332 20383
rect 14280 20340 14332 20349
rect 2780 20272 2832 20324
rect 3332 20272 3384 20324
rect 4160 20204 4212 20256
rect 14924 20272 14976 20324
rect 19064 20476 19116 20528
rect 19340 20476 19392 20528
rect 23756 20476 23808 20528
rect 16764 20408 16816 20460
rect 22192 20408 22244 20460
rect 23388 20451 23440 20460
rect 23388 20417 23397 20451
rect 23397 20417 23431 20451
rect 23431 20417 23440 20451
rect 23388 20408 23440 20417
rect 25688 20544 25740 20596
rect 25780 20544 25832 20596
rect 26332 20544 26384 20596
rect 25228 20408 25280 20460
rect 16856 20340 16908 20392
rect 20444 20340 20496 20392
rect 21180 20383 21232 20392
rect 21180 20349 21189 20383
rect 21189 20349 21223 20383
rect 21223 20349 21232 20383
rect 21180 20340 21232 20349
rect 16488 20272 16540 20324
rect 19064 20315 19116 20324
rect 19064 20281 19073 20315
rect 19073 20281 19107 20315
rect 19107 20281 19116 20315
rect 19064 20272 19116 20281
rect 22468 20383 22520 20392
rect 22468 20349 22477 20383
rect 22477 20349 22511 20383
rect 22511 20349 22520 20383
rect 22468 20340 22520 20349
rect 22560 20383 22612 20392
rect 22560 20349 22569 20383
rect 22569 20349 22603 20383
rect 22603 20349 22612 20383
rect 22560 20340 22612 20349
rect 24216 20340 24268 20392
rect 26976 20476 27028 20528
rect 25504 20408 25556 20460
rect 30840 20544 30892 20596
rect 31484 20544 31536 20596
rect 32496 20544 32548 20596
rect 27804 20476 27856 20528
rect 29828 20519 29880 20528
rect 29828 20485 29837 20519
rect 29837 20485 29871 20519
rect 29871 20485 29880 20519
rect 29828 20476 29880 20485
rect 31116 20476 31168 20528
rect 31852 20476 31904 20528
rect 32128 20476 32180 20528
rect 28908 20408 28960 20460
rect 25596 20383 25648 20392
rect 25596 20349 25605 20383
rect 25605 20349 25639 20383
rect 25639 20349 25648 20383
rect 25596 20340 25648 20349
rect 25780 20340 25832 20392
rect 25872 20340 25924 20392
rect 29276 20340 29328 20392
rect 29460 20340 29512 20392
rect 30196 20408 30248 20460
rect 30288 20408 30340 20460
rect 31024 20340 31076 20392
rect 31944 20408 31996 20460
rect 31300 20383 31352 20392
rect 31300 20349 31309 20383
rect 31309 20349 31343 20383
rect 31343 20349 31352 20383
rect 31300 20340 31352 20349
rect 32312 20383 32364 20392
rect 32312 20349 32321 20383
rect 32321 20349 32355 20383
rect 32355 20349 32364 20383
rect 32312 20340 32364 20349
rect 32588 20340 32640 20392
rect 36176 20544 36228 20596
rect 36636 20544 36688 20596
rect 13360 20204 13412 20256
rect 15568 20204 15620 20256
rect 17040 20204 17092 20256
rect 17132 20204 17184 20256
rect 19616 20204 19668 20256
rect 21456 20204 21508 20256
rect 22008 20247 22060 20256
rect 22008 20213 22017 20247
rect 22017 20213 22051 20247
rect 22051 20213 22060 20247
rect 22008 20204 22060 20213
rect 22652 20272 22704 20324
rect 26148 20272 26200 20324
rect 28632 20272 28684 20324
rect 30932 20272 30984 20324
rect 31392 20272 31444 20324
rect 25412 20204 25464 20256
rect 26240 20247 26292 20256
rect 26240 20213 26249 20247
rect 26249 20213 26283 20247
rect 26283 20213 26292 20247
rect 26240 20204 26292 20213
rect 26332 20204 26384 20256
rect 27252 20204 27304 20256
rect 30288 20204 30340 20256
rect 30840 20204 30892 20256
rect 31116 20204 31168 20256
rect 32772 20272 32824 20324
rect 34520 20340 34572 20392
rect 36360 20476 36412 20528
rect 37096 20476 37148 20528
rect 38476 20476 38528 20528
rect 34796 20383 34848 20392
rect 34796 20349 34805 20383
rect 34805 20349 34839 20383
rect 34839 20349 34848 20383
rect 34796 20340 34848 20349
rect 35072 20408 35124 20460
rect 37188 20408 37240 20460
rect 39580 20408 39632 20460
rect 40408 20544 40460 20596
rect 49148 20544 49200 20596
rect 40592 20476 40644 20528
rect 35348 20340 35400 20392
rect 34888 20272 34940 20324
rect 34980 20272 35032 20324
rect 36636 20340 36688 20392
rect 37464 20340 37516 20392
rect 37648 20340 37700 20392
rect 40132 20383 40184 20392
rect 40132 20349 40141 20383
rect 40141 20349 40175 20383
rect 40175 20349 40184 20383
rect 40132 20340 40184 20349
rect 36084 20315 36136 20324
rect 36084 20281 36093 20315
rect 36093 20281 36127 20315
rect 36127 20281 36136 20315
rect 36084 20272 36136 20281
rect 36544 20272 36596 20324
rect 35716 20247 35768 20256
rect 35716 20213 35725 20247
rect 35725 20213 35759 20247
rect 35759 20213 35768 20247
rect 35716 20204 35768 20213
rect 36820 20204 36872 20256
rect 37740 20247 37792 20256
rect 37740 20213 37749 20247
rect 37749 20213 37783 20247
rect 37783 20213 37792 20247
rect 37740 20204 37792 20213
rect 48780 20408 48832 20460
rect 49424 20408 49476 20460
rect 40684 20247 40736 20256
rect 40684 20213 40693 20247
rect 40693 20213 40727 20247
rect 40727 20213 40736 20247
rect 40684 20204 40736 20213
rect 48412 20247 48464 20256
rect 48412 20213 48421 20247
rect 48421 20213 48455 20247
rect 48455 20213 48464 20247
rect 48412 20204 48464 20213
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 4804 20000 4856 20052
rect 9956 19975 10008 19984
rect 9956 19941 9965 19975
rect 9965 19941 9999 19975
rect 9999 19941 10008 19975
rect 9956 19932 10008 19941
rect 10600 19975 10652 19984
rect 10600 19941 10609 19975
rect 10609 19941 10643 19975
rect 10643 19941 10652 19975
rect 10600 19932 10652 19941
rect 4252 19907 4304 19916
rect 4252 19873 4261 19907
rect 4261 19873 4295 19907
rect 4295 19873 4304 19907
rect 4252 19864 4304 19873
rect 5724 19864 5776 19916
rect 11980 20000 12032 20052
rect 12808 20000 12860 20052
rect 14464 20043 14516 20052
rect 14464 20009 14473 20043
rect 14473 20009 14507 20043
rect 14507 20009 14516 20043
rect 14464 20000 14516 20009
rect 3332 19796 3384 19848
rect 5264 19839 5316 19848
rect 5264 19805 5273 19839
rect 5273 19805 5307 19839
rect 5307 19805 5316 19839
rect 5264 19796 5316 19805
rect 1492 19728 1544 19780
rect 9588 19796 9640 19848
rect 11980 19907 12032 19916
rect 11980 19873 11989 19907
rect 11989 19873 12023 19907
rect 12023 19873 12032 19907
rect 11980 19864 12032 19873
rect 14924 19975 14976 19984
rect 14924 19941 14933 19975
rect 14933 19941 14967 19975
rect 14967 19941 14976 19975
rect 14924 19932 14976 19941
rect 13636 19864 13688 19916
rect 16304 19907 16356 19916
rect 16304 19873 16313 19907
rect 16313 19873 16347 19907
rect 16347 19873 16356 19907
rect 16304 19864 16356 19873
rect 10968 19796 11020 19848
rect 11428 19771 11480 19780
rect 11428 19737 11437 19771
rect 11437 19737 11471 19771
rect 11471 19737 11480 19771
rect 11428 19728 11480 19737
rect 13360 19796 13412 19848
rect 14188 19796 14240 19848
rect 14280 19839 14332 19848
rect 14280 19805 14289 19839
rect 14289 19805 14323 19839
rect 14323 19805 14332 19839
rect 14280 19796 14332 19805
rect 15568 19796 15620 19848
rect 18880 19932 18932 19984
rect 19524 19932 19576 19984
rect 19984 20000 20036 20052
rect 22008 20000 22060 20052
rect 22468 20000 22520 20052
rect 26792 20043 26844 20052
rect 26792 20009 26801 20043
rect 26801 20009 26835 20043
rect 26835 20009 26844 20043
rect 26792 20000 26844 20009
rect 27068 20000 27120 20052
rect 34980 20000 35032 20052
rect 35440 20000 35492 20052
rect 37004 20000 37056 20052
rect 38384 20000 38436 20052
rect 38844 20000 38896 20052
rect 13820 19728 13872 19780
rect 19892 19864 19944 19916
rect 19524 19796 19576 19848
rect 17868 19728 17920 19780
rect 20536 19796 20588 19848
rect 22836 19864 22888 19916
rect 23388 19907 23440 19916
rect 23388 19873 23397 19907
rect 23397 19873 23431 19907
rect 23431 19873 23440 19907
rect 23388 19864 23440 19873
rect 23940 19932 23992 19984
rect 27620 19932 27672 19984
rect 27988 19932 28040 19984
rect 29828 19932 29880 19984
rect 24584 19907 24636 19916
rect 24584 19873 24593 19907
rect 24593 19873 24627 19907
rect 24627 19873 24636 19907
rect 24584 19864 24636 19873
rect 25044 19864 25096 19916
rect 22744 19796 22796 19848
rect 25228 19796 25280 19848
rect 26976 19864 27028 19916
rect 28356 19864 28408 19916
rect 29000 19864 29052 19916
rect 33324 19932 33376 19984
rect 27252 19796 27304 19848
rect 30196 19839 30248 19848
rect 30196 19805 30205 19839
rect 30205 19805 30239 19839
rect 30239 19805 30248 19839
rect 30196 19796 30248 19805
rect 30564 19796 30616 19848
rect 31300 19796 31352 19848
rect 13636 19660 13688 19712
rect 15936 19660 15988 19712
rect 17132 19660 17184 19712
rect 17224 19703 17276 19712
rect 17224 19669 17233 19703
rect 17233 19669 17267 19703
rect 17267 19669 17276 19703
rect 17224 19660 17276 19669
rect 18328 19660 18380 19712
rect 18420 19660 18472 19712
rect 20352 19728 20404 19780
rect 21548 19728 21600 19780
rect 22100 19728 22152 19780
rect 26700 19728 26752 19780
rect 30012 19728 30064 19780
rect 30104 19771 30156 19780
rect 30104 19737 30113 19771
rect 30113 19737 30147 19771
rect 30147 19737 30156 19771
rect 30104 19728 30156 19737
rect 19340 19703 19392 19712
rect 19340 19669 19349 19703
rect 19349 19669 19383 19703
rect 19383 19669 19392 19703
rect 19340 19660 19392 19669
rect 20260 19703 20312 19712
rect 20260 19669 20269 19703
rect 20269 19669 20303 19703
rect 20303 19669 20312 19703
rect 20260 19660 20312 19669
rect 20444 19660 20496 19712
rect 22652 19703 22704 19712
rect 22652 19669 22661 19703
rect 22661 19669 22695 19703
rect 22695 19669 22704 19703
rect 22652 19660 22704 19669
rect 23388 19660 23440 19712
rect 23480 19660 23532 19712
rect 26332 19660 26384 19712
rect 27068 19660 27120 19712
rect 27252 19703 27304 19712
rect 27252 19669 27261 19703
rect 27261 19669 27295 19703
rect 27295 19669 27304 19703
rect 27252 19660 27304 19669
rect 27620 19660 27672 19712
rect 28632 19660 28684 19712
rect 28908 19660 28960 19712
rect 29736 19703 29788 19712
rect 29736 19669 29745 19703
rect 29745 19669 29779 19703
rect 29779 19669 29788 19703
rect 29736 19660 29788 19669
rect 30932 19660 30984 19712
rect 31116 19660 31168 19712
rect 31576 19660 31628 19712
rect 32220 19728 32272 19780
rect 32128 19703 32180 19712
rect 32128 19669 32137 19703
rect 32137 19669 32171 19703
rect 32171 19669 32180 19703
rect 32128 19660 32180 19669
rect 34060 19864 34112 19916
rect 35072 19907 35124 19916
rect 35072 19873 35081 19907
rect 35081 19873 35115 19907
rect 35115 19873 35124 19907
rect 35072 19864 35124 19873
rect 35716 19864 35768 19916
rect 35808 19864 35860 19916
rect 36452 19864 36504 19916
rect 37648 19864 37700 19916
rect 38476 19932 38528 19984
rect 39212 19864 39264 19916
rect 39396 19864 39448 19916
rect 41052 20043 41104 20052
rect 41052 20009 41061 20043
rect 41061 20009 41095 20043
rect 41095 20009 41104 20043
rect 41052 20000 41104 20009
rect 48780 20043 48832 20052
rect 48780 20009 48789 20043
rect 48789 20009 48823 20043
rect 48823 20009 48832 20043
rect 48780 20000 48832 20009
rect 40960 19932 41012 19984
rect 33784 19839 33836 19848
rect 33784 19805 33793 19839
rect 33793 19805 33827 19839
rect 33827 19805 33836 19839
rect 33784 19796 33836 19805
rect 34152 19796 34204 19848
rect 35532 19796 35584 19848
rect 37372 19796 37424 19848
rect 40868 19796 40920 19848
rect 34888 19728 34940 19780
rect 34980 19728 35032 19780
rect 36268 19728 36320 19780
rect 40040 19728 40092 19780
rect 41052 19728 41104 19780
rect 49332 19728 49384 19780
rect 33416 19660 33468 19712
rect 34152 19703 34204 19712
rect 34152 19669 34161 19703
rect 34161 19669 34195 19703
rect 34195 19669 34204 19703
rect 34152 19660 34204 19669
rect 35992 19660 36044 19712
rect 36544 19703 36596 19712
rect 36544 19669 36553 19703
rect 36553 19669 36587 19703
rect 36587 19669 36596 19703
rect 36544 19660 36596 19669
rect 37556 19703 37608 19712
rect 37556 19669 37565 19703
rect 37565 19669 37599 19703
rect 37599 19669 37608 19703
rect 37556 19660 37608 19669
rect 38384 19660 38436 19712
rect 40776 19703 40828 19712
rect 40776 19669 40785 19703
rect 40785 19669 40819 19703
rect 40819 19669 40828 19703
rect 40776 19660 40828 19669
rect 49148 19703 49200 19712
rect 49148 19669 49157 19703
rect 49157 19669 49191 19703
rect 49191 19669 49200 19703
rect 49148 19660 49200 19669
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 7840 19456 7892 19508
rect 13452 19456 13504 19508
rect 3424 19388 3476 19440
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 9220 19388 9272 19440
rect 12808 19388 12860 19440
rect 14188 19388 14240 19440
rect 3884 19252 3936 19304
rect 5908 19320 5960 19372
rect 9128 19320 9180 19372
rect 6828 19252 6880 19304
rect 9864 19295 9916 19304
rect 9864 19261 9873 19295
rect 9873 19261 9907 19295
rect 9907 19261 9916 19295
rect 9864 19252 9916 19261
rect 11152 19363 11204 19372
rect 11152 19329 11161 19363
rect 11161 19329 11195 19363
rect 11195 19329 11204 19363
rect 11152 19320 11204 19329
rect 12164 19363 12216 19372
rect 12164 19329 12173 19363
rect 12173 19329 12207 19363
rect 12207 19329 12216 19363
rect 12164 19320 12216 19329
rect 15016 19456 15068 19508
rect 19432 19456 19484 19508
rect 20812 19456 20864 19508
rect 21272 19456 21324 19508
rect 16212 19431 16264 19440
rect 16212 19397 16221 19431
rect 16221 19397 16255 19431
rect 16255 19397 16264 19431
rect 16212 19388 16264 19397
rect 19064 19388 19116 19440
rect 20260 19388 20312 19440
rect 23480 19456 23532 19508
rect 22652 19388 22704 19440
rect 23388 19388 23440 19440
rect 24492 19388 24544 19440
rect 24860 19388 24912 19440
rect 15384 19320 15436 19372
rect 15476 19363 15528 19372
rect 15476 19329 15485 19363
rect 15485 19329 15519 19363
rect 15519 19329 15528 19363
rect 15476 19320 15528 19329
rect 17040 19320 17092 19372
rect 18420 19320 18472 19372
rect 7564 19184 7616 19236
rect 12072 19184 12124 19236
rect 12716 19252 12768 19304
rect 15200 19252 15252 19304
rect 15752 19252 15804 19304
rect 16028 19295 16080 19304
rect 16028 19261 16037 19295
rect 16037 19261 16071 19295
rect 16071 19261 16080 19295
rect 16028 19252 16080 19261
rect 16120 19252 16172 19304
rect 15476 19184 15528 19236
rect 19432 19252 19484 19304
rect 19800 19295 19852 19304
rect 19800 19261 19809 19295
rect 19809 19261 19843 19295
rect 19843 19261 19852 19295
rect 19800 19252 19852 19261
rect 5908 19159 5960 19168
rect 5908 19125 5917 19159
rect 5917 19125 5951 19159
rect 5951 19125 5960 19159
rect 5908 19116 5960 19125
rect 8300 19116 8352 19168
rect 11888 19116 11940 19168
rect 12440 19116 12492 19168
rect 12716 19159 12768 19168
rect 12716 19125 12725 19159
rect 12725 19125 12759 19159
rect 12759 19125 12768 19159
rect 12716 19116 12768 19125
rect 15108 19116 15160 19168
rect 16488 19116 16540 19168
rect 19064 19116 19116 19168
rect 19616 19116 19668 19168
rect 22192 19363 22244 19372
rect 22192 19329 22201 19363
rect 22201 19329 22235 19363
rect 22235 19329 22244 19363
rect 22192 19320 22244 19329
rect 25688 19320 25740 19372
rect 22284 19252 22336 19304
rect 22836 19252 22888 19304
rect 24860 19252 24912 19304
rect 24952 19295 25004 19304
rect 24952 19261 24961 19295
rect 24961 19261 24995 19295
rect 24995 19261 25004 19295
rect 24952 19252 25004 19261
rect 25596 19252 25648 19304
rect 26148 19499 26200 19508
rect 26148 19465 26157 19499
rect 26157 19465 26191 19499
rect 26191 19465 26200 19499
rect 26148 19456 26200 19465
rect 26240 19499 26292 19508
rect 26240 19465 26249 19499
rect 26249 19465 26283 19499
rect 26283 19465 26292 19499
rect 26240 19456 26292 19465
rect 27344 19456 27396 19508
rect 27436 19456 27488 19508
rect 28356 19456 28408 19508
rect 28724 19456 28776 19508
rect 30196 19456 30248 19508
rect 31852 19456 31904 19508
rect 32496 19456 32548 19508
rect 34980 19456 35032 19508
rect 36544 19456 36596 19508
rect 37004 19456 37056 19508
rect 27436 19252 27488 19304
rect 28448 19320 28500 19372
rect 21180 19116 21232 19168
rect 23848 19116 23900 19168
rect 25780 19159 25832 19168
rect 25780 19125 25789 19159
rect 25789 19125 25823 19159
rect 25823 19125 25832 19159
rect 25780 19116 25832 19125
rect 27252 19159 27304 19168
rect 27252 19125 27261 19159
rect 27261 19125 27295 19159
rect 27295 19125 27304 19159
rect 27252 19116 27304 19125
rect 28080 19252 28132 19304
rect 28632 19252 28684 19304
rect 28540 19184 28592 19236
rect 29276 19252 29328 19304
rect 30380 19320 30432 19372
rect 31484 19431 31536 19440
rect 31484 19397 31493 19431
rect 31493 19397 31527 19431
rect 31527 19397 31536 19431
rect 31484 19388 31536 19397
rect 31760 19388 31812 19440
rect 32864 19388 32916 19440
rect 34704 19388 34756 19440
rect 34796 19388 34848 19440
rect 35348 19388 35400 19440
rect 35900 19388 35952 19440
rect 34244 19320 34296 19372
rect 31668 19252 31720 19304
rect 32404 19295 32456 19304
rect 32404 19261 32413 19295
rect 32413 19261 32447 19295
rect 32447 19261 32456 19295
rect 32404 19252 32456 19261
rect 34888 19320 34940 19372
rect 34980 19363 35032 19372
rect 34980 19329 34989 19363
rect 34989 19329 35023 19363
rect 35023 19329 35032 19363
rect 34980 19320 35032 19329
rect 35532 19320 35584 19372
rect 36728 19320 36780 19372
rect 37372 19320 37424 19372
rect 38476 19456 38528 19508
rect 40040 19456 40092 19508
rect 40408 19456 40460 19508
rect 39396 19431 39448 19440
rect 39396 19397 39405 19431
rect 39405 19397 39439 19431
rect 39439 19397 39448 19431
rect 39396 19388 39448 19397
rect 48412 19388 48464 19440
rect 39672 19363 39724 19372
rect 39672 19329 39681 19363
rect 39681 19329 39715 19363
rect 39715 19329 39724 19363
rect 39672 19320 39724 19329
rect 49240 19363 49292 19372
rect 49240 19329 49249 19363
rect 49249 19329 49283 19363
rect 49283 19329 49292 19363
rect 49240 19320 49292 19329
rect 29920 19184 29972 19236
rect 34428 19184 34480 19236
rect 28908 19116 28960 19168
rect 30012 19116 30064 19168
rect 30380 19159 30432 19168
rect 30380 19125 30389 19159
rect 30389 19125 30423 19159
rect 30423 19125 30432 19159
rect 30380 19116 30432 19125
rect 35900 19252 35952 19304
rect 36084 19252 36136 19304
rect 40316 19252 40368 19304
rect 37740 19184 37792 19236
rect 36636 19159 36688 19168
rect 36636 19125 36645 19159
rect 36645 19125 36679 19159
rect 36679 19125 36688 19159
rect 36636 19116 36688 19125
rect 36820 19116 36872 19168
rect 37832 19116 37884 19168
rect 40868 19184 40920 19236
rect 41052 19116 41104 19168
rect 42064 19116 42116 19168
rect 49424 19116 49476 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 6828 18912 6880 18964
rect 10876 18912 10928 18964
rect 11888 18955 11940 18964
rect 11888 18921 11897 18955
rect 11897 18921 11931 18955
rect 11931 18921 11940 18955
rect 11888 18912 11940 18921
rect 12348 18912 12400 18964
rect 3516 18776 3568 18828
rect 11060 18844 11112 18896
rect 1400 18640 1452 18692
rect 5356 18751 5408 18760
rect 5356 18717 5365 18751
rect 5365 18717 5399 18751
rect 5399 18717 5408 18751
rect 5356 18708 5408 18717
rect 12532 18776 12584 18828
rect 12440 18708 12492 18760
rect 4344 18640 4396 18692
rect 10140 18640 10192 18692
rect 10232 18640 10284 18692
rect 10416 18572 10468 18624
rect 10692 18683 10744 18692
rect 10692 18649 10701 18683
rect 10701 18649 10735 18683
rect 10735 18649 10744 18683
rect 10692 18640 10744 18649
rect 12164 18640 12216 18692
rect 15108 18912 15160 18964
rect 15200 18912 15252 18964
rect 16120 18912 16172 18964
rect 13360 18844 13412 18896
rect 13820 18844 13872 18896
rect 15660 18844 15712 18896
rect 17868 18912 17920 18964
rect 19524 18912 19576 18964
rect 20720 18912 20772 18964
rect 23112 18912 23164 18964
rect 27620 18912 27672 18964
rect 27712 18912 27764 18964
rect 30196 18912 30248 18964
rect 30472 18912 30524 18964
rect 12716 18776 12768 18828
rect 13176 18776 13228 18828
rect 16948 18776 17000 18828
rect 17500 18819 17552 18828
rect 17500 18785 17509 18819
rect 17509 18785 17543 18819
rect 17543 18785 17552 18819
rect 17500 18776 17552 18785
rect 19708 18776 19760 18828
rect 20628 18844 20680 18896
rect 20444 18819 20496 18828
rect 20444 18785 20453 18819
rect 20453 18785 20487 18819
rect 20487 18785 20496 18819
rect 20444 18776 20496 18785
rect 21364 18776 21416 18828
rect 23020 18776 23072 18828
rect 25596 18776 25648 18828
rect 25688 18776 25740 18828
rect 28908 18844 28960 18896
rect 29000 18887 29052 18896
rect 29000 18853 29009 18887
rect 29009 18853 29043 18887
rect 29043 18853 29052 18887
rect 29000 18844 29052 18853
rect 29184 18844 29236 18896
rect 30748 18844 30800 18896
rect 30932 18887 30984 18896
rect 30932 18853 30941 18887
rect 30941 18853 30975 18887
rect 30975 18853 30984 18887
rect 30932 18844 30984 18853
rect 27068 18776 27120 18828
rect 12808 18708 12860 18760
rect 18512 18751 18564 18760
rect 18512 18717 18521 18751
rect 18521 18717 18555 18751
rect 18555 18717 18564 18751
rect 18512 18708 18564 18717
rect 21088 18708 21140 18760
rect 21824 18708 21876 18760
rect 24124 18708 24176 18760
rect 27436 18776 27488 18828
rect 27988 18776 28040 18828
rect 28448 18819 28500 18828
rect 28448 18785 28457 18819
rect 28457 18785 28491 18819
rect 28491 18785 28500 18819
rect 28448 18776 28500 18785
rect 28080 18708 28132 18760
rect 29276 18776 29328 18828
rect 29552 18776 29604 18828
rect 33324 18912 33376 18964
rect 33968 18912 34020 18964
rect 34336 18912 34388 18964
rect 34428 18912 34480 18964
rect 31024 18708 31076 18760
rect 31116 18708 31168 18760
rect 11520 18615 11572 18624
rect 11520 18581 11529 18615
rect 11529 18581 11563 18615
rect 11563 18581 11572 18615
rect 11520 18572 11572 18581
rect 14096 18572 14148 18624
rect 14556 18683 14608 18692
rect 14556 18649 14565 18683
rect 14565 18649 14599 18683
rect 14599 18649 14608 18683
rect 14556 18640 14608 18649
rect 14832 18640 14884 18692
rect 16304 18683 16356 18692
rect 16304 18649 16313 18683
rect 16313 18649 16347 18683
rect 16347 18649 16356 18683
rect 16304 18640 16356 18649
rect 17408 18683 17460 18692
rect 17408 18649 17417 18683
rect 17417 18649 17451 18683
rect 17451 18649 17460 18683
rect 17408 18640 17460 18649
rect 19340 18683 19392 18692
rect 19340 18649 19349 18683
rect 19349 18649 19383 18683
rect 19383 18649 19392 18683
rect 19340 18640 19392 18649
rect 19432 18640 19484 18692
rect 15568 18572 15620 18624
rect 16672 18615 16724 18624
rect 16672 18581 16681 18615
rect 16681 18581 16715 18615
rect 16715 18581 16724 18615
rect 16672 18572 16724 18581
rect 19616 18615 19668 18624
rect 19616 18581 19625 18615
rect 19625 18581 19659 18615
rect 19659 18581 19668 18615
rect 19616 18572 19668 18581
rect 21456 18572 21508 18624
rect 22008 18572 22060 18624
rect 22100 18572 22152 18624
rect 22376 18572 22428 18624
rect 23296 18640 23348 18692
rect 23480 18640 23532 18692
rect 23848 18640 23900 18692
rect 24860 18572 24912 18624
rect 25044 18615 25096 18624
rect 25044 18581 25053 18615
rect 25053 18581 25087 18615
rect 25087 18581 25096 18615
rect 25044 18572 25096 18581
rect 26332 18572 26384 18624
rect 29368 18640 29420 18692
rect 27620 18572 27672 18624
rect 28080 18572 28132 18624
rect 28632 18615 28684 18624
rect 28632 18581 28641 18615
rect 28641 18581 28675 18615
rect 28675 18581 28684 18615
rect 28632 18572 28684 18581
rect 29184 18572 29236 18624
rect 29644 18572 29696 18624
rect 31300 18640 31352 18692
rect 31668 18708 31720 18760
rect 33048 18844 33100 18896
rect 39396 18912 39448 18964
rect 42064 18955 42116 18964
rect 42064 18921 42073 18955
rect 42073 18921 42107 18955
rect 42107 18921 42116 18955
rect 42064 18912 42116 18921
rect 34336 18776 34388 18828
rect 34520 18776 34572 18828
rect 36544 18776 36596 18828
rect 35256 18708 35308 18760
rect 38568 18819 38620 18828
rect 38568 18785 38577 18819
rect 38577 18785 38611 18819
rect 38611 18785 38620 18819
rect 38568 18776 38620 18785
rect 48780 18708 48832 18760
rect 49424 18708 49476 18760
rect 35624 18640 35676 18692
rect 37372 18640 37424 18692
rect 30472 18615 30524 18624
rect 30472 18581 30481 18615
rect 30481 18581 30515 18615
rect 30515 18581 30524 18615
rect 30472 18572 30524 18581
rect 30656 18572 30708 18624
rect 31576 18572 31628 18624
rect 33416 18572 33468 18624
rect 34244 18615 34296 18624
rect 34244 18581 34253 18615
rect 34253 18581 34287 18615
rect 34287 18581 34296 18615
rect 34244 18572 34296 18581
rect 34704 18572 34756 18624
rect 34888 18572 34940 18624
rect 37280 18572 37332 18624
rect 37556 18572 37608 18624
rect 39764 18640 39816 18692
rect 41052 18640 41104 18692
rect 38476 18615 38528 18624
rect 38476 18581 38485 18615
rect 38485 18581 38519 18615
rect 38519 18581 38528 18615
rect 38476 18572 38528 18581
rect 40132 18572 40184 18624
rect 40224 18572 40276 18624
rect 48412 18615 48464 18624
rect 48412 18581 48421 18615
rect 48421 18581 48455 18615
rect 48455 18581 48464 18615
rect 48412 18572 48464 18581
rect 48504 18572 48556 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 3608 18411 3660 18420
rect 3608 18377 3617 18411
rect 3617 18377 3651 18411
rect 3651 18377 3660 18411
rect 3608 18368 3660 18377
rect 9864 18368 9916 18420
rect 12440 18368 12492 18420
rect 4160 18300 4212 18352
rect 5632 18300 5684 18352
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 4068 18232 4120 18284
rect 4252 18164 4304 18216
rect 9772 18300 9824 18352
rect 11244 18300 11296 18352
rect 11520 18300 11572 18352
rect 13176 18343 13228 18352
rect 13176 18309 13185 18343
rect 13185 18309 13219 18343
rect 13219 18309 13228 18343
rect 13176 18300 13228 18309
rect 13912 18300 13964 18352
rect 16764 18300 16816 18352
rect 11796 18232 11848 18284
rect 12164 18232 12216 18284
rect 13452 18275 13504 18284
rect 13452 18241 13461 18275
rect 13461 18241 13495 18275
rect 13495 18241 13504 18275
rect 13452 18232 13504 18241
rect 10048 18096 10100 18148
rect 10968 18207 11020 18216
rect 10968 18173 10977 18207
rect 10977 18173 11011 18207
rect 11011 18173 11020 18207
rect 10968 18164 11020 18173
rect 14832 18232 14884 18284
rect 14556 18207 14608 18216
rect 14556 18173 14565 18207
rect 14565 18173 14599 18207
rect 14599 18173 14608 18207
rect 14556 18164 14608 18173
rect 9680 18028 9732 18080
rect 12072 18096 12124 18148
rect 13728 18096 13780 18148
rect 17868 18232 17920 18284
rect 16488 18164 16540 18216
rect 13636 18028 13688 18080
rect 15108 18028 15160 18080
rect 15292 18096 15344 18148
rect 16304 18028 16356 18080
rect 16948 18071 17000 18080
rect 16948 18037 16957 18071
rect 16957 18037 16991 18071
rect 16991 18037 17000 18071
rect 16948 18028 17000 18037
rect 18696 18368 18748 18420
rect 19156 18300 19208 18352
rect 21180 18300 21232 18352
rect 21640 18300 21692 18352
rect 25780 18368 25832 18420
rect 27252 18368 27304 18420
rect 27712 18368 27764 18420
rect 29736 18368 29788 18420
rect 31208 18368 31260 18420
rect 35532 18368 35584 18420
rect 36912 18411 36964 18420
rect 36912 18377 36921 18411
rect 36921 18377 36955 18411
rect 36955 18377 36964 18411
rect 36912 18368 36964 18377
rect 37372 18368 37424 18420
rect 38200 18368 38252 18420
rect 40776 18368 40828 18420
rect 48780 18411 48832 18420
rect 48780 18377 48789 18411
rect 48789 18377 48823 18411
rect 48823 18377 48832 18411
rect 48780 18368 48832 18377
rect 22652 18300 22704 18352
rect 23296 18343 23348 18352
rect 23296 18309 23305 18343
rect 23305 18309 23339 18343
rect 23339 18309 23348 18343
rect 23296 18300 23348 18309
rect 24124 18343 24176 18352
rect 24124 18309 24133 18343
rect 24133 18309 24167 18343
rect 24167 18309 24176 18343
rect 24124 18300 24176 18309
rect 24768 18300 24820 18352
rect 25228 18300 25280 18352
rect 32128 18300 32180 18352
rect 19432 18232 19484 18284
rect 23112 18232 23164 18284
rect 25044 18275 25096 18284
rect 25044 18241 25053 18275
rect 25053 18241 25087 18275
rect 25087 18241 25096 18275
rect 25044 18232 25096 18241
rect 19156 18164 19208 18216
rect 19616 18207 19668 18216
rect 19616 18173 19625 18207
rect 19625 18173 19659 18207
rect 19659 18173 19668 18207
rect 19616 18164 19668 18173
rect 21548 18164 21600 18216
rect 26332 18275 26384 18284
rect 26332 18241 26341 18275
rect 26341 18241 26375 18275
rect 26375 18241 26384 18275
rect 26332 18232 26384 18241
rect 29092 18232 29144 18284
rect 29368 18232 29420 18284
rect 21272 18028 21324 18080
rect 21456 18028 21508 18080
rect 26516 18207 26568 18216
rect 26516 18173 26525 18207
rect 26525 18173 26559 18207
rect 26559 18173 26568 18207
rect 26516 18164 26568 18173
rect 26608 18164 26660 18216
rect 23756 18096 23808 18148
rect 26056 18096 26108 18148
rect 25044 18028 25096 18080
rect 27160 18071 27212 18080
rect 27160 18037 27169 18071
rect 27169 18037 27203 18071
rect 27203 18037 27212 18071
rect 27160 18028 27212 18037
rect 27528 18028 27580 18080
rect 30104 18164 30156 18216
rect 32680 18275 32732 18284
rect 32680 18241 32689 18275
rect 32689 18241 32723 18275
rect 32723 18241 32732 18275
rect 32680 18232 32732 18241
rect 28540 18096 28592 18148
rect 31944 18164 31996 18216
rect 33600 18300 33652 18352
rect 34336 18300 34388 18352
rect 37004 18300 37056 18352
rect 37740 18300 37792 18352
rect 38752 18300 38804 18352
rect 40040 18300 40092 18352
rect 41052 18300 41104 18352
rect 35716 18232 35768 18284
rect 36360 18275 36412 18284
rect 36360 18241 36369 18275
rect 36369 18241 36403 18275
rect 36403 18241 36412 18275
rect 36360 18232 36412 18241
rect 33600 18207 33652 18216
rect 33600 18173 33609 18207
rect 33609 18173 33643 18207
rect 33643 18173 33652 18207
rect 33600 18164 33652 18173
rect 34612 18164 34664 18216
rect 36452 18164 36504 18216
rect 37280 18207 37332 18216
rect 37280 18173 37289 18207
rect 37289 18173 37323 18207
rect 37323 18173 37332 18207
rect 37280 18164 37332 18173
rect 37464 18232 37516 18284
rect 38016 18232 38068 18284
rect 39764 18275 39816 18284
rect 39764 18241 39773 18275
rect 39773 18241 39807 18275
rect 39807 18241 39816 18275
rect 39764 18232 39816 18241
rect 48412 18232 48464 18284
rect 49332 18275 49384 18284
rect 49332 18241 49341 18275
rect 49341 18241 49375 18275
rect 49375 18241 49384 18275
rect 49332 18232 49384 18241
rect 37740 18164 37792 18216
rect 37832 18164 37884 18216
rect 31024 18096 31076 18148
rect 29368 18028 29420 18080
rect 30104 18028 30156 18080
rect 32588 18028 32640 18080
rect 38016 18139 38068 18148
rect 38016 18105 38025 18139
rect 38025 18105 38059 18139
rect 38059 18105 38068 18139
rect 38016 18096 38068 18105
rect 35624 18028 35676 18080
rect 36360 18028 36412 18080
rect 37096 18028 37148 18080
rect 37280 18028 37332 18080
rect 40224 18028 40276 18080
rect 48320 18028 48372 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 10140 17867 10192 17876
rect 10140 17833 10149 17867
rect 10149 17833 10183 17867
rect 10183 17833 10192 17867
rect 10140 17824 10192 17833
rect 10968 17824 11020 17876
rect 9864 17756 9916 17808
rect 12348 17824 12400 17876
rect 12624 17824 12676 17876
rect 14556 17824 14608 17876
rect 15200 17824 15252 17876
rect 15752 17824 15804 17876
rect 17224 17824 17276 17876
rect 19340 17824 19392 17876
rect 19616 17824 19668 17876
rect 21364 17824 21416 17876
rect 21548 17824 21600 17876
rect 11428 17688 11480 17740
rect 12532 17688 12584 17740
rect 13452 17688 13504 17740
rect 10232 17620 10284 17672
rect 13360 17620 13412 17672
rect 940 17552 992 17604
rect 10140 17552 10192 17604
rect 12072 17595 12124 17604
rect 12072 17561 12081 17595
rect 12081 17561 12115 17595
rect 12115 17561 12124 17595
rect 12072 17552 12124 17561
rect 14740 17688 14792 17740
rect 15384 17688 15436 17740
rect 16028 17731 16080 17740
rect 16028 17697 16037 17731
rect 16037 17697 16071 17731
rect 16071 17697 16080 17731
rect 16028 17688 16080 17697
rect 11152 17484 11204 17536
rect 13636 17484 13688 17536
rect 16212 17552 16264 17604
rect 20720 17756 20772 17808
rect 22284 17756 22336 17808
rect 23572 17756 23624 17808
rect 16856 17731 16908 17740
rect 16856 17697 16865 17731
rect 16865 17697 16899 17731
rect 16899 17697 16908 17731
rect 16856 17688 16908 17697
rect 16948 17688 17000 17740
rect 19708 17688 19760 17740
rect 20352 17688 20404 17740
rect 21732 17731 21784 17740
rect 21732 17697 21741 17731
rect 21741 17697 21775 17731
rect 21775 17697 21784 17731
rect 21732 17688 21784 17697
rect 22100 17688 22152 17740
rect 24952 17688 25004 17740
rect 25044 17731 25096 17740
rect 25044 17697 25053 17731
rect 25053 17697 25087 17731
rect 25087 17697 25096 17731
rect 25044 17688 25096 17697
rect 16488 17620 16540 17672
rect 18604 17552 18656 17604
rect 16488 17527 16540 17536
rect 16488 17493 16497 17527
rect 16497 17493 16531 17527
rect 16531 17493 16540 17527
rect 16488 17484 16540 17493
rect 17408 17484 17460 17536
rect 18880 17484 18932 17536
rect 20352 17484 20404 17536
rect 23480 17620 23532 17672
rect 30932 17824 30984 17876
rect 31392 17824 31444 17876
rect 26332 17799 26384 17808
rect 26332 17765 26341 17799
rect 26341 17765 26375 17799
rect 26375 17765 26384 17799
rect 26332 17756 26384 17765
rect 29828 17756 29880 17808
rect 26424 17688 26476 17740
rect 31392 17688 31444 17740
rect 31484 17731 31536 17740
rect 31484 17697 31493 17731
rect 31493 17697 31527 17731
rect 31527 17697 31536 17731
rect 31484 17688 31536 17697
rect 27436 17620 27488 17672
rect 28908 17620 28960 17672
rect 33692 17824 33744 17876
rect 33876 17867 33928 17876
rect 33876 17833 33885 17867
rect 33885 17833 33919 17867
rect 33919 17833 33928 17867
rect 33876 17824 33928 17833
rect 32864 17756 32916 17808
rect 34336 17756 34388 17808
rect 38476 17824 38528 17876
rect 32956 17731 33008 17740
rect 32956 17697 32965 17731
rect 32965 17697 32999 17731
rect 32999 17697 33008 17731
rect 32956 17688 33008 17697
rect 33508 17688 33560 17740
rect 34612 17688 34664 17740
rect 21640 17552 21692 17604
rect 21824 17552 21876 17604
rect 24492 17552 24544 17604
rect 26516 17552 26568 17604
rect 22192 17484 22244 17536
rect 23756 17527 23808 17536
rect 23756 17493 23765 17527
rect 23765 17493 23799 17527
rect 23799 17493 23808 17527
rect 23756 17484 23808 17493
rect 24676 17484 24728 17536
rect 25044 17484 25096 17536
rect 26976 17484 27028 17536
rect 27068 17527 27120 17536
rect 27068 17493 27077 17527
rect 27077 17493 27111 17527
rect 27111 17493 27120 17527
rect 27068 17484 27120 17493
rect 27528 17484 27580 17536
rect 28632 17552 28684 17604
rect 29920 17595 29972 17604
rect 29920 17561 29929 17595
rect 29929 17561 29963 17595
rect 29963 17561 29972 17595
rect 29920 17552 29972 17561
rect 31484 17552 31536 17604
rect 33876 17620 33928 17672
rect 29000 17484 29052 17536
rect 29184 17527 29236 17536
rect 29184 17493 29193 17527
rect 29193 17493 29227 17527
rect 29227 17493 29236 17527
rect 29184 17484 29236 17493
rect 30012 17484 30064 17536
rect 33232 17552 33284 17604
rect 35072 17620 35124 17672
rect 35256 17620 35308 17672
rect 36728 17688 36780 17740
rect 37280 17688 37332 17740
rect 37556 17663 37608 17672
rect 37556 17629 37565 17663
rect 37565 17629 37599 17663
rect 37599 17629 37608 17663
rect 37556 17620 37608 17629
rect 40868 17756 40920 17808
rect 40684 17688 40736 17740
rect 41052 17731 41104 17740
rect 41052 17697 41061 17731
rect 41061 17697 41095 17731
rect 41095 17697 41104 17731
rect 41052 17688 41104 17697
rect 43444 17756 43496 17808
rect 49332 17663 49384 17672
rect 49332 17629 49341 17663
rect 49341 17629 49375 17663
rect 49375 17629 49384 17663
rect 49332 17620 49384 17629
rect 37004 17552 37056 17604
rect 37372 17552 37424 17604
rect 48412 17552 48464 17604
rect 32128 17484 32180 17536
rect 32312 17484 32364 17536
rect 32680 17484 32732 17536
rect 33324 17484 33376 17536
rect 34520 17527 34572 17536
rect 34520 17493 34529 17527
rect 34529 17493 34563 17527
rect 34563 17493 34572 17527
rect 34520 17484 34572 17493
rect 35072 17527 35124 17536
rect 35072 17493 35081 17527
rect 35081 17493 35115 17527
rect 35115 17493 35124 17527
rect 35072 17484 35124 17493
rect 35532 17484 35584 17536
rect 36636 17484 36688 17536
rect 38936 17484 38988 17536
rect 40040 17484 40092 17536
rect 48688 17527 48740 17536
rect 48688 17493 48697 17527
rect 48697 17493 48731 17527
rect 48731 17493 48740 17527
rect 48688 17484 48740 17493
rect 49148 17527 49200 17536
rect 49148 17493 49157 17527
rect 49157 17493 49191 17527
rect 49191 17493 49200 17527
rect 49148 17484 49200 17493
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 13820 17323 13872 17332
rect 1032 17076 1084 17128
rect 2136 17008 2188 17060
rect 13820 17289 13829 17323
rect 13829 17289 13863 17323
rect 13863 17289 13872 17323
rect 13820 17280 13872 17289
rect 14004 17280 14056 17332
rect 15568 17323 15620 17332
rect 15568 17289 15577 17323
rect 15577 17289 15611 17323
rect 15611 17289 15620 17323
rect 15568 17280 15620 17289
rect 10416 17212 10468 17264
rect 4344 17144 4396 17196
rect 5908 17144 5960 17196
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 9956 17144 10008 17196
rect 11428 17212 11480 17264
rect 11888 17255 11940 17264
rect 11888 17221 11897 17255
rect 11897 17221 11931 17255
rect 11931 17221 11940 17255
rect 11888 17212 11940 17221
rect 12348 17212 12400 17264
rect 13268 17212 13320 17264
rect 14096 17212 14148 17264
rect 14740 17212 14792 17264
rect 15752 17212 15804 17264
rect 16028 17212 16080 17264
rect 17960 17255 18012 17264
rect 17960 17221 17969 17255
rect 17969 17221 18003 17255
rect 18003 17221 18012 17255
rect 17960 17212 18012 17221
rect 18696 17255 18748 17264
rect 18696 17221 18705 17255
rect 18705 17221 18739 17255
rect 18739 17221 18748 17255
rect 18696 17212 18748 17221
rect 19156 17323 19208 17332
rect 19156 17289 19165 17323
rect 19165 17289 19199 17323
rect 19199 17289 19208 17323
rect 19156 17280 19208 17289
rect 20260 17280 20312 17332
rect 21732 17280 21784 17332
rect 22008 17280 22060 17332
rect 23480 17280 23532 17332
rect 24032 17280 24084 17332
rect 27712 17323 27764 17332
rect 27712 17289 27721 17323
rect 27721 17289 27755 17323
rect 27755 17289 27764 17323
rect 27712 17280 27764 17289
rect 27804 17280 27856 17332
rect 32312 17280 32364 17332
rect 20536 17212 20588 17264
rect 20996 17212 21048 17264
rect 21456 17212 21508 17264
rect 23664 17212 23716 17264
rect 24124 17212 24176 17264
rect 11980 17144 12032 17196
rect 10600 17076 10652 17128
rect 12348 17076 12400 17128
rect 12716 17008 12768 17060
rect 9496 16983 9548 16992
rect 9496 16949 9505 16983
rect 9505 16949 9539 16983
rect 9539 16949 9548 16983
rect 9496 16940 9548 16949
rect 10508 16940 10560 16992
rect 10600 16940 10652 16992
rect 11980 16940 12032 16992
rect 12808 16940 12860 16992
rect 15108 17187 15160 17196
rect 15108 17153 15117 17187
rect 15117 17153 15151 17187
rect 15151 17153 15160 17187
rect 15108 17144 15160 17153
rect 14280 17076 14332 17128
rect 16856 17144 16908 17196
rect 19340 17144 19392 17196
rect 22100 17144 22152 17196
rect 22744 17144 22796 17196
rect 25780 17212 25832 17264
rect 25964 17212 26016 17264
rect 26148 17212 26200 17264
rect 27620 17212 27672 17264
rect 25596 17144 25648 17196
rect 26332 17144 26384 17196
rect 27712 17144 27764 17196
rect 28816 17212 28868 17264
rect 29828 17212 29880 17264
rect 16120 17119 16172 17128
rect 16120 17085 16129 17119
rect 16129 17085 16163 17119
rect 16163 17085 16172 17119
rect 16120 17076 16172 17085
rect 16396 17076 16448 17128
rect 21180 17076 21232 17128
rect 21640 17119 21692 17128
rect 21640 17085 21649 17119
rect 21649 17085 21683 17119
rect 21683 17085 21692 17119
rect 21640 17076 21692 17085
rect 22008 17076 22060 17128
rect 23388 17076 23440 17128
rect 24492 17076 24544 17128
rect 25504 17119 25556 17128
rect 25504 17085 25513 17119
rect 25513 17085 25547 17119
rect 25547 17085 25556 17119
rect 25504 17076 25556 17085
rect 28448 17144 28500 17196
rect 29276 17144 29328 17196
rect 30288 17212 30340 17264
rect 33600 17280 33652 17332
rect 35072 17280 35124 17332
rect 16488 17008 16540 17060
rect 13452 16983 13504 16992
rect 13452 16949 13461 16983
rect 13461 16949 13495 16983
rect 13495 16949 13504 16983
rect 13452 16940 13504 16949
rect 14188 16983 14240 16992
rect 14188 16949 14197 16983
rect 14197 16949 14231 16983
rect 14231 16949 14240 16983
rect 14188 16940 14240 16949
rect 15936 16940 15988 16992
rect 17408 16983 17460 16992
rect 17408 16949 17417 16983
rect 17417 16949 17451 16983
rect 17451 16949 17460 16983
rect 17408 16940 17460 16949
rect 21640 16940 21692 16992
rect 25136 17008 25188 17060
rect 26516 17008 26568 17060
rect 27528 17008 27580 17060
rect 29000 17076 29052 17128
rect 29460 17076 29512 17128
rect 30564 17144 30616 17196
rect 31392 17187 31444 17196
rect 31392 17153 31401 17187
rect 31401 17153 31435 17187
rect 31435 17153 31444 17187
rect 31392 17144 31444 17153
rect 31484 17144 31536 17196
rect 32220 17144 32272 17196
rect 33048 17212 33100 17264
rect 35532 17255 35584 17264
rect 35532 17221 35541 17255
rect 35541 17221 35575 17255
rect 35575 17221 35584 17255
rect 35532 17212 35584 17221
rect 48320 17280 48372 17332
rect 48412 17323 48464 17332
rect 48412 17289 48421 17323
rect 48421 17289 48455 17323
rect 48455 17289 48464 17323
rect 48412 17280 48464 17289
rect 35164 17144 35216 17196
rect 36360 17187 36412 17196
rect 36360 17153 36369 17187
rect 36369 17153 36403 17187
rect 36403 17153 36412 17187
rect 36360 17144 36412 17153
rect 30288 17076 30340 17128
rect 30748 17076 30800 17128
rect 32588 17119 32640 17128
rect 32588 17085 32597 17119
rect 32597 17085 32631 17119
rect 32631 17085 32640 17119
rect 32588 17076 32640 17085
rect 32956 17076 33008 17128
rect 34796 17119 34848 17128
rect 34796 17085 34805 17119
rect 34805 17085 34839 17119
rect 34839 17085 34848 17119
rect 34796 17076 34848 17085
rect 36176 17119 36228 17128
rect 36176 17085 36185 17119
rect 36185 17085 36219 17119
rect 36219 17085 36228 17119
rect 36176 17076 36228 17085
rect 32312 17008 32364 17060
rect 33692 17008 33744 17060
rect 36084 17008 36136 17060
rect 39948 17212 40000 17264
rect 40132 17212 40184 17264
rect 40960 17255 41012 17264
rect 40960 17221 40969 17255
rect 40969 17221 41003 17255
rect 41003 17221 41012 17255
rect 40960 17212 41012 17221
rect 48228 17212 48280 17264
rect 48688 17212 48740 17264
rect 38936 17144 38988 17196
rect 48780 17144 48832 17196
rect 37832 17076 37884 17128
rect 40684 17119 40736 17128
rect 40684 17085 40693 17119
rect 40693 17085 40727 17119
rect 40727 17085 40736 17119
rect 40684 17076 40736 17085
rect 49056 17119 49108 17128
rect 49056 17085 49065 17119
rect 49065 17085 49099 17119
rect 49099 17085 49108 17119
rect 49056 17076 49108 17085
rect 29460 16940 29512 16992
rect 30564 16983 30616 16992
rect 30564 16949 30573 16983
rect 30573 16949 30607 16983
rect 30607 16949 30616 16983
rect 30564 16940 30616 16949
rect 33784 16940 33836 16992
rect 35624 16940 35676 16992
rect 37188 17008 37240 17060
rect 36728 16983 36780 16992
rect 36728 16949 36737 16983
rect 36737 16949 36771 16983
rect 36771 16949 36780 16983
rect 36728 16940 36780 16949
rect 38752 16940 38804 16992
rect 38844 16940 38896 16992
rect 41052 17008 41104 17060
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 14188 16736 14240 16788
rect 14648 16736 14700 16788
rect 4436 16668 4488 16720
rect 5448 16668 5500 16720
rect 10232 16668 10284 16720
rect 12440 16668 12492 16720
rect 13820 16668 13872 16720
rect 10876 16600 10928 16652
rect 9036 16532 9088 16584
rect 1032 16464 1084 16516
rect 7840 16464 7892 16516
rect 9680 16464 9732 16516
rect 10508 16507 10560 16516
rect 10508 16473 10517 16507
rect 10517 16473 10551 16507
rect 10551 16473 10560 16507
rect 10508 16464 10560 16473
rect 12624 16464 12676 16516
rect 12808 16532 12860 16584
rect 13544 16532 13596 16584
rect 15384 16600 15436 16652
rect 16672 16668 16724 16720
rect 14924 16532 14976 16584
rect 16672 16532 16724 16584
rect 9036 16439 9088 16448
rect 9036 16405 9045 16439
rect 9045 16405 9079 16439
rect 9079 16405 9088 16439
rect 9036 16396 9088 16405
rect 11336 16439 11388 16448
rect 11336 16405 11345 16439
rect 11345 16405 11379 16439
rect 11379 16405 11388 16439
rect 11336 16396 11388 16405
rect 11980 16396 12032 16448
rect 12900 16396 12952 16448
rect 13544 16396 13596 16448
rect 13636 16396 13688 16448
rect 14188 16439 14240 16448
rect 14188 16405 14197 16439
rect 14197 16405 14231 16439
rect 14231 16405 14240 16439
rect 14188 16396 14240 16405
rect 14740 16439 14792 16448
rect 14740 16405 14749 16439
rect 14749 16405 14783 16439
rect 14783 16405 14792 16439
rect 14740 16396 14792 16405
rect 14832 16439 14884 16448
rect 14832 16405 14841 16439
rect 14841 16405 14875 16439
rect 14875 16405 14884 16439
rect 14832 16396 14884 16405
rect 15476 16396 15528 16448
rect 15660 16439 15712 16448
rect 15660 16405 15669 16439
rect 15669 16405 15703 16439
rect 15703 16405 15712 16439
rect 15660 16396 15712 16405
rect 16396 16396 16448 16448
rect 17132 16439 17184 16448
rect 17132 16405 17141 16439
rect 17141 16405 17175 16439
rect 17175 16405 17184 16439
rect 17132 16396 17184 16405
rect 18880 16736 18932 16788
rect 20996 16779 21048 16788
rect 20996 16745 21005 16779
rect 21005 16745 21039 16779
rect 21039 16745 21048 16779
rect 20996 16736 21048 16745
rect 21180 16736 21232 16788
rect 20168 16668 20220 16720
rect 17960 16600 18012 16652
rect 19156 16600 19208 16652
rect 20628 16600 20680 16652
rect 22376 16600 22428 16652
rect 22836 16668 22888 16720
rect 23296 16736 23348 16788
rect 27620 16736 27672 16788
rect 28632 16736 28684 16788
rect 28816 16779 28868 16788
rect 28816 16745 28825 16779
rect 28825 16745 28859 16779
rect 28859 16745 28868 16779
rect 28816 16736 28868 16745
rect 22744 16643 22796 16652
rect 22744 16609 22753 16643
rect 22753 16609 22787 16643
rect 22787 16609 22796 16643
rect 22744 16600 22796 16609
rect 17500 16532 17552 16584
rect 26056 16668 26108 16720
rect 27804 16668 27856 16720
rect 31116 16736 31168 16788
rect 25872 16600 25924 16652
rect 26424 16600 26476 16652
rect 27068 16643 27120 16652
rect 27068 16609 27077 16643
rect 27077 16609 27111 16643
rect 27111 16609 27120 16643
rect 27068 16600 27120 16609
rect 27436 16600 27488 16652
rect 27988 16643 28040 16652
rect 27988 16609 27997 16643
rect 27997 16609 28031 16643
rect 28031 16609 28040 16643
rect 27988 16600 28040 16609
rect 18788 16396 18840 16448
rect 20536 16396 20588 16448
rect 20812 16396 20864 16448
rect 22008 16464 22060 16516
rect 24584 16507 24636 16516
rect 24584 16473 24593 16507
rect 24593 16473 24627 16507
rect 24627 16473 24636 16507
rect 24584 16464 24636 16473
rect 27804 16532 27856 16584
rect 26792 16464 26844 16516
rect 22836 16396 22888 16448
rect 22928 16396 22980 16448
rect 23664 16439 23716 16448
rect 23664 16405 23673 16439
rect 23673 16405 23707 16439
rect 23707 16405 23716 16439
rect 23664 16396 23716 16405
rect 25136 16396 25188 16448
rect 28264 16600 28316 16652
rect 29276 16643 29328 16652
rect 29276 16609 29285 16643
rect 29285 16609 29319 16643
rect 29319 16609 29328 16643
rect 29276 16600 29328 16609
rect 30104 16600 30156 16652
rect 30196 16600 30248 16652
rect 34612 16736 34664 16788
rect 36360 16736 36412 16788
rect 36452 16736 36504 16788
rect 36636 16736 36688 16788
rect 37188 16736 37240 16788
rect 37464 16736 37516 16788
rect 40224 16736 40276 16788
rect 40960 16736 41012 16788
rect 41328 16736 41380 16788
rect 34060 16668 34112 16720
rect 31944 16600 31996 16652
rect 32220 16643 32272 16652
rect 32220 16609 32229 16643
rect 32229 16609 32263 16643
rect 32263 16609 32272 16643
rect 32220 16600 32272 16609
rect 33692 16600 33744 16652
rect 37556 16668 37608 16720
rect 35348 16600 35400 16652
rect 28356 16575 28408 16584
rect 28356 16541 28365 16575
rect 28365 16541 28399 16575
rect 28399 16541 28408 16575
rect 28356 16532 28408 16541
rect 28632 16464 28684 16516
rect 29000 16464 29052 16516
rect 29092 16464 29144 16516
rect 29736 16396 29788 16448
rect 31944 16464 31996 16516
rect 35532 16532 35584 16584
rect 36820 16643 36872 16652
rect 36820 16609 36829 16643
rect 36829 16609 36863 16643
rect 36863 16609 36872 16643
rect 36820 16600 36872 16609
rect 37464 16600 37516 16652
rect 38844 16600 38896 16652
rect 40316 16600 40368 16652
rect 41236 16711 41288 16720
rect 41236 16677 41245 16711
rect 41245 16677 41279 16711
rect 41279 16677 41288 16711
rect 41236 16668 41288 16677
rect 46020 16736 46072 16788
rect 48780 16779 48832 16788
rect 48780 16745 48789 16779
rect 48789 16745 48823 16779
rect 48823 16745 48832 16779
rect 48780 16736 48832 16745
rect 39488 16575 39540 16584
rect 39488 16541 39497 16575
rect 39497 16541 39531 16575
rect 39531 16541 39540 16575
rect 39488 16532 39540 16541
rect 40684 16532 40736 16584
rect 49424 16532 49476 16584
rect 32772 16464 32824 16516
rect 32956 16464 33008 16516
rect 35900 16464 35952 16516
rect 36084 16464 36136 16516
rect 36820 16464 36872 16516
rect 38752 16464 38804 16516
rect 39948 16464 40000 16516
rect 40224 16464 40276 16516
rect 41236 16464 41288 16516
rect 31208 16439 31260 16448
rect 31208 16405 31217 16439
rect 31217 16405 31251 16439
rect 31251 16405 31260 16439
rect 31208 16396 31260 16405
rect 31300 16439 31352 16448
rect 31300 16405 31309 16439
rect 31309 16405 31343 16439
rect 31343 16405 31352 16439
rect 31300 16396 31352 16405
rect 31668 16439 31720 16448
rect 31668 16405 31677 16439
rect 31677 16405 31711 16439
rect 31711 16405 31720 16439
rect 31668 16396 31720 16405
rect 32680 16396 32732 16448
rect 33416 16396 33468 16448
rect 33968 16439 34020 16448
rect 33968 16405 33977 16439
rect 33977 16405 34011 16439
rect 34011 16405 34020 16439
rect 33968 16396 34020 16405
rect 34612 16396 34664 16448
rect 35808 16396 35860 16448
rect 37188 16396 37240 16448
rect 38568 16396 38620 16448
rect 40960 16396 41012 16448
rect 49148 16439 49200 16448
rect 49148 16405 49157 16439
rect 49157 16405 49191 16439
rect 49191 16405 49200 16439
rect 49148 16396 49200 16405
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 8300 16235 8352 16244
rect 8300 16201 8309 16235
rect 8309 16201 8343 16235
rect 8343 16201 8352 16235
rect 8300 16192 8352 16201
rect 9220 16235 9272 16244
rect 9220 16201 9229 16235
rect 9229 16201 9263 16235
rect 9263 16201 9272 16235
rect 9220 16192 9272 16201
rect 9772 16192 9824 16244
rect 11060 16192 11112 16244
rect 11336 16192 11388 16244
rect 13636 16235 13688 16244
rect 13636 16201 13645 16235
rect 13645 16201 13679 16235
rect 13679 16201 13688 16235
rect 13636 16192 13688 16201
rect 10876 16124 10928 16176
rect 4252 16056 4304 16108
rect 1032 15988 1084 16040
rect 9036 15988 9088 16040
rect 12164 16056 12216 16108
rect 15844 16192 15896 16244
rect 15016 16124 15068 16176
rect 18328 16192 18380 16244
rect 18696 16192 18748 16244
rect 21272 16192 21324 16244
rect 21456 16192 21508 16244
rect 22652 16192 22704 16244
rect 23388 16192 23440 16244
rect 24676 16192 24728 16244
rect 24768 16192 24820 16244
rect 26608 16192 26660 16244
rect 26792 16192 26844 16244
rect 26976 16192 27028 16244
rect 27436 16192 27488 16244
rect 28356 16192 28408 16244
rect 30564 16192 30616 16244
rect 32036 16192 32088 16244
rect 32956 16192 33008 16244
rect 33692 16192 33744 16244
rect 33784 16235 33836 16244
rect 33784 16201 33793 16235
rect 33793 16201 33827 16235
rect 33827 16201 33836 16235
rect 33784 16192 33836 16201
rect 34796 16192 34848 16244
rect 17132 16124 17184 16176
rect 14464 16056 14516 16108
rect 9772 15920 9824 15972
rect 9864 15852 9916 15904
rect 10600 15852 10652 15904
rect 11520 15852 11572 15904
rect 13636 15988 13688 16040
rect 14280 15988 14332 16040
rect 13544 15920 13596 15972
rect 15292 16056 15344 16108
rect 15384 16056 15436 16108
rect 14924 16031 14976 16040
rect 14924 15997 14933 16031
rect 14933 15997 14967 16031
rect 14967 15997 14976 16031
rect 14924 15988 14976 15997
rect 16120 16056 16172 16108
rect 15844 16031 15896 16040
rect 15844 15997 15853 16031
rect 15853 15997 15887 16031
rect 15887 15997 15896 16031
rect 15844 15988 15896 15997
rect 17132 15988 17184 16040
rect 15936 15920 15988 15972
rect 17592 15920 17644 15972
rect 16396 15852 16448 15904
rect 16948 15895 17000 15904
rect 16948 15861 16957 15895
rect 16957 15861 16991 15895
rect 16991 15861 17000 15895
rect 16948 15852 17000 15861
rect 17224 15852 17276 15904
rect 20812 16124 20864 16176
rect 20904 16124 20956 16176
rect 19156 16099 19208 16108
rect 19156 16065 19165 16099
rect 19165 16065 19199 16099
rect 19199 16065 19208 16099
rect 19156 16056 19208 16065
rect 21548 16124 21600 16176
rect 21916 16124 21968 16176
rect 25780 16124 25832 16176
rect 27804 16124 27856 16176
rect 22928 16056 22980 16108
rect 23480 16099 23532 16108
rect 23480 16065 23489 16099
rect 23489 16065 23523 16099
rect 23523 16065 23532 16099
rect 23480 16056 23532 16065
rect 28908 16124 28960 16176
rect 29184 16124 29236 16176
rect 29920 16124 29972 16176
rect 30656 16124 30708 16176
rect 30840 16167 30892 16176
rect 30840 16133 30849 16167
rect 30849 16133 30883 16167
rect 30883 16133 30892 16167
rect 30840 16124 30892 16133
rect 31668 16124 31720 16176
rect 19984 15988 20036 16040
rect 20996 15988 21048 16040
rect 21916 15988 21968 16040
rect 20444 15920 20496 15972
rect 22100 15920 22152 15972
rect 23388 16031 23440 16040
rect 23388 15997 23397 16031
rect 23397 15997 23431 16031
rect 23431 15997 23440 16031
rect 23388 15988 23440 15997
rect 24492 15988 24544 16040
rect 26056 16031 26108 16040
rect 26056 15997 26065 16031
rect 26065 15997 26099 16031
rect 26099 15997 26108 16031
rect 26056 15988 26108 15997
rect 26884 15988 26936 16040
rect 28632 16031 28684 16040
rect 28632 15997 28641 16031
rect 28641 15997 28675 16031
rect 28675 15997 28684 16031
rect 28632 15988 28684 15997
rect 29828 15988 29880 16040
rect 31208 15988 31260 16040
rect 18420 15852 18472 15904
rect 20812 15852 20864 15904
rect 22008 15852 22060 15904
rect 26700 15852 26752 15904
rect 27252 15852 27304 15904
rect 32036 15920 32088 15972
rect 30748 15852 30800 15904
rect 31208 15852 31260 15904
rect 31484 15852 31536 15904
rect 32404 16031 32456 16040
rect 32404 15997 32413 16031
rect 32413 15997 32447 16031
rect 32447 15997 32456 16031
rect 32404 15988 32456 15997
rect 33324 16056 33376 16108
rect 35532 16056 35584 16108
rect 37096 16192 37148 16244
rect 40960 16235 41012 16244
rect 40960 16201 40969 16235
rect 40969 16201 41003 16235
rect 41003 16201 41012 16235
rect 40960 16192 41012 16201
rect 41420 16192 41472 16244
rect 38568 16124 38620 16176
rect 39948 16124 40000 16176
rect 37372 16056 37424 16108
rect 48688 16056 48740 16108
rect 49332 16099 49384 16108
rect 49332 16065 49341 16099
rect 49341 16065 49375 16099
rect 49375 16065 49384 16099
rect 49332 16056 49384 16065
rect 32772 15988 32824 16040
rect 34428 15988 34480 16040
rect 35164 16031 35216 16040
rect 35164 15997 35173 16031
rect 35173 15997 35207 16031
rect 35207 15997 35216 16031
rect 35164 15988 35216 15997
rect 36084 15988 36136 16040
rect 37004 15988 37056 16040
rect 39212 15988 39264 16040
rect 41788 15988 41840 16040
rect 32772 15852 32824 15904
rect 32864 15852 32916 15904
rect 37280 15920 37332 15972
rect 49148 15963 49200 15972
rect 49148 15929 49157 15963
rect 49157 15929 49191 15963
rect 49191 15929 49200 15963
rect 49148 15920 49200 15929
rect 38568 15852 38620 15904
rect 40316 15852 40368 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 10692 15648 10744 15700
rect 11520 15648 11572 15700
rect 15292 15648 15344 15700
rect 16764 15691 16816 15700
rect 16764 15657 16773 15691
rect 16773 15657 16807 15691
rect 16807 15657 16816 15691
rect 16764 15648 16816 15657
rect 17316 15648 17368 15700
rect 20812 15648 20864 15700
rect 22468 15691 22520 15700
rect 22468 15657 22477 15691
rect 22477 15657 22511 15691
rect 22511 15657 22520 15691
rect 22468 15648 22520 15657
rect 22560 15648 22612 15700
rect 11060 15512 11112 15564
rect 14280 15580 14332 15632
rect 17500 15580 17552 15632
rect 18604 15580 18656 15632
rect 18972 15623 19024 15632
rect 18972 15589 18981 15623
rect 18981 15589 19015 15623
rect 19015 15589 19024 15623
rect 18972 15580 19024 15589
rect 19340 15580 19392 15632
rect 12532 15555 12584 15564
rect 12532 15521 12541 15555
rect 12541 15521 12575 15555
rect 12575 15521 12584 15555
rect 12532 15512 12584 15521
rect 14096 15512 14148 15564
rect 14924 15555 14976 15564
rect 14924 15521 14933 15555
rect 14933 15521 14967 15555
rect 14967 15521 14976 15555
rect 14924 15512 14976 15521
rect 16120 15555 16172 15564
rect 16120 15521 16129 15555
rect 16129 15521 16163 15555
rect 16163 15521 16172 15555
rect 16120 15512 16172 15521
rect 16212 15512 16264 15564
rect 16488 15512 16540 15564
rect 19524 15512 19576 15564
rect 22100 15580 22152 15632
rect 24032 15580 24084 15632
rect 29184 15580 29236 15632
rect 21272 15512 21324 15564
rect 21456 15512 21508 15564
rect 22008 15512 22060 15564
rect 24768 15512 24820 15564
rect 25320 15512 25372 15564
rect 26608 15512 26660 15564
rect 28724 15555 28776 15564
rect 28724 15521 28733 15555
rect 28733 15521 28767 15555
rect 28767 15521 28776 15555
rect 28724 15512 28776 15521
rect 31116 15512 31168 15564
rect 32588 15648 32640 15700
rect 33692 15648 33744 15700
rect 35532 15648 35584 15700
rect 37280 15648 37332 15700
rect 37740 15691 37792 15700
rect 37740 15657 37749 15691
rect 37749 15657 37783 15691
rect 37783 15657 37792 15691
rect 37740 15648 37792 15657
rect 41420 15648 41472 15700
rect 48688 15648 48740 15700
rect 31852 15580 31904 15632
rect 41788 15623 41840 15632
rect 41788 15589 41797 15623
rect 41797 15589 41831 15623
rect 41831 15589 41840 15623
rect 41788 15580 41840 15589
rect 10232 15444 10284 15496
rect 11152 15444 11204 15496
rect 12716 15444 12768 15496
rect 13452 15444 13504 15496
rect 18420 15444 18472 15496
rect 20904 15444 20956 15496
rect 21180 15444 21232 15496
rect 22468 15444 22520 15496
rect 27344 15444 27396 15496
rect 27712 15444 27764 15496
rect 940 15376 992 15428
rect 4160 15376 4212 15428
rect 9036 15351 9088 15360
rect 9036 15317 9045 15351
rect 9045 15317 9079 15351
rect 9079 15317 9088 15351
rect 9036 15308 9088 15317
rect 15936 15419 15988 15428
rect 15936 15385 15945 15419
rect 15945 15385 15979 15419
rect 15979 15385 15988 15419
rect 15936 15376 15988 15385
rect 16396 15376 16448 15428
rect 11888 15308 11940 15360
rect 12808 15308 12860 15360
rect 13544 15308 13596 15360
rect 13912 15308 13964 15360
rect 14648 15351 14700 15360
rect 14648 15317 14657 15351
rect 14657 15317 14691 15351
rect 14691 15317 14700 15351
rect 14648 15308 14700 15317
rect 15568 15351 15620 15360
rect 15568 15317 15577 15351
rect 15577 15317 15611 15351
rect 15611 15317 15620 15351
rect 15568 15308 15620 15317
rect 16120 15308 16172 15360
rect 17132 15351 17184 15360
rect 17132 15317 17141 15351
rect 17141 15317 17175 15351
rect 17175 15317 17184 15351
rect 17132 15308 17184 15317
rect 17316 15308 17368 15360
rect 18512 15376 18564 15428
rect 21456 15376 21508 15428
rect 19800 15308 19852 15360
rect 20260 15351 20312 15360
rect 20260 15317 20269 15351
rect 20269 15317 20303 15351
rect 20303 15317 20312 15351
rect 20260 15308 20312 15317
rect 21088 15308 21140 15360
rect 22100 15376 22152 15428
rect 22284 15351 22336 15360
rect 22284 15317 22293 15351
rect 22293 15317 22327 15351
rect 22327 15317 22336 15351
rect 22284 15308 22336 15317
rect 25688 15376 25740 15428
rect 26332 15419 26384 15428
rect 26332 15385 26341 15419
rect 26341 15385 26375 15419
rect 26375 15385 26384 15419
rect 26332 15376 26384 15385
rect 26976 15376 27028 15428
rect 30288 15376 30340 15428
rect 30748 15419 30800 15428
rect 30748 15385 30757 15419
rect 30757 15385 30791 15419
rect 30791 15385 30800 15419
rect 30748 15376 30800 15385
rect 31208 15376 31260 15428
rect 34796 15512 34848 15564
rect 35900 15512 35952 15564
rect 37372 15512 37424 15564
rect 39488 15555 39540 15564
rect 39488 15521 39497 15555
rect 39497 15521 39531 15555
rect 39531 15521 39540 15555
rect 39488 15512 39540 15521
rect 40316 15555 40368 15564
rect 40316 15521 40325 15555
rect 40325 15521 40359 15555
rect 40359 15521 40368 15555
rect 40316 15512 40368 15521
rect 34060 15444 34112 15496
rect 49332 15487 49384 15496
rect 49332 15453 49341 15487
rect 49341 15453 49375 15487
rect 49375 15453 49384 15487
rect 49332 15444 49384 15453
rect 34612 15376 34664 15428
rect 35624 15376 35676 15428
rect 38752 15376 38804 15428
rect 39212 15419 39264 15428
rect 39212 15385 39221 15419
rect 39221 15385 39255 15419
rect 39255 15385 39264 15419
rect 39212 15376 39264 15385
rect 39948 15376 40000 15428
rect 25136 15351 25188 15360
rect 25136 15317 25145 15351
rect 25145 15317 25179 15351
rect 25179 15317 25188 15351
rect 25136 15308 25188 15317
rect 25872 15351 25924 15360
rect 25872 15317 25881 15351
rect 25881 15317 25915 15351
rect 25915 15317 25924 15351
rect 25872 15308 25924 15317
rect 26240 15351 26292 15360
rect 26240 15317 26249 15351
rect 26249 15317 26283 15351
rect 26283 15317 26292 15351
rect 26240 15308 26292 15317
rect 26792 15308 26844 15360
rect 27160 15351 27212 15360
rect 27160 15317 27169 15351
rect 27169 15317 27203 15351
rect 27203 15317 27212 15351
rect 27160 15308 27212 15317
rect 29000 15351 29052 15360
rect 29000 15317 29009 15351
rect 29009 15317 29043 15351
rect 29043 15317 29052 15351
rect 29000 15308 29052 15317
rect 31024 15308 31076 15360
rect 32312 15308 32364 15360
rect 32680 15308 32732 15360
rect 33324 15308 33376 15360
rect 33692 15308 33744 15360
rect 33876 15351 33928 15360
rect 33876 15317 33885 15351
rect 33885 15317 33919 15351
rect 33919 15317 33928 15351
rect 33876 15308 33928 15317
rect 36452 15308 36504 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 9680 15147 9732 15156
rect 9680 15113 9689 15147
rect 9689 15113 9723 15147
rect 9723 15113 9732 15147
rect 9680 15104 9732 15113
rect 9772 15147 9824 15156
rect 9772 15113 9781 15147
rect 9781 15113 9815 15147
rect 9815 15113 9824 15147
rect 9772 15104 9824 15113
rect 11336 15104 11388 15156
rect 11796 15104 11848 15156
rect 10876 15079 10928 15088
rect 10876 15045 10885 15079
rect 10885 15045 10919 15079
rect 10919 15045 10928 15079
rect 10876 15036 10928 15045
rect 11060 15079 11112 15088
rect 11060 15045 11069 15079
rect 11069 15045 11103 15079
rect 11103 15045 11112 15079
rect 11060 15036 11112 15045
rect 11152 15036 11204 15088
rect 19340 15104 19392 15156
rect 19432 15104 19484 15156
rect 14832 15079 14884 15088
rect 14832 15045 14841 15079
rect 14841 15045 14875 15079
rect 14875 15045 14884 15079
rect 14832 15036 14884 15045
rect 15660 15036 15712 15088
rect 16120 15036 16172 15088
rect 21548 15104 21600 15156
rect 22836 15104 22888 15156
rect 23756 15104 23808 15156
rect 24676 15104 24728 15156
rect 20812 15036 20864 15088
rect 21640 15036 21692 15088
rect 25872 15036 25924 15088
rect 940 14968 992 15020
rect 4160 14968 4212 15020
rect 12256 15011 12308 15020
rect 12256 14977 12265 15011
rect 12265 14977 12299 15011
rect 12299 14977 12308 15011
rect 12256 14968 12308 14977
rect 13728 14968 13780 15020
rect 15108 15011 15160 15020
rect 15108 14977 15117 15011
rect 15117 14977 15151 15011
rect 15151 14977 15160 15011
rect 15108 14968 15160 14977
rect 15292 14968 15344 15020
rect 17500 14968 17552 15020
rect 18512 14968 18564 15020
rect 9772 14900 9824 14952
rect 12348 14943 12400 14952
rect 12348 14909 12357 14943
rect 12357 14909 12391 14943
rect 12391 14909 12400 14943
rect 12348 14900 12400 14909
rect 11060 14832 11112 14884
rect 10692 14764 10744 14816
rect 12072 14832 12124 14884
rect 13820 14900 13872 14952
rect 14188 14900 14240 14952
rect 14280 14900 14332 14952
rect 15384 14900 15436 14952
rect 17316 14943 17368 14952
rect 17316 14909 17325 14943
rect 17325 14909 17359 14943
rect 17359 14909 17368 14943
rect 17316 14900 17368 14909
rect 17408 14943 17460 14952
rect 17408 14909 17417 14943
rect 17417 14909 17451 14943
rect 17451 14909 17460 14943
rect 17408 14900 17460 14909
rect 18052 14943 18104 14952
rect 18052 14909 18061 14943
rect 18061 14909 18095 14943
rect 18095 14909 18104 14943
rect 20904 14968 20956 15020
rect 18052 14900 18104 14909
rect 20168 14943 20220 14952
rect 20168 14909 20177 14943
rect 20177 14909 20211 14943
rect 20211 14909 20220 14943
rect 20168 14900 20220 14909
rect 20536 14900 20588 14952
rect 21456 14968 21508 15020
rect 23296 15011 23348 15020
rect 23296 14977 23305 15011
rect 23305 14977 23339 15011
rect 23339 14977 23348 15011
rect 23296 14968 23348 14977
rect 25044 14968 25096 15020
rect 25136 14968 25188 15020
rect 25412 14968 25464 15020
rect 25688 14968 25740 15020
rect 29644 15104 29696 15156
rect 31300 15104 31352 15156
rect 27068 15079 27120 15088
rect 27068 15045 27077 15079
rect 27077 15045 27111 15079
rect 27111 15045 27120 15079
rect 27068 15036 27120 15045
rect 27896 15036 27948 15088
rect 28540 15036 28592 15088
rect 29276 15036 29328 15088
rect 29552 15036 29604 15088
rect 27252 15011 27304 15020
rect 27252 14977 27261 15011
rect 27261 14977 27295 15011
rect 27295 14977 27304 15011
rect 27252 14968 27304 14977
rect 27804 14968 27856 15020
rect 21364 14900 21416 14952
rect 23572 14943 23624 14952
rect 23572 14909 23581 14943
rect 23581 14909 23615 14943
rect 23615 14909 23624 14943
rect 23572 14900 23624 14909
rect 24216 14900 24268 14952
rect 24768 14900 24820 14952
rect 27344 14900 27396 14952
rect 30196 14968 30248 15020
rect 30564 15011 30616 15020
rect 30564 14977 30573 15011
rect 30573 14977 30607 15011
rect 30607 14977 30616 15011
rect 30564 14968 30616 14977
rect 29828 14900 29880 14952
rect 30012 14900 30064 14952
rect 30656 14943 30708 14952
rect 30656 14909 30665 14943
rect 30665 14909 30699 14943
rect 30699 14909 30708 14943
rect 30656 14900 30708 14909
rect 30932 15036 30984 15088
rect 33876 15147 33928 15156
rect 33876 15113 33885 15147
rect 33885 15113 33919 15147
rect 33919 15113 33928 15147
rect 33876 15104 33928 15113
rect 37004 15104 37056 15156
rect 37648 15104 37700 15156
rect 40132 15147 40184 15156
rect 40132 15113 40141 15147
rect 40141 15113 40175 15147
rect 40175 15113 40184 15147
rect 40132 15104 40184 15113
rect 35992 15036 36044 15088
rect 36268 15079 36320 15088
rect 36268 15045 36277 15079
rect 36277 15045 36311 15079
rect 36311 15045 36320 15079
rect 36268 15036 36320 15045
rect 37740 15079 37792 15088
rect 37740 15045 37749 15079
rect 37749 15045 37783 15079
rect 37783 15045 37792 15079
rect 37740 15036 37792 15045
rect 38752 15036 38804 15088
rect 48412 15036 48464 15088
rect 31760 14968 31812 15020
rect 35900 14968 35952 15020
rect 31852 14943 31904 14952
rect 31852 14909 31861 14943
rect 31861 14909 31895 14943
rect 31895 14909 31904 14943
rect 31852 14900 31904 14909
rect 32312 14900 32364 14952
rect 17960 14832 18012 14884
rect 12808 14764 12860 14816
rect 14280 14764 14332 14816
rect 14464 14764 14516 14816
rect 15936 14764 15988 14816
rect 18604 14764 18656 14816
rect 25044 14764 25096 14816
rect 25688 14764 25740 14816
rect 27712 14832 27764 14884
rect 33784 14943 33836 14952
rect 33784 14909 33793 14943
rect 33793 14909 33827 14943
rect 33827 14909 33836 14943
rect 33784 14900 33836 14909
rect 34888 14943 34940 14952
rect 34888 14909 34897 14943
rect 34897 14909 34931 14943
rect 34931 14909 34940 14943
rect 34888 14900 34940 14909
rect 37372 14968 37424 15020
rect 40868 15011 40920 15020
rect 40868 14977 40877 15011
rect 40877 14977 40911 15011
rect 40911 14977 40920 15011
rect 40868 14968 40920 14977
rect 49332 15011 49384 15020
rect 49332 14977 49341 15011
rect 49341 14977 49375 15011
rect 49375 14977 49384 15011
rect 49332 14968 49384 14977
rect 36084 14943 36136 14952
rect 36084 14909 36093 14943
rect 36093 14909 36127 14943
rect 36127 14909 36136 14943
rect 36084 14900 36136 14909
rect 36268 14900 36320 14952
rect 37096 14900 37148 14952
rect 30196 14807 30248 14816
rect 30196 14773 30205 14807
rect 30205 14773 30239 14807
rect 30239 14773 30248 14807
rect 30196 14764 30248 14773
rect 33968 14832 34020 14884
rect 36544 14832 36596 14884
rect 33324 14764 33376 14816
rect 33508 14764 33560 14816
rect 37464 14764 37516 14816
rect 39672 14875 39724 14884
rect 39672 14841 39681 14875
rect 39681 14841 39715 14875
rect 39715 14841 39724 14875
rect 39672 14832 39724 14841
rect 39764 14832 39816 14884
rect 38752 14764 38804 14816
rect 45652 14764 45704 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 11244 14560 11296 14612
rect 12624 14560 12676 14612
rect 14004 14560 14056 14612
rect 14648 14560 14700 14612
rect 16764 14560 16816 14612
rect 17408 14560 17460 14612
rect 18420 14560 18472 14612
rect 18512 14560 18564 14612
rect 10232 14535 10284 14544
rect 10232 14501 10241 14535
rect 10241 14501 10275 14535
rect 10275 14501 10284 14535
rect 10232 14492 10284 14501
rect 940 14424 992 14476
rect 10416 14399 10468 14408
rect 10416 14365 10425 14399
rect 10425 14365 10459 14399
rect 10459 14365 10468 14399
rect 10416 14356 10468 14365
rect 9956 14288 10008 14340
rect 10692 14424 10744 14476
rect 12256 14424 12308 14476
rect 13268 14424 13320 14476
rect 13636 14467 13688 14476
rect 13636 14433 13645 14467
rect 13645 14433 13679 14467
rect 13679 14433 13688 14467
rect 13636 14424 13688 14433
rect 14832 14424 14884 14476
rect 13820 14356 13872 14408
rect 20720 14535 20772 14544
rect 20720 14501 20729 14535
rect 20729 14501 20763 14535
rect 20763 14501 20772 14535
rect 20720 14492 20772 14501
rect 22744 14492 22796 14544
rect 24676 14535 24728 14544
rect 24676 14501 24685 14535
rect 24685 14501 24719 14535
rect 24719 14501 24728 14535
rect 24676 14492 24728 14501
rect 25504 14560 25556 14612
rect 26332 14560 26384 14612
rect 26516 14560 26568 14612
rect 30012 14560 30064 14612
rect 33784 14560 33836 14612
rect 36636 14603 36688 14612
rect 36636 14569 36645 14603
rect 36645 14569 36679 14603
rect 36679 14569 36688 14603
rect 36636 14560 36688 14569
rect 37096 14603 37148 14612
rect 37096 14569 37105 14603
rect 37105 14569 37139 14603
rect 37139 14569 37148 14603
rect 37096 14560 37148 14569
rect 38568 14560 38620 14612
rect 27436 14492 27488 14544
rect 15384 14424 15436 14476
rect 17408 14424 17460 14476
rect 19340 14424 19392 14476
rect 21364 14424 21416 14476
rect 21732 14424 21784 14476
rect 17224 14356 17276 14408
rect 17684 14356 17736 14408
rect 18604 14399 18656 14408
rect 18604 14365 18613 14399
rect 18613 14365 18647 14399
rect 18647 14365 18656 14399
rect 18604 14356 18656 14365
rect 19892 14399 19944 14408
rect 19892 14365 19901 14399
rect 19901 14365 19935 14399
rect 19935 14365 19944 14399
rect 19892 14356 19944 14365
rect 20444 14356 20496 14408
rect 22652 14356 22704 14408
rect 23020 14356 23072 14408
rect 27344 14399 27396 14408
rect 27344 14365 27353 14399
rect 27353 14365 27387 14399
rect 27387 14365 27396 14399
rect 27344 14356 27396 14365
rect 27896 14467 27948 14476
rect 27896 14433 27905 14467
rect 27905 14433 27939 14467
rect 27939 14433 27948 14467
rect 27896 14424 27948 14433
rect 29368 14424 29420 14476
rect 29736 14424 29788 14476
rect 30012 14467 30064 14476
rect 30012 14433 30021 14467
rect 30021 14433 30055 14467
rect 30055 14433 30064 14467
rect 30012 14424 30064 14433
rect 28632 14356 28684 14408
rect 31668 14535 31720 14544
rect 31668 14501 31677 14535
rect 31677 14501 31711 14535
rect 31711 14501 31720 14535
rect 31668 14492 31720 14501
rect 32496 14492 32548 14544
rect 30748 14424 30800 14476
rect 31576 14424 31628 14476
rect 11244 14331 11296 14340
rect 11244 14297 11253 14331
rect 11253 14297 11287 14331
rect 11287 14297 11296 14331
rect 11244 14288 11296 14297
rect 12808 14288 12860 14340
rect 10508 14220 10560 14272
rect 12716 14220 12768 14272
rect 14004 14220 14056 14272
rect 14188 14220 14240 14272
rect 16948 14288 17000 14340
rect 17316 14288 17368 14340
rect 19432 14288 19484 14340
rect 17500 14220 17552 14272
rect 17960 14220 18012 14272
rect 18052 14220 18104 14272
rect 18420 14220 18472 14272
rect 18972 14220 19024 14272
rect 19524 14263 19576 14272
rect 19524 14229 19533 14263
rect 19533 14229 19567 14263
rect 19567 14229 19576 14263
rect 19524 14220 19576 14229
rect 19800 14220 19852 14272
rect 20536 14263 20588 14272
rect 20536 14229 20545 14263
rect 20545 14229 20579 14263
rect 20579 14229 20588 14263
rect 20536 14220 20588 14229
rect 21272 14288 21324 14340
rect 24492 14288 24544 14340
rect 21732 14220 21784 14272
rect 23848 14263 23900 14272
rect 23848 14229 23857 14263
rect 23857 14229 23891 14263
rect 23891 14229 23900 14263
rect 23848 14220 23900 14229
rect 24400 14263 24452 14272
rect 24400 14229 24409 14263
rect 24409 14229 24443 14263
rect 24443 14229 24452 14263
rect 24400 14220 24452 14229
rect 25136 14263 25188 14272
rect 25136 14229 25145 14263
rect 25145 14229 25179 14263
rect 25179 14229 25188 14263
rect 25136 14220 25188 14229
rect 25780 14288 25832 14340
rect 27068 14331 27120 14340
rect 27068 14297 27077 14331
rect 27077 14297 27111 14331
rect 27111 14297 27120 14331
rect 27068 14288 27120 14297
rect 27712 14220 27764 14272
rect 28448 14220 28500 14272
rect 31852 14356 31904 14408
rect 34796 14424 34848 14476
rect 36360 14492 36412 14544
rect 37096 14424 37148 14476
rect 37372 14424 37424 14476
rect 32956 14356 33008 14408
rect 39948 14603 40000 14612
rect 39948 14569 39957 14603
rect 39957 14569 39991 14603
rect 39991 14569 40000 14603
rect 39948 14560 40000 14569
rect 49056 14399 49108 14408
rect 49056 14365 49065 14399
rect 49065 14365 49099 14399
rect 49099 14365 49108 14399
rect 49056 14356 49108 14365
rect 49240 14399 49292 14408
rect 49240 14365 49249 14399
rect 49249 14365 49283 14399
rect 49283 14365 49292 14399
rect 49240 14356 49292 14365
rect 33508 14288 33560 14340
rect 34612 14288 34664 14340
rect 35164 14331 35216 14340
rect 35164 14297 35173 14331
rect 35173 14297 35207 14331
rect 35207 14297 35216 14331
rect 35164 14288 35216 14297
rect 35624 14288 35676 14340
rect 36820 14288 36872 14340
rect 29000 14263 29052 14272
rect 29000 14229 29009 14263
rect 29009 14229 29043 14263
rect 29043 14229 29052 14263
rect 29000 14220 29052 14229
rect 29644 14220 29696 14272
rect 30012 14220 30064 14272
rect 30288 14220 30340 14272
rect 31024 14220 31076 14272
rect 32772 14220 32824 14272
rect 33416 14220 33468 14272
rect 34888 14220 34940 14272
rect 37556 14220 37608 14272
rect 37648 14220 37700 14272
rect 39488 14263 39540 14272
rect 39488 14229 39497 14263
rect 39497 14229 39531 14263
rect 39531 14229 39540 14263
rect 39488 14220 39540 14229
rect 48320 14220 48372 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 9864 14016 9916 14068
rect 9956 14059 10008 14068
rect 9956 14025 9965 14059
rect 9965 14025 9999 14059
rect 9999 14025 10008 14059
rect 9956 14016 10008 14025
rect 10416 14059 10468 14068
rect 10416 14025 10425 14059
rect 10425 14025 10459 14059
rect 10459 14025 10468 14059
rect 10416 14016 10468 14025
rect 11888 14016 11940 14068
rect 12900 14016 12952 14068
rect 14188 14016 14240 14068
rect 14280 14016 14332 14068
rect 15936 14059 15988 14068
rect 15936 14025 15945 14059
rect 15945 14025 15979 14059
rect 15979 14025 15988 14059
rect 15936 14016 15988 14025
rect 16580 14016 16632 14068
rect 17500 14059 17552 14068
rect 17500 14025 17509 14059
rect 17509 14025 17543 14059
rect 17543 14025 17552 14059
rect 17500 14016 17552 14025
rect 17592 14059 17644 14068
rect 17592 14025 17601 14059
rect 17601 14025 17635 14059
rect 17635 14025 17644 14059
rect 17592 14016 17644 14025
rect 18328 14059 18380 14068
rect 18328 14025 18337 14059
rect 18337 14025 18371 14059
rect 18371 14025 18380 14059
rect 18328 14016 18380 14025
rect 18788 14016 18840 14068
rect 19892 14016 19944 14068
rect 21272 14016 21324 14068
rect 21548 14016 21600 14068
rect 24492 14016 24544 14068
rect 25320 14016 25372 14068
rect 25504 14016 25556 14068
rect 1032 13948 1084 14000
rect 10508 13948 10560 14000
rect 11244 13948 11296 14000
rect 13268 13991 13320 14000
rect 13268 13957 13277 13991
rect 13277 13957 13311 13991
rect 13311 13957 13320 13991
rect 13268 13948 13320 13957
rect 13728 13948 13780 14000
rect 15016 13991 15068 14000
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 12256 13812 12308 13864
rect 12348 13744 12400 13796
rect 10784 13676 10836 13728
rect 13728 13812 13780 13864
rect 14464 13812 14516 13864
rect 15016 13957 15025 13991
rect 15025 13957 15059 13991
rect 15059 13957 15068 13991
rect 15016 13948 15068 13957
rect 15292 13991 15344 14000
rect 15292 13957 15301 13991
rect 15301 13957 15335 13991
rect 15335 13957 15344 13991
rect 15292 13948 15344 13957
rect 19524 13948 19576 14000
rect 20720 13948 20772 14000
rect 23020 13948 23072 14000
rect 25780 13948 25832 14000
rect 27620 14059 27672 14068
rect 27620 14025 27629 14059
rect 27629 14025 27663 14059
rect 27663 14025 27672 14059
rect 27620 14016 27672 14025
rect 27068 13948 27120 14000
rect 27528 13948 27580 14000
rect 30012 14016 30064 14068
rect 31116 14016 31168 14068
rect 41328 14016 41380 14068
rect 47032 14016 47084 14068
rect 48412 14059 48464 14068
rect 48412 14025 48421 14059
rect 48421 14025 48455 14059
rect 48455 14025 48464 14059
rect 48412 14016 48464 14025
rect 49148 14059 49200 14068
rect 49148 14025 49157 14059
rect 49157 14025 49191 14059
rect 49191 14025 49200 14059
rect 49148 14016 49200 14025
rect 31208 13948 31260 14000
rect 33692 13948 33744 14000
rect 35164 13948 35216 14000
rect 16488 13880 16540 13932
rect 17040 13880 17092 13932
rect 17592 13880 17644 13932
rect 19432 13880 19484 13932
rect 16212 13855 16264 13864
rect 16212 13821 16221 13855
rect 16221 13821 16255 13855
rect 16255 13821 16264 13855
rect 16212 13812 16264 13821
rect 13636 13676 13688 13728
rect 14648 13676 14700 13728
rect 15292 13744 15344 13796
rect 17132 13744 17184 13796
rect 18880 13855 18932 13864
rect 18880 13821 18889 13855
rect 18889 13821 18923 13855
rect 18923 13821 18932 13855
rect 18880 13812 18932 13821
rect 18972 13812 19024 13864
rect 20720 13812 20772 13864
rect 22008 13855 22060 13864
rect 17960 13744 18012 13796
rect 21088 13744 21140 13796
rect 19800 13676 19852 13728
rect 19984 13719 20036 13728
rect 19984 13685 20014 13719
rect 20014 13685 20036 13719
rect 22008 13821 22017 13855
rect 22017 13821 22051 13855
rect 22051 13821 22060 13855
rect 22008 13812 22060 13821
rect 24308 13880 24360 13932
rect 28908 13923 28960 13932
rect 28908 13889 28917 13923
rect 28917 13889 28951 13923
rect 28951 13889 28960 13923
rect 28908 13880 28960 13889
rect 29276 13880 29328 13932
rect 31116 13923 31168 13932
rect 31116 13889 31125 13923
rect 31125 13889 31159 13923
rect 31159 13889 31168 13923
rect 31116 13880 31168 13889
rect 31944 13880 31996 13932
rect 32496 13880 32548 13932
rect 34152 13880 34204 13932
rect 21916 13744 21968 13796
rect 23940 13812 23992 13864
rect 27344 13812 27396 13864
rect 30288 13812 30340 13864
rect 32312 13855 32364 13864
rect 24584 13744 24636 13796
rect 29736 13744 29788 13796
rect 32312 13821 32321 13855
rect 32321 13821 32355 13855
rect 32355 13821 32364 13855
rect 32312 13812 32364 13821
rect 34060 13855 34112 13864
rect 34060 13821 34069 13855
rect 34069 13821 34103 13855
rect 34103 13821 34112 13855
rect 34060 13812 34112 13821
rect 34704 13744 34756 13796
rect 36084 13880 36136 13932
rect 36728 13948 36780 14000
rect 38660 13948 38712 14000
rect 39488 13948 39540 14000
rect 49240 13991 49292 14000
rect 49240 13957 49249 13991
rect 49249 13957 49283 13991
rect 49283 13957 49292 13991
rect 49240 13948 49292 13957
rect 45652 13923 45704 13932
rect 45652 13889 45661 13923
rect 45661 13889 45695 13923
rect 45695 13889 45704 13923
rect 45652 13880 45704 13889
rect 48228 13880 48280 13932
rect 35992 13855 36044 13864
rect 35992 13821 36001 13855
rect 36001 13821 36035 13855
rect 36035 13821 36044 13855
rect 35992 13812 36044 13821
rect 36636 13744 36688 13796
rect 46296 13812 46348 13864
rect 38200 13744 38252 13796
rect 19984 13676 20036 13685
rect 22836 13676 22888 13728
rect 26332 13676 26384 13728
rect 30840 13676 30892 13728
rect 36360 13676 36412 13728
rect 36728 13719 36780 13728
rect 36728 13685 36737 13719
rect 36737 13685 36771 13719
rect 36771 13685 36780 13719
rect 36728 13676 36780 13685
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 1768 13379 1820 13388
rect 1768 13345 1777 13379
rect 1777 13345 1811 13379
rect 1811 13345 1820 13379
rect 1768 13336 1820 13345
rect 10508 13447 10560 13456
rect 10508 13413 10517 13447
rect 10517 13413 10551 13447
rect 10551 13413 10560 13447
rect 12256 13472 12308 13524
rect 12992 13472 13044 13524
rect 13728 13515 13780 13524
rect 13728 13481 13737 13515
rect 13737 13481 13771 13515
rect 13771 13481 13780 13515
rect 13728 13472 13780 13481
rect 14188 13472 14240 13524
rect 10508 13404 10560 13413
rect 10784 13379 10836 13388
rect 10784 13345 10793 13379
rect 10793 13345 10827 13379
rect 10827 13345 10836 13379
rect 10784 13336 10836 13345
rect 15016 13472 15068 13524
rect 15200 13404 15252 13456
rect 11152 13336 11204 13388
rect 12900 13336 12952 13388
rect 13820 13336 13872 13388
rect 14832 13336 14884 13388
rect 17960 13472 18012 13524
rect 18420 13472 18472 13524
rect 20260 13472 20312 13524
rect 20904 13515 20956 13524
rect 20904 13481 20913 13515
rect 20913 13481 20947 13515
rect 20947 13481 20956 13515
rect 20904 13472 20956 13481
rect 22192 13472 22244 13524
rect 17868 13404 17920 13456
rect 22560 13404 22612 13456
rect 15476 13379 15528 13388
rect 15476 13345 15485 13379
rect 15485 13345 15519 13379
rect 15519 13345 15528 13379
rect 15476 13336 15528 13345
rect 15752 13336 15804 13388
rect 18972 13336 19024 13388
rect 19984 13336 20036 13388
rect 21364 13336 21416 13388
rect 22744 13472 22796 13524
rect 23664 13472 23716 13524
rect 25596 13515 25648 13524
rect 25596 13481 25605 13515
rect 25605 13481 25639 13515
rect 25639 13481 25648 13515
rect 25596 13472 25648 13481
rect 25780 13472 25832 13524
rect 27436 13515 27488 13524
rect 27436 13481 27445 13515
rect 27445 13481 27479 13515
rect 27479 13481 27488 13515
rect 27436 13472 27488 13481
rect 27804 13515 27856 13524
rect 27804 13481 27813 13515
rect 27813 13481 27847 13515
rect 27847 13481 27856 13515
rect 27804 13472 27856 13481
rect 28356 13472 28408 13524
rect 28908 13472 28960 13524
rect 33784 13472 33836 13524
rect 35716 13472 35768 13524
rect 38200 13515 38252 13524
rect 38200 13481 38209 13515
rect 38209 13481 38243 13515
rect 38243 13481 38252 13515
rect 38200 13472 38252 13481
rect 38660 13472 38712 13524
rect 38844 13472 38896 13524
rect 24492 13404 24544 13456
rect 22836 13336 22888 13388
rect 24400 13336 24452 13388
rect 27068 13336 27120 13388
rect 29920 13404 29972 13456
rect 30380 13404 30432 13456
rect 29828 13379 29880 13388
rect 29828 13345 29837 13379
rect 29837 13345 29871 13379
rect 29871 13345 29880 13379
rect 29828 13336 29880 13345
rect 30472 13336 30524 13388
rect 31392 13336 31444 13388
rect 33876 13379 33928 13388
rect 33876 13345 33885 13379
rect 33885 13345 33919 13379
rect 33919 13345 33928 13379
rect 33876 13336 33928 13345
rect 14556 13268 14608 13320
rect 18328 13268 18380 13320
rect 9036 13200 9088 13252
rect 10968 13132 11020 13184
rect 11152 13200 11204 13252
rect 12992 13200 13044 13252
rect 14924 13200 14976 13252
rect 16212 13200 16264 13252
rect 16304 13200 16356 13252
rect 17132 13200 17184 13252
rect 21456 13200 21508 13252
rect 21640 13200 21692 13252
rect 22836 13200 22888 13252
rect 13820 13132 13872 13184
rect 14096 13132 14148 13184
rect 15108 13132 15160 13184
rect 15568 13175 15620 13184
rect 15568 13141 15577 13175
rect 15577 13141 15611 13175
rect 15611 13141 15620 13175
rect 15568 13132 15620 13141
rect 15936 13175 15988 13184
rect 15936 13141 15945 13175
rect 15945 13141 15979 13175
rect 15979 13141 15988 13175
rect 15936 13132 15988 13141
rect 16764 13132 16816 13184
rect 18512 13132 18564 13184
rect 19340 13175 19392 13184
rect 19340 13141 19349 13175
rect 19349 13141 19383 13175
rect 19383 13141 19392 13175
rect 19340 13132 19392 13141
rect 19984 13175 20036 13184
rect 19984 13141 19993 13175
rect 19993 13141 20027 13175
rect 20027 13141 20036 13175
rect 19984 13132 20036 13141
rect 21548 13132 21600 13184
rect 21824 13132 21876 13184
rect 24032 13200 24084 13252
rect 23664 13175 23716 13184
rect 23664 13141 23673 13175
rect 23673 13141 23707 13175
rect 23707 13141 23716 13175
rect 23664 13132 23716 13141
rect 23848 13132 23900 13184
rect 24400 13132 24452 13184
rect 25136 13268 25188 13320
rect 29000 13268 29052 13320
rect 30196 13268 30248 13320
rect 31208 13268 31260 13320
rect 34060 13268 34112 13320
rect 24860 13200 24912 13252
rect 25780 13200 25832 13252
rect 26056 13243 26108 13252
rect 26056 13209 26065 13243
rect 26065 13209 26099 13243
rect 26099 13209 26108 13243
rect 26056 13200 26108 13209
rect 28632 13200 28684 13252
rect 26516 13132 26568 13184
rect 28724 13175 28776 13184
rect 28724 13141 28733 13175
rect 28733 13141 28767 13175
rect 28767 13141 28776 13175
rect 28724 13132 28776 13141
rect 33600 13200 33652 13252
rect 33692 13243 33744 13252
rect 33692 13209 33701 13243
rect 33701 13209 33735 13243
rect 33735 13209 33744 13243
rect 39212 13336 39264 13388
rect 34888 13268 34940 13320
rect 33692 13200 33744 13209
rect 35164 13243 35216 13252
rect 35164 13209 35173 13243
rect 35173 13209 35207 13243
rect 35207 13209 35216 13243
rect 35164 13200 35216 13209
rect 36360 13200 36412 13252
rect 31668 13132 31720 13184
rect 34428 13132 34480 13184
rect 35624 13132 35676 13184
rect 41328 13311 41380 13320
rect 41328 13277 41337 13311
rect 41337 13277 41371 13311
rect 41371 13277 41380 13311
rect 41328 13268 41380 13277
rect 46296 13268 46348 13320
rect 49148 13311 49200 13320
rect 49148 13277 49157 13311
rect 49157 13277 49191 13311
rect 49191 13277 49200 13311
rect 49148 13268 49200 13277
rect 36636 13200 36688 13252
rect 38844 13200 38896 13252
rect 37464 13132 37516 13184
rect 37648 13132 37700 13184
rect 39580 13132 39632 13184
rect 45928 13132 45980 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 5448 12928 5500 12980
rect 10968 12971 11020 12980
rect 10968 12937 10977 12971
rect 10977 12937 11011 12971
rect 11011 12937 11020 12971
rect 10968 12928 11020 12937
rect 11152 12971 11204 12980
rect 11152 12937 11161 12971
rect 11161 12937 11195 12971
rect 11195 12937 11204 12971
rect 11152 12928 11204 12937
rect 11336 12928 11388 12980
rect 12440 12928 12492 12980
rect 13268 12928 13320 12980
rect 13636 12928 13688 12980
rect 1308 12860 1360 12912
rect 14464 12860 14516 12912
rect 1216 12792 1268 12844
rect 9496 12724 9548 12776
rect 11796 12767 11848 12776
rect 11796 12733 11805 12767
rect 11805 12733 11839 12767
rect 11839 12733 11848 12767
rect 11796 12724 11848 12733
rect 13912 12724 13964 12776
rect 14556 12767 14608 12776
rect 14556 12733 14565 12767
rect 14565 12733 14599 12767
rect 14599 12733 14608 12767
rect 14556 12724 14608 12733
rect 15292 12971 15344 12980
rect 15292 12937 15301 12971
rect 15301 12937 15335 12971
rect 15335 12937 15344 12971
rect 15292 12928 15344 12937
rect 18328 12928 18380 12980
rect 19064 12928 19116 12980
rect 22928 12971 22980 12980
rect 22928 12937 22937 12971
rect 22937 12937 22971 12971
rect 22971 12937 22980 12971
rect 22928 12928 22980 12937
rect 23388 12971 23440 12980
rect 23388 12937 23397 12971
rect 23397 12937 23431 12971
rect 23431 12937 23440 12971
rect 23388 12928 23440 12937
rect 24308 12928 24360 12980
rect 24584 12928 24636 12980
rect 16396 12860 16448 12912
rect 18972 12860 19024 12912
rect 15476 12724 15528 12776
rect 16304 12792 16356 12844
rect 16856 12792 16908 12844
rect 17776 12792 17828 12844
rect 18604 12792 18656 12844
rect 19064 12792 19116 12844
rect 19892 12860 19944 12912
rect 24860 12860 24912 12912
rect 25320 12903 25372 12912
rect 25320 12869 25329 12903
rect 25329 12869 25363 12903
rect 25363 12869 25372 12903
rect 25320 12860 25372 12869
rect 19524 12792 19576 12844
rect 21916 12792 21968 12844
rect 22192 12792 22244 12844
rect 23020 12835 23072 12844
rect 23020 12801 23029 12835
rect 23029 12801 23063 12835
rect 23063 12801 23072 12835
rect 23020 12792 23072 12801
rect 25780 12928 25832 12980
rect 26240 12971 26292 12980
rect 26240 12937 26249 12971
rect 26249 12937 26283 12971
rect 26283 12937 26292 12971
rect 26240 12928 26292 12937
rect 26516 12928 26568 12980
rect 27896 12928 27948 12980
rect 27436 12860 27488 12912
rect 29644 12903 29696 12912
rect 29644 12869 29653 12903
rect 29653 12869 29687 12903
rect 29687 12869 29696 12903
rect 29644 12860 29696 12869
rect 30196 12860 30248 12912
rect 31300 12860 31352 12912
rect 31852 12928 31904 12980
rect 32404 12928 32456 12980
rect 33508 12928 33560 12980
rect 33692 12928 33744 12980
rect 34060 12928 34112 12980
rect 26424 12835 26476 12844
rect 26424 12801 26433 12835
rect 26433 12801 26467 12835
rect 26467 12801 26476 12835
rect 27160 12835 27212 12844
rect 26424 12792 26476 12801
rect 27160 12801 27169 12835
rect 27169 12801 27203 12835
rect 27203 12801 27212 12835
rect 27160 12792 27212 12801
rect 30012 12835 30064 12844
rect 30012 12801 30021 12835
rect 30021 12801 30055 12835
rect 30055 12801 30064 12835
rect 30012 12792 30064 12801
rect 19708 12767 19760 12776
rect 19708 12733 19717 12767
rect 19717 12733 19751 12767
rect 19751 12733 19760 12767
rect 19708 12724 19760 12733
rect 20260 12724 20312 12776
rect 11244 12631 11296 12640
rect 11244 12597 11253 12631
rect 11253 12597 11287 12631
rect 11287 12597 11296 12631
rect 11244 12588 11296 12597
rect 12532 12588 12584 12640
rect 17316 12656 17368 12708
rect 17776 12656 17828 12708
rect 21272 12767 21324 12776
rect 21272 12733 21281 12767
rect 21281 12733 21315 12767
rect 21315 12733 21324 12767
rect 21272 12724 21324 12733
rect 21732 12724 21784 12776
rect 22744 12767 22796 12776
rect 22744 12733 22753 12767
rect 22753 12733 22787 12767
rect 22787 12733 22796 12767
rect 22744 12724 22796 12733
rect 23572 12724 23624 12776
rect 24952 12724 25004 12776
rect 28908 12767 28960 12776
rect 28908 12733 28917 12767
rect 28917 12733 28951 12767
rect 28951 12733 28960 12767
rect 28908 12724 28960 12733
rect 32680 12724 32732 12776
rect 16764 12631 16816 12640
rect 16764 12597 16773 12631
rect 16773 12597 16807 12631
rect 16807 12597 16816 12631
rect 16764 12588 16816 12597
rect 16856 12631 16908 12640
rect 16856 12597 16865 12631
rect 16865 12597 16899 12631
rect 16899 12597 16908 12631
rect 16856 12588 16908 12597
rect 17132 12588 17184 12640
rect 19340 12588 19392 12640
rect 21180 12588 21232 12640
rect 23848 12588 23900 12640
rect 25688 12588 25740 12640
rect 25964 12631 26016 12640
rect 25964 12597 25973 12631
rect 25973 12597 26007 12631
rect 26007 12597 26016 12631
rect 25964 12588 26016 12597
rect 27804 12588 27856 12640
rect 33876 12860 33928 12912
rect 35164 12928 35216 12980
rect 40316 12928 40368 12980
rect 34888 12860 34940 12912
rect 34060 12835 34112 12844
rect 34060 12801 34069 12835
rect 34069 12801 34103 12835
rect 34103 12801 34112 12835
rect 34060 12792 34112 12801
rect 34336 12792 34388 12844
rect 37004 12860 37056 12912
rect 37188 12860 37240 12912
rect 37648 12860 37700 12912
rect 33232 12724 33284 12776
rect 34796 12656 34848 12708
rect 35256 12724 35308 12776
rect 35624 12767 35676 12776
rect 35624 12733 35633 12767
rect 35633 12733 35667 12767
rect 35667 12733 35676 12767
rect 35624 12724 35676 12733
rect 37464 12835 37516 12844
rect 37464 12801 37473 12835
rect 37473 12801 37507 12835
rect 37507 12801 37516 12835
rect 37464 12792 37516 12801
rect 38844 12792 38896 12844
rect 40040 12835 40092 12844
rect 40040 12801 40049 12835
rect 40049 12801 40083 12835
rect 40083 12801 40092 12835
rect 40040 12792 40092 12801
rect 45928 12835 45980 12844
rect 45928 12801 45937 12835
rect 45937 12801 45971 12835
rect 45971 12801 45980 12835
rect 45928 12792 45980 12801
rect 47032 12792 47084 12844
rect 49148 12835 49200 12844
rect 49148 12801 49157 12835
rect 49157 12801 49191 12835
rect 49191 12801 49200 12835
rect 49148 12792 49200 12801
rect 38292 12724 38344 12776
rect 39304 12724 39356 12776
rect 37280 12656 37332 12708
rect 42708 12656 42760 12708
rect 33324 12588 33376 12640
rect 35624 12588 35676 12640
rect 39304 12588 39356 12640
rect 47952 12588 48004 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 11796 12384 11848 12436
rect 14096 12384 14148 12436
rect 14556 12384 14608 12436
rect 15292 12384 15344 12436
rect 16028 12384 16080 12436
rect 16304 12384 16356 12436
rect 13820 12316 13872 12368
rect 14740 12316 14792 12368
rect 1308 12248 1360 12300
rect 10784 12248 10836 12300
rect 15476 12248 15528 12300
rect 15752 12248 15804 12300
rect 5908 12180 5960 12232
rect 17408 12291 17460 12300
rect 17408 12257 17417 12291
rect 17417 12257 17451 12291
rect 17451 12257 17460 12291
rect 17408 12248 17460 12257
rect 19892 12248 19944 12300
rect 21180 12291 21232 12300
rect 21180 12257 21189 12291
rect 21189 12257 21223 12291
rect 21223 12257 21232 12291
rect 21180 12248 21232 12257
rect 22100 12316 22152 12368
rect 22560 12384 22612 12436
rect 23480 12316 23532 12368
rect 9772 12155 9824 12164
rect 9772 12121 9781 12155
rect 9781 12121 9815 12155
rect 9815 12121 9824 12155
rect 9772 12112 9824 12121
rect 10508 12112 10560 12164
rect 11060 12112 11112 12164
rect 13636 12112 13688 12164
rect 14464 12112 14516 12164
rect 15844 12155 15896 12164
rect 15844 12121 15853 12155
rect 15853 12121 15887 12155
rect 15887 12121 15896 12155
rect 15844 12112 15896 12121
rect 12256 12044 12308 12096
rect 13452 12044 13504 12096
rect 16764 12087 16816 12096
rect 16764 12053 16773 12087
rect 16773 12053 16807 12087
rect 16807 12053 16816 12087
rect 16764 12044 16816 12053
rect 17224 12087 17276 12096
rect 17224 12053 17233 12087
rect 17233 12053 17267 12087
rect 17267 12053 17276 12087
rect 17224 12044 17276 12053
rect 17592 12112 17644 12164
rect 18788 12112 18840 12164
rect 18880 12155 18932 12164
rect 18880 12121 18889 12155
rect 18889 12121 18923 12155
rect 18923 12121 18932 12155
rect 18880 12112 18932 12121
rect 19800 12223 19852 12232
rect 19800 12189 19809 12223
rect 19809 12189 19843 12223
rect 19843 12189 19852 12223
rect 19800 12180 19852 12189
rect 20536 12180 20588 12232
rect 20904 12180 20956 12232
rect 21456 12180 21508 12232
rect 22284 12291 22336 12300
rect 22284 12257 22293 12291
rect 22293 12257 22327 12291
rect 22327 12257 22336 12291
rect 22284 12248 22336 12257
rect 26700 12384 26752 12436
rect 27896 12384 27948 12436
rect 32036 12384 32088 12436
rect 34612 12384 34664 12436
rect 26332 12359 26384 12368
rect 26332 12325 26341 12359
rect 26341 12325 26375 12359
rect 26375 12325 26384 12359
rect 26332 12316 26384 12325
rect 26884 12316 26936 12368
rect 29460 12316 29512 12368
rect 34520 12316 34572 12368
rect 35624 12384 35676 12436
rect 36636 12427 36688 12436
rect 36636 12393 36645 12427
rect 36645 12393 36679 12427
rect 36679 12393 36688 12427
rect 36636 12384 36688 12393
rect 39212 12384 39264 12436
rect 39304 12427 39356 12436
rect 39304 12393 39313 12427
rect 39313 12393 39347 12427
rect 39347 12393 39356 12427
rect 39304 12384 39356 12393
rect 24400 12248 24452 12300
rect 24952 12248 25004 12300
rect 27160 12291 27212 12300
rect 27160 12257 27169 12291
rect 27169 12257 27203 12291
rect 27203 12257 27212 12291
rect 27160 12248 27212 12257
rect 27344 12248 27396 12300
rect 30012 12248 30064 12300
rect 31300 12248 31352 12300
rect 31760 12291 31812 12300
rect 31760 12257 31769 12291
rect 31769 12257 31803 12291
rect 31803 12257 31812 12291
rect 31760 12248 31812 12257
rect 33600 12248 33652 12300
rect 38384 12291 38436 12300
rect 38384 12257 38393 12291
rect 38393 12257 38427 12291
rect 38427 12257 38436 12291
rect 38384 12248 38436 12257
rect 38752 12248 38804 12300
rect 47124 12316 47176 12368
rect 22744 12180 22796 12232
rect 24584 12223 24636 12232
rect 24584 12189 24593 12223
rect 24593 12189 24627 12223
rect 24627 12189 24636 12223
rect 24584 12180 24636 12189
rect 26516 12180 26568 12232
rect 27528 12180 27580 12232
rect 27620 12180 27672 12232
rect 28816 12180 28868 12232
rect 31484 12180 31536 12232
rect 32128 12223 32180 12232
rect 32128 12189 32137 12223
rect 32137 12189 32171 12223
rect 32171 12189 32180 12223
rect 32128 12180 32180 12189
rect 34888 12223 34940 12232
rect 34888 12189 34897 12223
rect 34897 12189 34931 12223
rect 34931 12189 34940 12223
rect 34888 12180 34940 12189
rect 37096 12180 37148 12232
rect 49148 12291 49200 12300
rect 49148 12257 49157 12291
rect 49157 12257 49191 12291
rect 49191 12257 49200 12291
rect 49148 12248 49200 12257
rect 20168 12112 20220 12164
rect 19800 12044 19852 12096
rect 20076 12044 20128 12096
rect 22192 12044 22244 12096
rect 22560 12044 22612 12096
rect 25504 12044 25556 12096
rect 27436 12112 27488 12164
rect 29920 12112 29972 12164
rect 32312 12112 32364 12164
rect 32404 12155 32456 12164
rect 32404 12121 32413 12155
rect 32413 12121 32447 12155
rect 32447 12121 32456 12155
rect 32404 12112 32456 12121
rect 27344 12087 27396 12096
rect 27344 12053 27353 12087
rect 27353 12053 27387 12087
rect 27387 12053 27396 12087
rect 27344 12044 27396 12053
rect 27620 12044 27672 12096
rect 31392 12044 31444 12096
rect 31760 12044 31812 12096
rect 33324 12044 33376 12096
rect 34244 12044 34296 12096
rect 34336 12087 34388 12096
rect 34336 12053 34345 12087
rect 34345 12053 34379 12087
rect 34379 12053 34388 12087
rect 34336 12044 34388 12053
rect 35440 12044 35492 12096
rect 36176 12044 36228 12096
rect 36636 12044 36688 12096
rect 37372 12044 37424 12096
rect 38844 12112 38896 12164
rect 40132 12155 40184 12164
rect 40132 12121 40141 12155
rect 40141 12121 40175 12155
rect 40175 12121 40184 12155
rect 40132 12112 40184 12121
rect 38660 12087 38712 12096
rect 38660 12053 38669 12087
rect 38669 12053 38703 12087
rect 38703 12053 38712 12087
rect 38660 12044 38712 12053
rect 40960 12087 41012 12096
rect 40960 12053 40969 12087
rect 40969 12053 41003 12087
rect 41003 12053 41012 12087
rect 40960 12044 41012 12053
rect 47952 12223 48004 12232
rect 47952 12189 47961 12223
rect 47961 12189 47995 12223
rect 47995 12189 48004 12223
rect 47952 12180 48004 12189
rect 46112 12087 46164 12096
rect 46112 12053 46121 12087
rect 46121 12053 46155 12087
rect 46155 12053 46164 12087
rect 46112 12044 46164 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 10508 11840 10560 11892
rect 11336 11840 11388 11892
rect 13544 11840 13596 11892
rect 14280 11883 14332 11892
rect 14280 11849 14289 11883
rect 14289 11849 14323 11883
rect 14323 11849 14332 11883
rect 14280 11840 14332 11849
rect 2504 11772 2556 11824
rect 14740 11772 14792 11824
rect 19340 11840 19392 11892
rect 19984 11840 20036 11892
rect 20720 11883 20772 11892
rect 20720 11849 20729 11883
rect 20729 11849 20763 11883
rect 20763 11849 20772 11883
rect 20720 11840 20772 11849
rect 21180 11883 21232 11892
rect 21180 11849 21189 11883
rect 21189 11849 21223 11883
rect 21223 11849 21232 11883
rect 21180 11840 21232 11849
rect 21640 11840 21692 11892
rect 22560 11840 22612 11892
rect 1216 11704 1268 11756
rect 1308 11636 1360 11688
rect 12348 11704 12400 11756
rect 14372 11704 14424 11756
rect 14648 11704 14700 11756
rect 15108 11704 15160 11756
rect 15292 11704 15344 11756
rect 17040 11772 17092 11824
rect 11796 11636 11848 11688
rect 11520 11568 11572 11620
rect 13452 11636 13504 11688
rect 13636 11679 13688 11688
rect 13636 11645 13645 11679
rect 13645 11645 13679 11679
rect 13679 11645 13688 11679
rect 13636 11636 13688 11645
rect 13912 11636 13964 11688
rect 13268 11568 13320 11620
rect 13544 11568 13596 11620
rect 13820 11568 13872 11620
rect 15568 11679 15620 11688
rect 15568 11645 15577 11679
rect 15577 11645 15611 11679
rect 15611 11645 15620 11679
rect 15568 11636 15620 11645
rect 16028 11704 16080 11756
rect 16856 11704 16908 11756
rect 20076 11772 20128 11824
rect 21732 11772 21784 11824
rect 19524 11704 19576 11756
rect 20628 11704 20680 11756
rect 20904 11704 20956 11756
rect 22468 11704 22520 11756
rect 24492 11772 24544 11824
rect 27344 11840 27396 11892
rect 27436 11840 27488 11892
rect 28724 11840 28776 11892
rect 31852 11840 31904 11892
rect 32220 11840 32272 11892
rect 32772 11840 32824 11892
rect 33784 11840 33836 11892
rect 34244 11840 34296 11892
rect 25504 11704 25556 11756
rect 25780 11704 25832 11756
rect 27068 11704 27120 11756
rect 27344 11704 27396 11756
rect 16120 11636 16172 11688
rect 17592 11636 17644 11688
rect 4160 11500 4212 11552
rect 12348 11543 12400 11552
rect 12348 11509 12357 11543
rect 12357 11509 12391 11543
rect 12391 11509 12400 11543
rect 12348 11500 12400 11509
rect 13360 11543 13412 11552
rect 13360 11509 13369 11543
rect 13369 11509 13403 11543
rect 13403 11509 13412 11543
rect 13360 11500 13412 11509
rect 14832 11500 14884 11552
rect 15476 11500 15528 11552
rect 16212 11500 16264 11552
rect 16488 11500 16540 11552
rect 18788 11636 18840 11688
rect 20076 11636 20128 11688
rect 20996 11568 21048 11620
rect 21364 11679 21416 11688
rect 21364 11645 21373 11679
rect 21373 11645 21407 11679
rect 21407 11645 21416 11679
rect 21364 11636 21416 11645
rect 22284 11636 22336 11688
rect 26332 11636 26384 11688
rect 27252 11679 27304 11688
rect 27252 11645 27261 11679
rect 27261 11645 27295 11679
rect 27295 11645 27304 11679
rect 27252 11636 27304 11645
rect 27620 11772 27672 11824
rect 31392 11772 31444 11824
rect 31116 11747 31168 11756
rect 31116 11713 31125 11747
rect 31125 11713 31159 11747
rect 31159 11713 31168 11747
rect 31116 11704 31168 11713
rect 31576 11772 31628 11824
rect 31760 11815 31812 11824
rect 31760 11781 31769 11815
rect 31769 11781 31803 11815
rect 31803 11781 31812 11815
rect 31760 11772 31812 11781
rect 32312 11772 32364 11824
rect 34796 11840 34848 11892
rect 34980 11840 35032 11892
rect 36084 11840 36136 11892
rect 38660 11883 38712 11892
rect 38660 11849 38669 11883
rect 38669 11849 38703 11883
rect 38703 11849 38712 11883
rect 38660 11840 38712 11849
rect 40132 11840 40184 11892
rect 35900 11772 35952 11824
rect 37280 11772 37332 11824
rect 40960 11772 41012 11824
rect 49148 11815 49200 11824
rect 49148 11781 49157 11815
rect 49157 11781 49191 11815
rect 49191 11781 49200 11815
rect 49148 11772 49200 11781
rect 27712 11636 27764 11688
rect 27344 11568 27396 11620
rect 29552 11636 29604 11688
rect 29644 11636 29696 11688
rect 30840 11679 30892 11688
rect 30840 11645 30849 11679
rect 30849 11645 30883 11679
rect 30883 11645 30892 11679
rect 30840 11636 30892 11645
rect 31852 11636 31904 11688
rect 32588 11636 32640 11688
rect 30472 11568 30524 11620
rect 33508 11636 33560 11688
rect 36820 11704 36872 11756
rect 34888 11636 34940 11688
rect 33876 11568 33928 11620
rect 35072 11568 35124 11620
rect 21272 11500 21324 11552
rect 22468 11500 22520 11552
rect 24032 11500 24084 11552
rect 24400 11500 24452 11552
rect 34612 11543 34664 11552
rect 34612 11509 34621 11543
rect 34621 11509 34655 11543
rect 34655 11509 34664 11543
rect 34612 11500 34664 11509
rect 35440 11679 35492 11688
rect 35440 11645 35449 11679
rect 35449 11645 35483 11679
rect 35483 11645 35492 11679
rect 35440 11636 35492 11645
rect 36636 11636 36688 11688
rect 38384 11704 38436 11756
rect 39028 11747 39080 11756
rect 39028 11713 39037 11747
rect 39037 11713 39071 11747
rect 39071 11713 39080 11747
rect 39028 11704 39080 11713
rect 39212 11679 39264 11688
rect 39212 11645 39221 11679
rect 39221 11645 39255 11679
rect 39255 11645 39264 11679
rect 39212 11636 39264 11645
rect 38016 11568 38068 11620
rect 46112 11704 46164 11756
rect 35624 11500 35676 11552
rect 40224 11500 40276 11552
rect 46756 11568 46808 11620
rect 47768 11500 47820 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 1216 11296 1268 11348
rect 14004 11296 14056 11348
rect 14464 11228 14516 11280
rect 11060 11160 11112 11212
rect 11796 11160 11848 11212
rect 12900 11160 12952 11212
rect 15568 11296 15620 11348
rect 16672 11296 16724 11348
rect 15108 11228 15160 11280
rect 18880 11296 18932 11348
rect 22468 11296 22520 11348
rect 23296 11339 23348 11348
rect 23296 11305 23305 11339
rect 23305 11305 23339 11339
rect 23339 11305 23348 11339
rect 23296 11296 23348 11305
rect 17592 11228 17644 11280
rect 19524 11271 19576 11280
rect 19524 11237 19533 11271
rect 19533 11237 19567 11271
rect 19567 11237 19576 11271
rect 19524 11228 19576 11237
rect 14832 11203 14884 11212
rect 14832 11169 14841 11203
rect 14841 11169 14875 11203
rect 14875 11169 14884 11203
rect 14832 11160 14884 11169
rect 15384 11160 15436 11212
rect 1584 11135 1636 11144
rect 1584 11101 1593 11135
rect 1593 11101 1627 11135
rect 1627 11101 1636 11135
rect 1584 11092 1636 11101
rect 11336 11092 11388 11144
rect 13636 11092 13688 11144
rect 15936 11160 15988 11212
rect 16396 11092 16448 11144
rect 16488 11092 16540 11144
rect 12900 11024 12952 11076
rect 13452 11024 13504 11076
rect 15844 11024 15896 11076
rect 16580 11024 16632 11076
rect 14740 10999 14792 11008
rect 14740 10965 14749 10999
rect 14749 10965 14783 10999
rect 14783 10965 14792 10999
rect 14740 10956 14792 10965
rect 16304 10999 16356 11008
rect 16304 10965 16313 10999
rect 16313 10965 16347 10999
rect 16347 10965 16356 10999
rect 16304 10956 16356 10965
rect 18328 11092 18380 11144
rect 18604 11203 18656 11212
rect 18604 11169 18613 11203
rect 18613 11169 18647 11203
rect 18647 11169 18656 11203
rect 18604 11160 18656 11169
rect 18696 11160 18748 11212
rect 20076 11228 20128 11280
rect 20168 11160 20220 11212
rect 21272 11160 21324 11212
rect 23756 11160 23808 11212
rect 25228 11296 25280 11348
rect 26608 11296 26660 11348
rect 28816 11296 28868 11348
rect 28908 11228 28960 11280
rect 30472 11271 30524 11280
rect 30472 11237 30481 11271
rect 30481 11237 30515 11271
rect 30515 11237 30524 11271
rect 30472 11228 30524 11237
rect 24400 11160 24452 11212
rect 27160 11203 27212 11212
rect 27160 11169 27169 11203
rect 27169 11169 27203 11203
rect 27203 11169 27212 11203
rect 27160 11160 27212 11169
rect 32036 11160 32088 11212
rect 32588 11160 32640 11212
rect 19524 11092 19576 11144
rect 24584 11135 24636 11144
rect 24584 11101 24593 11135
rect 24593 11101 24627 11135
rect 24627 11101 24636 11135
rect 24584 11092 24636 11101
rect 26884 11135 26936 11144
rect 26884 11101 26893 11135
rect 26893 11101 26927 11135
rect 26927 11101 26936 11135
rect 26884 11092 26936 11101
rect 29644 11092 29696 11144
rect 34060 11296 34112 11348
rect 34612 11296 34664 11348
rect 35072 11296 35124 11348
rect 33508 11228 33560 11280
rect 35992 11228 36044 11280
rect 35900 11160 35952 11212
rect 33968 11092 34020 11144
rect 36912 11160 36964 11212
rect 37464 11160 37516 11212
rect 38844 11296 38896 11348
rect 39580 11339 39632 11348
rect 39580 11305 39589 11339
rect 39589 11305 39623 11339
rect 39623 11305 39632 11339
rect 39580 11296 39632 11305
rect 44088 11296 44140 11348
rect 17132 11067 17184 11076
rect 17132 11033 17141 11067
rect 17141 11033 17175 11067
rect 17175 11033 17184 11067
rect 17132 11024 17184 11033
rect 20536 11024 20588 11076
rect 21180 11024 21232 11076
rect 23940 11024 23992 11076
rect 25504 11024 25556 11076
rect 27620 11024 27672 11076
rect 18788 10956 18840 11008
rect 19984 10956 20036 11008
rect 22376 10956 22428 11008
rect 22652 10999 22704 11008
rect 22652 10965 22661 10999
rect 22661 10965 22695 10999
rect 22695 10965 22704 10999
rect 22652 10956 22704 10965
rect 24032 10956 24084 11008
rect 24676 10956 24728 11008
rect 29184 10999 29236 11008
rect 29184 10965 29193 10999
rect 29193 10965 29227 10999
rect 29227 10965 29236 10999
rect 29184 10956 29236 10965
rect 29368 10956 29420 11008
rect 30012 10999 30064 11008
rect 30012 10965 30021 10999
rect 30021 10965 30055 10999
rect 30055 10965 30064 10999
rect 30012 10956 30064 10965
rect 31392 11067 31444 11076
rect 31392 11033 31401 11067
rect 31401 11033 31435 11067
rect 31435 11033 31444 11067
rect 31392 11024 31444 11033
rect 31484 11024 31536 11076
rect 39580 11092 39632 11144
rect 40224 11092 40276 11144
rect 42708 11160 42760 11212
rect 49148 11203 49200 11212
rect 49148 11169 49157 11203
rect 49157 11169 49191 11203
rect 49191 11169 49200 11203
rect 49148 11160 49200 11169
rect 30748 10999 30800 11008
rect 30748 10965 30757 10999
rect 30757 10965 30791 10999
rect 30791 10965 30800 10999
rect 30748 10956 30800 10965
rect 30840 10956 30892 11008
rect 32036 10956 32088 11008
rect 32128 10956 32180 11008
rect 35900 11024 35952 11076
rect 38384 11024 38436 11076
rect 45744 11024 45796 11076
rect 46940 11024 46992 11076
rect 32956 10956 33008 11008
rect 38936 10956 38988 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 2504 10795 2556 10804
rect 2504 10761 2513 10795
rect 2513 10761 2547 10795
rect 2547 10761 2556 10795
rect 2504 10752 2556 10761
rect 11336 10752 11388 10804
rect 12808 10752 12860 10804
rect 14372 10795 14424 10804
rect 14372 10761 14381 10795
rect 14381 10761 14415 10795
rect 14415 10761 14424 10795
rect 14372 10752 14424 10761
rect 15568 10795 15620 10804
rect 15568 10761 15577 10795
rect 15577 10761 15611 10795
rect 15611 10761 15620 10795
rect 15568 10752 15620 10761
rect 19708 10752 19760 10804
rect 22652 10752 22704 10804
rect 22928 10752 22980 10804
rect 25504 10752 25556 10804
rect 26700 10752 26752 10804
rect 27712 10752 27764 10804
rect 1216 10684 1268 10736
rect 1308 10616 1360 10668
rect 14556 10684 14608 10736
rect 12256 10616 12308 10668
rect 15752 10684 15804 10736
rect 15844 10684 15896 10736
rect 13452 10548 13504 10600
rect 16764 10616 16816 10668
rect 20352 10684 20404 10736
rect 22284 10684 22336 10736
rect 23940 10684 23992 10736
rect 27620 10684 27672 10736
rect 18696 10659 18748 10668
rect 18696 10625 18705 10659
rect 18705 10625 18739 10659
rect 18739 10625 18748 10659
rect 18696 10616 18748 10625
rect 13820 10591 13872 10600
rect 13820 10557 13829 10591
rect 13829 10557 13863 10591
rect 13863 10557 13872 10591
rect 13820 10548 13872 10557
rect 14924 10591 14976 10600
rect 14924 10557 14933 10591
rect 14933 10557 14967 10591
rect 14967 10557 14976 10591
rect 14924 10548 14976 10557
rect 16028 10591 16080 10600
rect 16028 10557 16037 10591
rect 16037 10557 16071 10591
rect 16071 10557 16080 10591
rect 16028 10548 16080 10557
rect 12256 10455 12308 10464
rect 12256 10421 12265 10455
rect 12265 10421 12299 10455
rect 12299 10421 12308 10455
rect 12256 10412 12308 10421
rect 12716 10412 12768 10464
rect 13912 10480 13964 10532
rect 16672 10548 16724 10600
rect 17684 10591 17736 10600
rect 17684 10557 17693 10591
rect 17693 10557 17727 10591
rect 17727 10557 17736 10591
rect 17684 10548 17736 10557
rect 18052 10548 18104 10600
rect 16212 10480 16264 10532
rect 14740 10412 14792 10464
rect 16580 10412 16632 10464
rect 17040 10412 17092 10464
rect 18512 10480 18564 10532
rect 20444 10616 20496 10668
rect 19984 10548 20036 10600
rect 21088 10548 21140 10600
rect 21272 10480 21324 10532
rect 26056 10659 26108 10668
rect 26056 10625 26065 10659
rect 26065 10625 26099 10659
rect 26099 10625 26108 10659
rect 26056 10616 26108 10625
rect 27252 10616 27304 10668
rect 28816 10727 28868 10736
rect 28816 10693 28825 10727
rect 28825 10693 28859 10727
rect 28859 10693 28868 10727
rect 31116 10752 31168 10804
rect 32956 10752 33008 10804
rect 28816 10684 28868 10693
rect 32036 10684 32088 10736
rect 32772 10684 32824 10736
rect 29920 10616 29972 10668
rect 22008 10591 22060 10600
rect 22008 10557 22017 10591
rect 22017 10557 22051 10591
rect 22051 10557 22060 10591
rect 22008 10548 22060 10557
rect 24124 10548 24176 10600
rect 24676 10591 24728 10600
rect 24676 10557 24685 10591
rect 24685 10557 24719 10591
rect 24719 10557 24728 10591
rect 24676 10548 24728 10557
rect 26608 10548 26660 10600
rect 23756 10523 23808 10532
rect 23756 10489 23765 10523
rect 23765 10489 23799 10523
rect 23799 10489 23808 10523
rect 23756 10480 23808 10489
rect 24768 10480 24820 10532
rect 22100 10412 22152 10464
rect 22376 10412 22428 10464
rect 25780 10480 25832 10532
rect 26240 10523 26292 10532
rect 26240 10489 26249 10523
rect 26249 10489 26283 10523
rect 26283 10489 26292 10523
rect 26240 10480 26292 10489
rect 29276 10548 29328 10600
rect 29644 10548 29696 10600
rect 29828 10548 29880 10600
rect 30472 10591 30524 10600
rect 30472 10557 30481 10591
rect 30481 10557 30515 10591
rect 30515 10557 30524 10591
rect 30472 10548 30524 10557
rect 30656 10548 30708 10600
rect 33324 10659 33376 10668
rect 33324 10625 33333 10659
rect 33333 10625 33367 10659
rect 33367 10625 33376 10659
rect 33324 10616 33376 10625
rect 32404 10591 32456 10600
rect 32404 10557 32413 10591
rect 32413 10557 32447 10591
rect 32447 10557 32456 10591
rect 32404 10548 32456 10557
rect 36636 10684 36688 10736
rect 36820 10795 36872 10804
rect 36820 10761 36829 10795
rect 36829 10761 36863 10795
rect 36863 10761 36872 10795
rect 36820 10752 36872 10761
rect 36912 10752 36964 10804
rect 38844 10752 38896 10804
rect 37372 10684 37424 10736
rect 49240 10684 49292 10736
rect 34244 10616 34296 10668
rect 35624 10659 35676 10668
rect 35624 10625 35633 10659
rect 35633 10625 35667 10659
rect 35667 10625 35676 10659
rect 35624 10616 35676 10625
rect 36452 10659 36504 10668
rect 36452 10625 36461 10659
rect 36461 10625 36495 10659
rect 36495 10625 36504 10659
rect 36452 10616 36504 10625
rect 30196 10412 30248 10464
rect 30840 10412 30892 10464
rect 31760 10412 31812 10464
rect 31852 10412 31904 10464
rect 32036 10412 32088 10464
rect 34704 10548 34756 10600
rect 36360 10591 36412 10600
rect 36360 10557 36369 10591
rect 36369 10557 36403 10591
rect 36403 10557 36412 10591
rect 36360 10548 36412 10557
rect 46940 10616 46992 10668
rect 35624 10480 35676 10532
rect 46940 10480 46992 10532
rect 33876 10412 33928 10464
rect 34796 10412 34848 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 16028 10208 16080 10260
rect 14740 10140 14792 10192
rect 2136 10115 2188 10124
rect 2136 10081 2145 10115
rect 2145 10081 2179 10115
rect 2179 10081 2188 10115
rect 2136 10072 2188 10081
rect 2412 10047 2464 10056
rect 2412 10013 2421 10047
rect 2421 10013 2455 10047
rect 2455 10013 2464 10047
rect 2412 10004 2464 10013
rect 15108 10072 15160 10124
rect 15200 10072 15252 10124
rect 18052 10208 18104 10260
rect 18328 10208 18380 10260
rect 20444 10208 20496 10260
rect 16580 10183 16632 10192
rect 16580 10149 16589 10183
rect 16589 10149 16623 10183
rect 16623 10149 16632 10183
rect 16580 10140 16632 10149
rect 17500 10140 17552 10192
rect 17316 10072 17368 10124
rect 17868 10140 17920 10192
rect 18512 10140 18564 10192
rect 18420 10072 18472 10124
rect 19156 10140 19208 10192
rect 19432 10072 19484 10124
rect 19616 10072 19668 10124
rect 14464 10004 14516 10056
rect 14648 10004 14700 10056
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 16672 10004 16724 10056
rect 21640 10208 21692 10260
rect 22192 10208 22244 10260
rect 24032 10208 24084 10260
rect 24308 10208 24360 10260
rect 26700 10251 26752 10260
rect 26700 10217 26709 10251
rect 26709 10217 26743 10251
rect 26743 10217 26752 10251
rect 26700 10208 26752 10217
rect 27620 10208 27672 10260
rect 23480 10140 23532 10192
rect 23940 10183 23992 10192
rect 23940 10149 23949 10183
rect 23949 10149 23983 10183
rect 23983 10149 23992 10183
rect 23940 10140 23992 10149
rect 21088 10072 21140 10124
rect 26608 10140 26660 10192
rect 29092 10208 29144 10260
rect 29828 10208 29880 10260
rect 31392 10208 31444 10260
rect 26884 10072 26936 10124
rect 29276 10072 29328 10124
rect 29368 10115 29420 10124
rect 29368 10081 29377 10115
rect 29377 10081 29411 10115
rect 29411 10081 29420 10115
rect 29368 10072 29420 10081
rect 30656 10072 30708 10124
rect 32864 10208 32916 10260
rect 32128 10115 32180 10124
rect 32128 10081 32137 10115
rect 32137 10081 32171 10115
rect 32171 10081 32180 10115
rect 32128 10072 32180 10081
rect 20628 10004 20680 10056
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12440 9868 12492 9877
rect 13912 9868 13964 9920
rect 15016 9868 15068 9920
rect 15108 9868 15160 9920
rect 17684 9936 17736 9988
rect 16948 9911 17000 9920
rect 16948 9877 16957 9911
rect 16957 9877 16991 9911
rect 16991 9877 17000 9911
rect 16948 9868 17000 9877
rect 17316 9911 17368 9920
rect 17316 9877 17325 9911
rect 17325 9877 17359 9911
rect 17359 9877 17368 9911
rect 17316 9868 17368 9877
rect 17500 9868 17552 9920
rect 19984 9936 20036 9988
rect 18512 9911 18564 9920
rect 18512 9877 18521 9911
rect 18521 9877 18555 9911
rect 18555 9877 18564 9911
rect 18512 9868 18564 9877
rect 21364 9868 21416 9920
rect 21456 9868 21508 9920
rect 22008 9868 22060 9920
rect 24032 10004 24084 10056
rect 22468 9979 22520 9988
rect 22468 9945 22477 9979
rect 22477 9945 22511 9979
rect 22511 9945 22520 9979
rect 22468 9936 22520 9945
rect 25504 9936 25556 9988
rect 27344 9936 27396 9988
rect 24124 9911 24176 9920
rect 24124 9877 24133 9911
rect 24133 9877 24167 9911
rect 24167 9877 24176 9911
rect 24124 9868 24176 9877
rect 26700 9868 26752 9920
rect 27712 9936 27764 9988
rect 29184 9936 29236 9988
rect 30380 9936 30432 9988
rect 31852 9979 31904 9988
rect 31852 9945 31861 9979
rect 31861 9945 31895 9979
rect 31895 9945 31904 9979
rect 31852 9936 31904 9945
rect 29736 9868 29788 9920
rect 34428 10140 34480 10192
rect 32772 10115 32824 10124
rect 32772 10081 32781 10115
rect 32781 10081 32815 10115
rect 32815 10081 32824 10115
rect 32772 10072 32824 10081
rect 34704 10072 34756 10124
rect 35164 10115 35216 10124
rect 35164 10081 35173 10115
rect 35173 10081 35207 10115
rect 35207 10081 35216 10115
rect 35164 10072 35216 10081
rect 32496 10004 32548 10056
rect 34888 10047 34940 10056
rect 34888 10013 34897 10047
rect 34897 10013 34931 10047
rect 34931 10013 34940 10047
rect 34888 10004 34940 10013
rect 36636 10251 36688 10260
rect 36636 10217 36645 10251
rect 36645 10217 36679 10251
rect 36679 10217 36688 10251
rect 36636 10208 36688 10217
rect 36912 10251 36964 10260
rect 36912 10217 36921 10251
rect 36921 10217 36955 10251
rect 36955 10217 36964 10251
rect 36912 10208 36964 10217
rect 47032 10072 47084 10124
rect 49148 10115 49200 10124
rect 49148 10081 49157 10115
rect 49157 10081 49191 10115
rect 49191 10081 49200 10115
rect 49148 10072 49200 10081
rect 38936 10004 38988 10056
rect 44088 10004 44140 10056
rect 45744 10004 45796 10056
rect 46756 10004 46808 10056
rect 32680 9936 32732 9988
rect 34244 9936 34296 9988
rect 35440 9936 35492 9988
rect 32404 9868 32456 9920
rect 35808 9868 35860 9920
rect 36084 9868 36136 9920
rect 36912 9936 36964 9988
rect 42708 9936 42760 9988
rect 46204 9936 46256 9988
rect 47308 9979 47360 9988
rect 47308 9945 47317 9979
rect 47317 9945 47351 9979
rect 47351 9945 47360 9979
rect 47308 9936 47360 9945
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 1308 9664 1360 9716
rect 2412 9664 2464 9716
rect 14464 9664 14516 9716
rect 15108 9664 15160 9716
rect 15752 9664 15804 9716
rect 13728 9596 13780 9648
rect 14648 9596 14700 9648
rect 14832 9596 14884 9648
rect 15384 9596 15436 9648
rect 16488 9664 16540 9716
rect 17224 9664 17276 9716
rect 16672 9596 16724 9648
rect 18328 9596 18380 9648
rect 19524 9596 19576 9648
rect 21088 9707 21140 9716
rect 21088 9673 21097 9707
rect 21097 9673 21131 9707
rect 21131 9673 21140 9707
rect 21088 9664 21140 9673
rect 21272 9596 21324 9648
rect 22284 9707 22336 9716
rect 22284 9673 22293 9707
rect 22293 9673 22327 9707
rect 22327 9673 22336 9707
rect 22284 9664 22336 9673
rect 26056 9664 26108 9716
rect 31760 9664 31812 9716
rect 1308 9528 1360 9580
rect 12348 9528 12400 9580
rect 20628 9528 20680 9580
rect 11060 9460 11112 9512
rect 1768 9435 1820 9444
rect 1768 9401 1777 9435
rect 1777 9401 1811 9435
rect 1811 9401 1820 9435
rect 1768 9392 1820 9401
rect 15108 9503 15160 9512
rect 15108 9469 15117 9503
rect 15117 9469 15151 9503
rect 15151 9469 15160 9503
rect 15108 9460 15160 9469
rect 12532 9392 12584 9444
rect 14096 9392 14148 9444
rect 13636 9324 13688 9376
rect 16028 9460 16080 9512
rect 17592 9460 17644 9512
rect 18604 9503 18656 9512
rect 18604 9469 18613 9503
rect 18613 9469 18647 9503
rect 18647 9469 18656 9503
rect 18604 9460 18656 9469
rect 18880 9503 18932 9512
rect 18880 9469 18889 9503
rect 18889 9469 18923 9503
rect 18923 9469 18932 9503
rect 18880 9460 18932 9469
rect 17316 9392 17368 9444
rect 23480 9596 23532 9648
rect 24676 9596 24728 9648
rect 22652 9571 22704 9580
rect 22652 9537 22661 9571
rect 22661 9537 22695 9571
rect 22695 9537 22704 9571
rect 22652 9528 22704 9537
rect 22008 9392 22060 9444
rect 15660 9367 15712 9376
rect 15660 9333 15669 9367
rect 15669 9333 15703 9367
rect 15703 9333 15712 9367
rect 15660 9324 15712 9333
rect 16212 9324 16264 9376
rect 16488 9324 16540 9376
rect 18512 9324 18564 9376
rect 21548 9324 21600 9376
rect 21824 9367 21876 9376
rect 21824 9333 21833 9367
rect 21833 9333 21867 9367
rect 21867 9333 21876 9367
rect 21824 9324 21876 9333
rect 24308 9460 24360 9512
rect 27344 9596 27396 9648
rect 27712 9596 27764 9648
rect 30104 9596 30156 9648
rect 30656 9596 30708 9648
rect 31944 9596 31996 9648
rect 32128 9596 32180 9648
rect 32496 9596 32548 9648
rect 34888 9664 34940 9716
rect 35164 9664 35216 9716
rect 36084 9707 36136 9716
rect 36084 9673 36093 9707
rect 36093 9673 36127 9707
rect 36127 9673 36136 9707
rect 36084 9664 36136 9673
rect 25964 9503 26016 9512
rect 25964 9469 25973 9503
rect 25973 9469 26007 9503
rect 26007 9469 26016 9503
rect 25964 9460 26016 9469
rect 23756 9324 23808 9376
rect 25688 9392 25740 9444
rect 31668 9528 31720 9580
rect 35992 9596 36044 9648
rect 49240 9596 49292 9648
rect 47124 9528 47176 9580
rect 27160 9392 27212 9444
rect 29276 9503 29328 9512
rect 29276 9469 29285 9503
rect 29285 9469 29319 9503
rect 29319 9469 29328 9503
rect 29276 9460 29328 9469
rect 30012 9503 30064 9512
rect 30012 9469 30021 9503
rect 30021 9469 30055 9503
rect 30055 9469 30064 9503
rect 30012 9460 30064 9469
rect 30104 9460 30156 9512
rect 31576 9460 31628 9512
rect 31760 9460 31812 9512
rect 31944 9460 31996 9512
rect 34152 9503 34204 9512
rect 34152 9469 34161 9503
rect 34161 9469 34195 9503
rect 34195 9469 34204 9503
rect 35900 9503 35952 9512
rect 34152 9460 34204 9469
rect 35900 9469 35909 9503
rect 35909 9469 35943 9503
rect 35943 9469 35952 9503
rect 35900 9460 35952 9469
rect 25412 9324 25464 9376
rect 32772 9392 32824 9444
rect 30472 9324 30524 9376
rect 30656 9324 30708 9376
rect 31576 9324 31628 9376
rect 31760 9324 31812 9376
rect 32864 9324 32916 9376
rect 35532 9324 35584 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 17224 9120 17276 9172
rect 17868 9163 17920 9172
rect 17868 9129 17889 9163
rect 17889 9129 17920 9163
rect 17868 9120 17920 9129
rect 19524 9120 19576 9172
rect 22100 9120 22152 9172
rect 22468 9120 22520 9172
rect 32404 9120 32456 9172
rect 36360 9120 36412 9172
rect 43720 9120 43772 9172
rect 16856 9052 16908 9104
rect 1216 8916 1268 8968
rect 15108 8984 15160 9036
rect 15476 9027 15528 9036
rect 15476 8993 15485 9027
rect 15485 8993 15519 9027
rect 15519 8993 15528 9027
rect 15476 8984 15528 8993
rect 16028 8984 16080 9036
rect 18880 8984 18932 9036
rect 19432 8984 19484 9036
rect 1308 8848 1360 8900
rect 11980 8916 12032 8968
rect 15568 8959 15620 8968
rect 15568 8925 15577 8959
rect 15577 8925 15611 8959
rect 15611 8925 15620 8959
rect 15568 8916 15620 8925
rect 18696 8959 18748 8968
rect 18696 8925 18705 8959
rect 18705 8925 18739 8959
rect 18739 8925 18748 8959
rect 18696 8916 18748 8925
rect 21456 8916 21508 8968
rect 22008 8916 22060 8968
rect 23388 8984 23440 9036
rect 23756 9027 23808 9036
rect 23756 8993 23765 9027
rect 23765 8993 23799 9027
rect 23799 8993 23808 9027
rect 23756 8984 23808 8993
rect 30012 9052 30064 9104
rect 28448 8984 28500 9036
rect 31760 8984 31812 9036
rect 33876 9052 33928 9104
rect 34244 9052 34296 9104
rect 36268 9052 36320 9104
rect 32496 9027 32548 9036
rect 32496 8993 32505 9027
rect 32505 8993 32539 9027
rect 32539 8993 32548 9027
rect 32496 8984 32548 8993
rect 33048 8984 33100 9036
rect 34152 8984 34204 9036
rect 34980 9027 35032 9036
rect 34980 8993 34989 9027
rect 34989 8993 35023 9027
rect 35023 8993 35032 9027
rect 34980 8984 35032 8993
rect 35072 8984 35124 9036
rect 24032 8959 24084 8968
rect 24032 8925 24041 8959
rect 24041 8925 24075 8959
rect 24075 8925 24084 8959
rect 24032 8916 24084 8925
rect 16120 8848 16172 8900
rect 16212 8848 16264 8900
rect 14924 8823 14976 8832
rect 14924 8789 14933 8823
rect 14933 8789 14967 8823
rect 14967 8789 14976 8823
rect 14924 8780 14976 8789
rect 15936 8823 15988 8832
rect 15936 8789 15945 8823
rect 15945 8789 15979 8823
rect 15979 8789 15988 8823
rect 15936 8780 15988 8789
rect 16396 8823 16448 8832
rect 16396 8789 16405 8823
rect 16405 8789 16439 8823
rect 16439 8789 16448 8823
rect 16396 8780 16448 8789
rect 17408 8848 17460 8900
rect 18328 8848 18380 8900
rect 20444 8848 20496 8900
rect 25964 8916 26016 8968
rect 30840 8916 30892 8968
rect 34796 8916 34848 8968
rect 35532 8984 35584 9036
rect 44180 8984 44232 9036
rect 49332 8984 49384 9036
rect 47676 8916 47728 8968
rect 47768 8916 47820 8968
rect 18788 8780 18840 8832
rect 18880 8780 18932 8832
rect 22192 8780 22244 8832
rect 30932 8848 30984 8900
rect 32772 8848 32824 8900
rect 36452 8848 36504 8900
rect 23480 8780 23532 8832
rect 25688 8823 25740 8832
rect 25688 8789 25697 8823
rect 25697 8789 25731 8823
rect 25731 8789 25740 8823
rect 25688 8780 25740 8789
rect 27804 8823 27856 8832
rect 27804 8789 27813 8823
rect 27813 8789 27847 8823
rect 27847 8789 27856 8823
rect 28448 8823 28500 8832
rect 27804 8780 27856 8789
rect 28448 8789 28457 8823
rect 28457 8789 28491 8823
rect 28491 8789 28500 8823
rect 28448 8780 28500 8789
rect 30380 8780 30432 8832
rect 30656 8780 30708 8832
rect 32864 8823 32916 8832
rect 32864 8789 32873 8823
rect 32873 8789 32907 8823
rect 32907 8789 32916 8823
rect 32864 8780 32916 8789
rect 33140 8780 33192 8832
rect 33600 8823 33652 8832
rect 33600 8789 33609 8823
rect 33609 8789 33643 8823
rect 33643 8789 33652 8823
rect 33600 8780 33652 8789
rect 34244 8780 34296 8832
rect 35256 8823 35308 8832
rect 35256 8789 35265 8823
rect 35265 8789 35299 8823
rect 35299 8789 35308 8823
rect 35256 8780 35308 8789
rect 35624 8823 35676 8832
rect 35624 8789 35633 8823
rect 35633 8789 35667 8823
rect 35667 8789 35676 8823
rect 35624 8780 35676 8789
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 13544 8576 13596 8628
rect 13728 8576 13780 8628
rect 13912 8551 13964 8560
rect 13912 8517 13921 8551
rect 13921 8517 13955 8551
rect 13955 8517 13964 8551
rect 13912 8508 13964 8517
rect 16396 8508 16448 8560
rect 16764 8508 16816 8560
rect 18604 8619 18656 8628
rect 18604 8585 18613 8619
rect 18613 8585 18647 8619
rect 18647 8585 18656 8619
rect 18604 8576 18656 8585
rect 19892 8576 19944 8628
rect 18880 8508 18932 8560
rect 20444 8508 20496 8560
rect 2688 8440 2740 8492
rect 14924 8440 14976 8492
rect 2412 8415 2464 8424
rect 2412 8381 2421 8415
rect 2421 8381 2455 8415
rect 2455 8381 2464 8415
rect 2412 8372 2464 8381
rect 13636 8415 13688 8424
rect 13636 8381 13645 8415
rect 13645 8381 13679 8415
rect 13679 8381 13688 8415
rect 13636 8372 13688 8381
rect 16028 8440 16080 8492
rect 18236 8440 18288 8492
rect 18512 8440 18564 8492
rect 15108 8372 15160 8424
rect 17132 8372 17184 8424
rect 21456 8415 21508 8424
rect 21456 8381 21465 8415
rect 21465 8381 21499 8415
rect 21499 8381 21508 8415
rect 21456 8372 21508 8381
rect 23480 8576 23532 8628
rect 32772 8576 32824 8628
rect 33876 8576 33928 8628
rect 34980 8576 35032 8628
rect 29092 8551 29144 8560
rect 29092 8517 29101 8551
rect 29101 8517 29135 8551
rect 29135 8517 29144 8551
rect 29092 8508 29144 8517
rect 30472 8508 30524 8560
rect 32036 8508 32088 8560
rect 32864 8508 32916 8560
rect 33140 8508 33192 8560
rect 35992 8576 36044 8628
rect 40040 8576 40092 8628
rect 42708 8576 42760 8628
rect 35624 8508 35676 8560
rect 22008 8440 22060 8492
rect 24032 8440 24084 8492
rect 30656 8440 30708 8492
rect 30932 8440 30984 8492
rect 31116 8440 31168 8492
rect 31760 8440 31812 8492
rect 32312 8483 32364 8492
rect 32312 8449 32321 8483
rect 32321 8449 32355 8483
rect 32355 8449 32364 8483
rect 32312 8440 32364 8449
rect 35808 8440 35860 8492
rect 40316 8551 40368 8560
rect 40316 8517 40325 8551
rect 40325 8517 40359 8551
rect 40359 8517 40368 8551
rect 40316 8508 40368 8517
rect 44180 8551 44232 8560
rect 44180 8517 44189 8551
rect 44189 8517 44223 8551
rect 44223 8517 44232 8551
rect 44180 8508 44232 8517
rect 45468 8576 45520 8628
rect 47584 8576 47636 8628
rect 45468 8440 45520 8492
rect 49148 8551 49200 8560
rect 49148 8517 49157 8551
rect 49157 8517 49191 8551
rect 49191 8517 49200 8551
rect 49148 8508 49200 8517
rect 46204 8440 46256 8492
rect 22100 8372 22152 8424
rect 28816 8415 28868 8424
rect 28816 8381 28825 8415
rect 28825 8381 28859 8415
rect 28859 8381 28868 8415
rect 28816 8372 28868 8381
rect 29184 8372 29236 8424
rect 31944 8372 31996 8424
rect 32220 8372 32272 8424
rect 32588 8415 32640 8424
rect 32588 8381 32597 8415
rect 32597 8381 32631 8415
rect 32631 8381 32640 8415
rect 32588 8372 32640 8381
rect 32956 8372 33008 8424
rect 38752 8372 38804 8424
rect 22468 8304 22520 8356
rect 31852 8304 31904 8356
rect 17316 8236 17368 8288
rect 31944 8236 31996 8288
rect 33048 8236 33100 8288
rect 33692 8236 33744 8288
rect 40224 8372 40276 8424
rect 44916 8304 44968 8356
rect 46848 8415 46900 8424
rect 46848 8381 46857 8415
rect 46857 8381 46891 8415
rect 46891 8381 46900 8415
rect 46848 8372 46900 8381
rect 47768 8304 47820 8356
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 1308 8032 1360 8084
rect 2412 8032 2464 8084
rect 18420 8032 18472 8084
rect 19432 8075 19484 8084
rect 19432 8041 19441 8075
rect 19441 8041 19475 8075
rect 19475 8041 19484 8075
rect 19432 8032 19484 8041
rect 21916 8032 21968 8084
rect 30564 8032 30616 8084
rect 35256 8032 35308 8084
rect 18880 7964 18932 8016
rect 21640 7964 21692 8016
rect 22652 7964 22704 8016
rect 32588 7964 32640 8016
rect 39028 7964 39080 8016
rect 16764 7939 16816 7948
rect 16764 7905 16773 7939
rect 16773 7905 16807 7939
rect 16807 7905 16816 7939
rect 16764 7896 16816 7905
rect 16948 7939 17000 7948
rect 16948 7905 16957 7939
rect 16957 7905 16991 7939
rect 16991 7905 17000 7939
rect 16948 7896 17000 7905
rect 18604 7896 18656 7948
rect 19892 7896 19944 7948
rect 23664 7896 23716 7948
rect 29920 7939 29972 7948
rect 29920 7905 29929 7939
rect 29929 7905 29963 7939
rect 29963 7905 29972 7939
rect 29920 7896 29972 7905
rect 32220 7896 32272 7948
rect 34520 7896 34572 7948
rect 49240 7896 49292 7948
rect 1308 7828 1360 7880
rect 14096 7828 14148 7880
rect 17040 7871 17092 7880
rect 17040 7837 17049 7871
rect 17049 7837 17083 7871
rect 17083 7837 17092 7871
rect 17040 7828 17092 7837
rect 13728 7760 13780 7812
rect 16304 7760 16356 7812
rect 19616 7760 19668 7812
rect 20444 7760 20496 7812
rect 20996 7760 21048 7812
rect 21456 7828 21508 7880
rect 22192 7828 22244 7880
rect 30564 7828 30616 7880
rect 32680 7871 32732 7880
rect 32680 7837 32689 7871
rect 32689 7837 32723 7871
rect 32723 7837 32732 7871
rect 32680 7828 32732 7837
rect 38752 7871 38804 7880
rect 38752 7837 38761 7871
rect 38761 7837 38795 7871
rect 38795 7837 38804 7871
rect 38752 7828 38804 7837
rect 46940 7828 46992 7880
rect 30472 7803 30524 7812
rect 30472 7769 30481 7803
rect 30481 7769 30515 7803
rect 30515 7769 30524 7803
rect 30472 7760 30524 7769
rect 21456 7735 21508 7744
rect 21456 7701 21465 7735
rect 21465 7701 21499 7735
rect 21499 7701 21508 7735
rect 21456 7692 21508 7701
rect 21640 7735 21692 7744
rect 21640 7701 21649 7735
rect 21649 7701 21683 7735
rect 21683 7701 21692 7735
rect 21640 7692 21692 7701
rect 22376 7692 22428 7744
rect 22468 7735 22520 7744
rect 22468 7701 22477 7735
rect 22477 7701 22511 7735
rect 22511 7701 22520 7735
rect 22468 7692 22520 7701
rect 25688 7692 25740 7744
rect 27528 7692 27580 7744
rect 40132 7760 40184 7812
rect 30656 7735 30708 7744
rect 30656 7701 30665 7735
rect 30665 7701 30699 7735
rect 30699 7701 30708 7735
rect 30656 7692 30708 7701
rect 31392 7735 31444 7744
rect 31392 7701 31401 7735
rect 31401 7701 31435 7735
rect 31435 7701 31444 7735
rect 31392 7692 31444 7701
rect 32588 7735 32640 7744
rect 32588 7701 32597 7735
rect 32597 7701 32631 7735
rect 32631 7701 32640 7735
rect 32588 7692 32640 7701
rect 38660 7692 38712 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 19800 7488 19852 7540
rect 22284 7488 22336 7540
rect 31116 7531 31168 7540
rect 31116 7497 31125 7531
rect 31125 7497 31159 7531
rect 31159 7497 31168 7531
rect 31116 7488 31168 7497
rect 31392 7488 31444 7540
rect 17868 7420 17920 7472
rect 18512 7420 18564 7472
rect 20444 7420 20496 7472
rect 31944 7463 31996 7472
rect 31944 7429 31953 7463
rect 31953 7429 31987 7463
rect 31987 7429 31996 7463
rect 31944 7420 31996 7429
rect 34428 7420 34480 7472
rect 38660 7420 38712 7472
rect 47308 7420 47360 7472
rect 49332 7420 49384 7472
rect 1308 7352 1360 7404
rect 22376 7395 22428 7404
rect 22376 7361 22385 7395
rect 22385 7361 22419 7395
rect 22419 7361 22428 7395
rect 22376 7352 22428 7361
rect 22560 7327 22612 7336
rect 22560 7293 22569 7327
rect 22569 7293 22603 7327
rect 22603 7293 22612 7327
rect 22560 7284 22612 7293
rect 19248 7216 19300 7268
rect 28632 7216 28684 7268
rect 44916 7395 44968 7404
rect 44916 7361 44925 7395
rect 44925 7361 44959 7395
rect 44959 7361 44968 7395
rect 44916 7352 44968 7361
rect 47032 7352 47084 7404
rect 21456 7148 21508 7200
rect 22008 7148 22060 7200
rect 32588 7148 32640 7200
rect 37280 7148 37332 7200
rect 37924 7191 37976 7200
rect 37924 7157 37933 7191
rect 37933 7157 37967 7191
rect 37967 7157 37976 7191
rect 37924 7148 37976 7157
rect 47860 7216 47912 7268
rect 45836 7148 45888 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 30472 6944 30524 6996
rect 38476 6944 38528 6996
rect 37924 6876 37976 6928
rect 46940 6876 46992 6928
rect 15660 6808 15712 6860
rect 22376 6808 22428 6860
rect 49148 6851 49200 6860
rect 49148 6817 49157 6851
rect 49157 6817 49191 6851
rect 49191 6817 49200 6851
rect 49148 6808 49200 6817
rect 1308 6740 1360 6792
rect 15936 6740 15988 6792
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 40132 6740 40184 6792
rect 47768 6740 47820 6792
rect 1216 6672 1268 6724
rect 1768 6647 1820 6656
rect 1768 6613 1777 6647
rect 1777 6613 1811 6647
rect 1811 6613 1820 6647
rect 1768 6604 1820 6613
rect 10600 6672 10652 6724
rect 48688 6672 48740 6724
rect 19248 6604 19300 6656
rect 21732 6604 21784 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 1216 6400 1268 6452
rect 1768 6332 1820 6384
rect 27804 6332 27856 6384
rect 30748 6332 30800 6384
rect 40040 6332 40092 6384
rect 49332 6332 49384 6384
rect 1308 6264 1360 6316
rect 16856 6264 16908 6316
rect 47676 6264 47728 6316
rect 18328 6196 18380 6248
rect 11244 6128 11296 6180
rect 47032 6128 47084 6180
rect 19432 6060 19484 6112
rect 37648 6103 37700 6112
rect 37648 6069 37657 6103
rect 37657 6069 37691 6103
rect 37691 6069 37700 6103
rect 37648 6060 37700 6069
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 37648 5856 37700 5908
rect 47216 5856 47268 5908
rect 13360 5788 13412 5840
rect 1308 5652 1360 5704
rect 49240 5720 49292 5772
rect 2780 5652 2832 5704
rect 43720 5695 43772 5704
rect 43720 5661 43729 5695
rect 43729 5661 43763 5695
rect 43763 5661 43772 5695
rect 43720 5652 43772 5661
rect 47584 5652 47636 5704
rect 16212 5584 16264 5636
rect 45744 5584 45796 5636
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 37280 5244 37332 5296
rect 38476 5287 38528 5296
rect 38476 5253 38485 5287
rect 38485 5253 38519 5287
rect 38519 5253 38528 5287
rect 38476 5244 38528 5253
rect 49148 5287 49200 5296
rect 49148 5253 49157 5287
rect 49157 5253 49191 5287
rect 49191 5253 49200 5287
rect 49148 5244 49200 5253
rect 12808 5176 12860 5228
rect 18880 5219 18932 5228
rect 18880 5185 18889 5219
rect 18889 5185 18923 5219
rect 18923 5185 18932 5219
rect 18880 5176 18932 5185
rect 45836 5219 45888 5228
rect 45836 5185 45845 5219
rect 45845 5185 45879 5219
rect 45879 5185 45888 5219
rect 45836 5176 45888 5185
rect 47860 5176 47912 5228
rect 1308 5108 1360 5160
rect 19064 5151 19116 5160
rect 19064 5117 19073 5151
rect 19073 5117 19107 5151
rect 19107 5117 19116 5151
rect 19064 5108 19116 5117
rect 48320 5108 48372 5160
rect 40040 5040 40092 5092
rect 20628 4972 20680 5024
rect 37832 5015 37884 5024
rect 37832 4981 37841 5015
rect 37841 4981 37875 5015
rect 37875 4981 37884 5015
rect 37832 4972 37884 4981
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 1308 4768 1360 4820
rect 24124 4768 24176 4820
rect 37832 4768 37884 4820
rect 47124 4768 47176 4820
rect 26148 4700 26200 4752
rect 37004 4700 37056 4752
rect 19248 4632 19300 4684
rect 21732 4632 21784 4684
rect 1308 4564 1360 4616
rect 19984 4564 20036 4616
rect 22928 4632 22980 4684
rect 23204 4632 23256 4684
rect 27252 4632 27304 4684
rect 40224 4700 40276 4752
rect 22100 4607 22152 4616
rect 22100 4573 22109 4607
rect 22109 4573 22143 4607
rect 22143 4573 22152 4607
rect 22100 4564 22152 4573
rect 19064 4496 19116 4548
rect 23572 4564 23624 4616
rect 32772 4564 32824 4616
rect 49424 4632 49476 4684
rect 47308 4564 47360 4616
rect 21272 4428 21324 4480
rect 21456 4428 21508 4480
rect 21824 4428 21876 4480
rect 27068 4496 27120 4548
rect 25872 4428 25924 4480
rect 37372 4471 37424 4480
rect 37372 4437 37381 4471
rect 37381 4437 37415 4471
rect 37415 4437 37424 4471
rect 37372 4428 37424 4437
rect 39764 4428 39816 4480
rect 47676 4496 47728 4548
rect 49792 4428 49844 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 1400 4156 1452 4208
rect 1308 3952 1360 4004
rect 37372 4224 37424 4276
rect 45652 4224 45704 4276
rect 22100 4156 22152 4208
rect 15660 4088 15712 4140
rect 17960 3952 18012 4004
rect 18328 3952 18380 4004
rect 22928 4131 22980 4140
rect 22928 4097 22972 4131
rect 22972 4097 22980 4131
rect 22928 4088 22980 4097
rect 23204 4088 23256 4140
rect 25872 4199 25924 4208
rect 25872 4165 25881 4199
rect 25881 4165 25915 4199
rect 25915 4165 25924 4199
rect 25872 4156 25924 4165
rect 27620 4088 27672 4140
rect 45836 4131 45888 4140
rect 45836 4097 45845 4131
rect 45845 4097 45879 4131
rect 45879 4097 45888 4131
rect 45836 4088 45888 4097
rect 46940 4088 46992 4140
rect 49332 4088 49384 4140
rect 23296 4020 23348 4072
rect 24860 4063 24912 4072
rect 24860 4029 24869 4063
rect 24869 4029 24903 4063
rect 24903 4029 24912 4063
rect 24860 4020 24912 4029
rect 25780 4020 25832 4072
rect 21640 3884 21692 3936
rect 22836 3884 22888 3936
rect 32864 4020 32916 4072
rect 46664 4063 46716 4072
rect 46664 4029 46673 4063
rect 46673 4029 46707 4063
rect 46707 4029 46716 4063
rect 46664 4020 46716 4029
rect 27528 3884 27580 3936
rect 47676 3927 47728 3936
rect 47676 3893 47685 3927
rect 47685 3893 47719 3927
rect 47719 3893 47728 3927
rect 47676 3884 47728 3893
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 7472 3680 7524 3732
rect 3332 3612 3384 3664
rect 12440 3544 12492 3596
rect 1308 3476 1360 3528
rect 22008 3680 22060 3732
rect 23572 3723 23624 3732
rect 23572 3689 23581 3723
rect 23581 3689 23615 3723
rect 23615 3689 23624 3723
rect 23572 3680 23624 3689
rect 25964 3680 26016 3732
rect 24952 3612 25004 3664
rect 26332 3612 26384 3664
rect 29644 3612 29696 3664
rect 33416 3612 33468 3664
rect 17960 3476 18012 3528
rect 20996 3519 21048 3528
rect 20996 3485 21005 3519
rect 21005 3485 21039 3519
rect 21039 3485 21048 3519
rect 20996 3476 21048 3485
rect 13912 3408 13964 3460
rect 19340 3408 19392 3460
rect 21364 3408 21416 3460
rect 22008 3408 22060 3460
rect 22836 3544 22888 3596
rect 29000 3544 29052 3596
rect 40040 3544 40092 3596
rect 24032 3519 24084 3528
rect 24032 3485 24041 3519
rect 24041 3485 24075 3519
rect 24075 3485 24084 3519
rect 24032 3476 24084 3485
rect 28356 3476 28408 3528
rect 39212 3476 39264 3528
rect 23940 3408 23992 3460
rect 21456 3340 21508 3392
rect 22744 3383 22796 3392
rect 22744 3349 22753 3383
rect 22753 3349 22787 3383
rect 22787 3349 22796 3383
rect 22744 3340 22796 3349
rect 23112 3340 23164 3392
rect 45836 3476 45888 3528
rect 49148 3587 49200 3596
rect 49148 3553 49157 3587
rect 49157 3553 49191 3587
rect 49191 3553 49200 3587
rect 49148 3544 49200 3553
rect 47032 3476 47084 3528
rect 45560 3451 45612 3460
rect 45560 3417 45569 3451
rect 45569 3417 45603 3451
rect 45603 3417 45612 3451
rect 45560 3408 45612 3417
rect 48688 3408 48740 3460
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 1308 3136 1360 3188
rect 1308 3000 1360 3052
rect 9680 3043 9732 3052
rect 9680 3009 9689 3043
rect 9689 3009 9723 3043
rect 9723 3009 9732 3043
rect 9680 3000 9732 3009
rect 19340 3136 19392 3188
rect 17868 3068 17920 3120
rect 13636 3000 13688 3052
rect 19064 3000 19116 3052
rect 21456 3179 21508 3188
rect 21456 3145 21465 3179
rect 21465 3145 21499 3179
rect 21499 3145 21508 3179
rect 21456 3136 21508 3145
rect 20628 3043 20680 3052
rect 20628 3009 20637 3043
rect 20637 3009 20671 3043
rect 20671 3009 20680 3043
rect 20628 3000 20680 3009
rect 21272 3043 21324 3052
rect 21272 3009 21281 3043
rect 21281 3009 21315 3043
rect 21315 3009 21324 3043
rect 21272 3000 21324 3009
rect 22192 3000 22244 3052
rect 24032 3068 24084 3120
rect 24952 3068 25004 3120
rect 26148 3000 26200 3052
rect 37740 3136 37792 3188
rect 29644 3068 29696 3120
rect 49240 3068 49292 3120
rect 28816 3000 28868 3052
rect 39764 3000 39816 3052
rect 45744 3000 45796 3052
rect 47216 3000 47268 3052
rect 18328 2975 18380 2984
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18328 2932 18380 2941
rect 20996 2932 21048 2984
rect 12716 2864 12768 2916
rect 22100 2864 22152 2916
rect 22192 2907 22244 2916
rect 22192 2873 22201 2907
rect 22201 2873 22235 2907
rect 22235 2873 22244 2907
rect 22192 2864 22244 2873
rect 22744 2864 22796 2916
rect 25964 2975 26016 2984
rect 25964 2941 25973 2975
rect 25973 2941 26007 2975
rect 26007 2941 26016 2975
rect 25964 2932 26016 2941
rect 29644 2932 29696 2984
rect 30656 2932 30708 2984
rect 46756 2932 46808 2984
rect 46848 2975 46900 2984
rect 46848 2941 46857 2975
rect 46857 2941 46891 2975
rect 46891 2941 46900 2975
rect 46848 2932 46900 2941
rect 2320 2839 2372 2848
rect 2320 2805 2329 2839
rect 2329 2805 2363 2839
rect 2363 2805 2372 2839
rect 2320 2796 2372 2805
rect 2780 2839 2832 2848
rect 2780 2805 2789 2839
rect 2789 2805 2823 2839
rect 2823 2805 2832 2839
rect 2780 2796 2832 2805
rect 17408 2839 17460 2848
rect 17408 2805 17417 2839
rect 17417 2805 17451 2839
rect 17451 2805 17460 2839
rect 17408 2796 17460 2805
rect 21364 2796 21416 2848
rect 23296 2839 23348 2848
rect 23296 2805 23305 2839
rect 23305 2805 23339 2839
rect 23339 2805 23348 2839
rect 23296 2796 23348 2805
rect 27528 2907 27580 2916
rect 27528 2873 27537 2907
rect 27537 2873 27571 2907
rect 27571 2873 27580 2907
rect 27528 2864 27580 2873
rect 27160 2796 27212 2848
rect 38292 2864 38344 2916
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 9680 2524 9732 2576
rect 24032 2635 24084 2644
rect 24032 2601 24041 2635
rect 24041 2601 24075 2635
rect 24075 2601 24084 2635
rect 24032 2592 24084 2601
rect 26332 2635 26384 2644
rect 26332 2601 26341 2635
rect 26341 2601 26375 2635
rect 26375 2601 26384 2635
rect 26332 2592 26384 2601
rect 27620 2592 27672 2644
rect 29000 2635 29052 2644
rect 29000 2601 29009 2635
rect 29009 2601 29043 2635
rect 29043 2601 29052 2635
rect 29000 2592 29052 2601
rect 32864 2592 32916 2644
rect 22468 2524 22520 2576
rect 32772 2524 32824 2576
rect 34428 2524 34480 2576
rect 1308 2388 1360 2440
rect 2780 2388 2832 2440
rect 1216 2320 1268 2372
rect 2320 2320 2372 2372
rect 1308 2252 1360 2304
rect 12256 2456 12308 2508
rect 9588 2388 9640 2440
rect 13912 2388 13964 2440
rect 17408 2388 17460 2440
rect 9588 2252 9640 2304
rect 11704 2320 11756 2372
rect 13820 2320 13872 2372
rect 15936 2320 15988 2372
rect 14740 2252 14792 2304
rect 19984 2456 20036 2508
rect 20168 2456 20220 2508
rect 22284 2456 22336 2508
rect 24400 2456 24452 2508
rect 26516 2456 26568 2508
rect 37740 2499 37792 2508
rect 37740 2465 37749 2499
rect 37749 2465 37783 2499
rect 37783 2465 37792 2499
rect 37740 2456 37792 2465
rect 41328 2456 41380 2508
rect 49148 2499 49200 2508
rect 49148 2465 49157 2499
rect 49157 2465 49191 2499
rect 49191 2465 49200 2499
rect 49148 2456 49200 2465
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 22100 2388 22152 2440
rect 21456 2320 21508 2372
rect 27160 2431 27212 2440
rect 27160 2397 27169 2431
rect 27169 2397 27203 2431
rect 27203 2397 27212 2431
rect 27160 2388 27212 2397
rect 29000 2388 29052 2440
rect 30748 2388 30800 2440
rect 33140 2431 33192 2440
rect 33140 2397 33149 2431
rect 33149 2397 33183 2431
rect 33183 2397 33192 2431
rect 33140 2388 33192 2397
rect 34980 2388 35032 2440
rect 38292 2388 38344 2440
rect 45652 2388 45704 2440
rect 47124 2388 47176 2440
rect 48504 2320 48556 2372
rect 37096 2295 37148 2304
rect 37096 2261 37105 2295
rect 37105 2261 37139 2295
rect 37139 2261 37148 2295
rect 37096 2252 37148 2261
rect 43444 2252 43496 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
<< metal2 >>
rect 1582 26200 1638 27000
rect 2226 26200 2282 27000
rect 2870 26330 2926 27000
rect 2870 26302 3372 26330
rect 2870 26200 2926 26302
rect 1596 22778 1624 26200
rect 1768 23044 1820 23050
rect 1768 22986 1820 22992
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 1032 21956 1084 21962
rect 1032 21898 1084 21904
rect 1044 20777 1072 21898
rect 1780 21593 1808 22986
rect 2240 22234 2268 26200
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2778 24440 2834 24449
rect 2950 24443 3258 24452
rect 2778 24375 2834 24384
rect 2792 23526 2820 24375
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 3054 23216 3110 23225
rect 3054 23151 3110 23160
rect 2870 22808 2926 22817
rect 2870 22743 2926 22752
rect 2780 22568 2832 22574
rect 2780 22510 2832 22516
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 1766 21584 1822 21593
rect 1766 21519 1822 21528
rect 1768 21480 1820 21486
rect 1768 21422 1820 21428
rect 1030 20768 1086 20777
rect 1030 20703 1086 20712
rect 1308 20528 1360 20534
rect 1308 20470 1360 20476
rect 1320 20369 1348 20470
rect 1306 20360 1362 20369
rect 1306 20295 1362 20304
rect 1780 19961 1808 21422
rect 2792 21185 2820 22510
rect 2884 22166 2912 22743
rect 3068 22438 3096 23151
rect 3056 22432 3108 22438
rect 3056 22374 3108 22380
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2872 22160 2924 22166
rect 2872 22102 2924 22108
rect 3238 21992 3294 22001
rect 3238 21927 3240 21936
rect 3292 21927 3294 21936
rect 3240 21898 3292 21904
rect 3344 21622 3372 26302
rect 3514 26200 3570 27000
rect 4158 26200 4214 27000
rect 4802 26200 4858 27000
rect 5446 26200 5502 27000
rect 6090 26200 6146 27000
rect 6734 26200 6790 27000
rect 7378 26200 7434 27000
rect 8022 26200 8078 27000
rect 8666 26200 8722 27000
rect 9310 26200 9366 27000
rect 9954 26200 10010 27000
rect 10598 26200 10654 27000
rect 11242 26200 11298 27000
rect 11886 26200 11942 27000
rect 12530 26330 12586 27000
rect 13174 26330 13230 27000
rect 12530 26302 12848 26330
rect 12530 26200 12586 26302
rect 3422 25664 3478 25673
rect 3422 25599 3478 25608
rect 3436 24886 3464 25599
rect 3424 24880 3476 24886
rect 3424 24822 3476 24828
rect 3528 24274 3556 26200
rect 3698 25256 3754 25265
rect 3698 25191 3754 25200
rect 3606 24848 3662 24857
rect 3606 24783 3608 24792
rect 3660 24783 3662 24792
rect 3608 24754 3660 24760
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3514 24032 3570 24041
rect 3514 23967 3570 23976
rect 3422 23624 3478 23633
rect 3422 23559 3424 23568
rect 3476 23559 3478 23568
rect 3424 23530 3476 23536
rect 3424 22772 3476 22778
rect 3424 22714 3476 22720
rect 3332 21616 3384 21622
rect 3332 21558 3384 21564
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2778 21176 2834 21185
rect 2950 21179 3258 21188
rect 2778 21111 2834 21120
rect 2872 21004 2924 21010
rect 2872 20946 2924 20952
rect 2780 20324 2832 20330
rect 2780 20266 2832 20272
rect 1766 19952 1822 19961
rect 1766 19887 1822 19896
rect 1492 19780 1544 19786
rect 1492 19722 1544 19728
rect 1504 18737 1532 19722
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1490 18728 1546 18737
rect 1400 18692 1452 18698
rect 1490 18663 1546 18672
rect 1400 18634 1452 18640
rect 1412 17921 1440 18634
rect 1780 18329 1808 19314
rect 2792 19145 2820 20266
rect 2884 19553 2912 20946
rect 3332 20324 3384 20330
rect 3332 20266 3384 20272
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 3344 19854 3372 20266
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 2870 19544 2926 19553
rect 2870 19479 2926 19488
rect 3436 19446 3464 22714
rect 3424 19440 3476 19446
rect 3424 19382 3476 19388
rect 2778 19136 2834 19145
rect 2778 19071 2834 19080
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 3528 18834 3556 23967
rect 3608 22772 3660 22778
rect 3608 22714 3660 22720
rect 3516 18828 3568 18834
rect 3516 18770 3568 18776
rect 3620 18426 3648 22714
rect 3712 22094 3740 25191
rect 3884 24200 3936 24206
rect 3884 24142 3936 24148
rect 3712 22066 3832 22094
rect 3804 21350 3832 22066
rect 3792 21344 3844 21350
rect 3792 21286 3844 21292
rect 3896 19310 3924 24142
rect 4068 23724 4120 23730
rect 4068 23666 4120 23672
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3988 19417 4016 20402
rect 3974 19408 4030 19417
rect 3974 19343 4030 19352
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 1766 18320 1822 18329
rect 4080 18290 4108 23666
rect 4172 23662 4200 26200
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 4632 23866 4660 24142
rect 4620 23860 4672 23866
rect 4620 23802 4672 23808
rect 4712 23724 4764 23730
rect 4712 23666 4764 23672
rect 4160 23656 4212 23662
rect 4160 23598 4212 23604
rect 4724 23322 4752 23666
rect 4712 23316 4764 23322
rect 4712 23258 4764 23264
rect 4436 23112 4488 23118
rect 4436 23054 4488 23060
rect 4158 22536 4214 22545
rect 4158 22471 4214 22480
rect 4172 21010 4200 22471
rect 4252 22228 4304 22234
rect 4252 22170 4304 22176
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 4172 18358 4200 20198
rect 4264 19922 4292 22170
rect 4252 19916 4304 19922
rect 4252 19858 4304 19864
rect 4344 18692 4396 18698
rect 4344 18634 4396 18640
rect 4160 18352 4212 18358
rect 4160 18294 4212 18300
rect 1766 18255 1822 18264
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 4252 18216 4304 18222
rect 4252 18158 4304 18164
rect 1398 17912 1454 17921
rect 1398 17847 1454 17856
rect 940 17604 992 17610
rect 940 17546 992 17552
rect 952 17105 980 17546
rect 1780 17513 1808 18158
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 1766 17504 1822 17513
rect 1766 17439 1822 17448
rect 1032 17128 1084 17134
rect 938 17096 994 17105
rect 1032 17070 1084 17076
rect 938 17031 994 17040
rect 1044 16697 1072 17070
rect 2136 17060 2188 17066
rect 2136 17002 2188 17008
rect 1030 16688 1086 16697
rect 1030 16623 1086 16632
rect 1032 16516 1084 16522
rect 1032 16458 1084 16464
rect 1044 16289 1072 16458
rect 1030 16280 1086 16289
rect 1030 16215 1086 16224
rect 1032 16040 1084 16046
rect 1032 15982 1084 15988
rect 1044 15881 1072 15982
rect 1030 15872 1086 15881
rect 1030 15807 1086 15816
rect 938 15464 994 15473
rect 938 15399 940 15408
rect 992 15399 994 15408
rect 940 15370 992 15376
rect 938 15056 994 15065
rect 938 14991 940 15000
rect 992 14991 994 15000
rect 940 14962 992 14968
rect 938 14648 994 14657
rect 938 14583 994 14592
rect 952 14482 980 14583
rect 940 14476 992 14482
rect 940 14418 992 14424
rect 1030 14240 1086 14249
rect 1030 14175 1086 14184
rect 1044 14006 1072 14175
rect 1032 14000 1084 14006
rect 1032 13942 1084 13948
rect 1766 13832 1822 13841
rect 1766 13767 1822 13776
rect 1780 13394 1808 13767
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1306 13016 1362 13025
rect 1306 12951 1362 12960
rect 1320 12918 1348 12951
rect 1308 12912 1360 12918
rect 1308 12854 1360 12860
rect 1216 12844 1268 12850
rect 1216 12786 1268 12792
rect 1228 12617 1256 12786
rect 1214 12608 1270 12617
rect 1214 12543 1270 12552
rect 1308 12300 1360 12306
rect 1308 12242 1360 12248
rect 1214 12200 1270 12209
rect 1214 12135 1270 12144
rect 1228 11762 1256 12135
rect 1320 11801 1348 12242
rect 1306 11792 1362 11801
rect 1216 11756 1268 11762
rect 1306 11727 1362 11736
rect 1216 11698 1268 11704
rect 1228 11354 1256 11698
rect 1308 11688 1360 11694
rect 1308 11630 1360 11636
rect 1320 11393 1348 11630
rect 1306 11384 1362 11393
rect 1216 11348 1268 11354
rect 1306 11319 1362 11328
rect 1216 11290 1268 11296
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1596 10985 1624 11086
rect 1582 10976 1638 10985
rect 1582 10911 1638 10920
rect 1216 10736 1268 10742
rect 1216 10678 1268 10684
rect 1228 10169 1256 10678
rect 1308 10668 1360 10674
rect 1308 10610 1360 10616
rect 1320 10577 1348 10610
rect 1306 10568 1362 10577
rect 1306 10503 1362 10512
rect 1214 10160 1270 10169
rect 2148 10130 2176 17002
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 4264 16114 4292 18158
rect 4356 17202 4384 18634
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4448 16726 4476 23054
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4632 21554 4660 22918
rect 4816 22710 4844 26200
rect 5460 23662 5488 26200
rect 5908 24812 5960 24818
rect 5908 24754 5960 24760
rect 5540 24064 5592 24070
rect 5540 24006 5592 24012
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5264 23248 5316 23254
rect 5264 23190 5316 23196
rect 4804 22704 4856 22710
rect 4804 22646 4856 22652
rect 4620 21548 4672 21554
rect 4620 21490 4672 21496
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 4816 20058 4844 20402
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 5276 19854 5304 23190
rect 5552 23118 5580 24006
rect 5816 23588 5868 23594
rect 5816 23530 5868 23536
rect 5724 23520 5776 23526
rect 5724 23462 5776 23468
rect 5632 23180 5684 23186
rect 5632 23122 5684 23128
rect 5356 23112 5408 23118
rect 5356 23054 5408 23060
rect 5540 23112 5592 23118
rect 5540 23054 5592 23060
rect 5368 22778 5396 23054
rect 5356 22772 5408 22778
rect 5356 22714 5408 22720
rect 5448 22500 5500 22506
rect 5448 22442 5500 22448
rect 5460 20466 5488 22442
rect 5644 21962 5672 23122
rect 5632 21956 5684 21962
rect 5632 21898 5684 21904
rect 5632 21480 5684 21486
rect 5632 21422 5684 21428
rect 5448 20460 5500 20466
rect 5448 20402 5500 20408
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 5354 18864 5410 18873
rect 5354 18799 5410 18808
rect 5368 18766 5396 18799
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 5644 18358 5672 21422
rect 5736 19922 5764 23462
rect 5828 21486 5856 23530
rect 5816 21480 5868 21486
rect 5816 21422 5868 21428
rect 5920 20398 5948 24754
rect 6000 23520 6052 23526
rect 6000 23462 6052 23468
rect 6012 22642 6040 23462
rect 6104 23186 6132 26200
rect 6748 24274 6776 26200
rect 6736 24268 6788 24274
rect 6736 24210 6788 24216
rect 7196 24200 7248 24206
rect 7196 24142 7248 24148
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 7208 22778 7236 24142
rect 7196 22772 7248 22778
rect 7196 22714 7248 22720
rect 7104 22704 7156 22710
rect 7104 22646 7156 22652
rect 6000 22636 6052 22642
rect 6000 22578 6052 22584
rect 6000 22432 6052 22438
rect 6000 22374 6052 22380
rect 6012 21010 6040 22374
rect 7116 22166 7144 22646
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 7104 22160 7156 22166
rect 7104 22102 7156 22108
rect 7208 22114 7236 22578
rect 7392 22574 7420 26200
rect 8036 24698 8064 26200
rect 7852 24670 8064 24698
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7484 22642 7512 24006
rect 7852 23186 7880 24670
rect 7930 24304 7986 24313
rect 8680 24274 8708 26200
rect 7930 24239 7986 24248
rect 8668 24268 8720 24274
rect 7944 24206 7972 24239
rect 8668 24210 8720 24216
rect 7932 24200 7984 24206
rect 7932 24142 7984 24148
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8484 23724 8536 23730
rect 8484 23666 8536 23672
rect 8392 23656 8444 23662
rect 8392 23598 8444 23604
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 7840 22160 7892 22166
rect 7208 22086 7328 22114
rect 7840 22102 7892 22108
rect 6736 22024 6788 22030
rect 6736 21966 6788 21972
rect 6748 21622 6776 21966
rect 6736 21616 6788 21622
rect 6550 21584 6606 21593
rect 6736 21558 6788 21564
rect 6550 21519 6552 21528
rect 6604 21519 6606 21528
rect 6644 21548 6696 21554
rect 6552 21490 6604 21496
rect 6644 21490 6696 21496
rect 6000 21004 6052 21010
rect 6000 20946 6052 20952
rect 6656 20602 6684 21490
rect 7300 20806 7328 22086
rect 7748 22024 7800 22030
rect 7748 21966 7800 21972
rect 7760 21010 7788 21966
rect 7748 21004 7800 21010
rect 7748 20946 7800 20952
rect 7288 20800 7340 20806
rect 7288 20742 7340 20748
rect 7564 20800 7616 20806
rect 7564 20742 7616 20748
rect 6644 20596 6696 20602
rect 6644 20538 6696 20544
rect 5908 20392 5960 20398
rect 5908 20334 5960 20340
rect 5724 19916 5776 19922
rect 5724 19858 5776 19864
rect 5908 19372 5960 19378
rect 5908 19314 5960 19320
rect 5920 19174 5948 19314
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 5632 18352 5684 18358
rect 5632 18294 5684 18300
rect 5920 17202 5948 19110
rect 6840 18970 6868 19246
rect 7576 19242 7604 20742
rect 7852 19514 7880 22102
rect 8404 21894 8432 23598
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8496 21298 8524 23666
rect 9140 23118 9168 24006
rect 9324 23746 9352 26200
rect 9772 24880 9824 24886
rect 9772 24822 9824 24828
rect 9588 24404 9640 24410
rect 9588 24346 9640 24352
rect 9232 23718 9352 23746
rect 9232 23662 9260 23718
rect 9220 23656 9272 23662
rect 9220 23598 9272 23604
rect 9128 23112 9180 23118
rect 9128 23054 9180 23060
rect 9220 22976 9272 22982
rect 9220 22918 9272 22924
rect 9128 22500 9180 22506
rect 9128 22442 9180 22448
rect 9140 22030 9168 22442
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 8956 21350 8984 21830
rect 9034 21584 9090 21593
rect 9034 21519 9036 21528
rect 9088 21519 9090 21528
rect 9036 21490 9088 21496
rect 8404 21270 8524 21298
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 8404 20942 8432 21270
rect 9232 21146 9260 22918
rect 9600 21690 9628 24346
rect 9784 22098 9812 24822
rect 9968 22710 9996 26200
rect 10140 24132 10192 24138
rect 10140 24074 10192 24080
rect 9956 22704 10008 22710
rect 9956 22646 10008 22652
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9772 22092 9824 22098
rect 10152 22094 10180 24074
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 10232 22160 10284 22166
rect 10232 22102 10284 22108
rect 9772 22034 9824 22040
rect 10060 22066 10180 22094
rect 9588 21684 9640 21690
rect 9588 21626 9640 21632
rect 9128 21140 9180 21146
rect 9128 21082 9180 21088
rect 9220 21140 9272 21146
rect 9220 21082 9272 21088
rect 8392 20936 8444 20942
rect 8390 20904 8392 20913
rect 8444 20904 8446 20913
rect 8390 20839 8446 20848
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 7564 19236 7616 19242
rect 7564 19178 7616 19184
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 4436 16720 4488 16726
rect 4436 16662 4488 16668
rect 5448 16720 5500 16726
rect 5448 16662 5500 16668
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 4160 15428 4212 15434
rect 4160 15370 4212 15376
rect 4172 15026 4200 15370
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 3528 13433 3556 13874
rect 3514 13424 3570 13433
rect 3514 13359 3570 13368
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 4264 12434 4292 16050
rect 5460 12986 5488 16662
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 4172 12406 4292 12434
rect 2504 11824 2556 11830
rect 2504 11766 2556 11772
rect 2686 11792 2742 11801
rect 2516 10810 2544 11766
rect 2686 11727 2742 11736
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 1214 10095 1270 10104
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 1306 9752 1362 9761
rect 2424 9722 2452 9998
rect 1306 9687 1308 9696
rect 1360 9687 1362 9696
rect 2412 9716 2464 9722
rect 1308 9658 1360 9664
rect 2412 9658 2464 9664
rect 1308 9580 1360 9586
rect 1308 9522 1360 9528
rect 1320 9353 1348 9522
rect 1766 9480 1822 9489
rect 1766 9415 1768 9424
rect 1820 9415 1822 9424
rect 1768 9386 1820 9392
rect 1306 9344 1362 9353
rect 1306 9279 1362 9288
rect 1216 8968 1268 8974
rect 1216 8910 1268 8916
rect 1306 8936 1362 8945
rect 1228 8537 1256 8910
rect 1306 8871 1308 8880
rect 1360 8871 1362 8880
rect 1308 8842 1360 8848
rect 1214 8528 1270 8537
rect 2700 8498 2728 11727
rect 4172 11558 4200 12406
rect 5920 12238 5948 17138
rect 7852 16522 7880 19450
rect 8312 19174 8340 20470
rect 9140 19378 9168 21082
rect 9692 20602 9720 22034
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9220 19440 9272 19446
rect 9220 19382 9272 19388
rect 9128 19372 9180 19378
rect 9128 19314 9180 19320
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 7840 16516 7892 16522
rect 7840 16458 7892 16464
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8312 16250 8340 19110
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 9048 16454 9076 16526
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 9048 16046 9076 16390
rect 9232 16250 9260 19382
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 9048 15366 9076 15982
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 9048 13258 9076 15302
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 9508 12782 9536 16934
rect 9600 16017 9628 19790
rect 9692 18086 9720 20402
rect 9968 19990 9996 21490
rect 9956 19984 10008 19990
rect 9956 19926 10008 19932
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9876 18426 9904 19246
rect 9864 18420 9916 18426
rect 9864 18362 9916 18368
rect 9772 18352 9824 18358
rect 9772 18294 9824 18300
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 9586 16008 9642 16017
rect 9586 15943 9642 15952
rect 9692 15162 9720 16458
rect 9784 16250 9812 18294
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9876 17202 9904 17750
rect 9968 17202 9996 19926
rect 10060 18154 10088 22066
rect 10244 21010 10272 22102
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 10336 20602 10364 23802
rect 10612 23662 10640 26200
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 10600 23656 10652 23662
rect 10600 23598 10652 23604
rect 11164 22642 11192 24006
rect 11256 23186 11284 26200
rect 11900 24342 11928 26200
rect 12348 24404 12400 24410
rect 12348 24346 12400 24352
rect 11888 24336 11940 24342
rect 11888 24278 11940 24284
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11808 23798 11836 24006
rect 11796 23792 11848 23798
rect 11796 23734 11848 23740
rect 12360 23730 12388 24346
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12348 23724 12400 23730
rect 12348 23666 12400 23672
rect 11244 23180 11296 23186
rect 11244 23122 11296 23128
rect 11888 23112 11940 23118
rect 11334 23080 11390 23089
rect 11888 23054 11940 23060
rect 11334 23015 11390 23024
rect 11152 22636 11204 22642
rect 11152 22578 11204 22584
rect 11060 22500 11112 22506
rect 11060 22442 11112 22448
rect 11072 22094 11100 22442
rect 11072 22066 11284 22094
rect 10968 21616 11020 21622
rect 10968 21558 11020 21564
rect 10876 21344 10928 21350
rect 10876 21286 10928 21292
rect 10600 20800 10652 20806
rect 10600 20742 10652 20748
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10612 19990 10640 20742
rect 10704 20641 10732 20742
rect 10690 20632 10746 20641
rect 10690 20567 10746 20576
rect 10888 20466 10916 21286
rect 10980 20534 11008 21558
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 10968 20528 11020 20534
rect 10968 20470 11020 20476
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10600 19984 10652 19990
rect 10600 19926 10652 19932
rect 10612 19689 10640 19926
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 10598 19680 10654 19689
rect 10598 19615 10654 19624
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 10140 18692 10192 18698
rect 10232 18692 10284 18698
rect 10192 18652 10232 18680
rect 10140 18634 10192 18640
rect 10232 18634 10284 18640
rect 10692 18692 10744 18698
rect 10692 18634 10744 18640
rect 10048 18148 10100 18154
rect 10048 18090 10100 18096
rect 10152 17882 10180 18634
rect 10416 18624 10468 18630
rect 10416 18566 10468 18572
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10152 17610 10180 17818
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 10140 17604 10192 17610
rect 10140 17546 10192 17552
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 10244 16726 10272 17614
rect 10428 17270 10456 18566
rect 10598 17776 10654 17785
rect 10598 17711 10654 17720
rect 10416 17264 10468 17270
rect 10416 17206 10468 17212
rect 10612 17134 10640 17711
rect 10600 17128 10652 17134
rect 10520 17076 10600 17082
rect 10520 17070 10652 17076
rect 10520 17054 10640 17070
rect 10520 16998 10548 17054
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10232 16720 10284 16726
rect 10232 16662 10284 16668
rect 10508 16516 10560 16522
rect 10508 16458 10560 16464
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 10520 16153 10548 16458
rect 10506 16144 10562 16153
rect 10506 16079 10562 16088
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9784 15162 9812 15914
rect 10612 15910 10640 16934
rect 10704 16266 10732 18634
rect 10888 16658 10916 18906
rect 10980 18222 11008 19790
rect 11072 18902 11100 20742
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 11060 18896 11112 18902
rect 11060 18838 11112 18844
rect 10968 18216 11020 18222
rect 11164 18193 11192 19314
rect 11256 18873 11284 22066
rect 11348 20942 11376 23015
rect 11796 22568 11848 22574
rect 11796 22510 11848 22516
rect 11808 22114 11836 22510
rect 11900 22234 11928 23054
rect 12072 22432 12124 22438
rect 12072 22374 12124 22380
rect 11888 22228 11940 22234
rect 11888 22170 11940 22176
rect 11886 22128 11942 22137
rect 11808 22086 11886 22114
rect 11886 22063 11888 22072
rect 11940 22063 11942 22072
rect 12084 22094 12112 22374
rect 12084 22066 12204 22094
rect 11888 22034 11940 22040
rect 12176 21554 12204 22066
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 11428 21480 11480 21486
rect 11704 21480 11756 21486
rect 11428 21422 11480 21428
rect 11702 21448 11704 21457
rect 11756 21448 11758 21457
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11440 19786 11468 21422
rect 11702 21383 11758 21392
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11808 20466 11836 21286
rect 12084 20874 12112 21490
rect 12176 21026 12204 21490
rect 12452 21434 12480 21626
rect 12360 21406 12480 21434
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12268 21146 12296 21286
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 12176 20998 12296 21026
rect 12072 20868 12124 20874
rect 12072 20810 12124 20816
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 11992 19922 12020 19994
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 12084 19825 12112 20810
rect 12070 19816 12126 19825
rect 11428 19780 11480 19786
rect 12070 19751 12126 19760
rect 11428 19722 11480 19728
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 12072 19236 12124 19242
rect 12072 19178 12124 19184
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11900 18970 11928 19110
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 11242 18864 11298 18873
rect 11242 18799 11298 18808
rect 11520 18624 11572 18630
rect 11520 18566 11572 18572
rect 11532 18358 11560 18566
rect 11244 18352 11296 18358
rect 11244 18294 11296 18300
rect 11520 18352 11572 18358
rect 11520 18294 11572 18300
rect 10968 18158 11020 18164
rect 11150 18184 11206 18193
rect 10980 17882 11008 18158
rect 11150 18119 11206 18128
rect 10968 17876 11020 17882
rect 10968 17818 11020 17824
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 10704 16250 11100 16266
rect 10704 16244 11112 16250
rect 10704 16238 11060 16244
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 9784 12170 9812 14894
rect 9876 14074 9904 15846
rect 10704 15706 10732 16238
rect 11060 16186 11112 16192
rect 10876 16176 10928 16182
rect 10876 16118 10928 16124
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10244 14550 10272 15438
rect 10888 15094 10916 16118
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 11072 15094 11100 15506
rect 11164 15502 11192 17478
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11164 15094 11192 15438
rect 10876 15088 10928 15094
rect 10876 15030 10928 15036
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 11072 14890 11100 15030
rect 11060 14884 11112 14890
rect 11060 14826 11112 14832
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10232 14544 10284 14550
rect 10232 14486 10284 14492
rect 10414 14512 10470 14521
rect 10704 14482 10732 14758
rect 10414 14447 10470 14456
rect 10692 14476 10744 14482
rect 10428 14414 10456 14447
rect 10692 14418 10744 14424
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 9968 14074 9996 14282
rect 10428 14074 10456 14350
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10520 14006 10548 14214
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10508 13456 10560 13462
rect 10508 13398 10560 13404
rect 10520 12170 10548 13398
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 10520 11898 10548 12106
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 1214 8463 1270 8472
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 1306 8120 1362 8129
rect 2424 8090 2452 8366
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 1306 8055 1308 8064
rect 1360 8055 1362 8064
rect 2412 8084 2464 8090
rect 1308 8026 1360 8032
rect 2412 8026 2464 8032
rect 1308 7880 1360 7886
rect 1308 7822 1360 7828
rect 1320 7721 1348 7822
rect 1306 7712 1362 7721
rect 1306 7647 1362 7656
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 1308 7404 1360 7410
rect 1308 7346 1360 7352
rect 1320 7313 1348 7346
rect 1306 7304 1362 7313
rect 1306 7239 1362 7248
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 10704 6914 10732 14418
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 10796 13394 10824 13670
rect 11164 13394 11192 15030
rect 11256 14618 11284 18294
rect 11796 18284 11848 18290
rect 12084 18272 12112 19178
rect 12176 18698 12204 19314
rect 12164 18692 12216 18698
rect 12164 18634 12216 18640
rect 12164 18284 12216 18290
rect 12084 18244 12164 18272
rect 11796 18226 11848 18232
rect 12164 18226 12216 18232
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11440 17270 11468 17682
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11336 16448 11388 16454
rect 11336 16390 11388 16396
rect 11348 16250 11376 16390
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11532 15706 11560 15846
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 11256 14006 11284 14282
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11256 13841 11284 13942
rect 11242 13832 11298 13841
rect 11242 13767 11298 13776
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 10796 12306 10824 13330
rect 11164 13258 11192 13330
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 11150 13152 11206 13161
rect 10980 12986 11008 13126
rect 11150 13087 11206 13096
rect 11164 12986 11192 13087
rect 11348 12986 11376 15098
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 11072 11218 11100 12106
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 11072 9518 11100 11154
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 1214 6896 1270 6905
rect 1214 6831 1270 6840
rect 10612 6886 10732 6914
rect 1228 6730 1256 6831
rect 1308 6792 1360 6798
rect 1308 6734 1360 6740
rect 1216 6724 1268 6730
rect 1216 6666 1268 6672
rect 1228 6458 1256 6666
rect 1320 6497 1348 6734
rect 10612 6730 10640 6886
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 1768 6656 1820 6662
rect 1768 6598 1820 6604
rect 1306 6488 1362 6497
rect 1216 6452 1268 6458
rect 1306 6423 1362 6432
rect 1216 6394 1268 6400
rect 1780 6390 1808 6598
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 1768 6384 1820 6390
rect 1768 6326 1820 6332
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 1320 6089 1348 6258
rect 11256 6186 11284 12582
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11348 11150 11376 11834
rect 11532 11626 11560 15642
rect 11808 15162 11836 18226
rect 12072 18148 12124 18154
rect 12072 18090 12124 18096
rect 12084 17610 12112 18090
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 11888 17264 11940 17270
rect 11888 17206 11940 17212
rect 11900 17105 11928 17206
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 11886 17096 11942 17105
rect 11886 17031 11942 17040
rect 11992 16998 12020 17138
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11900 14074 11928 15302
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11808 12442 11836 12718
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11808 11694 11836 12378
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11808 11218 11836 11630
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11348 10810 11376 11086
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11992 8974 12020 16390
rect 12084 14890 12112 17546
rect 12268 17241 12296 20998
rect 12360 20534 12388 21406
rect 12348 20528 12400 20534
rect 12348 20470 12400 20476
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 12360 19938 12388 20334
rect 12360 19910 12480 19938
rect 12452 19258 12480 19910
rect 12360 19230 12480 19258
rect 12360 18970 12388 19230
rect 12544 19224 12572 21966
rect 12636 21622 12664 24074
rect 12716 23724 12768 23730
rect 12716 23666 12768 23672
rect 12624 21616 12676 21622
rect 12624 21558 12676 21564
rect 12624 21480 12676 21486
rect 12624 21422 12676 21428
rect 12636 21049 12664 21422
rect 12622 21040 12678 21049
rect 12728 21010 12756 23666
rect 12820 22710 12848 26302
rect 13174 26302 13400 26330
rect 13174 26200 13230 26302
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13372 23186 13400 26302
rect 13818 26200 13874 27000
rect 14462 26200 14518 27000
rect 15106 26200 15162 27000
rect 15750 26200 15806 27000
rect 16394 26200 16450 27000
rect 17038 26200 17094 27000
rect 17682 26200 17738 27000
rect 18326 26200 18382 27000
rect 18970 26200 19026 27000
rect 19614 26200 19670 27000
rect 20258 26200 20314 27000
rect 20902 26200 20958 27000
rect 21546 26200 21602 27000
rect 22190 26200 22246 27000
rect 22834 26200 22890 27000
rect 23478 26200 23534 27000
rect 24122 26200 24178 27000
rect 24766 26200 24822 27000
rect 25410 26200 25466 27000
rect 26054 26330 26110 27000
rect 26698 26330 26754 27000
rect 26054 26302 26188 26330
rect 26054 26200 26110 26302
rect 13832 24274 13860 26200
rect 14476 24290 14504 26200
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 14384 24262 14504 24290
rect 14280 24200 14332 24206
rect 14280 24142 14332 24148
rect 14188 23792 14240 23798
rect 14188 23734 14240 23740
rect 14200 23254 14228 23734
rect 14188 23248 14240 23254
rect 14188 23190 14240 23196
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 12808 22704 12860 22710
rect 12808 22646 12860 22652
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12808 21480 12860 21486
rect 12808 21422 12860 21428
rect 12820 21146 12848 21422
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12808 21140 12860 21146
rect 12808 21082 12860 21088
rect 12622 20975 12678 20984
rect 12716 21004 12768 21010
rect 12716 20946 12768 20952
rect 12624 20936 12676 20942
rect 12676 20884 12756 20890
rect 12624 20878 12756 20884
rect 12636 20862 12756 20878
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12636 19334 12664 20742
rect 12728 20602 12756 20862
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12820 20058 12848 21082
rect 12898 21040 12954 21049
rect 12898 20975 12954 20984
rect 12912 20466 12940 20975
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 13360 20256 13412 20262
rect 13360 20198 13412 20204
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12808 20052 12860 20058
rect 12808 19994 12860 20000
rect 13372 19854 13400 20198
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13464 19666 13492 22578
rect 13832 21690 13860 23054
rect 13912 22500 13964 22506
rect 13912 22442 13964 22448
rect 13820 21684 13872 21690
rect 13820 21626 13872 21632
rect 13924 21486 13952 22442
rect 14188 22160 14240 22166
rect 14188 22102 14240 22108
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13912 21480 13964 21486
rect 13912 21422 13964 21428
rect 13728 21412 13780 21418
rect 13728 21354 13780 21360
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13372 19638 13492 19666
rect 12808 19440 12860 19446
rect 12808 19382 12860 19388
rect 12636 19310 12756 19334
rect 12636 19306 12768 19310
rect 12716 19304 12768 19306
rect 12716 19246 12768 19252
rect 12544 19196 12664 19224
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 12452 18850 12480 19110
rect 12360 18822 12480 18850
rect 12532 18828 12584 18834
rect 12360 18034 12388 18822
rect 12532 18770 12584 18776
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12452 18426 12480 18702
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12360 18006 12480 18034
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12360 17270 12388 17818
rect 12348 17264 12400 17270
rect 12254 17232 12310 17241
rect 12348 17206 12400 17212
rect 12254 17167 12310 17176
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12360 16232 12388 17070
rect 12452 16726 12480 18006
rect 12544 17746 12572 18770
rect 12636 17882 12664 19196
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12728 18834 12756 19110
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12820 18766 12848 19382
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 13372 18902 13400 19638
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 13360 18896 13412 18902
rect 13360 18838 13412 18844
rect 13176 18828 13228 18834
rect 13176 18770 13228 18776
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 13188 18358 13216 18770
rect 13176 18352 13228 18358
rect 13176 18294 13228 18300
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 13372 17762 13400 18838
rect 13464 18290 13492 19450
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 13280 17734 13400 17762
rect 13464 17746 13492 18226
rect 13452 17740 13504 17746
rect 12440 16720 12492 16726
rect 12440 16662 12492 16668
rect 12360 16204 12480 16232
rect 12164 16108 12216 16114
rect 12164 16050 12216 16056
rect 12072 14884 12124 14890
rect 12072 14826 12124 14832
rect 12176 12753 12204 16050
rect 12256 15020 12308 15026
rect 12256 14962 12308 14968
rect 12268 14482 12296 14962
rect 12348 14952 12400 14958
rect 12346 14920 12348 14929
rect 12400 14920 12402 14929
rect 12346 14855 12402 14864
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12268 13530 12296 13806
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12162 12744 12218 12753
rect 12162 12679 12218 12688
rect 12268 12102 12296 13466
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12360 11762 12388 13738
rect 12452 12986 12480 16204
rect 12544 15570 12572 17682
rect 13280 17270 13308 17734
rect 13452 17682 13504 17688
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 12716 17060 12768 17066
rect 12716 17002 12768 17008
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12636 14618 12664 16458
rect 12728 15502 12756 17002
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12820 16674 12848 16934
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12820 16646 12940 16674
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 12820 15366 12848 16526
rect 12912 16454 12940 16646
rect 12900 16448 12952 16454
rect 12900 16390 12952 16396
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 13372 15042 13400 17614
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13464 15502 13492 16934
rect 13556 16590 13584 20742
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 13648 19718 13676 19858
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13740 18154 13768 21354
rect 13912 20528 13964 20534
rect 13912 20470 13964 20476
rect 13820 19780 13872 19786
rect 13820 19722 13872 19728
rect 13832 18902 13860 19722
rect 13820 18896 13872 18902
rect 13820 18838 13872 18844
rect 13924 18358 13952 20470
rect 13912 18352 13964 18358
rect 13912 18294 13964 18300
rect 13728 18148 13780 18154
rect 13728 18090 13780 18096
rect 13636 18080 13688 18086
rect 13636 18022 13688 18028
rect 13648 17542 13676 18022
rect 13636 17536 13688 17542
rect 13688 17496 13768 17524
rect 13636 17478 13688 17484
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13544 16448 13596 16454
rect 13542 16416 13544 16425
rect 13636 16448 13688 16454
rect 13596 16416 13598 16425
rect 13636 16390 13688 16396
rect 13542 16351 13598 16360
rect 13648 16250 13676 16390
rect 13636 16244 13688 16250
rect 13636 16186 13688 16192
rect 13636 16040 13688 16046
rect 13542 16008 13598 16017
rect 13636 15982 13688 15988
rect 13542 15943 13544 15952
rect 13596 15943 13598 15952
rect 13544 15914 13596 15920
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13372 15014 13492 15042
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12624 14612 12676 14618
rect 12820 14600 12848 14758
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 12820 14572 12940 14600
rect 12624 14554 12676 14560
rect 12808 14340 12860 14346
rect 12808 14282 12860 14288
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12728 13172 12756 14214
rect 12820 13376 12848 14282
rect 12912 14074 12940 14572
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 13280 14006 13308 14418
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13280 13818 13308 13942
rect 13280 13790 13400 13818
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 12900 13388 12952 13394
rect 12820 13348 12900 13376
rect 12900 13330 12952 13336
rect 13004 13258 13032 13466
rect 12992 13252 13044 13258
rect 12992 13194 13044 13200
rect 12728 13144 12848 13172
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12452 12209 12480 12922
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12438 12200 12494 12209
rect 12438 12135 12494 12144
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12268 10470 12296 10610
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11244 6180 11296 6186
rect 11244 6122 11296 6128
rect 1306 6080 1362 6089
rect 1306 6015 1362 6024
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 1308 5704 1360 5710
rect 1306 5672 1308 5681
rect 2780 5704 2832 5710
rect 1360 5672 1362 5681
rect 2780 5646 2832 5652
rect 1306 5607 1362 5616
rect 2792 5273 2820 5646
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 2778 5264 2834 5273
rect 2778 5199 2834 5208
rect 1308 5160 1360 5166
rect 1308 5102 1360 5108
rect 1320 4865 1348 5102
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 1306 4856 1362 4865
rect 2950 4859 3258 4868
rect 1306 4791 1308 4800
rect 1360 4791 1362 4800
rect 1308 4762 1360 4768
rect 1308 4616 1360 4622
rect 1308 4558 1360 4564
rect 1320 4457 1348 4558
rect 1306 4448 1362 4457
rect 1306 4383 1362 4392
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 1400 4208 1452 4214
rect 1400 4150 1452 4156
rect 1412 4049 1440 4150
rect 1398 4040 1454 4049
rect 1308 4004 1360 4010
rect 1398 3975 1454 3984
rect 5354 4040 5410 4049
rect 5354 3975 5410 3984
rect 1308 3946 1360 3952
rect 1320 3641 1348 3946
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 3332 3664 3384 3670
rect 1306 3632 1362 3641
rect 3332 3606 3384 3612
rect 1306 3567 1362 3576
rect 1308 3528 1360 3534
rect 1122 3496 1178 3505
rect 1308 3470 1360 3476
rect 1122 3431 1178 3440
rect 1136 800 1164 3431
rect 1320 3233 1348 3470
rect 1306 3224 1362 3233
rect 1306 3159 1308 3168
rect 1360 3159 1362 3168
rect 1308 3130 1360 3136
rect 1308 3052 1360 3058
rect 1308 2994 1360 3000
rect 1320 2825 1348 2994
rect 2320 2848 2372 2854
rect 1306 2816 1362 2825
rect 2320 2790 2372 2796
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 1306 2751 1362 2760
rect 1308 2440 1360 2446
rect 1306 2408 1308 2417
rect 1360 2408 1362 2417
rect 1216 2372 1268 2378
rect 2332 2378 2360 2790
rect 2792 2446 2820 2790
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 1306 2343 1362 2352
rect 2320 2372 2372 2378
rect 1216 2314 1268 2320
rect 2320 2314 2372 2320
rect 1228 2009 1256 2314
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1214 2000 1270 2009
rect 1214 1935 1270 1944
rect 1320 1601 1348 2246
rect 3344 1850 3372 3606
rect 3252 1822 3372 1850
rect 1306 1592 1362 1601
rect 1306 1527 1362 1536
rect 3252 800 3280 1822
rect 5368 800 5396 3975
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7484 800 7512 3674
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9692 2582 9720 2994
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 12268 2514 12296 10406
rect 12360 9586 12388 11494
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12452 3602 12480 9862
rect 12544 9450 12572 12582
rect 12820 10810 12848 13144
rect 13372 13138 13400 13790
rect 13280 13110 13400 13138
rect 13280 12986 13308 13110
rect 13268 12980 13320 12986
rect 13464 12968 13492 15014
rect 13268 12922 13320 12928
rect 13372 12940 13492 12968
rect 13372 12730 13400 12940
rect 13372 12702 13492 12730
rect 13358 12608 13414 12617
rect 12950 12540 13258 12549
rect 13358 12543 13414 12552
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13372 12434 13400 12543
rect 13280 12406 13400 12434
rect 13280 11626 13308 12406
rect 13464 12102 13492 12702
rect 13452 12096 13504 12102
rect 13358 12064 13414 12073
rect 13452 12038 13504 12044
rect 13358 11999 13414 12008
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13372 11558 13400 11999
rect 13556 11898 13584 15302
rect 13648 14482 13676 15982
rect 13740 15144 13768 17496
rect 14016 17338 14044 21490
rect 14094 20632 14150 20641
rect 14094 20567 14096 20576
rect 14148 20567 14150 20576
rect 14096 20538 14148 20544
rect 14200 19854 14228 22102
rect 14292 22098 14320 24142
rect 14384 23798 14412 24262
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 14372 23792 14424 23798
rect 14372 23734 14424 23740
rect 14372 22976 14424 22982
rect 14372 22918 14424 22924
rect 14384 22438 14412 22918
rect 14372 22432 14424 22438
rect 14372 22374 14424 22380
rect 14384 22166 14412 22374
rect 14372 22160 14424 22166
rect 14372 22102 14424 22108
rect 14280 22092 14332 22098
rect 14280 22034 14332 22040
rect 14280 21616 14332 21622
rect 14280 21558 14332 21564
rect 14292 21146 14320 21558
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14384 21146 14412 21490
rect 14280 21140 14332 21146
rect 14280 21082 14332 21088
rect 14372 21140 14424 21146
rect 14372 21082 14424 21088
rect 14292 20398 14320 21082
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14476 20058 14504 24142
rect 14924 24132 14976 24138
rect 14924 24074 14976 24080
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14660 22642 14688 22918
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14200 19446 14228 19790
rect 14188 19440 14240 19446
rect 14188 19382 14240 19388
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14108 18329 14136 18566
rect 14094 18320 14150 18329
rect 14094 18255 14150 18264
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 13832 16726 13860 17274
rect 14108 17270 14136 18255
rect 14096 17264 14148 17270
rect 14096 17206 14148 17212
rect 14292 17134 14320 19790
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14568 18222 14596 18634
rect 14556 18216 14608 18222
rect 14556 18158 14608 18164
rect 14568 17882 14596 18158
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14200 16794 14228 16934
rect 14660 16794 14688 21898
rect 14936 20602 14964 24074
rect 15120 22710 15148 26200
rect 15476 24336 15528 24342
rect 15476 24278 15528 24284
rect 15108 22704 15160 22710
rect 15108 22646 15160 22652
rect 15200 22704 15252 22710
rect 15200 22646 15252 22652
rect 15108 22160 15160 22166
rect 15108 22102 15160 22108
rect 15120 21978 15148 22102
rect 15212 22098 15240 22646
rect 15200 22092 15252 22098
rect 15200 22034 15252 22040
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 15120 21950 15240 21978
rect 15212 21486 15240 21950
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 15212 20874 15240 21422
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15200 20868 15252 20874
rect 15200 20810 15252 20816
rect 14924 20596 14976 20602
rect 14924 20538 14976 20544
rect 15016 20460 15068 20466
rect 15016 20402 15068 20408
rect 14924 20324 14976 20330
rect 14924 20266 14976 20272
rect 14936 19990 14964 20266
rect 14924 19984 14976 19990
rect 14924 19926 14976 19932
rect 15028 19514 15056 20402
rect 15016 19508 15068 19514
rect 15016 19450 15068 19456
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 15120 18970 15148 19110
rect 15212 18970 15240 19246
rect 15108 18964 15160 18970
rect 15108 18906 15160 18912
rect 15200 18964 15252 18970
rect 15200 18906 15252 18912
rect 14830 18728 14886 18737
rect 14752 18672 14830 18680
rect 14752 18652 14832 18672
rect 14752 17746 14780 18652
rect 14884 18663 14886 18672
rect 14832 18634 14884 18640
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14740 17264 14792 17270
rect 14740 17206 14792 17212
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 13820 16720 13872 16726
rect 13820 16662 13872 16668
rect 14752 16454 14780 17206
rect 14844 16454 14872 18226
rect 15014 18184 15070 18193
rect 15304 18154 15332 21082
rect 15396 19378 15424 22034
rect 15488 20602 15516 24278
rect 15764 23186 15792 26200
rect 16028 24336 16080 24342
rect 16028 24278 16080 24284
rect 15844 23316 15896 23322
rect 15844 23258 15896 23264
rect 15752 23180 15804 23186
rect 15752 23122 15804 23128
rect 15752 22772 15804 22778
rect 15752 22714 15804 22720
rect 15660 22160 15712 22166
rect 15660 22102 15712 22108
rect 15566 21584 15622 21593
rect 15566 21519 15622 21528
rect 15476 20596 15528 20602
rect 15476 20538 15528 20544
rect 15580 20262 15608 21519
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15474 19952 15530 19961
rect 15474 19887 15530 19896
rect 15488 19378 15516 19887
rect 15580 19854 15608 20198
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15476 19372 15528 19378
rect 15476 19314 15528 19320
rect 15014 18119 15070 18128
rect 15292 18148 15344 18154
rect 14924 16584 14976 16590
rect 14924 16526 14976 16532
rect 14188 16448 14240 16454
rect 14002 16416 14058 16425
rect 14188 16390 14240 16396
rect 14740 16448 14792 16454
rect 14832 16448 14884 16454
rect 14740 16390 14792 16396
rect 14830 16416 14832 16425
rect 14884 16416 14886 16425
rect 14002 16351 14058 16360
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 13740 15116 13860 15144
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13740 14006 13768 14962
rect 13832 14958 13860 15116
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13728 14000 13780 14006
rect 13728 13942 13780 13948
rect 13740 13870 13768 13942
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13648 12986 13676 13670
rect 13728 13524 13780 13530
rect 13832 13512 13860 14350
rect 13780 13484 13860 13512
rect 13728 13466 13780 13472
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13740 12617 13768 13466
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13832 13190 13860 13330
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13726 12608 13782 12617
rect 13726 12543 13782 12552
rect 13832 12458 13860 13126
rect 13924 12782 13952 15302
rect 14016 14618 14044 16351
rect 14200 16153 14228 16390
rect 14830 16351 14886 16360
rect 14186 16144 14242 16153
rect 14554 16144 14610 16153
rect 14186 16079 14242 16088
rect 14464 16108 14516 16114
rect 14554 16079 14610 16088
rect 14464 16050 14516 16056
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14292 15638 14320 15982
rect 14280 15632 14332 15638
rect 14280 15574 14332 15580
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 13740 12430 13860 12458
rect 13636 12164 13688 12170
rect 13636 12106 13688 12112
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13648 11694 13676 12106
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12912 11082 12940 11154
rect 12900 11076 12952 11082
rect 12900 11018 12952 11024
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12912 10690 12940 11018
rect 12820 10662 12940 10690
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 12728 2922 12756 10406
rect 12820 5234 12848 10662
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 13372 5846 13400 11494
rect 13464 11082 13492 11630
rect 13544 11620 13596 11626
rect 13544 11562 13596 11568
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13464 10985 13492 11018
rect 13450 10976 13506 10985
rect 13450 10911 13506 10920
rect 13452 10600 13504 10606
rect 13450 10568 13452 10577
rect 13504 10568 13506 10577
rect 13450 10503 13506 10512
rect 13556 8634 13584 11562
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13648 9382 13676 11086
rect 13740 9654 13768 12430
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13832 11626 13860 12310
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 13832 10606 13860 11562
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13924 10538 13952 11630
rect 14016 11354 14044 14214
rect 14108 13190 14136 15506
rect 14292 14958 14320 15574
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14200 14278 14228 14894
rect 14292 14822 14320 14894
rect 14476 14822 14504 16050
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14568 14498 14596 16079
rect 14936 16046 14964 16526
rect 15028 16182 15056 18119
rect 15292 18090 15344 18096
rect 15108 18080 15160 18086
rect 15160 18040 15240 18068
rect 15108 18022 15160 18028
rect 15212 17882 15240 18040
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15396 17746 15424 19314
rect 15488 19242 15516 19314
rect 15476 19236 15528 19242
rect 15476 19178 15528 19184
rect 15672 18902 15700 22102
rect 15764 19310 15792 22714
rect 15856 20602 15884 23258
rect 16040 20602 16068 24278
rect 16408 23662 16436 26200
rect 16396 23656 16448 23662
rect 16396 23598 16448 23604
rect 16580 23044 16632 23050
rect 16580 22986 16632 22992
rect 16120 21956 16172 21962
rect 16120 21898 16172 21904
rect 16132 21622 16160 21898
rect 16120 21616 16172 21622
rect 16120 21558 16172 21564
rect 16304 21140 16356 21146
rect 16304 21082 16356 21088
rect 16120 20868 16172 20874
rect 16120 20810 16172 20816
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 15936 19712 15988 19718
rect 15842 19680 15898 19689
rect 16132 19666 16160 20810
rect 16210 20360 16266 20369
rect 16210 20295 16266 20304
rect 15988 19660 16160 19666
rect 15936 19654 16160 19660
rect 15948 19638 16160 19654
rect 15842 19615 15898 19624
rect 15752 19304 15804 19310
rect 15752 19246 15804 19252
rect 15660 18896 15712 18902
rect 15660 18838 15712 18844
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15384 17740 15436 17746
rect 15304 17700 15384 17728
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15120 16697 15148 17138
rect 15106 16688 15162 16697
rect 15106 16623 15162 16632
rect 15304 16436 15332 17700
rect 15384 17682 15436 17688
rect 15580 17338 15608 18566
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15764 17270 15792 17818
rect 15752 17264 15804 17270
rect 15752 17206 15804 17212
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15120 16408 15332 16436
rect 15016 16176 15068 16182
rect 15016 16118 15068 16124
rect 14924 16040 14976 16046
rect 14844 16000 14924 16028
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14660 14618 14688 15302
rect 14844 15094 14872 16000
rect 14924 15982 14976 15988
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 14832 15088 14884 15094
rect 14752 15056 14832 15076
rect 14884 15056 14886 15065
rect 14752 15048 14830 15056
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14384 14470 14596 14498
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14200 13530 14228 14010
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14108 12442 14136 13126
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 14292 11898 14320 14010
rect 14280 11892 14332 11898
rect 14384 11880 14412 14470
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14476 12918 14504 13806
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 14554 13424 14610 13433
rect 14554 13359 14610 13368
rect 14568 13326 14596 13359
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14568 13161 14596 13262
rect 14554 13152 14610 13161
rect 14554 13087 14610 13096
rect 14464 12912 14516 12918
rect 14464 12854 14516 12860
rect 14476 12170 14504 12854
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14568 12442 14596 12718
rect 14556 12436 14608 12442
rect 14556 12378 14608 12384
rect 14660 12288 14688 13670
rect 14752 12374 14780 15048
rect 14830 14991 14886 15000
rect 14832 14476 14884 14482
rect 14832 14418 14884 14424
rect 14844 13394 14872 14418
rect 14832 13388 14884 13394
rect 14832 13330 14884 13336
rect 14844 13025 14872 13330
rect 14936 13258 14964 15506
rect 15120 15026 15148 16408
rect 15396 16114 15424 16594
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 15384 16108 15436 16114
rect 15384 16050 15436 16056
rect 15304 15706 15332 16050
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 15304 15026 15332 15642
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15304 14006 15332 14962
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15396 14482 15424 14894
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15016 14000 15068 14006
rect 15016 13942 15068 13948
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15028 13530 15056 13942
rect 15120 13802 15332 13818
rect 15120 13796 15344 13802
rect 15120 13790 15292 13796
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 15120 13410 15148 13790
rect 15292 13738 15344 13744
rect 15028 13382 15148 13410
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 14830 13016 14886 13025
rect 14830 12951 14886 12960
rect 14740 12368 14792 12374
rect 14740 12310 14792 12316
rect 14568 12260 14688 12288
rect 14464 12164 14516 12170
rect 14464 12106 14516 12112
rect 14384 11852 14504 11880
rect 14280 11834 14332 11840
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 14384 10810 14412 11698
rect 14476 11286 14504 11852
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14568 10742 14596 12260
rect 14752 11830 14780 12310
rect 14740 11824 14792 11830
rect 14740 11766 14792 11772
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14556 10736 14608 10742
rect 14556 10678 14608 10684
rect 14660 10554 14688 11698
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14844 11218 14872 11494
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14830 10976 14886 10985
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 14476 10526 14688 10554
rect 13924 9926 13952 10474
rect 14476 10062 14504 10526
rect 14752 10470 14780 10950
rect 14830 10911 14886 10920
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 10198 14780 10406
rect 14740 10192 14792 10198
rect 14740 10134 14792 10140
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13648 8430 13676 9318
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13648 3058 13676 8366
rect 13740 7818 13768 8570
rect 13924 8566 13952 9862
rect 14476 9722 14504 9998
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14660 9654 14688 9998
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 14096 9444 14148 9450
rect 14096 9386 14148 9392
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 14108 7886 14136 9386
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13912 3460 13964 3466
rect 13912 3402 13964 3408
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 13924 2446 13952 3402
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 9600 2310 9628 2382
rect 11704 2372 11756 2378
rect 11704 2314 11756 2320
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 9600 800 9628 2246
rect 11716 800 11744 2314
rect 13832 800 13860 2314
rect 14752 2310 14780 10134
rect 14844 9654 14872 10911
rect 14936 10606 14964 13194
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 15028 9926 15056 13382
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15120 11762 15148 13126
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15108 11280 15160 11286
rect 15108 11222 15160 11228
rect 15120 10130 15148 11222
rect 15212 10130 15240 13398
rect 15290 13016 15346 13025
rect 15290 12951 15292 12960
rect 15344 12951 15346 12960
rect 15292 12922 15344 12928
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15304 11762 15332 12378
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15304 11098 15332 11698
rect 15396 11218 15424 14418
rect 15488 13394 15516 16390
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 15580 13190 15608 15302
rect 15672 15094 15700 16390
rect 15660 15088 15712 15094
rect 15660 15030 15712 15036
rect 15764 14906 15792 17206
rect 15856 16250 15884 19615
rect 16132 19310 16160 19638
rect 16224 19446 16252 20295
rect 16316 19922 16344 21082
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16212 19440 16264 19446
rect 16212 19382 16264 19388
rect 16028 19304 16080 19310
rect 16026 19272 16028 19281
rect 16120 19304 16172 19310
rect 16080 19272 16082 19281
rect 16120 19246 16172 19252
rect 16026 19207 16082 19216
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 16040 17270 16068 17682
rect 16028 17264 16080 17270
rect 16028 17206 16080 17212
rect 16132 17134 16160 18906
rect 16302 18728 16358 18737
rect 16302 18663 16304 18672
rect 16356 18663 16358 18672
rect 16304 18634 16356 18640
rect 16316 18086 16344 18634
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 16212 17604 16264 17610
rect 16212 17546 16264 17552
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15842 16144 15898 16153
rect 15842 16079 15898 16088
rect 15856 16046 15884 16079
rect 15844 16040 15896 16046
rect 15844 15982 15896 15988
rect 15856 15473 15884 15982
rect 15948 15978 15976 16934
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16026 16008 16082 16017
rect 15936 15972 15988 15978
rect 16026 15943 16082 15952
rect 15936 15914 15988 15920
rect 15842 15464 15898 15473
rect 15948 15434 15976 15914
rect 15842 15399 15898 15408
rect 15936 15428 15988 15434
rect 15936 15370 15988 15376
rect 15672 14878 15792 14906
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15488 12306 15516 12718
rect 15672 12434 15700 14878
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15948 14074 15976 14758
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15580 12406 15700 12434
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15580 11694 15608 12406
rect 15764 12306 15792 13330
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15842 12200 15898 12209
rect 15842 12135 15844 12144
rect 15896 12135 15898 12144
rect 15844 12106 15896 12112
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15304 11070 15424 11098
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15120 9722 15148 9862
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 15396 9654 15424 11070
rect 14832 9648 14884 9654
rect 14832 9590 14884 9596
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 14844 8820 14872 9590
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15120 9042 15148 9454
rect 15488 9042 15516 11494
rect 15580 11354 15608 11630
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15948 11218 15976 13126
rect 16040 12442 16068 15943
rect 16132 15570 16160 16050
rect 16224 15570 16252 17546
rect 16316 16697 16344 18022
rect 16408 17134 16436 20538
rect 16488 20324 16540 20330
rect 16488 20266 16540 20272
rect 16500 19174 16528 20266
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16500 17678 16528 18158
rect 16592 18057 16620 22986
rect 16764 22568 16816 22574
rect 16764 22510 16816 22516
rect 16672 21956 16724 21962
rect 16672 21898 16724 21904
rect 16684 21486 16712 21898
rect 16672 21480 16724 21486
rect 16672 21422 16724 21428
rect 16776 21418 16804 22510
rect 17052 22166 17080 26200
rect 17224 24812 17276 24818
rect 17224 24754 17276 24760
rect 17236 24410 17264 24754
rect 17224 24404 17276 24410
rect 17224 24346 17276 24352
rect 17696 24274 17724 26200
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18340 23662 18368 26200
rect 18880 24744 18932 24750
rect 18880 24686 18932 24692
rect 18604 24404 18656 24410
rect 18604 24346 18656 24352
rect 18420 24064 18472 24070
rect 18420 24006 18472 24012
rect 18328 23656 18380 23662
rect 18328 23598 18380 23604
rect 17868 23044 17920 23050
rect 17868 22986 17920 22992
rect 17132 22976 17184 22982
rect 17132 22918 17184 22924
rect 17040 22160 17092 22166
rect 17040 22102 17092 22108
rect 17144 22030 17172 22918
rect 17880 22710 17908 22986
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17868 22704 17920 22710
rect 17868 22646 17920 22652
rect 17880 22574 17908 22646
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 16948 21616 17000 21622
rect 16948 21558 17000 21564
rect 16764 21412 16816 21418
rect 16764 21354 16816 21360
rect 16776 20942 16804 21354
rect 16960 21350 16988 21558
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16764 20936 16816 20942
rect 16764 20878 16816 20884
rect 16776 20466 16804 20878
rect 17144 20602 17172 21966
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 17500 21480 17552 21486
rect 17500 21422 17552 21428
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16856 20392 16908 20398
rect 16856 20334 16908 20340
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16578 18048 16634 18057
rect 16578 17983 16634 17992
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16396 17128 16448 17134
rect 16396 17070 16448 17076
rect 16302 16688 16358 16697
rect 16302 16623 16358 16632
rect 16408 16454 16436 17070
rect 16500 17066 16528 17478
rect 16488 17060 16540 17066
rect 16488 17002 16540 17008
rect 16684 16726 16712 18566
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 16672 16720 16724 16726
rect 16672 16662 16724 16668
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16120 15564 16172 15570
rect 16120 15506 16172 15512
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16132 15450 16160 15506
rect 16132 15422 16344 15450
rect 16408 15434 16436 15846
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 16132 15094 16160 15302
rect 16120 15088 16172 15094
rect 16120 15030 16172 15036
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16224 13258 16252 13806
rect 16316 13258 16344 15422
rect 16396 15428 16448 15434
rect 16396 15370 16448 15376
rect 16212 13252 16264 13258
rect 16212 13194 16264 13200
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 16316 12850 16344 13194
rect 16408 12918 16436 15370
rect 16500 13938 16528 15506
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 16486 13696 16542 13705
rect 16486 13631 16542 13640
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16302 12744 16358 12753
rect 16302 12679 16358 12688
rect 16210 12472 16266 12481
rect 16028 12436 16080 12442
rect 16316 12442 16344 12679
rect 16210 12407 16266 12416
rect 16304 12436 16356 12442
rect 16028 12378 16080 12384
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 14924 8832 14976 8838
rect 14844 8792 14924 8820
rect 14924 8774 14976 8780
rect 14936 8498 14964 8774
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 15120 8430 15148 8978
rect 15580 8974 15608 10746
rect 15856 10742 15884 11018
rect 16040 10985 16068 11698
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16026 10976 16082 10985
rect 16026 10911 16082 10920
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 15844 10736 15896 10742
rect 15844 10678 15896 10684
rect 15764 9722 15792 10678
rect 16028 10600 16080 10606
rect 16028 10542 16080 10548
rect 16040 10266 16068 10542
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 16040 9518 16068 9998
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 15672 6866 15700 9318
rect 16040 9042 16068 9454
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15672 4146 15700 6802
rect 15948 6798 15976 8774
rect 16040 8498 16068 8978
rect 16132 8906 16160 11630
rect 16224 11558 16252 12407
rect 16500 12434 16528 13631
rect 16304 12378 16356 12384
rect 16408 12406 16528 12434
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16408 11234 16436 12406
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16224 11206 16436 11234
rect 16224 10538 16252 11206
rect 16500 11150 16528 11494
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 16212 10532 16264 10538
rect 16212 10474 16264 10480
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16224 8906 16252 9318
rect 16120 8900 16172 8906
rect 16120 8842 16172 8848
rect 16212 8900 16264 8906
rect 16212 8842 16264 8848
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 16224 5642 16252 8842
rect 16316 7818 16344 10950
rect 16408 8838 16436 11086
rect 16592 11082 16620 14010
rect 16684 11354 16712 16526
rect 16776 15706 16804 18294
rect 16868 17746 16896 20334
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17052 19378 17080 20198
rect 17144 19718 17172 20198
rect 17132 19712 17184 19718
rect 17132 19654 17184 19660
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16960 18086 16988 18770
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16960 17746 16988 18022
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16776 13190 16804 14554
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16776 12646 16804 13126
rect 16868 12850 16896 17138
rect 16948 15904 17000 15910
rect 17052 15892 17080 19314
rect 17236 17882 17264 19654
rect 17512 18834 17540 21422
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17880 20874 17908 21286
rect 17868 20868 17920 20874
rect 17868 20810 17920 20816
rect 17880 20584 17908 20810
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17960 20596 18012 20602
rect 17880 20556 17960 20584
rect 17960 20538 18012 20544
rect 17868 19780 17920 19786
rect 17868 19722 17920 19728
rect 17880 18970 17908 19722
rect 18340 19718 18368 21490
rect 18432 19718 18460 24006
rect 18616 23050 18644 24346
rect 18892 24206 18920 24686
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 18788 23520 18840 23526
rect 18788 23462 18840 23468
rect 18604 23044 18656 23050
rect 18604 22986 18656 22992
rect 18616 22778 18644 22986
rect 18604 22772 18656 22778
rect 18604 22714 18656 22720
rect 18800 22642 18828 23462
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 18800 21622 18828 22578
rect 18892 22574 18920 22918
rect 18880 22568 18932 22574
rect 18880 22510 18932 22516
rect 18984 22098 19012 26200
rect 19628 24342 19656 26200
rect 20272 24342 20300 26200
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 19616 24336 19668 24342
rect 19616 24278 19668 24284
rect 20260 24336 20312 24342
rect 20260 24278 20312 24284
rect 20548 24206 20576 24550
rect 20916 24274 20944 26200
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20536 24200 20588 24206
rect 20536 24142 20588 24148
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 20628 24132 20680 24138
rect 20628 24074 20680 24080
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 20260 24064 20312 24070
rect 20260 24006 20312 24012
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19352 22778 19380 23054
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19352 22506 19380 22714
rect 19340 22500 19392 22506
rect 19340 22442 19392 22448
rect 18972 22092 19024 22098
rect 18972 22034 19024 22040
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 18788 21616 18840 21622
rect 18788 21558 18840 21564
rect 19156 21616 19208 21622
rect 19156 21558 19208 21564
rect 18880 21480 18932 21486
rect 18602 21448 18658 21457
rect 18880 21422 18932 21428
rect 18602 21383 18658 21392
rect 18512 20800 18564 20806
rect 18512 20742 18564 20748
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 17868 18964 17920 18970
rect 17868 18906 17920 18912
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17406 18728 17462 18737
rect 17406 18663 17408 18672
rect 17460 18663 17462 18672
rect 17408 18634 17460 18640
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17868 18284 17920 18290
rect 17868 18226 17920 18232
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17420 16998 17448 17478
rect 17408 16992 17460 16998
rect 17406 16960 17408 16969
rect 17460 16960 17462 16969
rect 17406 16895 17462 16904
rect 17498 16688 17554 16697
rect 17498 16623 17554 16632
rect 17512 16590 17540 16623
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 17144 16182 17172 16390
rect 17132 16176 17184 16182
rect 17132 16118 17184 16124
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 17000 15864 17080 15892
rect 16948 15846 17000 15852
rect 16960 14346 16988 15846
rect 17144 15366 17172 15982
rect 17592 15972 17644 15978
rect 17592 15914 17644 15920
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17236 15609 17264 15846
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 17222 15600 17278 15609
rect 17222 15535 17278 15544
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 16948 14340 17000 14346
rect 16948 14282 17000 14288
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16776 12209 16804 12582
rect 16762 12200 16818 12209
rect 16762 12135 16818 12144
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16776 10674 16804 12038
rect 16868 11762 16896 12582
rect 16960 11801 16988 14282
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17052 11830 17080 13874
rect 17144 13802 17172 15302
rect 17236 14414 17264 15535
rect 17328 15366 17356 15642
rect 17500 15632 17552 15638
rect 17500 15574 17552 15580
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17512 15026 17540 15574
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17328 14346 17356 14894
rect 17420 14618 17448 14894
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 17132 13796 17184 13802
rect 17132 13738 17184 13744
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 17144 12646 17172 13194
rect 17420 13025 17448 14418
rect 17500 14272 17552 14278
rect 17500 14214 17552 14220
rect 17512 14074 17540 14214
rect 17604 14074 17632 15914
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17592 13932 17644 13938
rect 17696 13920 17724 14350
rect 17644 13892 17724 13920
rect 17592 13874 17644 13880
rect 17880 13462 17908 18226
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17972 16658 18000 17206
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 17960 14884 18012 14890
rect 17960 14826 18012 14832
rect 17972 14278 18000 14826
rect 18064 14278 18092 14894
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 18340 14074 18368 16186
rect 18432 15910 18460 19314
rect 18524 18766 18552 20742
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18616 18442 18644 21383
rect 18892 20602 18920 21422
rect 19168 21060 19196 21558
rect 19260 21486 19288 21966
rect 19248 21480 19300 21486
rect 19248 21422 19300 21428
rect 19352 21350 19380 22442
rect 19444 22030 19472 24006
rect 19616 23860 19668 23866
rect 19616 23802 19668 23808
rect 19628 23254 19656 23802
rect 20272 23798 20300 24006
rect 20260 23792 20312 23798
rect 20260 23734 20312 23740
rect 20272 23322 20300 23734
rect 19892 23316 19944 23322
rect 19892 23258 19944 23264
rect 20260 23316 20312 23322
rect 20260 23258 20312 23264
rect 19616 23248 19668 23254
rect 19616 23190 19668 23196
rect 19524 23180 19576 23186
rect 19524 23122 19576 23128
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19248 21072 19300 21078
rect 19168 21032 19248 21060
rect 19248 21014 19300 21020
rect 19260 20754 19288 21014
rect 19352 20942 19380 21286
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19432 20868 19484 20874
rect 19432 20810 19484 20816
rect 19340 20800 19392 20806
rect 19260 20748 19340 20754
rect 19260 20742 19392 20748
rect 19260 20726 19380 20742
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18892 19990 18920 20538
rect 19352 20534 19380 20726
rect 19444 20602 19472 20810
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19064 20528 19116 20534
rect 19064 20470 19116 20476
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19076 20330 19104 20470
rect 19064 20324 19116 20330
rect 19064 20266 19116 20272
rect 18880 19984 18932 19990
rect 18880 19926 18932 19932
rect 19076 19446 19104 20266
rect 19536 19990 19564 23122
rect 19800 23044 19852 23050
rect 19800 22986 19852 22992
rect 19812 22681 19840 22986
rect 19798 22672 19854 22681
rect 19798 22607 19854 22616
rect 19708 22568 19760 22574
rect 19708 22510 19760 22516
rect 19616 22228 19668 22234
rect 19616 22170 19668 22176
rect 19628 22137 19656 22170
rect 19614 22128 19670 22137
rect 19614 22063 19670 22072
rect 19616 21344 19668 21350
rect 19616 21286 19668 21292
rect 19628 21078 19656 21286
rect 19720 21146 19748 22510
rect 19708 21140 19760 21146
rect 19708 21082 19760 21088
rect 19616 21072 19668 21078
rect 19616 21014 19668 21020
rect 19800 20936 19852 20942
rect 19800 20878 19852 20884
rect 19616 20800 19668 20806
rect 19616 20742 19668 20748
rect 19628 20262 19656 20742
rect 19708 20596 19760 20602
rect 19708 20538 19760 20544
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 19524 19984 19576 19990
rect 19524 19926 19576 19932
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19352 19530 19380 19654
rect 19352 19514 19472 19530
rect 19352 19508 19484 19514
rect 19352 19502 19432 19508
rect 19064 19440 19116 19446
rect 19352 19417 19380 19502
rect 19432 19450 19484 19456
rect 19064 19382 19116 19388
rect 19338 19408 19394 19417
rect 19338 19343 19394 19352
rect 19432 19304 19484 19310
rect 19432 19246 19484 19252
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 18524 18414 18644 18442
rect 18696 18420 18748 18426
rect 18524 15960 18552 18414
rect 18696 18362 18748 18368
rect 18604 17604 18656 17610
rect 18708 17592 18736 18362
rect 18656 17564 18736 17592
rect 18604 17546 18656 17552
rect 18708 17270 18736 17564
rect 18880 17536 18932 17542
rect 18880 17478 18932 17484
rect 18696 17264 18748 17270
rect 18696 17206 18748 17212
rect 18708 16250 18736 17206
rect 18892 16794 18920 17478
rect 18970 17232 19026 17241
rect 18970 17167 19026 17176
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 18524 15932 18644 15960
rect 18420 15904 18472 15910
rect 18472 15864 18552 15892
rect 18420 15846 18472 15852
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18432 14618 18460 15438
rect 18524 15434 18552 15864
rect 18616 15638 18644 15932
rect 18604 15632 18656 15638
rect 18604 15574 18656 15580
rect 18512 15428 18564 15434
rect 18512 15370 18564 15376
rect 18510 15056 18566 15065
rect 18510 14991 18512 15000
rect 18564 14991 18566 15000
rect 18512 14962 18564 14968
rect 18510 14920 18566 14929
rect 18510 14855 18566 14864
rect 18524 14618 18552 14855
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18616 14414 18644 14758
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18420 14272 18472 14278
rect 18472 14232 18552 14260
rect 18420 14214 18472 14220
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 17972 13530 18000 13738
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 17868 13456 17920 13462
rect 17868 13398 17920 13404
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17406 13016 17462 13025
rect 17950 13019 18258 13028
rect 18340 12986 18368 13262
rect 17406 12951 17462 12960
rect 18328 12980 18380 12986
rect 17316 12708 17368 12714
rect 17316 12650 17368 12656
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 17222 12336 17278 12345
rect 17222 12271 17278 12280
rect 17236 12102 17264 12271
rect 17224 12096 17276 12102
rect 17222 12064 17224 12073
rect 17276 12064 17278 12073
rect 17222 11999 17278 12008
rect 17040 11824 17092 11830
rect 16946 11792 17002 11801
rect 16856 11756 16908 11762
rect 17040 11766 17092 11772
rect 16946 11727 17002 11736
rect 16856 11698 16908 11704
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16592 10198 16620 10406
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 16684 10062 16712 10542
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16488 9716 16540 9722
rect 16488 9658 16540 9664
rect 16500 9382 16528 9658
rect 16684 9654 16712 9998
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16856 9104 16908 9110
rect 16856 9046 16908 9052
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16408 8566 16436 8774
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 16776 7954 16804 8502
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16304 7812 16356 7818
rect 16304 7754 16356 7760
rect 16868 6322 16896 9046
rect 16960 7954 16988 9862
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 17052 7886 17080 10406
rect 17144 8430 17172 11018
rect 17328 10130 17356 12650
rect 17420 12306 17448 12951
rect 18328 12922 18380 12928
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17788 12714 17816 12786
rect 17776 12708 17828 12714
rect 17776 12650 17828 12656
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17592 12164 17644 12170
rect 17592 12106 17644 12112
rect 17604 11694 17632 12106
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 18432 11370 18460 13466
rect 18524 13297 18552 14232
rect 18510 13288 18566 13297
rect 18510 13223 18566 13232
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18524 12730 18552 13126
rect 18604 12844 18656 12850
rect 18708 12832 18736 16186
rect 18800 14074 18828 16390
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18892 13870 18920 16730
rect 18984 15638 19012 17167
rect 18972 15632 19024 15638
rect 18972 15574 19024 15580
rect 18984 14278 19012 15574
rect 18972 14272 19024 14278
rect 18972 14214 19024 14220
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 18984 13394 19012 13806
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18984 12918 19012 13330
rect 19076 12986 19104 19110
rect 19338 18728 19394 18737
rect 19444 18698 19472 19246
rect 19536 18970 19564 19790
rect 19628 19174 19656 20198
rect 19616 19168 19668 19174
rect 19616 19110 19668 19116
rect 19524 18964 19576 18970
rect 19524 18906 19576 18912
rect 19338 18663 19340 18672
rect 19392 18663 19394 18672
rect 19432 18692 19484 18698
rect 19340 18634 19392 18640
rect 19432 18634 19484 18640
rect 19444 18442 19472 18634
rect 19628 18630 19656 19110
rect 19720 18834 19748 20538
rect 19812 19310 19840 20878
rect 19904 19922 19932 23258
rect 20168 22160 20220 22166
rect 20168 22102 20220 22108
rect 20180 20602 20208 22102
rect 20640 21622 20668 24074
rect 21468 23866 21496 24142
rect 21456 23860 21508 23866
rect 21456 23802 21508 23808
rect 21270 23760 21326 23769
rect 21270 23695 21272 23704
rect 21324 23695 21326 23704
rect 21272 23666 21324 23672
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 20812 22976 20864 22982
rect 20812 22918 20864 22924
rect 20824 22642 20852 22918
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 20824 22438 20852 22578
rect 20812 22432 20864 22438
rect 20812 22374 20864 22380
rect 21008 21690 21036 23462
rect 21560 22982 21588 26200
rect 21640 23792 21692 23798
rect 21640 23734 21692 23740
rect 21652 23032 21680 23734
rect 21732 23656 21784 23662
rect 21732 23598 21784 23604
rect 21744 23202 21772 23598
rect 21744 23186 21956 23202
rect 21732 23180 21956 23186
rect 21784 23174 21956 23180
rect 21732 23122 21784 23128
rect 21732 23044 21784 23050
rect 21652 23004 21732 23032
rect 21548 22976 21600 22982
rect 21548 22918 21600 22924
rect 21364 22772 21416 22778
rect 21364 22714 21416 22720
rect 21270 22128 21326 22137
rect 21270 22063 21326 22072
rect 21284 21894 21312 22063
rect 21272 21888 21324 21894
rect 21272 21830 21324 21836
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 20628 21616 20680 21622
rect 20628 21558 20680 21564
rect 21088 21412 21140 21418
rect 21088 21354 21140 21360
rect 21100 20602 21128 21354
rect 20168 20596 20220 20602
rect 20168 20538 20220 20544
rect 21088 20596 21140 20602
rect 21088 20538 21140 20544
rect 20444 20392 20496 20398
rect 20444 20334 20496 20340
rect 21180 20392 21232 20398
rect 21180 20334 21232 20340
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 19892 19916 19944 19922
rect 19892 19858 19944 19864
rect 19800 19304 19852 19310
rect 19800 19246 19852 19252
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19616 18624 19668 18630
rect 19616 18566 19668 18572
rect 19444 18414 19564 18442
rect 19156 18352 19208 18358
rect 19156 18294 19208 18300
rect 19168 18222 19196 18294
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19156 18216 19208 18222
rect 19156 18158 19208 18164
rect 19168 17338 19196 18158
rect 19338 18048 19394 18057
rect 19338 17983 19394 17992
rect 19352 17882 19380 17983
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19156 17332 19208 17338
rect 19156 17274 19208 17280
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 19156 16652 19208 16658
rect 19156 16594 19208 16600
rect 19168 16114 19196 16594
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 19352 15638 19380 17138
rect 19340 15632 19392 15638
rect 19154 15600 19210 15609
rect 19340 15574 19392 15580
rect 19154 15535 19210 15544
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 18972 12912 19024 12918
rect 18972 12854 19024 12860
rect 18656 12804 18736 12832
rect 19064 12844 19116 12850
rect 18604 12786 18656 12792
rect 19064 12786 19116 12792
rect 18524 12702 18644 12730
rect 18432 11342 18552 11370
rect 17592 11280 17644 11286
rect 17592 11222 17644 11228
rect 17500 10192 17552 10198
rect 17500 10134 17552 10140
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17512 9926 17540 10134
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17236 9178 17264 9658
rect 17328 9450 17356 9862
rect 17604 9518 17632 11222
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 17696 9994 17724 10542
rect 18064 10266 18092 10542
rect 18340 10266 18368 11086
rect 18524 10538 18552 11342
rect 18616 11218 18644 12702
rect 19076 12434 19104 12786
rect 18892 12406 19104 12434
rect 18892 12170 18920 12406
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 18880 12164 18932 12170
rect 18880 12106 18932 12112
rect 18800 11694 18828 12106
rect 18788 11688 18840 11694
rect 18788 11630 18840 11636
rect 18800 11234 18828 11630
rect 18892 11354 18920 12106
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18696 11212 18748 11218
rect 18800 11206 18920 11234
rect 18696 11154 18748 11160
rect 18708 11098 18736 11154
rect 18708 11070 18828 11098
rect 18800 11014 18828 11070
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18524 10198 18552 10474
rect 17868 10192 17920 10198
rect 17868 10134 17920 10140
rect 18512 10192 18564 10198
rect 18512 10134 18564 10140
rect 17684 9988 17736 9994
rect 17684 9930 17736 9936
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17316 9444 17368 9450
rect 17316 9386 17368 9392
rect 17880 9178 17908 10134
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 18328 9648 18380 9654
rect 18328 9590 18380 9596
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 18340 8906 18368 9590
rect 17408 8900 17460 8906
rect 17408 8842 17460 8848
rect 18328 8900 18380 8906
rect 18328 8842 18380 8848
rect 17132 8424 17184 8430
rect 17420 8412 17448 8842
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 18340 8514 18368 8842
rect 18248 8498 18368 8514
rect 18236 8492 18368 8498
rect 18288 8486 18368 8492
rect 18236 8434 18288 8440
rect 17132 8366 17184 8372
rect 17328 8384 17448 8412
rect 17328 8294 17356 8384
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 18432 8090 18460 10066
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18524 9382 18552 9862
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18616 8634 18644 9454
rect 18708 8974 18736 10610
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18800 8838 18828 10950
rect 18892 9518 18920 11206
rect 19168 10198 19196 15535
rect 19444 15162 19472 18226
rect 19536 15570 19564 18414
rect 19628 18222 19656 18566
rect 19616 18216 19668 18222
rect 19616 18158 19668 18164
rect 19628 17882 19656 18158
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19628 17728 19656 17818
rect 19708 17740 19760 17746
rect 19628 17700 19708 17728
rect 19708 17682 19760 17688
rect 19996 16046 20024 19994
rect 20352 19780 20404 19786
rect 20352 19722 20404 19728
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 20272 19446 20300 19654
rect 20260 19440 20312 19446
rect 20260 19382 20312 19388
rect 20272 17338 20300 19382
rect 20364 18873 20392 19722
rect 20456 19718 20484 20334
rect 20536 19848 20588 19854
rect 20588 19796 20760 19802
rect 20536 19790 20760 19796
rect 20548 19774 20760 19790
rect 20444 19712 20496 19718
rect 20444 19654 20496 19660
rect 20350 18864 20406 18873
rect 20456 18834 20484 19654
rect 20626 19272 20682 19281
rect 20626 19207 20682 19216
rect 20640 18902 20668 19207
rect 20732 18970 20760 19774
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20628 18896 20680 18902
rect 20628 18838 20680 18844
rect 20350 18799 20406 18808
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20350 18048 20406 18057
rect 20350 17983 20406 17992
rect 20364 17746 20392 17983
rect 20824 17898 20852 19450
rect 21192 19334 21220 20334
rect 21270 19544 21326 19553
rect 21270 19479 21272 19488
rect 21324 19479 21326 19488
rect 21272 19450 21324 19456
rect 21192 19306 21312 19334
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21088 18760 21140 18766
rect 21088 18702 21140 18708
rect 20732 17870 20852 17898
rect 20732 17814 20760 17870
rect 20720 17808 20772 17814
rect 20720 17750 20772 17756
rect 20352 17740 20404 17746
rect 20352 17682 20404 17688
rect 20364 17542 20392 17682
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20536 17264 20588 17270
rect 20536 17206 20588 17212
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 20168 16720 20220 16726
rect 20168 16662 20220 16668
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19524 15564 19576 15570
rect 19524 15506 19576 15512
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19352 15042 19380 15098
rect 19536 15042 19564 15506
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19352 15014 19564 15042
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 19246 13288 19302 13297
rect 19246 13223 19302 13232
rect 19156 10192 19208 10198
rect 19156 10134 19208 10140
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18892 9042 18920 9454
rect 18880 9036 18932 9042
rect 18880 8978 18932 8984
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18512 8492 18564 8498
rect 18512 8434 18564 8440
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18524 7478 18552 8434
rect 18616 7954 18644 8570
rect 18892 8566 18920 8774
rect 18880 8560 18932 8566
rect 18880 8502 18932 8508
rect 18880 8016 18932 8022
rect 18880 7958 18932 7964
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 17868 7472 17920 7478
rect 17868 7414 17920 7420
rect 18512 7472 18564 7478
rect 18512 7414 18564 7420
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16212 5636 16264 5642
rect 16212 5578 16264 5584
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 17880 3126 17908 7414
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18340 4010 18368 6190
rect 18892 5234 18920 7958
rect 19260 7274 19288 13223
rect 19352 13190 19380 14418
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 19444 13938 19472 14282
rect 19812 14278 19840 15302
rect 20180 14958 20208 16662
rect 20548 16454 20576 17206
rect 21008 16794 21036 17206
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20536 16448 20588 16454
rect 20536 16390 20588 16396
rect 20444 15972 20496 15978
rect 20444 15914 20496 15920
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 20074 14376 20130 14385
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19536 14006 19564 14214
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19352 11898 19380 12582
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19444 11744 19472 13874
rect 19812 13734 19840 14214
rect 19904 14074 19932 14350
rect 20074 14311 20130 14320
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 20088 13841 20116 14311
rect 20074 13832 20130 13841
rect 20074 13767 20130 13776
rect 19800 13728 19852 13734
rect 19800 13670 19852 13676
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19996 13394 20024 13670
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19892 12912 19944 12918
rect 19892 12854 19944 12860
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19536 12288 19564 12786
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 19536 12260 19656 12288
rect 19524 11756 19576 11762
rect 19444 11716 19524 11744
rect 19524 11698 19576 11704
rect 19536 11286 19564 11698
rect 19524 11280 19576 11286
rect 19524 11222 19576 11228
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 19444 9042 19472 10066
rect 19536 9654 19564 11086
rect 19628 10130 19656 12260
rect 19720 10810 19748 12718
rect 19904 12458 19932 12854
rect 19812 12430 19932 12458
rect 19812 12238 19840 12430
rect 19996 12424 20024 13126
rect 19983 12396 20024 12424
rect 20088 12434 20116 13767
rect 20272 13530 20300 15302
rect 20456 14414 20484 15914
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20548 14278 20576 14894
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20272 12434 20300 12718
rect 20088 12406 20208 12434
rect 20272 12406 20484 12434
rect 19892 12300 19944 12306
rect 19983 12288 20011 12396
rect 20180 12356 20208 12406
rect 20180 12328 20392 12356
rect 19983 12260 20024 12288
rect 19892 12242 19944 12248
rect 19800 12232 19852 12238
rect 19800 12174 19852 12180
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19708 10804 19760 10810
rect 19708 10746 19760 10752
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19536 9178 19564 9590
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19444 8090 19472 8978
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19616 7812 19668 7818
rect 19616 7754 19668 7760
rect 19248 7268 19300 7274
rect 19248 7210 19300 7216
rect 19628 6798 19656 7754
rect 19812 7546 19840 12038
rect 19904 8634 19932 12242
rect 19996 11898 20024 12260
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 20088 11830 20116 12038
rect 20076 11824 20128 11830
rect 20076 11766 20128 11772
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 20088 11286 20116 11630
rect 20076 11280 20128 11286
rect 20076 11222 20128 11228
rect 20180 11218 20208 12106
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 19984 11008 20036 11014
rect 19984 10950 20036 10956
rect 19996 10606 20024 10950
rect 20364 10742 20392 12328
rect 20352 10736 20404 10742
rect 20352 10678 20404 10684
rect 20456 10674 20484 12406
rect 20548 12238 20576 14214
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20640 12084 20668 16594
rect 20812 16448 20864 16454
rect 20812 16390 20864 16396
rect 20824 16182 20852 16390
rect 20812 16176 20864 16182
rect 20812 16118 20864 16124
rect 20904 16176 20956 16182
rect 20904 16118 20956 16124
rect 20824 15910 20852 16118
rect 20812 15904 20864 15910
rect 20732 15864 20812 15892
rect 20732 14550 20760 15864
rect 20812 15846 20864 15852
rect 20810 15736 20866 15745
rect 20810 15671 20812 15680
rect 20864 15671 20866 15680
rect 20812 15642 20864 15648
rect 20916 15502 20944 16118
rect 20996 16040 21048 16046
rect 20996 15982 21048 15988
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 20732 14006 20760 14486
rect 20720 14000 20772 14006
rect 20720 13942 20772 13948
rect 20732 13870 20760 13942
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20824 13682 20852 15030
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20548 12056 20668 12084
rect 20732 13654 20852 13682
rect 20548 11082 20576 12056
rect 20732 11898 20760 13654
rect 20916 13530 20944 14962
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20626 11792 20682 11801
rect 20916 11762 20944 12174
rect 20626 11727 20628 11736
rect 20680 11727 20682 11736
rect 20904 11756 20956 11762
rect 20628 11698 20680 11704
rect 20904 11698 20956 11704
rect 21008 11626 21036 15982
rect 21100 15366 21128 18702
rect 21192 18358 21220 19110
rect 21180 18352 21232 18358
rect 21180 18294 21232 18300
rect 21284 18086 21312 19306
rect 21376 18834 21404 22714
rect 21652 22438 21680 23004
rect 21732 22986 21784 22992
rect 21824 23044 21876 23050
rect 21824 22986 21876 22992
rect 21836 22778 21864 22986
rect 21824 22772 21876 22778
rect 21824 22714 21876 22720
rect 21836 22506 21864 22714
rect 21928 22642 21956 23174
rect 21916 22636 21968 22642
rect 21968 22596 22140 22624
rect 21916 22578 21968 22584
rect 21824 22500 21876 22506
rect 21824 22442 21876 22448
rect 21640 22432 21692 22438
rect 21640 22374 21692 22380
rect 21548 21956 21600 21962
rect 21548 21898 21600 21904
rect 21456 21888 21508 21894
rect 21456 21830 21508 21836
rect 21468 20262 21496 21830
rect 21560 21486 21588 21898
rect 21548 21480 21600 21486
rect 21548 21422 21600 21428
rect 21652 21350 21680 22374
rect 22112 22094 22140 22596
rect 22204 22234 22232 26200
rect 22560 24676 22612 24682
rect 22560 24618 22612 24624
rect 22376 24268 22428 24274
rect 22376 24210 22428 24216
rect 22192 22228 22244 22234
rect 22192 22170 22244 22176
rect 22388 22094 22416 24210
rect 22572 23662 22600 24618
rect 22560 23656 22612 23662
rect 22560 23598 22612 23604
rect 22848 23322 22876 26200
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23492 23730 23520 26200
rect 24032 24812 24084 24818
rect 24032 24754 24084 24760
rect 23848 24064 23900 24070
rect 23848 24006 23900 24012
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23664 23724 23716 23730
rect 23664 23666 23716 23672
rect 23388 23588 23440 23594
rect 23388 23530 23440 23536
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22836 23316 22888 23322
rect 22836 23258 22888 23264
rect 23400 23254 23428 23530
rect 23480 23520 23532 23526
rect 23480 23462 23532 23468
rect 23388 23248 23440 23254
rect 23388 23190 23440 23196
rect 23294 23080 23350 23089
rect 22560 23044 22612 23050
rect 23294 23015 23350 23024
rect 22560 22986 22612 22992
rect 22112 22066 22232 22094
rect 22388 22066 22508 22094
rect 21916 21888 21968 21894
rect 21916 21830 21968 21836
rect 21928 21690 21956 21830
rect 21916 21684 21968 21690
rect 21916 21626 21968 21632
rect 22204 21486 22232 22066
rect 22282 21856 22338 21865
rect 22282 21791 22338 21800
rect 22296 21554 22324 21791
rect 22284 21548 22336 21554
rect 22284 21490 22336 21496
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 21640 21344 21692 21350
rect 21560 21304 21640 21332
rect 21456 20256 21508 20262
rect 21456 20198 21508 20204
rect 21560 19786 21588 21304
rect 21640 21286 21692 21292
rect 21914 21040 21970 21049
rect 21914 20975 21970 20984
rect 21732 20596 21784 20602
rect 21732 20538 21784 20544
rect 21548 19780 21600 19786
rect 21548 19722 21600 19728
rect 21364 18828 21416 18834
rect 21364 18770 21416 18776
rect 21456 18624 21508 18630
rect 21454 18592 21456 18601
rect 21508 18592 21510 18601
rect 21454 18527 21510 18536
rect 21640 18352 21692 18358
rect 21640 18294 21692 18300
rect 21548 18216 21600 18222
rect 21548 18158 21600 18164
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 21192 16794 21220 17070
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 21284 16250 21312 18022
rect 21364 17876 21416 17882
rect 21364 17818 21416 17824
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 21178 15600 21234 15609
rect 21178 15535 21234 15544
rect 21272 15564 21324 15570
rect 21192 15502 21220 15535
rect 21272 15506 21324 15512
rect 21180 15496 21232 15502
rect 21180 15438 21232 15444
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 21284 14346 21312 15506
rect 21376 14958 21404 17818
rect 21468 17270 21496 18022
rect 21560 17882 21588 18158
rect 21548 17876 21600 17882
rect 21548 17818 21600 17824
rect 21652 17610 21680 18294
rect 21744 17746 21772 20538
rect 21824 18760 21876 18766
rect 21824 18702 21876 18708
rect 21732 17740 21784 17746
rect 21732 17682 21784 17688
rect 21836 17610 21864 18702
rect 21640 17604 21692 17610
rect 21640 17546 21692 17552
rect 21824 17604 21876 17610
rect 21824 17546 21876 17552
rect 21456 17264 21508 17270
rect 21456 17206 21508 17212
rect 21652 17134 21680 17546
rect 21732 17332 21784 17338
rect 21732 17274 21784 17280
rect 21640 17128 21692 17134
rect 21640 17070 21692 17076
rect 21640 16992 21692 16998
rect 21744 16980 21772 17274
rect 21692 16952 21772 16980
rect 21836 16969 21864 17546
rect 21822 16960 21878 16969
rect 21640 16934 21692 16940
rect 21456 16244 21508 16250
rect 21456 16186 21508 16192
rect 21468 15570 21496 16186
rect 21548 16176 21600 16182
rect 21548 16118 21600 16124
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21456 15428 21508 15434
rect 21456 15370 21508 15376
rect 21468 15026 21496 15370
rect 21560 15314 21588 16118
rect 21652 15450 21680 16934
rect 21822 16895 21878 16904
rect 21652 15422 21772 15450
rect 21560 15286 21680 15314
rect 21548 15156 21600 15162
rect 21548 15098 21600 15104
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 21364 14952 21416 14958
rect 21364 14894 21416 14900
rect 21376 14482 21404 14894
rect 21454 14512 21510 14521
rect 21364 14476 21416 14482
rect 21454 14447 21510 14456
rect 21364 14418 21416 14424
rect 21272 14340 21324 14346
rect 21272 14282 21324 14288
rect 21284 14074 21312 14282
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21088 13796 21140 13802
rect 21088 13738 21140 13744
rect 20996 11620 21048 11626
rect 20996 11562 21048 11568
rect 20536 11076 20588 11082
rect 21100 11064 21128 13738
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 21272 12776 21324 12782
rect 21272 12718 21324 12724
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 21192 12306 21220 12582
rect 21180 12300 21232 12306
rect 21180 12242 21232 12248
rect 21192 11898 21220 12242
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21284 11558 21312 12718
rect 21376 11694 21404 13330
rect 21468 13258 21496 14447
rect 21560 14074 21588 15098
rect 21652 15094 21680 15286
rect 21640 15088 21692 15094
rect 21640 15030 21692 15036
rect 21744 14906 21772 15422
rect 21652 14878 21772 14906
rect 21652 14385 21680 14878
rect 21732 14476 21784 14482
rect 21732 14418 21784 14424
rect 21638 14376 21694 14385
rect 21638 14311 21694 14320
rect 21744 14278 21772 14418
rect 21732 14272 21784 14278
rect 21732 14214 21784 14220
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 21456 13252 21508 13258
rect 21456 13194 21508 13200
rect 21640 13252 21692 13258
rect 21640 13194 21692 13200
rect 21548 13184 21600 13190
rect 21454 13152 21510 13161
rect 21548 13126 21600 13132
rect 21454 13087 21510 13096
rect 21468 12238 21496 13087
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21284 11218 21312 11494
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21180 11076 21232 11082
rect 21100 11036 21180 11064
rect 20536 11018 20588 11024
rect 21180 11018 21232 11024
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19996 9994 20024 10542
rect 20456 10266 20484 10610
rect 21088 10600 21140 10606
rect 21088 10542 21140 10548
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 21100 10130 21128 10542
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 21088 10124 21140 10130
rect 21088 10066 21140 10072
rect 20628 10056 20680 10062
rect 20628 9998 20680 10004
rect 19984 9988 20036 9994
rect 19984 9930 20036 9936
rect 20640 9586 20668 9998
rect 21100 9722 21128 10066
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21284 9654 21312 10474
rect 21362 10160 21418 10169
rect 21362 10095 21418 10104
rect 21376 9926 21404 10095
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21456 9920 21508 9926
rect 21456 9862 21508 9868
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 21468 8974 21496 9862
rect 21560 9382 21588 13126
rect 21652 11898 21680 13194
rect 21836 13190 21864 16895
rect 21928 16182 21956 20975
rect 22204 20466 22232 21422
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22008 20256 22060 20262
rect 22008 20198 22060 20204
rect 22020 20058 22048 20198
rect 22008 20052 22060 20058
rect 22008 19994 22060 20000
rect 22100 19780 22152 19786
rect 22100 19722 22152 19728
rect 22112 18630 22140 19722
rect 22204 19378 22232 20402
rect 22296 20210 22324 21490
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22388 20874 22416 21286
rect 22376 20868 22428 20874
rect 22376 20810 22428 20816
rect 22480 20516 22508 22066
rect 22572 22030 22600 22986
rect 23308 22982 23336 23015
rect 23204 22976 23256 22982
rect 23204 22918 23256 22924
rect 23296 22976 23348 22982
rect 23296 22918 23348 22924
rect 23216 22778 23244 22918
rect 23204 22772 23256 22778
rect 23204 22714 23256 22720
rect 23296 22568 23348 22574
rect 23296 22510 23348 22516
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 22744 22092 22796 22098
rect 22744 22034 22796 22040
rect 22560 22024 22612 22030
rect 22560 21966 22612 21972
rect 22652 21888 22704 21894
rect 22652 21830 22704 21836
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 22572 21350 22600 21626
rect 22560 21344 22612 21350
rect 22560 21286 22612 21292
rect 22560 21140 22612 21146
rect 22560 21082 22612 21088
rect 22572 20874 22600 21082
rect 22664 21010 22692 21830
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22756 20874 22784 22034
rect 22928 21956 22980 21962
rect 22928 21898 22980 21904
rect 22940 21690 22968 21898
rect 23112 21888 23164 21894
rect 23110 21856 23112 21865
rect 23164 21856 23166 21865
rect 23110 21791 23166 21800
rect 22928 21684 22980 21690
rect 22928 21626 22980 21632
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23308 21078 23336 22510
rect 23492 22012 23520 23462
rect 23572 22568 23624 22574
rect 23572 22510 23624 22516
rect 23584 22098 23612 22510
rect 23676 22098 23704 23666
rect 23860 23662 23888 24006
rect 23848 23656 23900 23662
rect 23848 23598 23900 23604
rect 23756 22976 23808 22982
rect 23756 22918 23808 22924
rect 23768 22273 23796 22918
rect 24044 22710 24072 24754
rect 24032 22704 24084 22710
rect 24032 22646 24084 22652
rect 23754 22264 23810 22273
rect 23754 22199 23810 22208
rect 23572 22092 23624 22098
rect 23572 22034 23624 22040
rect 23664 22092 23716 22098
rect 23664 22034 23716 22040
rect 23400 21984 23520 22012
rect 24032 22024 24084 22030
rect 23296 21072 23348 21078
rect 23296 21014 23348 21020
rect 22928 20936 22980 20942
rect 22928 20878 22980 20884
rect 22560 20868 22612 20874
rect 22560 20810 22612 20816
rect 22744 20868 22796 20874
rect 22744 20810 22796 20816
rect 22940 20602 22968 20878
rect 22744 20596 22796 20602
rect 22928 20596 22980 20602
rect 22744 20538 22796 20544
rect 22848 20556 22928 20584
rect 22480 20488 22692 20516
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22296 20182 22416 20210
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22388 19334 22416 20182
rect 22480 20058 22508 20334
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22008 18624 22060 18630
rect 22008 18566 22060 18572
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22020 17338 22048 18566
rect 22100 17740 22152 17746
rect 22204 17728 22232 19314
rect 22284 19304 22336 19310
rect 22388 19306 22508 19334
rect 22284 19246 22336 19252
rect 22296 17814 22324 19246
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22388 18465 22416 18566
rect 22374 18456 22430 18465
rect 22374 18391 22430 18400
rect 22284 17808 22336 17814
rect 22284 17750 22336 17756
rect 22152 17700 22232 17728
rect 22100 17682 22152 17688
rect 22008 17332 22060 17338
rect 22008 17274 22060 17280
rect 22112 17202 22140 17682
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 22100 17196 22152 17202
rect 22100 17138 22152 17144
rect 22008 17128 22060 17134
rect 22008 17070 22060 17076
rect 22098 17096 22154 17105
rect 22020 16522 22048 17070
rect 22098 17031 22154 17040
rect 22008 16516 22060 16522
rect 22008 16458 22060 16464
rect 21916 16176 21968 16182
rect 21916 16118 21968 16124
rect 21916 16040 21968 16046
rect 21916 15982 21968 15988
rect 21928 13802 21956 15982
rect 22020 15910 22048 16458
rect 22112 15978 22140 17031
rect 22100 15972 22152 15978
rect 22100 15914 22152 15920
rect 22008 15904 22060 15910
rect 22008 15846 22060 15852
rect 22100 15632 22152 15638
rect 22100 15574 22152 15580
rect 22008 15564 22060 15570
rect 22008 15506 22060 15512
rect 22020 13870 22048 15506
rect 22112 15434 22140 15574
rect 22100 15428 22152 15434
rect 22100 15370 22152 15376
rect 22008 13864 22060 13870
rect 22008 13806 22060 13812
rect 21916 13796 21968 13802
rect 21916 13738 21968 13744
rect 22204 13530 22232 17478
rect 22480 17377 22508 19306
rect 22572 18057 22600 20334
rect 22664 20330 22692 20488
rect 22652 20324 22704 20330
rect 22652 20266 22704 20272
rect 22756 19854 22784 20538
rect 22848 19922 22876 20556
rect 22928 20538 22980 20544
rect 23400 20466 23428 21984
rect 24032 21966 24084 21972
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23768 20913 23796 21830
rect 23848 21548 23900 21554
rect 23848 21490 23900 21496
rect 23860 21078 23888 21490
rect 23848 21072 23900 21078
rect 23848 21014 23900 21020
rect 23754 20904 23810 20913
rect 23572 20868 23624 20874
rect 23754 20839 23810 20848
rect 23572 20810 23624 20816
rect 23388 20460 23440 20466
rect 23388 20402 23440 20408
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 23388 19916 23440 19922
rect 23388 19858 23440 19864
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 23400 19718 23428 19858
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 23388 19712 23440 19718
rect 23388 19654 23440 19660
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 22664 19446 22692 19654
rect 23400 19446 23428 19654
rect 23492 19514 23520 19654
rect 23480 19508 23532 19514
rect 23480 19450 23532 19456
rect 22652 19440 22704 19446
rect 22652 19382 22704 19388
rect 23388 19440 23440 19446
rect 23388 19382 23440 19388
rect 22664 18358 22692 19382
rect 22836 19304 22888 19310
rect 22836 19246 22888 19252
rect 22652 18352 22704 18358
rect 22652 18294 22704 18300
rect 22558 18048 22614 18057
rect 22558 17983 22614 17992
rect 22466 17368 22522 17377
rect 22466 17303 22522 17312
rect 22376 16652 22428 16658
rect 22480 16640 22508 17303
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 22756 16658 22784 17138
rect 22848 16726 22876 19246
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23112 18964 23164 18970
rect 23112 18906 23164 18912
rect 23020 18828 23072 18834
rect 23020 18770 23072 18776
rect 23032 18601 23060 18770
rect 23018 18592 23074 18601
rect 23018 18527 23074 18536
rect 23124 18290 23152 18906
rect 23296 18692 23348 18698
rect 23480 18692 23532 18698
rect 23348 18652 23428 18680
rect 23296 18634 23348 18640
rect 23296 18352 23348 18358
rect 23296 18294 23348 18300
rect 23112 18284 23164 18290
rect 23112 18226 23164 18232
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23308 16794 23336 18294
rect 23400 17218 23428 18652
rect 23480 18634 23532 18640
rect 23492 17678 23520 18634
rect 23584 17814 23612 20810
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23768 18154 23796 20470
rect 23938 20088 23994 20097
rect 23938 20023 23994 20032
rect 23952 19990 23980 20023
rect 23940 19984 23992 19990
rect 23940 19926 23992 19932
rect 23848 19168 23900 19174
rect 23848 19110 23900 19116
rect 23860 18698 23888 19110
rect 23848 18692 23900 18698
rect 23848 18634 23900 18640
rect 23756 18148 23808 18154
rect 23756 18090 23808 18096
rect 23572 17808 23624 17814
rect 23572 17750 23624 17756
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23492 17338 23520 17614
rect 23756 17536 23808 17542
rect 23756 17478 23808 17484
rect 23480 17332 23532 17338
rect 23480 17274 23532 17280
rect 23664 17264 23716 17270
rect 23400 17212 23664 17218
rect 23400 17206 23716 17212
rect 23400 17190 23704 17206
rect 23400 17134 23428 17190
rect 23388 17128 23440 17134
rect 23388 17070 23440 17076
rect 23296 16788 23348 16794
rect 23296 16730 23348 16736
rect 22836 16720 22888 16726
rect 22836 16662 22888 16668
rect 22428 16612 22508 16640
rect 22744 16652 22796 16658
rect 22376 16594 22428 16600
rect 22744 16594 22796 16600
rect 22466 16552 22522 16561
rect 22848 16538 22876 16662
rect 22466 16487 22522 16496
rect 22756 16510 22876 16538
rect 22480 15706 22508 16487
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22558 15736 22614 15745
rect 22468 15700 22520 15706
rect 22558 15671 22560 15680
rect 22468 15642 22520 15648
rect 22612 15671 22614 15680
rect 22560 15642 22612 15648
rect 22480 15502 22508 15642
rect 22468 15496 22520 15502
rect 22468 15438 22520 15444
rect 22284 15360 22336 15366
rect 22284 15302 22336 15308
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 21824 13184 21876 13190
rect 21824 13126 21876 13132
rect 22098 13016 22154 13025
rect 22098 12951 22154 12960
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21732 12776 21784 12782
rect 21732 12718 21784 12724
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 21652 10266 21680 11834
rect 21744 11830 21772 12718
rect 21732 11824 21784 11830
rect 21732 11766 21784 11772
rect 21640 10260 21692 10266
rect 21640 10202 21692 10208
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21824 9376 21876 9382
rect 21824 9318 21876 9324
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 20444 8900 20496 8906
rect 20444 8842 20496 8848
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19904 7954 19932 8570
rect 20456 8566 20484 8842
rect 20444 8560 20496 8566
rect 20444 8502 20496 8508
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 20456 7818 20484 8502
rect 21468 8430 21496 8910
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21468 7886 21496 8366
rect 21640 8016 21692 8022
rect 21640 7958 21692 7964
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20996 7812 21048 7818
rect 20996 7754 21048 7760
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 20456 7478 20484 7754
rect 20444 7472 20496 7478
rect 20444 7414 20496 7420
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 19076 4554 19104 5102
rect 19260 4690 19288 6598
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 19064 4548 19116 4554
rect 19064 4490 19116 4496
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 18328 4004 18380 4010
rect 18328 3946 18380 3952
rect 17972 3534 18000 3946
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 19076 3058 19104 4490
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 19352 3194 19380 3402
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 17420 2446 17448 2790
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 15948 800 15976 2314
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 1122 0 1178 800
rect 3238 0 3294 800
rect 5354 0 5410 800
rect 7470 0 7526 800
rect 9586 0 9642 800
rect 11702 0 11758 800
rect 13818 0 13874 800
rect 15934 0 15990 800
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18340 762 18368 2926
rect 19444 2446 19472 6054
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19996 2514 20024 4558
rect 20640 3058 20668 4966
rect 21008 3534 21036 7754
rect 21652 7750 21680 7958
rect 21456 7744 21508 7750
rect 21456 7686 21508 7692
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21468 7206 21496 7686
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21272 4480 21324 4486
rect 21272 4422 21324 4428
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 21008 2990 21036 3470
rect 21284 3058 21312 4422
rect 21364 3460 21416 3466
rect 21364 3402 21416 3408
rect 21272 3052 21324 3058
rect 21272 2994 21324 3000
rect 20996 2984 21048 2990
rect 20996 2926 21048 2932
rect 21376 2854 21404 3402
rect 21468 3398 21496 4422
rect 21652 3942 21680 7686
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 21744 4690 21772 6598
rect 21732 4684 21784 4690
rect 21732 4626 21784 4632
rect 21836 4486 21864 9318
rect 21928 8090 21956 12786
rect 22112 12374 22140 12951
rect 22192 12844 22244 12850
rect 22296 12832 22324 15302
rect 22664 14414 22692 16186
rect 22756 14550 22784 16510
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 22928 16448 22980 16454
rect 22928 16390 22980 16396
rect 22848 15162 22876 16390
rect 22940 16114 22968 16390
rect 23400 16250 23428 17070
rect 23676 16833 23704 17190
rect 23662 16824 23718 16833
rect 23662 16759 23718 16768
rect 23664 16448 23716 16454
rect 23664 16390 23716 16396
rect 23388 16244 23440 16250
rect 23388 16186 23440 16192
rect 22928 16108 22980 16114
rect 22928 16050 22980 16056
rect 23480 16108 23532 16114
rect 23480 16050 23532 16056
rect 23388 16040 23440 16046
rect 23388 15982 23440 15988
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22836 15156 22888 15162
rect 22836 15098 22888 15104
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22744 14544 22796 14550
rect 22744 14486 22796 14492
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 22756 13530 22784 14486
rect 23020 14408 23072 14414
rect 23020 14350 23072 14356
rect 23032 14006 23060 14350
rect 23020 14000 23072 14006
rect 23020 13942 23072 13948
rect 22836 13728 22888 13734
rect 22836 13670 22888 13676
rect 22744 13524 22796 13530
rect 22744 13466 22796 13472
rect 22560 13456 22612 13462
rect 22560 13398 22612 13404
rect 22244 12804 22324 12832
rect 22192 12786 22244 12792
rect 22100 12368 22152 12374
rect 22100 12310 22152 12316
rect 22204 12102 22232 12786
rect 22572 12442 22600 13398
rect 22848 13394 22876 13670
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22836 13388 22888 13394
rect 22836 13330 22888 13336
rect 22836 13252 22888 13258
rect 22836 13194 22888 13200
rect 22742 12880 22798 12889
rect 22742 12815 22798 12824
rect 22756 12782 22784 12815
rect 22744 12776 22796 12782
rect 22744 12718 22796 12724
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 22558 12336 22614 12345
rect 22284 12300 22336 12306
rect 22558 12271 22614 12280
rect 22284 12242 22336 12248
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 22296 11694 22324 12242
rect 22572 12102 22600 12271
rect 22756 12238 22784 12718
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22560 12096 22612 12102
rect 22560 12038 22612 12044
rect 22572 11898 22600 12038
rect 22560 11892 22612 11898
rect 22560 11834 22612 11840
rect 22468 11756 22520 11762
rect 22468 11698 22520 11704
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22480 11558 22508 11698
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22480 11354 22508 11494
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22376 11008 22428 11014
rect 22376 10950 22428 10956
rect 22284 10736 22336 10742
rect 22284 10678 22336 10684
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 22020 9926 22048 10542
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 22008 9444 22060 9450
rect 22008 9386 22060 9392
rect 22020 8974 22048 9386
rect 22112 9178 22140 10406
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 22020 8498 22048 8910
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 22020 7206 22048 8434
rect 22112 8430 22140 9114
rect 22204 8922 22232 10202
rect 22296 9722 22324 10678
rect 22388 10470 22416 10950
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 22480 9994 22508 11290
rect 22652 11008 22704 11014
rect 22652 10950 22704 10956
rect 22664 10810 22692 10950
rect 22848 10826 22876 13194
rect 22926 13016 22982 13025
rect 22926 12951 22928 12960
rect 22980 12951 22982 12960
rect 22928 12922 22980 12928
rect 23020 12844 23072 12850
rect 23020 12786 23072 12792
rect 23032 12753 23060 12786
rect 23018 12744 23074 12753
rect 23018 12679 23074 12688
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23308 11354 23336 14962
rect 23400 12986 23428 15982
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23492 12374 23520 16050
rect 23572 14952 23624 14958
rect 23572 14894 23624 14900
rect 23584 12782 23612 14894
rect 23676 13530 23704 16390
rect 23768 15162 23796 17478
rect 24044 17338 24072 21966
rect 24136 21146 24164 26200
rect 24780 24818 24808 26200
rect 24768 24812 24820 24818
rect 24768 24754 24820 24760
rect 25424 24206 25452 26200
rect 25780 24336 25832 24342
rect 25778 24304 25780 24313
rect 25832 24304 25834 24313
rect 26160 24290 26188 26302
rect 26698 26302 27016 26330
rect 26698 26200 26754 26302
rect 26332 24676 26384 24682
rect 26332 24618 26384 24624
rect 26424 24676 26476 24682
rect 26424 24618 26476 24624
rect 26160 24262 26280 24290
rect 25778 24239 25834 24248
rect 26252 24206 26280 24262
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 26240 24200 26292 24206
rect 26240 24142 26292 24148
rect 26344 24154 26372 24618
rect 26436 24410 26464 24618
rect 26424 24404 26476 24410
rect 26424 24346 26476 24352
rect 26606 24168 26662 24177
rect 25320 24132 25372 24138
rect 25320 24074 25372 24080
rect 24676 24064 24728 24070
rect 24676 24006 24728 24012
rect 24400 23520 24452 23526
rect 24400 23462 24452 23468
rect 24412 22642 24440 23462
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24216 22500 24268 22506
rect 24216 22442 24268 22448
rect 24124 21140 24176 21146
rect 24124 21082 24176 21088
rect 24136 20942 24164 21082
rect 24124 20936 24176 20942
rect 24124 20878 24176 20884
rect 24124 20800 24176 20806
rect 24124 20742 24176 20748
rect 24136 19553 24164 20742
rect 24228 20398 24256 22442
rect 24492 22432 24544 22438
rect 24492 22374 24544 22380
rect 24504 22137 24532 22374
rect 24688 22234 24716 24006
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 24872 23186 24900 23462
rect 25136 23316 25188 23322
rect 25136 23258 25188 23264
rect 24860 23180 24912 23186
rect 24860 23122 24912 23128
rect 24768 23044 24820 23050
rect 24768 22986 24820 22992
rect 24780 22545 24808 22986
rect 24860 22704 24912 22710
rect 24860 22646 24912 22652
rect 24766 22536 24822 22545
rect 24766 22471 24822 22480
rect 24676 22228 24728 22234
rect 24676 22170 24728 22176
rect 24872 22166 24900 22646
rect 24952 22500 25004 22506
rect 24952 22442 25004 22448
rect 24964 22166 24992 22442
rect 25148 22409 25176 23258
rect 25332 22982 25360 24074
rect 25424 23322 25452 24142
rect 26344 24126 26556 24154
rect 25872 23792 25924 23798
rect 25872 23734 25924 23740
rect 25412 23316 25464 23322
rect 25412 23258 25464 23264
rect 25688 23112 25740 23118
rect 25688 23054 25740 23060
rect 25320 22976 25372 22982
rect 25318 22944 25320 22953
rect 25412 22976 25464 22982
rect 25372 22944 25374 22953
rect 25412 22918 25464 22924
rect 25318 22879 25374 22888
rect 25134 22400 25190 22409
rect 25134 22335 25190 22344
rect 24860 22160 24912 22166
rect 24490 22128 24546 22137
rect 24860 22102 24912 22108
rect 24952 22160 25004 22166
rect 24952 22102 25004 22108
rect 25424 22098 25452 22918
rect 25504 22772 25556 22778
rect 25504 22714 25556 22720
rect 24490 22063 24546 22072
rect 25412 22092 25464 22098
rect 24504 21486 24532 22063
rect 25412 22034 25464 22040
rect 25320 22024 25372 22030
rect 25320 21966 25372 21972
rect 24584 21956 24636 21962
rect 24584 21898 24636 21904
rect 24952 21956 25004 21962
rect 24952 21898 25004 21904
rect 24492 21480 24544 21486
rect 24492 21422 24544 21428
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 24122 19544 24178 19553
rect 24122 19479 24178 19488
rect 24124 18760 24176 18766
rect 24124 18702 24176 18708
rect 24136 18358 24164 18702
rect 24124 18352 24176 18358
rect 24124 18294 24176 18300
rect 24032 17332 24084 17338
rect 24032 17274 24084 17280
rect 24136 17270 24164 18294
rect 24124 17264 24176 17270
rect 24124 17206 24176 17212
rect 24032 15632 24084 15638
rect 24032 15574 24084 15580
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23860 13274 23888 14214
rect 23940 13864 23992 13870
rect 23940 13806 23992 13812
rect 23676 13246 23888 13274
rect 23676 13190 23704 13246
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 23848 13184 23900 13190
rect 23848 13126 23900 13132
rect 23572 12776 23624 12782
rect 23572 12718 23624 12724
rect 23860 12646 23888 13126
rect 23848 12640 23900 12646
rect 23848 12582 23900 12588
rect 23480 12368 23532 12374
rect 23480 12310 23532 12316
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23756 11212 23808 11218
rect 23756 11154 23808 11160
rect 22848 10810 22968 10826
rect 22652 10804 22704 10810
rect 22848 10804 22980 10810
rect 22848 10798 22928 10804
rect 22652 10746 22704 10752
rect 22928 10746 22980 10752
rect 23768 10538 23796 11154
rect 23756 10532 23808 10538
rect 23756 10474 23808 10480
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23480 10192 23532 10198
rect 23480 10134 23532 10140
rect 22468 9988 22520 9994
rect 22468 9930 22520 9936
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22480 9178 22508 9930
rect 23492 9654 23520 10134
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 22652 9580 22704 9586
rect 22652 9522 22704 9528
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 22204 8894 22324 8922
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 22204 7886 22232 8774
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 22296 7546 22324 8894
rect 22468 8356 22520 8362
rect 22520 8316 22600 8344
rect 22468 8298 22520 8304
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 22388 7410 22416 7686
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 21824 4480 21876 4486
rect 21824 4422 21876 4428
rect 21640 3936 21692 3942
rect 21640 3878 21692 3884
rect 22020 3738 22048 7142
rect 22388 6866 22416 7346
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 22112 4214 22140 4558
rect 22100 4208 22152 4214
rect 22100 4150 22152 4156
rect 22008 3732 22060 3738
rect 22008 3674 22060 3680
rect 22020 3466 22048 3674
rect 22008 3460 22060 3466
rect 22008 3402 22060 3408
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 21456 3188 21508 3194
rect 21456 3130 21508 3136
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 20180 800 20208 2450
rect 21468 2378 21496 3130
rect 22112 3040 22140 4150
rect 22192 3052 22244 3058
rect 22112 3012 22192 3040
rect 22192 2994 22244 3000
rect 22204 2922 22232 2994
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 22112 2446 22140 2858
rect 22480 2774 22508 7686
rect 22572 7342 22600 8316
rect 22664 8022 22692 9522
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 23388 9036 23440 9042
rect 23492 9024 23520 9590
rect 23768 9466 23796 10474
rect 23860 9704 23888 12582
rect 23952 11082 23980 13806
rect 24044 13258 24072 15574
rect 24228 14958 24256 20334
rect 24490 20224 24546 20233
rect 24490 20159 24546 20168
rect 24504 19446 24532 20159
rect 24596 19922 24624 21898
rect 24964 21457 24992 21898
rect 25044 21616 25096 21622
rect 25044 21558 25096 21564
rect 24950 21448 25006 21457
rect 24688 21406 24900 21434
rect 24688 21350 24716 21406
rect 24676 21344 24728 21350
rect 24872 21332 24900 21406
rect 24950 21383 25006 21392
rect 25056 21332 25084 21558
rect 25136 21412 25188 21418
rect 25136 21354 25188 21360
rect 24872 21304 25084 21332
rect 24676 21286 24728 21292
rect 24584 19916 24636 19922
rect 24584 19858 24636 19864
rect 25044 19916 25096 19922
rect 25044 19858 25096 19864
rect 25056 19689 25084 19858
rect 25042 19680 25098 19689
rect 25042 19615 25098 19624
rect 24492 19440 24544 19446
rect 24492 19382 24544 19388
rect 24860 19440 24912 19446
rect 24860 19382 24912 19388
rect 24872 19310 24900 19382
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 24952 19304 25004 19310
rect 24952 19246 25004 19252
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 24768 18352 24820 18358
rect 24768 18294 24820 18300
rect 24492 17604 24544 17610
rect 24492 17546 24544 17552
rect 24504 17134 24532 17546
rect 24676 17536 24728 17542
rect 24676 17478 24728 17484
rect 24492 17128 24544 17134
rect 24492 17070 24544 17076
rect 24504 16046 24532 17070
rect 24582 16824 24638 16833
rect 24582 16759 24638 16768
rect 24596 16522 24624 16759
rect 24584 16516 24636 16522
rect 24584 16458 24636 16464
rect 24688 16250 24716 17478
rect 24780 17241 24808 18294
rect 24872 17524 24900 18566
rect 24964 17746 24992 19246
rect 25056 18630 25084 19615
rect 25044 18624 25096 18630
rect 25044 18566 25096 18572
rect 25042 18320 25098 18329
rect 25042 18255 25044 18264
rect 25096 18255 25098 18264
rect 25044 18226 25096 18232
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 25056 17746 25084 18022
rect 24952 17740 25004 17746
rect 24952 17682 25004 17688
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 25044 17536 25096 17542
rect 24872 17496 25044 17524
rect 24766 17232 24822 17241
rect 24766 17167 24822 17176
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24492 16040 24544 16046
rect 24492 15982 24544 15988
rect 24780 15570 24808 16186
rect 24872 16017 24900 17496
rect 25044 17478 25096 17484
rect 25148 17066 25176 21354
rect 25228 21072 25280 21078
rect 25228 21014 25280 21020
rect 25240 20466 25268 21014
rect 25228 20460 25280 20466
rect 25228 20402 25280 20408
rect 25240 20233 25268 20402
rect 25226 20224 25282 20233
rect 25226 20159 25282 20168
rect 25228 19848 25280 19854
rect 25228 19790 25280 19796
rect 25240 18358 25268 19790
rect 25332 19334 25360 21966
rect 25412 21480 25464 21486
rect 25412 21422 25464 21428
rect 25424 20262 25452 21422
rect 25516 21146 25544 22714
rect 25504 21140 25556 21146
rect 25504 21082 25556 21088
rect 25516 20466 25544 21082
rect 25700 20602 25728 23054
rect 25884 22710 25912 23734
rect 26056 23180 26108 23186
rect 26056 23122 26108 23128
rect 26068 22982 26096 23122
rect 26240 23044 26292 23050
rect 26240 22986 26292 22992
rect 26056 22976 26108 22982
rect 26056 22918 26108 22924
rect 25872 22704 25924 22710
rect 25792 22664 25872 22692
rect 25792 22574 25820 22664
rect 25872 22646 25924 22652
rect 25780 22568 25832 22574
rect 25780 22510 25832 22516
rect 25792 21078 25820 22510
rect 26056 21956 26108 21962
rect 26056 21898 26108 21904
rect 25964 21888 26016 21894
rect 25964 21830 26016 21836
rect 25872 21548 25924 21554
rect 25872 21490 25924 21496
rect 25884 21350 25912 21490
rect 25872 21344 25924 21350
rect 25872 21286 25924 21292
rect 25780 21072 25832 21078
rect 25780 21014 25832 21020
rect 25884 20913 25912 21286
rect 25870 20904 25926 20913
rect 25976 20874 26004 21830
rect 26068 21593 26096 21898
rect 26148 21888 26200 21894
rect 26148 21830 26200 21836
rect 26054 21584 26110 21593
rect 26054 21519 26056 21528
rect 26108 21519 26110 21528
rect 26056 21490 26108 21496
rect 26160 21434 26188 21830
rect 26068 21406 26188 21434
rect 25870 20839 25926 20848
rect 25964 20868 26016 20874
rect 25964 20810 26016 20816
rect 25688 20596 25740 20602
rect 25688 20538 25740 20544
rect 25780 20596 25832 20602
rect 25780 20538 25832 20544
rect 25504 20460 25556 20466
rect 25504 20402 25556 20408
rect 25596 20392 25648 20398
rect 25596 20334 25648 20340
rect 25412 20256 25464 20262
rect 25412 20198 25464 20204
rect 25332 19306 25452 19334
rect 25608 19310 25636 20334
rect 25700 19378 25728 20538
rect 25792 20398 25820 20538
rect 25780 20392 25832 20398
rect 25780 20334 25832 20340
rect 25872 20392 25924 20398
rect 25872 20334 25924 20340
rect 25688 19372 25740 19378
rect 25688 19314 25740 19320
rect 25228 18352 25280 18358
rect 25228 18294 25280 18300
rect 25424 18057 25452 19306
rect 25596 19304 25648 19310
rect 25596 19246 25648 19252
rect 25594 19000 25650 19009
rect 25594 18935 25650 18944
rect 25608 18834 25636 18935
rect 25700 18834 25728 19314
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25596 18828 25648 18834
rect 25596 18770 25648 18776
rect 25688 18828 25740 18834
rect 25688 18770 25740 18776
rect 25608 18465 25636 18770
rect 25594 18456 25650 18465
rect 25792 18426 25820 19110
rect 25594 18391 25650 18400
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 25410 18048 25466 18057
rect 25410 17983 25466 17992
rect 25780 17264 25832 17270
rect 25778 17232 25780 17241
rect 25832 17232 25834 17241
rect 25596 17196 25648 17202
rect 25778 17167 25834 17176
rect 25596 17138 25648 17144
rect 25504 17128 25556 17134
rect 25504 17070 25556 17076
rect 25136 17060 25188 17066
rect 25136 17002 25188 17008
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 24858 16008 24914 16017
rect 24858 15943 24914 15952
rect 24768 15564 24820 15570
rect 24596 15524 24768 15552
rect 24216 14952 24268 14958
rect 24216 14894 24268 14900
rect 24492 14340 24544 14346
rect 24492 14282 24544 14288
rect 24400 14272 24452 14278
rect 24400 14214 24452 14220
rect 24308 13932 24360 13938
rect 24308 13874 24360 13880
rect 24032 13252 24084 13258
rect 24032 13194 24084 13200
rect 24320 12986 24348 13874
rect 24412 13394 24440 14214
rect 24504 14074 24532 14282
rect 24492 14068 24544 14074
rect 24492 14010 24544 14016
rect 24596 13802 24624 15524
rect 24768 15506 24820 15512
rect 25148 15366 25176 16390
rect 25320 15564 25372 15570
rect 25320 15506 25372 15512
rect 25136 15360 25188 15366
rect 25136 15302 25188 15308
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 24688 14550 24716 15098
rect 25148 15026 25176 15302
rect 25044 15020 25096 15026
rect 25044 14962 25096 14968
rect 25136 15020 25188 15026
rect 25136 14962 25188 14968
rect 24768 14952 24820 14958
rect 24768 14894 24820 14900
rect 24676 14544 24728 14550
rect 24676 14486 24728 14492
rect 24584 13796 24636 13802
rect 24584 13738 24636 13744
rect 24492 13456 24544 13462
rect 24688 13433 24716 14486
rect 24492 13398 24544 13404
rect 24674 13424 24730 13433
rect 24400 13388 24452 13394
rect 24400 13330 24452 13336
rect 24412 13190 24440 13330
rect 24400 13184 24452 13190
rect 24400 13126 24452 13132
rect 24308 12980 24360 12986
rect 24308 12922 24360 12928
rect 24504 12434 24532 13398
rect 24674 13359 24730 13368
rect 24584 12980 24636 12986
rect 24584 12922 24636 12928
rect 24320 12406 24532 12434
rect 24032 11552 24084 11558
rect 24032 11494 24084 11500
rect 24044 11121 24072 11494
rect 24030 11112 24086 11121
rect 23940 11076 23992 11082
rect 24030 11047 24086 11056
rect 23940 11018 23992 11024
rect 24044 11014 24072 11047
rect 24032 11008 24084 11014
rect 24032 10950 24084 10956
rect 23940 10736 23992 10742
rect 23940 10678 23992 10684
rect 23952 10198 23980 10678
rect 24044 10266 24072 10950
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24032 10260 24084 10266
rect 24032 10202 24084 10208
rect 23940 10192 23992 10198
rect 23940 10134 23992 10140
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 23860 9676 23980 9704
rect 23440 8996 23520 9024
rect 23388 8978 23440 8984
rect 23492 8838 23520 8996
rect 23676 9438 23796 9466
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23492 8634 23520 8774
rect 23480 8628 23532 8634
rect 23480 8570 23532 8576
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22652 8016 22704 8022
rect 22652 7958 22704 7964
rect 23676 7954 23704 9438
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23768 9042 23796 9318
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 22560 7336 22612 7342
rect 22560 7278 22612 7284
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22928 4684 22980 4690
rect 22928 4626 22980 4632
rect 23204 4684 23256 4690
rect 23204 4626 23256 4632
rect 22940 4146 22968 4626
rect 23216 4146 23244 4626
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 22928 4140 22980 4146
rect 22928 4082 22980 4088
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23296 4072 23348 4078
rect 23296 4014 23348 4020
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22848 3602 22876 3878
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22836 3596 22888 3602
rect 22836 3538 22888 3544
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 23112 3392 23164 3398
rect 23112 3334 23164 3340
rect 22756 2922 22784 3334
rect 23124 2938 23152 3334
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 22848 2910 23152 2938
rect 22848 2774 22876 2910
rect 23308 2854 23336 4014
rect 23584 3738 23612 4558
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 23952 3466 23980 9676
rect 24044 8974 24072 9998
rect 24136 9926 24164 10542
rect 24320 10266 24348 12406
rect 24400 12300 24452 12306
rect 24400 12242 24452 12248
rect 24412 11558 24440 12242
rect 24596 12238 24624 12922
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24492 11824 24544 11830
rect 24596 11812 24624 12174
rect 24544 11784 24624 11812
rect 24492 11766 24544 11772
rect 24400 11552 24452 11558
rect 24400 11494 24452 11500
rect 24412 11218 24440 11494
rect 24400 11212 24452 11218
rect 24400 11154 24452 11160
rect 24596 11150 24624 11784
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24308 10260 24360 10266
rect 24308 10202 24360 10208
rect 24124 9920 24176 9926
rect 24124 9862 24176 9868
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 24044 8498 24072 8910
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 24136 4826 24164 9862
rect 24320 9518 24348 10202
rect 24596 9636 24624 11086
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 24688 10606 24716 10950
rect 24676 10600 24728 10606
rect 24676 10542 24728 10548
rect 24780 10538 24808 14894
rect 25056 14822 25084 14962
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 24860 13252 24912 13258
rect 24860 13194 24912 13200
rect 24872 12918 24900 13194
rect 24860 12912 24912 12918
rect 24860 12854 24912 12860
rect 24952 12776 25004 12782
rect 24952 12718 25004 12724
rect 24964 12306 24992 12718
rect 24952 12300 25004 12306
rect 24952 12242 25004 12248
rect 25056 12186 25084 14758
rect 25136 14272 25188 14278
rect 25136 14214 25188 14220
rect 25148 13326 25176 14214
rect 25332 14074 25360 15506
rect 25412 15020 25464 15026
rect 25412 14962 25464 14968
rect 25320 14068 25372 14074
rect 25320 14010 25372 14016
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 25332 12918 25360 14010
rect 25320 12912 25372 12918
rect 25320 12854 25372 12860
rect 25332 12322 25360 12854
rect 24872 12158 25084 12186
rect 25240 12294 25360 12322
rect 24872 11801 24900 12158
rect 24858 11792 24914 11801
rect 24858 11727 24914 11736
rect 24768 10532 24820 10538
rect 24768 10474 24820 10480
rect 24676 9648 24728 9654
rect 24596 9608 24676 9636
rect 24676 9590 24728 9596
rect 24308 9512 24360 9518
rect 24308 9454 24360 9460
rect 24124 4820 24176 4826
rect 24124 4762 24176 4768
rect 24872 4078 24900 11727
rect 25240 11354 25268 12294
rect 25228 11348 25280 11354
rect 25228 11290 25280 11296
rect 25424 9382 25452 14962
rect 25516 14618 25544 17070
rect 25504 14612 25556 14618
rect 25504 14554 25556 14560
rect 25516 14074 25544 14554
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25608 13530 25636 17138
rect 25778 16824 25834 16833
rect 25778 16759 25834 16768
rect 25792 16182 25820 16759
rect 25884 16658 25912 20334
rect 26068 19281 26096 21406
rect 26252 21350 26280 22986
rect 26332 22976 26384 22982
rect 26332 22918 26384 22924
rect 26344 22710 26372 22918
rect 26332 22704 26384 22710
rect 26332 22646 26384 22652
rect 26528 22522 26556 24126
rect 26606 24103 26608 24112
rect 26660 24103 26662 24112
rect 26608 24074 26660 24080
rect 26988 24070 27016 26302
rect 27342 26200 27398 27000
rect 27986 26330 28042 27000
rect 27986 26302 28396 26330
rect 27986 26200 28042 26302
rect 27252 24744 27304 24750
rect 27252 24686 27304 24692
rect 27264 24410 27292 24686
rect 27252 24404 27304 24410
rect 27252 24346 27304 24352
rect 27356 24274 27384 26200
rect 27344 24268 27396 24274
rect 27344 24210 27396 24216
rect 27252 24132 27304 24138
rect 27252 24074 27304 24080
rect 27344 24132 27396 24138
rect 27344 24074 27396 24080
rect 26976 24064 27028 24070
rect 26976 24006 27028 24012
rect 26608 23656 26660 23662
rect 26608 23598 26660 23604
rect 26620 22778 26648 23598
rect 27264 23050 27292 24074
rect 27252 23044 27304 23050
rect 27252 22986 27304 22992
rect 26608 22772 26660 22778
rect 26608 22714 26660 22720
rect 26620 22642 26648 22714
rect 27264 22710 27292 22986
rect 27252 22704 27304 22710
rect 27252 22646 27304 22652
rect 26608 22636 26660 22642
rect 26608 22578 26660 22584
rect 27264 22574 27292 22646
rect 27252 22568 27304 22574
rect 26528 22494 26924 22522
rect 27252 22510 27304 22516
rect 27356 22506 27384 24074
rect 27804 24064 27856 24070
rect 27804 24006 27856 24012
rect 27712 23792 27764 23798
rect 27712 23734 27764 23740
rect 27620 22704 27672 22710
rect 27620 22646 27672 22652
rect 27632 22574 27660 22646
rect 27724 22574 27752 23734
rect 27816 23730 27844 24006
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 27896 23860 27948 23866
rect 27896 23802 27948 23808
rect 27804 23724 27856 23730
rect 27804 23666 27856 23672
rect 27804 23520 27856 23526
rect 27804 23462 27856 23468
rect 27620 22568 27672 22574
rect 27620 22510 27672 22516
rect 27712 22568 27764 22574
rect 27712 22510 27764 22516
rect 26332 22432 26384 22438
rect 26332 22374 26384 22380
rect 26608 22432 26660 22438
rect 26608 22374 26660 22380
rect 26344 22098 26372 22374
rect 26332 22092 26384 22098
rect 26332 22034 26384 22040
rect 26620 22030 26648 22374
rect 26700 22160 26752 22166
rect 26700 22102 26752 22108
rect 26608 22024 26660 22030
rect 26608 21966 26660 21972
rect 26332 21956 26384 21962
rect 26384 21916 26464 21944
rect 26332 21898 26384 21904
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 26148 21072 26200 21078
rect 26148 21014 26200 21020
rect 26160 20806 26188 21014
rect 26240 21004 26292 21010
rect 26240 20946 26292 20952
rect 26332 21004 26384 21010
rect 26332 20946 26384 20952
rect 26148 20800 26200 20806
rect 26148 20742 26200 20748
rect 26252 20346 26280 20946
rect 26344 20602 26372 20946
rect 26332 20596 26384 20602
rect 26332 20538 26384 20544
rect 26148 20324 26200 20330
rect 26252 20318 26372 20346
rect 26148 20266 26200 20272
rect 26160 19961 26188 20266
rect 26344 20262 26372 20318
rect 26240 20256 26292 20262
rect 26240 20198 26292 20204
rect 26332 20256 26384 20262
rect 26332 20198 26384 20204
rect 26146 19952 26202 19961
rect 26146 19887 26202 19896
rect 26160 19514 26188 19887
rect 26252 19514 26280 20198
rect 26330 19952 26386 19961
rect 26330 19887 26386 19896
rect 26344 19718 26372 19887
rect 26332 19712 26384 19718
rect 26332 19654 26384 19660
rect 26148 19508 26200 19514
rect 26148 19450 26200 19456
rect 26240 19508 26292 19514
rect 26240 19450 26292 19456
rect 26054 19272 26110 19281
rect 26054 19207 26110 19216
rect 26332 18624 26384 18630
rect 26332 18566 26384 18572
rect 25962 18320 26018 18329
rect 26344 18290 26372 18566
rect 25962 18255 26018 18264
rect 26332 18284 26384 18290
rect 25976 17270 26004 18255
rect 26332 18226 26384 18232
rect 26330 18184 26386 18193
rect 26056 18148 26108 18154
rect 26330 18119 26386 18128
rect 26056 18090 26108 18096
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 26068 16726 26096 18090
rect 26344 17814 26372 18119
rect 26332 17808 26384 17814
rect 26332 17750 26384 17756
rect 26148 17264 26200 17270
rect 26148 17206 26200 17212
rect 26056 16720 26108 16726
rect 26056 16662 26108 16668
rect 25872 16652 25924 16658
rect 25872 16594 25924 16600
rect 25780 16176 25832 16182
rect 25686 16144 25742 16153
rect 25780 16118 25832 16124
rect 25686 16079 25742 16088
rect 25700 15434 25728 16079
rect 25688 15428 25740 15434
rect 25688 15370 25740 15376
rect 25700 15026 25728 15370
rect 25688 15020 25740 15026
rect 25688 14962 25740 14968
rect 25688 14816 25740 14822
rect 25688 14758 25740 14764
rect 25596 13524 25648 13530
rect 25596 13466 25648 13472
rect 25700 12646 25728 14758
rect 25792 14346 25820 16118
rect 26056 16040 26108 16046
rect 26160 16028 26188 17206
rect 26344 17202 26372 17750
rect 26436 17746 26464 21916
rect 26712 19786 26740 22102
rect 26792 20868 26844 20874
rect 26792 20810 26844 20816
rect 26804 20058 26832 20810
rect 26896 20806 26924 22494
rect 27344 22500 27396 22506
rect 27344 22442 27396 22448
rect 27620 22092 27672 22098
rect 27620 22034 27672 22040
rect 27712 22092 27764 22098
rect 27712 22034 27764 22040
rect 27632 22001 27660 22034
rect 27618 21992 27674 22001
rect 27618 21927 27674 21936
rect 27724 21876 27752 22034
rect 27816 22030 27844 23462
rect 27908 23322 27936 23802
rect 28264 23792 28316 23798
rect 28264 23734 28316 23740
rect 27896 23316 27948 23322
rect 27896 23258 27948 23264
rect 28276 23254 28304 23734
rect 28368 23662 28396 26302
rect 28630 26200 28686 27000
rect 29274 26330 29330 27000
rect 29274 26302 29868 26330
rect 29274 26200 29330 26302
rect 28644 24342 28672 26200
rect 29840 24614 29868 26302
rect 29918 26200 29974 27000
rect 30562 26200 30618 27000
rect 31206 26200 31262 27000
rect 31850 26200 31906 27000
rect 32494 26200 32550 27000
rect 33138 26200 33194 27000
rect 33782 26330 33838 27000
rect 33782 26302 34008 26330
rect 33782 26200 33838 26302
rect 29932 24750 29960 26200
rect 30576 25294 30604 26200
rect 30564 25288 30616 25294
rect 30564 25230 30616 25236
rect 30380 24812 30432 24818
rect 30380 24754 30432 24760
rect 29920 24744 29972 24750
rect 29920 24686 29972 24692
rect 29736 24608 29788 24614
rect 29736 24550 29788 24556
rect 29828 24608 29880 24614
rect 29828 24550 29880 24556
rect 29748 24410 29776 24550
rect 30392 24410 30420 24754
rect 29736 24404 29788 24410
rect 29736 24346 29788 24352
rect 30380 24404 30432 24410
rect 30380 24346 30432 24352
rect 28632 24336 28684 24342
rect 28632 24278 28684 24284
rect 30392 24206 30420 24346
rect 31116 24268 31168 24274
rect 31116 24210 31168 24216
rect 30380 24200 30432 24206
rect 30380 24142 30432 24148
rect 28540 24064 28592 24070
rect 28540 24006 28592 24012
rect 28724 24064 28776 24070
rect 28724 24006 28776 24012
rect 30564 24064 30616 24070
rect 30564 24006 30616 24012
rect 30932 24064 30984 24070
rect 30932 24006 30984 24012
rect 28448 23860 28500 23866
rect 28448 23802 28500 23808
rect 28460 23769 28488 23802
rect 28446 23760 28502 23769
rect 28446 23695 28502 23704
rect 28356 23656 28408 23662
rect 28356 23598 28408 23604
rect 28356 23316 28408 23322
rect 28356 23258 28408 23264
rect 28264 23248 28316 23254
rect 28264 23190 28316 23196
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 27896 22704 27948 22710
rect 27896 22646 27948 22652
rect 28264 22704 28316 22710
rect 28368 22692 28396 23258
rect 28316 22664 28396 22692
rect 28264 22646 28316 22652
rect 27804 22024 27856 22030
rect 27804 21966 27856 21972
rect 27908 21876 27936 22646
rect 28080 22568 28132 22574
rect 28080 22510 28132 22516
rect 28356 22568 28408 22574
rect 28356 22510 28408 22516
rect 28092 22098 28120 22510
rect 28262 22264 28318 22273
rect 28262 22199 28264 22208
rect 28316 22199 28318 22208
rect 28264 22170 28316 22176
rect 28080 22092 28132 22098
rect 28080 22034 28132 22040
rect 27540 21848 27752 21876
rect 27816 21848 27936 21876
rect 27068 21684 27120 21690
rect 27068 21626 27120 21632
rect 27436 21684 27488 21690
rect 27436 21626 27488 21632
rect 27080 21146 27108 21626
rect 27068 21140 27120 21146
rect 27068 21082 27120 21088
rect 27448 21049 27476 21626
rect 27434 21040 27490 21049
rect 27434 20975 27490 20984
rect 26976 20936 27028 20942
rect 26976 20878 27028 20884
rect 26884 20800 26936 20806
rect 26884 20742 26936 20748
rect 26988 20534 27016 20878
rect 27448 20874 27476 20975
rect 27436 20868 27488 20874
rect 27436 20810 27488 20816
rect 27160 20800 27212 20806
rect 27160 20742 27212 20748
rect 26976 20528 27028 20534
rect 26976 20470 27028 20476
rect 26792 20052 26844 20058
rect 26792 19994 26844 20000
rect 26988 19922 27016 20470
rect 27068 20052 27120 20058
rect 27068 19994 27120 20000
rect 26976 19916 27028 19922
rect 26976 19858 27028 19864
rect 26700 19780 26752 19786
rect 26700 19722 26752 19728
rect 26712 19553 26740 19722
rect 27080 19718 27108 19994
rect 27068 19712 27120 19718
rect 27068 19654 27120 19660
rect 27172 19700 27200 20742
rect 27252 20256 27304 20262
rect 27252 20198 27304 20204
rect 27264 19854 27292 20198
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 27252 19712 27304 19718
rect 27172 19672 27252 19700
rect 26698 19544 26754 19553
rect 26698 19479 26754 19488
rect 27080 18834 27108 19654
rect 27068 18828 27120 18834
rect 27068 18770 27120 18776
rect 27172 18306 27200 19672
rect 27252 19654 27304 19660
rect 27344 19508 27396 19514
rect 27344 19450 27396 19456
rect 27436 19508 27488 19514
rect 27436 19450 27488 19456
rect 27252 19168 27304 19174
rect 27252 19110 27304 19116
rect 27264 18426 27292 19110
rect 27252 18420 27304 18426
rect 27252 18362 27304 18368
rect 27172 18278 27292 18306
rect 26516 18216 26568 18222
rect 26516 18158 26568 18164
rect 26608 18216 26660 18222
rect 26608 18158 26660 18164
rect 26424 17740 26476 17746
rect 26424 17682 26476 17688
rect 26528 17610 26556 18158
rect 26516 17604 26568 17610
rect 26516 17546 26568 17552
rect 26332 17196 26384 17202
rect 26332 17138 26384 17144
rect 26516 17060 26568 17066
rect 26516 17002 26568 17008
rect 26424 16652 26476 16658
rect 26424 16594 26476 16600
rect 26108 16000 26188 16028
rect 26056 15982 26108 15988
rect 25872 15360 25924 15366
rect 26068 15337 26096 15982
rect 26332 15428 26384 15434
rect 26332 15370 26384 15376
rect 26240 15360 26292 15366
rect 25872 15302 25924 15308
rect 26054 15328 26110 15337
rect 25884 15094 25912 15302
rect 26240 15302 26292 15308
rect 26054 15263 26110 15272
rect 25872 15088 25924 15094
rect 25872 15030 25924 15036
rect 25780 14340 25832 14346
rect 25780 14282 25832 14288
rect 25792 14006 25820 14282
rect 25780 14000 25832 14006
rect 25780 13942 25832 13948
rect 25792 13530 25820 13942
rect 25780 13524 25832 13530
rect 25780 13466 25832 13472
rect 25792 13258 25820 13466
rect 25780 13252 25832 13258
rect 25780 13194 25832 13200
rect 26056 13252 26108 13258
rect 26056 13194 26108 13200
rect 25792 12986 25820 13194
rect 26068 13161 26096 13194
rect 26054 13152 26110 13161
rect 26054 13087 26110 13096
rect 26252 13025 26280 15302
rect 26344 14618 26372 15370
rect 26332 14612 26384 14618
rect 26332 14554 26384 14560
rect 26436 14498 26464 16594
rect 26528 14618 26556 17002
rect 26620 16250 26648 18158
rect 27160 18080 27212 18086
rect 27160 18022 27212 18028
rect 26976 17536 27028 17542
rect 26976 17478 27028 17484
rect 27068 17536 27120 17542
rect 27068 17478 27120 17484
rect 26790 16824 26846 16833
rect 26790 16759 26846 16768
rect 26804 16522 26832 16759
rect 26792 16516 26844 16522
rect 26792 16458 26844 16464
rect 26804 16250 26832 16458
rect 26988 16250 27016 17478
rect 27080 16658 27108 17478
rect 27068 16652 27120 16658
rect 27068 16594 27120 16600
rect 26608 16244 26660 16250
rect 26608 16186 26660 16192
rect 26792 16244 26844 16250
rect 26792 16186 26844 16192
rect 26976 16244 27028 16250
rect 26976 16186 27028 16192
rect 26884 16040 26936 16046
rect 26884 15982 26936 15988
rect 26700 15904 26752 15910
rect 26700 15846 26752 15852
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26516 14612 26568 14618
rect 26516 14554 26568 14560
rect 26344 14470 26464 14498
rect 26344 13734 26372 14470
rect 26332 13728 26384 13734
rect 26332 13670 26384 13676
rect 26516 13184 26568 13190
rect 26516 13126 26568 13132
rect 26238 13016 26294 13025
rect 25780 12980 25832 12986
rect 26528 12986 26556 13126
rect 26238 12951 26240 12960
rect 25780 12922 25832 12928
rect 26292 12951 26294 12960
rect 26516 12980 26568 12986
rect 26240 12922 26292 12928
rect 26516 12922 26568 12928
rect 26422 12880 26478 12889
rect 26422 12815 26424 12824
rect 26476 12815 26478 12824
rect 26424 12786 26476 12792
rect 25962 12744 26018 12753
rect 25962 12679 26018 12688
rect 25976 12646 26004 12679
rect 25688 12640 25740 12646
rect 25688 12582 25740 12588
rect 25964 12640 26016 12646
rect 25964 12582 26016 12588
rect 25504 12096 25556 12102
rect 25504 12038 25556 12044
rect 25516 11762 25544 12038
rect 25504 11756 25556 11762
rect 25504 11698 25556 11704
rect 25780 11756 25832 11762
rect 25780 11698 25832 11704
rect 25516 11082 25544 11698
rect 25504 11076 25556 11082
rect 25504 11018 25556 11024
rect 25516 10810 25544 11018
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 25516 9994 25544 10746
rect 25792 10538 25820 11698
rect 25780 10532 25832 10538
rect 25780 10474 25832 10480
rect 25504 9988 25556 9994
rect 25504 9930 25556 9936
rect 25976 9602 26004 12582
rect 26332 12368 26384 12374
rect 26332 12310 26384 12316
rect 26344 11694 26372 12310
rect 26528 12238 26556 12922
rect 26516 12232 26568 12238
rect 26516 12174 26568 12180
rect 26332 11688 26384 11694
rect 26332 11630 26384 11636
rect 26620 11354 26648 15506
rect 26712 12442 26740 15846
rect 26790 15600 26846 15609
rect 26790 15535 26846 15544
rect 26804 15366 26832 15535
rect 26792 15360 26844 15366
rect 26792 15302 26844 15308
rect 26700 12436 26752 12442
rect 26700 12378 26752 12384
rect 26896 12374 26924 15982
rect 27172 15620 27200 18022
rect 27264 15910 27292 18278
rect 27252 15904 27304 15910
rect 27252 15846 27304 15852
rect 27356 15858 27384 19450
rect 27448 19310 27476 19450
rect 27436 19304 27488 19310
rect 27436 19246 27488 19252
rect 27540 19009 27568 21848
rect 27816 21185 27844 21848
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 27896 21548 27948 21554
rect 27896 21490 27948 21496
rect 27802 21176 27858 21185
rect 27802 21111 27858 21120
rect 27620 20800 27672 20806
rect 27620 20742 27672 20748
rect 27632 19990 27660 20742
rect 27816 20534 27844 21111
rect 27908 21010 27936 21490
rect 27896 21004 27948 21010
rect 27896 20946 27948 20952
rect 28368 20874 28396 22510
rect 28552 21026 28580 24006
rect 28736 22234 28764 24006
rect 30380 23724 30432 23730
rect 30380 23666 30432 23672
rect 29368 23656 29420 23662
rect 29368 23598 29420 23604
rect 30194 23624 30250 23633
rect 29092 23520 29144 23526
rect 29092 23462 29144 23468
rect 28724 22228 28776 22234
rect 28724 22170 28776 22176
rect 28908 22092 28960 22098
rect 28908 22034 28960 22040
rect 28920 21486 28948 22034
rect 28816 21480 28868 21486
rect 28814 21448 28816 21457
rect 28908 21480 28960 21486
rect 28868 21448 28870 21457
rect 28908 21422 28960 21428
rect 28814 21383 28870 21392
rect 28460 20998 28580 21026
rect 28356 20868 28408 20874
rect 28356 20810 28408 20816
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 27804 20528 27856 20534
rect 27804 20470 27856 20476
rect 27620 19984 27672 19990
rect 27620 19926 27672 19932
rect 27620 19712 27672 19718
rect 27620 19654 27672 19660
rect 27526 19000 27582 19009
rect 27632 18970 27660 19654
rect 27710 19544 27766 19553
rect 27710 19479 27766 19488
rect 27816 19496 27844 20470
rect 28460 20074 28488 20998
rect 28724 20800 28776 20806
rect 28724 20742 28776 20748
rect 28632 20324 28684 20330
rect 28632 20266 28684 20272
rect 28460 20046 28580 20074
rect 27988 19984 28040 19990
rect 27986 19952 27988 19961
rect 28040 19952 28042 19961
rect 28446 19952 28502 19961
rect 27986 19887 28042 19896
rect 28356 19916 28408 19922
rect 28446 19887 28502 19896
rect 28356 19858 28408 19864
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 28368 19514 28396 19858
rect 28356 19508 28408 19514
rect 27724 19428 27752 19479
rect 27816 19468 28028 19496
rect 27724 19400 27844 19428
rect 27526 18935 27582 18944
rect 27620 18964 27672 18970
rect 27620 18906 27672 18912
rect 27712 18964 27764 18970
rect 27712 18906 27764 18912
rect 27436 18828 27488 18834
rect 27436 18770 27488 18776
rect 27448 17678 27476 18770
rect 27620 18624 27672 18630
rect 27620 18566 27672 18572
rect 27528 18080 27580 18086
rect 27528 18022 27580 18028
rect 27436 17672 27488 17678
rect 27436 17614 27488 17620
rect 27448 16833 27476 17614
rect 27540 17542 27568 18022
rect 27528 17536 27580 17542
rect 27528 17478 27580 17484
rect 27632 17270 27660 18566
rect 27724 18426 27752 18906
rect 27712 18420 27764 18426
rect 27712 18362 27764 18368
rect 27710 17368 27766 17377
rect 27816 17338 27844 19400
rect 28000 18834 28028 19468
rect 28356 19450 28408 19456
rect 28354 19408 28410 19417
rect 28460 19378 28488 19887
rect 28354 19343 28410 19352
rect 28448 19372 28500 19378
rect 28080 19304 28132 19310
rect 28080 19246 28132 19252
rect 27988 18828 28040 18834
rect 27988 18770 28040 18776
rect 28092 18766 28120 19246
rect 28080 18760 28132 18766
rect 28080 18702 28132 18708
rect 28092 18630 28120 18702
rect 28080 18624 28132 18630
rect 28080 18566 28132 18572
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 27710 17303 27712 17312
rect 27764 17303 27766 17312
rect 27804 17332 27856 17338
rect 27712 17274 27764 17280
rect 27804 17274 27856 17280
rect 27620 17264 27672 17270
rect 27620 17206 27672 17212
rect 28262 17232 28318 17241
rect 27712 17196 27764 17202
rect 28262 17167 28318 17176
rect 27712 17138 27764 17144
rect 27724 17105 27752 17138
rect 27710 17096 27766 17105
rect 27528 17060 27580 17066
rect 27710 17031 27766 17040
rect 27528 17002 27580 17008
rect 27434 16824 27490 16833
rect 27434 16759 27490 16768
rect 27436 16652 27488 16658
rect 27436 16594 27488 16600
rect 27448 16250 27476 16594
rect 27436 16244 27488 16250
rect 27436 16186 27488 16192
rect 27356 15830 27476 15858
rect 27172 15592 27384 15620
rect 27356 15502 27384 15592
rect 27344 15496 27396 15502
rect 27066 15464 27122 15473
rect 26988 15434 27066 15450
rect 26976 15428 27066 15434
rect 27028 15422 27066 15428
rect 27344 15438 27396 15444
rect 27066 15399 27122 15408
rect 26976 15370 27028 15376
rect 27080 15094 27108 15399
rect 27160 15360 27212 15366
rect 27158 15328 27160 15337
rect 27212 15328 27214 15337
rect 27158 15263 27214 15272
rect 27068 15088 27120 15094
rect 27068 15030 27120 15036
rect 27068 14340 27120 14346
rect 27068 14282 27120 14288
rect 27080 14006 27108 14282
rect 27068 14000 27120 14006
rect 27068 13942 27120 13948
rect 27080 13394 27108 13942
rect 27068 13388 27120 13394
rect 27068 13330 27120 13336
rect 27172 12850 27200 15263
rect 27250 15056 27306 15065
rect 27250 14991 27252 15000
rect 27304 14991 27306 15000
rect 27252 14962 27304 14968
rect 27344 14952 27396 14958
rect 27264 14900 27344 14906
rect 27264 14894 27396 14900
rect 27264 14878 27384 14894
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 26884 12368 26936 12374
rect 26884 12310 26936 12316
rect 27160 12300 27212 12306
rect 27160 12242 27212 12248
rect 27068 11756 27120 11762
rect 27068 11698 27120 11704
rect 26608 11348 26660 11354
rect 26608 11290 26660 11296
rect 26056 10668 26108 10674
rect 26056 10610 26108 10616
rect 26068 9722 26096 10610
rect 26620 10606 26648 11290
rect 26884 11144 26936 11150
rect 26884 11086 26936 11092
rect 26700 10804 26752 10810
rect 26700 10746 26752 10752
rect 26608 10600 26660 10606
rect 26608 10542 26660 10548
rect 26240 10532 26292 10538
rect 26240 10474 26292 10480
rect 26252 10169 26280 10474
rect 26620 10198 26648 10542
rect 26712 10266 26740 10746
rect 26700 10260 26752 10266
rect 26700 10202 26752 10208
rect 26608 10192 26660 10198
rect 26238 10160 26294 10169
rect 26608 10134 26660 10140
rect 26238 10095 26294 10104
rect 26712 9926 26740 10202
rect 26896 10130 26924 11086
rect 26884 10124 26936 10130
rect 26884 10066 26936 10072
rect 26700 9920 26752 9926
rect 26700 9862 26752 9868
rect 26056 9716 26108 9722
rect 26056 9658 26108 9664
rect 25792 9574 26004 9602
rect 25688 9444 25740 9450
rect 25688 9386 25740 9392
rect 25412 9376 25464 9382
rect 25412 9318 25464 9324
rect 25700 8838 25728 9386
rect 25688 8832 25740 8838
rect 25688 8774 25740 8780
rect 25700 7750 25728 8774
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25792 4078 25820 9574
rect 25964 9512 26016 9518
rect 25964 9454 26016 9460
rect 25976 8974 26004 9454
rect 25964 8968 26016 8974
rect 25964 8910 26016 8916
rect 26148 4752 26200 4758
rect 26148 4694 26200 4700
rect 25872 4480 25924 4486
rect 25872 4422 25924 4428
rect 25884 4214 25912 4422
rect 25872 4208 25924 4214
rect 25872 4150 25924 4156
rect 24860 4072 24912 4078
rect 24858 4040 24860 4049
rect 25780 4072 25832 4078
rect 24912 4040 24914 4049
rect 25780 4014 25832 4020
rect 24858 3975 24914 3984
rect 24952 3664 25004 3670
rect 24952 3606 25004 3612
rect 24032 3528 24084 3534
rect 24032 3470 24084 3476
rect 23940 3460 23992 3466
rect 23940 3402 23992 3408
rect 24044 3126 24072 3470
rect 24964 3126 24992 3606
rect 25792 3505 25820 4014
rect 25964 3732 26016 3738
rect 25964 3674 26016 3680
rect 25778 3496 25834 3505
rect 25778 3431 25834 3440
rect 24032 3120 24084 3126
rect 24032 3062 24084 3068
rect 24952 3120 25004 3126
rect 24952 3062 25004 3068
rect 23296 2848 23348 2854
rect 23296 2790 23348 2796
rect 22480 2746 22876 2774
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 22480 2582 22508 2746
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 24044 2650 24072 3062
rect 25976 2990 26004 3674
rect 26160 3058 26188 4694
rect 27080 4554 27108 11698
rect 27172 11218 27200 12242
rect 27264 11694 27292 14878
rect 27448 14550 27476 15830
rect 27436 14544 27488 14550
rect 27436 14486 27488 14492
rect 27344 14408 27396 14414
rect 27344 14350 27396 14356
rect 27356 13870 27384 14350
rect 27540 14006 27568 17002
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27632 14074 27660 16730
rect 27724 15502 27752 17031
rect 27802 16824 27858 16833
rect 27802 16759 27858 16768
rect 27816 16726 27844 16759
rect 27804 16720 27856 16726
rect 27804 16662 27856 16668
rect 27986 16688 28042 16697
rect 28276 16658 28304 17167
rect 27986 16623 27988 16632
rect 28040 16623 28042 16632
rect 28264 16652 28316 16658
rect 27988 16594 28040 16600
rect 28264 16594 28316 16600
rect 28368 16590 28396 19343
rect 28448 19314 28500 19320
rect 28460 18834 28488 19314
rect 28552 19242 28580 20046
rect 28644 19718 28672 20266
rect 28632 19712 28684 19718
rect 28632 19654 28684 19660
rect 28736 19514 28764 20742
rect 28908 20460 28960 20466
rect 28908 20402 28960 20408
rect 28920 19718 28948 20402
rect 29000 19916 29052 19922
rect 29000 19858 29052 19864
rect 28908 19712 28960 19718
rect 28814 19680 28870 19689
rect 28908 19654 28960 19660
rect 28814 19615 28870 19624
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 28632 19304 28684 19310
rect 28632 19246 28684 19252
rect 28540 19236 28592 19242
rect 28540 19178 28592 19184
rect 28448 18828 28500 18834
rect 28448 18770 28500 18776
rect 28552 18154 28580 19178
rect 28644 18630 28672 19246
rect 28722 18728 28778 18737
rect 28722 18663 28778 18672
rect 28632 18624 28684 18630
rect 28632 18566 28684 18572
rect 28540 18148 28592 18154
rect 28540 18090 28592 18096
rect 28446 18048 28502 18057
rect 28446 17983 28502 17992
rect 28460 17202 28488 17983
rect 28644 17728 28672 18566
rect 28736 18193 28764 18663
rect 28722 18184 28778 18193
rect 28722 18119 28778 18128
rect 28552 17700 28672 17728
rect 28448 17196 28500 17202
rect 28448 17138 28500 17144
rect 28552 16810 28580 17700
rect 28632 17604 28684 17610
rect 28632 17546 28684 17552
rect 28460 16782 28580 16810
rect 28644 16794 28672 17546
rect 28632 16788 28684 16794
rect 27804 16584 27856 16590
rect 27804 16526 27856 16532
rect 28356 16584 28408 16590
rect 28356 16526 28408 16532
rect 27816 16182 27844 16526
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 28368 16250 28396 16526
rect 28356 16244 28408 16250
rect 28356 16186 28408 16192
rect 27804 16176 27856 16182
rect 27804 16118 27856 16124
rect 27712 15496 27764 15502
rect 27712 15438 27764 15444
rect 27816 15026 27844 16118
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 27896 15088 27948 15094
rect 27896 15030 27948 15036
rect 27804 15020 27856 15026
rect 27804 14962 27856 14968
rect 27712 14884 27764 14890
rect 27712 14826 27764 14832
rect 27724 14278 27752 14826
rect 27908 14482 27936 15030
rect 27896 14476 27948 14482
rect 27816 14436 27896 14464
rect 27712 14272 27764 14278
rect 27712 14214 27764 14220
rect 27620 14068 27672 14074
rect 27620 14010 27672 14016
rect 27528 14000 27580 14006
rect 27528 13942 27580 13948
rect 27344 13864 27396 13870
rect 27344 13806 27396 13812
rect 27356 12306 27384 13806
rect 27436 13524 27488 13530
rect 27436 13466 27488 13472
rect 27448 12918 27476 13466
rect 27436 12912 27488 12918
rect 27436 12854 27488 12860
rect 27344 12300 27396 12306
rect 27344 12242 27396 12248
rect 27448 12170 27476 12854
rect 27632 12238 27660 14010
rect 27816 13530 27844 14436
rect 27896 14418 27948 14424
rect 28460 14278 28488 16782
rect 28632 16730 28684 16736
rect 28632 16516 28684 16522
rect 28632 16458 28684 16464
rect 28644 16046 28672 16458
rect 28632 16040 28684 16046
rect 28552 16000 28632 16028
rect 28552 15094 28580 16000
rect 28632 15982 28684 15988
rect 28736 15570 28764 18119
rect 28828 17270 28856 19615
rect 28920 19174 28948 19654
rect 28908 19168 28960 19174
rect 28908 19110 28960 19116
rect 29012 18986 29040 19858
rect 28920 18958 29040 18986
rect 28920 18902 28948 18958
rect 28908 18896 28960 18902
rect 29000 18896 29052 18902
rect 28908 18838 28960 18844
rect 28998 18864 29000 18873
rect 29052 18864 29054 18873
rect 28920 18748 28948 18838
rect 28998 18799 29054 18808
rect 28920 18720 29040 18748
rect 28908 17672 28960 17678
rect 28908 17614 28960 17620
rect 28816 17264 28868 17270
rect 28816 17206 28868 17212
rect 28828 16794 28856 17206
rect 28816 16788 28868 16794
rect 28816 16730 28868 16736
rect 28920 16182 28948 17614
rect 29012 17542 29040 18720
rect 29104 18290 29132 23462
rect 29184 22568 29236 22574
rect 29184 22510 29236 22516
rect 29196 22094 29224 22510
rect 29196 22066 29316 22094
rect 29288 20398 29316 22066
rect 29380 21622 29408 23598
rect 29644 23588 29696 23594
rect 30194 23559 30250 23568
rect 29644 23530 29696 23536
rect 29656 23186 29684 23530
rect 30208 23186 30236 23559
rect 30288 23520 30340 23526
rect 30288 23462 30340 23468
rect 30300 23186 30328 23462
rect 30392 23322 30420 23666
rect 30380 23316 30432 23322
rect 30380 23258 30432 23264
rect 29644 23180 29696 23186
rect 29644 23122 29696 23128
rect 30196 23180 30248 23186
rect 30196 23122 30248 23128
rect 30288 23180 30340 23186
rect 30288 23122 30340 23128
rect 30104 23112 30156 23118
rect 30156 23060 30328 23066
rect 30104 23054 30328 23060
rect 29920 23044 29972 23050
rect 30116 23038 30328 23054
rect 29920 22986 29972 22992
rect 29642 22672 29698 22681
rect 29642 22607 29698 22616
rect 29552 22092 29604 22098
rect 29552 22034 29604 22040
rect 29564 21894 29592 22034
rect 29552 21888 29604 21894
rect 29552 21830 29604 21836
rect 29368 21616 29420 21622
rect 29368 21558 29420 21564
rect 29276 20392 29328 20398
rect 29276 20334 29328 20340
rect 29276 19304 29328 19310
rect 29276 19246 29328 19252
rect 29184 18896 29236 18902
rect 29184 18838 29236 18844
rect 29196 18630 29224 18838
rect 29288 18834 29316 19246
rect 29276 18828 29328 18834
rect 29276 18770 29328 18776
rect 29380 18698 29408 21558
rect 29656 21350 29684 22607
rect 29932 22574 29960 22986
rect 30104 22976 30156 22982
rect 30104 22918 30156 22924
rect 29920 22568 29972 22574
rect 29920 22510 29972 22516
rect 29734 22400 29790 22409
rect 29734 22335 29790 22344
rect 29748 21894 29776 22335
rect 29828 22024 29880 22030
rect 29828 21966 29880 21972
rect 29736 21888 29788 21894
rect 29736 21830 29788 21836
rect 29736 21480 29788 21486
rect 29736 21422 29788 21428
rect 29552 21344 29604 21350
rect 29552 21286 29604 21292
rect 29644 21344 29696 21350
rect 29644 21286 29696 21292
rect 29460 21140 29512 21146
rect 29460 21082 29512 21088
rect 29472 20398 29500 21082
rect 29564 21078 29592 21286
rect 29552 21072 29604 21078
rect 29552 21014 29604 21020
rect 29642 21040 29698 21049
rect 29642 20975 29698 20984
rect 29460 20392 29512 20398
rect 29460 20334 29512 20340
rect 29368 18692 29420 18698
rect 29368 18634 29420 18640
rect 29184 18624 29236 18630
rect 29184 18566 29236 18572
rect 29092 18284 29144 18290
rect 29092 18226 29144 18232
rect 29368 18284 29420 18290
rect 29368 18226 29420 18232
rect 29000 17536 29052 17542
rect 29000 17478 29052 17484
rect 29000 17128 29052 17134
rect 29000 17070 29052 17076
rect 29012 16522 29040 17070
rect 29104 16522 29132 18226
rect 29380 18086 29408 18226
rect 29368 18080 29420 18086
rect 29368 18022 29420 18028
rect 29184 17536 29236 17542
rect 29184 17478 29236 17484
rect 29000 16516 29052 16522
rect 29000 16458 29052 16464
rect 29092 16516 29144 16522
rect 29092 16458 29144 16464
rect 29196 16182 29224 17478
rect 29276 17196 29328 17202
rect 29276 17138 29328 17144
rect 29288 16658 29316 17138
rect 29276 16652 29328 16658
rect 29276 16594 29328 16600
rect 28908 16176 28960 16182
rect 28908 16118 28960 16124
rect 29184 16176 29236 16182
rect 29184 16118 29236 16124
rect 29196 15638 29224 16118
rect 29184 15632 29236 15638
rect 29184 15574 29236 15580
rect 28724 15564 28776 15570
rect 28724 15506 28776 15512
rect 29000 15360 29052 15366
rect 29196 15337 29224 15574
rect 29000 15302 29052 15308
rect 29182 15328 29238 15337
rect 29012 15201 29040 15302
rect 29182 15263 29238 15272
rect 28998 15192 29054 15201
rect 28998 15127 29054 15136
rect 28540 15088 28592 15094
rect 29196 15076 29224 15263
rect 29276 15088 29328 15094
rect 29196 15048 29276 15076
rect 28540 15030 28592 15036
rect 29276 15030 29328 15036
rect 28632 14408 28684 14414
rect 28632 14350 28684 14356
rect 28448 14272 28500 14278
rect 28448 14214 28500 14220
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 27804 13524 27856 13530
rect 27804 13466 27856 13472
rect 28356 13524 28408 13530
rect 28356 13466 28408 13472
rect 27816 12646 27844 13466
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 27896 12980 27948 12986
rect 27896 12922 27948 12928
rect 27804 12640 27856 12646
rect 27804 12582 27856 12588
rect 27908 12442 27936 12922
rect 27896 12436 27948 12442
rect 27896 12378 27948 12384
rect 27528 12232 27580 12238
rect 27528 12174 27580 12180
rect 27620 12232 27672 12238
rect 27620 12174 27672 12180
rect 27436 12164 27488 12170
rect 27436 12106 27488 12112
rect 27344 12096 27396 12102
rect 27344 12038 27396 12044
rect 27356 11898 27384 12038
rect 27344 11892 27396 11898
rect 27344 11834 27396 11840
rect 27436 11892 27488 11898
rect 27436 11834 27488 11840
rect 27448 11778 27476 11834
rect 27356 11762 27476 11778
rect 27344 11756 27476 11762
rect 27396 11750 27476 11756
rect 27344 11698 27396 11704
rect 27252 11688 27304 11694
rect 27252 11630 27304 11636
rect 27344 11620 27396 11626
rect 27344 11562 27396 11568
rect 27160 11212 27212 11218
rect 27160 11154 27212 11160
rect 27172 9450 27200 11154
rect 27252 10668 27304 10674
rect 27252 10610 27304 10616
rect 27264 10169 27292 10610
rect 27250 10160 27306 10169
rect 27250 10095 27306 10104
rect 27160 9444 27212 9450
rect 27160 9386 27212 9392
rect 27264 4690 27292 10095
rect 27356 9994 27384 11562
rect 27344 9988 27396 9994
rect 27344 9930 27396 9936
rect 27356 9654 27384 9930
rect 27344 9648 27396 9654
rect 27344 9590 27396 9596
rect 27540 7750 27568 12174
rect 27620 12096 27672 12102
rect 27620 12038 27672 12044
rect 27632 11830 27660 12038
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 27620 11824 27672 11830
rect 27620 11766 27672 11772
rect 27632 11082 27660 11766
rect 27712 11688 27764 11694
rect 27712 11630 27764 11636
rect 27620 11076 27672 11082
rect 27620 11018 27672 11024
rect 27724 10810 27752 11630
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27712 10804 27764 10810
rect 27712 10746 27764 10752
rect 27620 10736 27672 10742
rect 27620 10678 27672 10684
rect 27632 10266 27660 10678
rect 27620 10260 27672 10266
rect 27620 10202 27672 10208
rect 27712 9988 27764 9994
rect 27712 9930 27764 9936
rect 27724 9654 27752 9930
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 27712 9648 27764 9654
rect 27712 9590 27764 9596
rect 27804 8832 27856 8838
rect 27804 8774 27856 8780
rect 27528 7744 27580 7750
rect 27528 7686 27580 7692
rect 27816 6390 27844 8774
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 27804 6384 27856 6390
rect 27804 6326 27856 6332
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 27252 4684 27304 4690
rect 27252 4626 27304 4632
rect 27068 4548 27120 4554
rect 27068 4490 27120 4496
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 27620 4140 27672 4146
rect 27620 4082 27672 4088
rect 27528 3936 27580 3942
rect 27528 3878 27580 3884
rect 26332 3664 26384 3670
rect 26332 3606 26384 3612
rect 26148 3052 26200 3058
rect 26148 2994 26200 3000
rect 25964 2984 26016 2990
rect 25964 2926 26016 2932
rect 26344 2650 26372 3606
rect 27540 2922 27568 3878
rect 27528 2916 27580 2922
rect 27528 2858 27580 2864
rect 27160 2848 27212 2854
rect 27160 2790 27212 2796
rect 24032 2644 24084 2650
rect 24032 2586 24084 2592
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 22468 2576 22520 2582
rect 22468 2518 22520 2524
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 24400 2508 24452 2514
rect 24400 2450 24452 2456
rect 26516 2508 26568 2514
rect 26516 2450 26568 2456
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 21456 2372 21508 2378
rect 21456 2314 21508 2320
rect 22296 800 22324 2450
rect 24412 800 24440 2450
rect 26528 800 26556 2450
rect 27172 2446 27200 2790
rect 27632 2650 27660 4082
rect 28368 3534 28396 13466
rect 28460 12889 28488 14214
rect 28644 13258 28672 14350
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 28908 13932 28960 13938
rect 28908 13874 28960 13880
rect 28920 13530 28948 13874
rect 28908 13524 28960 13530
rect 28908 13466 28960 13472
rect 29012 13326 29040 14214
rect 29288 13938 29316 15030
rect 29380 14482 29408 18022
rect 29472 17134 29500 20334
rect 29552 18828 29604 18834
rect 29552 18770 29604 18776
rect 29460 17128 29512 17134
rect 29460 17070 29512 17076
rect 29460 16992 29512 16998
rect 29460 16934 29512 16940
rect 29368 14476 29420 14482
rect 29368 14418 29420 14424
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 29000 13320 29052 13326
rect 29000 13262 29052 13268
rect 28632 13252 28684 13258
rect 28632 13194 28684 13200
rect 28446 12880 28502 12889
rect 28446 12815 28502 12824
rect 28644 11121 28672 13194
rect 28724 13184 28776 13190
rect 28724 13126 28776 13132
rect 28736 11898 28764 13126
rect 28908 12776 28960 12782
rect 28908 12718 28960 12724
rect 28816 12232 28868 12238
rect 28816 12174 28868 12180
rect 28724 11892 28776 11898
rect 28724 11834 28776 11840
rect 28828 11354 28856 12174
rect 28816 11348 28868 11354
rect 28816 11290 28868 11296
rect 28630 11112 28686 11121
rect 28630 11047 28686 11056
rect 28448 9036 28500 9042
rect 28448 8978 28500 8984
rect 28460 8838 28488 8978
rect 28448 8832 28500 8838
rect 28448 8774 28500 8780
rect 28644 7274 28672 11047
rect 28828 10742 28856 11290
rect 28920 11286 28948 12718
rect 28908 11280 28960 11286
rect 28908 11222 28960 11228
rect 29380 11014 29408 14418
rect 29472 12374 29500 16934
rect 29564 15094 29592 18770
rect 29656 18630 29684 20975
rect 29748 20942 29776 21422
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 29840 20534 29868 21966
rect 29920 21344 29972 21350
rect 29920 21286 29972 21292
rect 29932 21146 29960 21286
rect 30010 21176 30066 21185
rect 29920 21140 29972 21146
rect 30010 21111 30012 21120
rect 29920 21082 29972 21088
rect 30064 21111 30066 21120
rect 30012 21082 30064 21088
rect 29920 20936 29972 20942
rect 29920 20878 29972 20884
rect 29828 20528 29880 20534
rect 29828 20470 29880 20476
rect 29828 19984 29880 19990
rect 29828 19926 29880 19932
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29644 18624 29696 18630
rect 29644 18566 29696 18572
rect 29642 18456 29698 18465
rect 29748 18426 29776 19654
rect 29840 19417 29868 19926
rect 29826 19408 29882 19417
rect 29826 19343 29882 19352
rect 29642 18391 29698 18400
rect 29736 18420 29788 18426
rect 29656 15162 29684 18391
rect 29736 18362 29788 18368
rect 29840 17814 29868 19343
rect 29932 19242 29960 20878
rect 30116 20806 30144 22918
rect 30196 22228 30248 22234
rect 30196 22170 30248 22176
rect 30208 22001 30236 22170
rect 30194 21992 30250 22001
rect 30194 21927 30250 21936
rect 30104 20800 30156 20806
rect 30104 20742 30156 20748
rect 30208 20466 30236 21927
rect 30300 20466 30328 23038
rect 30380 22976 30432 22982
rect 30380 22918 30432 22924
rect 30392 22438 30420 22918
rect 30472 22636 30524 22642
rect 30472 22578 30524 22584
rect 30380 22432 30432 22438
rect 30380 22374 30432 22380
rect 30484 21962 30512 22578
rect 30576 22098 30604 24006
rect 30746 22808 30802 22817
rect 30746 22743 30802 22752
rect 30760 22710 30788 22743
rect 30656 22704 30708 22710
rect 30654 22672 30656 22681
rect 30748 22704 30800 22710
rect 30708 22672 30710 22681
rect 30748 22646 30800 22652
rect 30654 22607 30710 22616
rect 30564 22092 30616 22098
rect 30564 22034 30616 22040
rect 30472 21956 30524 21962
rect 30472 21898 30524 21904
rect 30380 21888 30432 21894
rect 30380 21830 30432 21836
rect 30392 21457 30420 21830
rect 30378 21448 30434 21457
rect 30576 21418 30604 22034
rect 30656 22024 30708 22030
rect 30656 21966 30708 21972
rect 30840 22024 30892 22030
rect 30840 21966 30892 21972
rect 30378 21383 30434 21392
rect 30472 21412 30524 21418
rect 30392 20641 30420 21383
rect 30472 21354 30524 21360
rect 30564 21412 30616 21418
rect 30564 21354 30616 21360
rect 30378 20632 30434 20641
rect 30378 20567 30434 20576
rect 30196 20460 30248 20466
rect 30196 20402 30248 20408
rect 30288 20460 30340 20466
rect 30288 20402 30340 20408
rect 30102 20360 30158 20369
rect 30102 20295 30158 20304
rect 30116 19786 30144 20295
rect 30288 20256 30340 20262
rect 30288 20198 30340 20204
rect 30196 19848 30248 19854
rect 30196 19790 30248 19796
rect 30012 19780 30064 19786
rect 30012 19722 30064 19728
rect 30104 19780 30156 19786
rect 30104 19722 30156 19728
rect 29920 19236 29972 19242
rect 29920 19178 29972 19184
rect 30024 19174 30052 19722
rect 30208 19514 30236 19790
rect 30196 19508 30248 19514
rect 30196 19450 30248 19456
rect 30012 19168 30064 19174
rect 30012 19110 30064 19116
rect 29828 17808 29880 17814
rect 29828 17750 29880 17756
rect 29840 17270 29868 17750
rect 29920 17604 29972 17610
rect 29920 17546 29972 17552
rect 29932 17513 29960 17546
rect 30024 17542 30052 19110
rect 30196 18964 30248 18970
rect 30196 18906 30248 18912
rect 30208 18601 30236 18906
rect 30194 18592 30250 18601
rect 30194 18527 30250 18536
rect 30104 18216 30156 18222
rect 30104 18158 30156 18164
rect 30116 18086 30144 18158
rect 30104 18080 30156 18086
rect 30104 18022 30156 18028
rect 30012 17536 30064 17542
rect 29918 17504 29974 17513
rect 30012 17478 30064 17484
rect 29918 17439 29974 17448
rect 29828 17264 29880 17270
rect 29828 17206 29880 17212
rect 30208 16658 30236 18527
rect 30300 17270 30328 20198
rect 30380 19372 30432 19378
rect 30380 19314 30432 19320
rect 30392 19174 30420 19314
rect 30380 19168 30432 19174
rect 30380 19110 30432 19116
rect 30392 17513 30420 19110
rect 30484 18970 30512 21354
rect 30668 20777 30696 21966
rect 30748 21548 30800 21554
rect 30748 21490 30800 21496
rect 30760 21457 30788 21490
rect 30746 21448 30802 21457
rect 30746 21383 30802 21392
rect 30748 21344 30800 21350
rect 30748 21286 30800 21292
rect 30654 20768 30710 20777
rect 30654 20703 30710 20712
rect 30564 19848 30616 19854
rect 30564 19790 30616 19796
rect 30472 18964 30524 18970
rect 30472 18906 30524 18912
rect 30472 18624 30524 18630
rect 30472 18566 30524 18572
rect 30378 17504 30434 17513
rect 30378 17439 30434 17448
rect 30288 17264 30340 17270
rect 30288 17206 30340 17212
rect 30288 17128 30340 17134
rect 30288 17070 30340 17076
rect 30104 16652 30156 16658
rect 30104 16594 30156 16600
rect 30196 16652 30248 16658
rect 30196 16594 30248 16600
rect 29736 16448 29788 16454
rect 29736 16390 29788 16396
rect 29644 15156 29696 15162
rect 29644 15098 29696 15104
rect 29552 15088 29604 15094
rect 29552 15030 29604 15036
rect 29460 12368 29512 12374
rect 29460 12310 29512 12316
rect 29564 11694 29592 15030
rect 29748 14482 29776 16390
rect 29920 16176 29972 16182
rect 29920 16118 29972 16124
rect 29828 16040 29880 16046
rect 29828 15982 29880 15988
rect 29840 14958 29868 15982
rect 29932 15745 29960 16118
rect 29918 15736 29974 15745
rect 29918 15671 29974 15680
rect 29828 14952 29880 14958
rect 29828 14894 29880 14900
rect 29736 14476 29788 14482
rect 29736 14418 29788 14424
rect 29644 14272 29696 14278
rect 29644 14214 29696 14220
rect 29840 14226 29868 14894
rect 29932 14464 29960 15671
rect 30012 14952 30064 14958
rect 30012 14894 30064 14900
rect 30024 14618 30052 14894
rect 30012 14612 30064 14618
rect 30012 14554 30064 14560
rect 30012 14476 30064 14482
rect 29932 14436 30012 14464
rect 30012 14418 30064 14424
rect 30024 14278 30052 14418
rect 30012 14272 30064 14278
rect 29656 12918 29684 14214
rect 29840 14198 29960 14226
rect 30012 14214 30064 14220
rect 29736 13796 29788 13802
rect 29736 13738 29788 13744
rect 29644 12912 29696 12918
rect 29644 12854 29696 12860
rect 29656 12209 29684 12854
rect 29748 12345 29776 13738
rect 29932 13462 29960 14198
rect 30012 14068 30064 14074
rect 30012 14010 30064 14016
rect 29920 13456 29972 13462
rect 29920 13398 29972 13404
rect 29828 13388 29880 13394
rect 29828 13330 29880 13336
rect 29734 12336 29790 12345
rect 29734 12271 29790 12280
rect 29642 12200 29698 12209
rect 29642 12135 29698 12144
rect 29552 11688 29604 11694
rect 29552 11630 29604 11636
rect 29644 11688 29696 11694
rect 29644 11630 29696 11636
rect 29656 11150 29684 11630
rect 29644 11144 29696 11150
rect 29644 11086 29696 11092
rect 29184 11008 29236 11014
rect 29184 10950 29236 10956
rect 29368 11008 29420 11014
rect 29368 10950 29420 10956
rect 28816 10736 28868 10742
rect 28816 10678 28868 10684
rect 29092 10260 29144 10266
rect 29092 10202 29144 10208
rect 29104 8566 29132 10202
rect 29196 9994 29224 10950
rect 29276 10600 29328 10606
rect 29276 10542 29328 10548
rect 29288 10130 29316 10542
rect 29380 10130 29408 10950
rect 29656 10606 29684 11086
rect 29644 10600 29696 10606
rect 29644 10542 29696 10548
rect 29276 10124 29328 10130
rect 29276 10066 29328 10072
rect 29368 10124 29420 10130
rect 29368 10066 29420 10072
rect 29184 9988 29236 9994
rect 29184 9930 29236 9936
rect 29288 9518 29316 10066
rect 29748 9926 29776 12271
rect 29840 10606 29868 13330
rect 29932 12170 29960 13398
rect 30024 12850 30052 14010
rect 30012 12844 30064 12850
rect 30012 12786 30064 12792
rect 30024 12306 30052 12786
rect 30012 12300 30064 12306
rect 30012 12242 30064 12248
rect 29920 12164 29972 12170
rect 29920 12106 29972 12112
rect 30010 11112 30066 11121
rect 30010 11047 30066 11056
rect 30024 11014 30052 11047
rect 30012 11008 30064 11014
rect 30012 10950 30064 10956
rect 29920 10668 29972 10674
rect 29920 10610 29972 10616
rect 29828 10600 29880 10606
rect 29828 10542 29880 10548
rect 29840 10266 29868 10542
rect 29828 10260 29880 10266
rect 29828 10202 29880 10208
rect 29736 9920 29788 9926
rect 29736 9862 29788 9868
rect 29276 9512 29328 9518
rect 29196 9472 29276 9500
rect 29092 8560 29144 8566
rect 29092 8502 29144 8508
rect 29196 8430 29224 9472
rect 29276 9454 29328 9460
rect 28816 8424 28868 8430
rect 28816 8366 28868 8372
rect 29184 8424 29236 8430
rect 29184 8366 29236 8372
rect 28632 7268 28684 7274
rect 28632 7210 28684 7216
rect 28356 3528 28408 3534
rect 28356 3470 28408 3476
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 28828 3058 28856 8366
rect 29932 7954 29960 10610
rect 30116 9976 30144 16594
rect 30300 15552 30328 17070
rect 30208 15524 30420 15552
rect 30208 15026 30236 15524
rect 30288 15428 30340 15434
rect 30288 15370 30340 15376
rect 30196 15020 30248 15026
rect 30196 14962 30248 14968
rect 30196 14816 30248 14822
rect 30196 14758 30248 14764
rect 30208 13326 30236 14758
rect 30300 14278 30328 15370
rect 30288 14272 30340 14278
rect 30288 14214 30340 14220
rect 30300 13870 30328 14214
rect 30288 13864 30340 13870
rect 30288 13806 30340 13812
rect 30392 13462 30420 15524
rect 30380 13456 30432 13462
rect 30380 13398 30432 13404
rect 30484 13394 30512 18566
rect 30576 17202 30604 19790
rect 30760 18902 30788 21286
rect 30852 20602 30880 21966
rect 30840 20596 30892 20602
rect 30840 20538 30892 20544
rect 30944 20330 30972 24006
rect 31024 22500 31076 22506
rect 31024 22442 31076 22448
rect 31036 21962 31064 22442
rect 31128 22438 31156 24210
rect 31220 22982 31248 26200
rect 31864 24614 31892 26200
rect 31942 24712 31998 24721
rect 31942 24647 31998 24656
rect 31576 24608 31628 24614
rect 31576 24550 31628 24556
rect 31852 24608 31904 24614
rect 31852 24550 31904 24556
rect 31588 24206 31616 24550
rect 31576 24200 31628 24206
rect 31576 24142 31628 24148
rect 31484 23316 31536 23322
rect 31588 23304 31616 24142
rect 31760 23656 31812 23662
rect 31760 23598 31812 23604
rect 31536 23276 31616 23304
rect 31484 23258 31536 23264
rect 31772 23186 31800 23598
rect 31760 23180 31812 23186
rect 31760 23122 31812 23128
rect 31392 23112 31444 23118
rect 31392 23054 31444 23060
rect 31208 22976 31260 22982
rect 31208 22918 31260 22924
rect 31404 22778 31432 23054
rect 31392 22772 31444 22778
rect 31392 22714 31444 22720
rect 31116 22432 31168 22438
rect 31116 22374 31168 22380
rect 31024 21956 31076 21962
rect 31024 21898 31076 21904
rect 31036 20398 31064 21898
rect 31128 20534 31156 22374
rect 31404 22094 31432 22714
rect 31482 22536 31538 22545
rect 31482 22471 31538 22480
rect 31496 22438 31524 22471
rect 31484 22432 31536 22438
rect 31484 22374 31536 22380
rect 31852 22228 31904 22234
rect 31852 22170 31904 22176
rect 31484 22094 31536 22098
rect 31404 22092 31536 22094
rect 31404 22066 31484 22092
rect 31484 22034 31536 22040
rect 31864 22094 31892 22170
rect 31956 22094 31984 24647
rect 32128 24064 32180 24070
rect 32128 24006 32180 24012
rect 32312 24064 32364 24070
rect 32312 24006 32364 24012
rect 32140 23905 32168 24006
rect 32126 23896 32182 23905
rect 32126 23831 32182 23840
rect 32140 23050 32168 23831
rect 32324 23594 32352 24006
rect 32404 23792 32456 23798
rect 32404 23734 32456 23740
rect 32312 23588 32364 23594
rect 32312 23530 32364 23536
rect 32128 23044 32180 23050
rect 32128 22986 32180 22992
rect 31864 22066 31984 22094
rect 31496 22003 31524 22034
rect 31392 21956 31444 21962
rect 31392 21898 31444 21904
rect 31206 21584 31262 21593
rect 31206 21519 31208 21528
rect 31260 21519 31262 21528
rect 31208 21490 31260 21496
rect 31404 21185 31432 21898
rect 31760 21684 31812 21690
rect 31760 21626 31812 21632
rect 31576 21480 31628 21486
rect 31576 21422 31628 21428
rect 31484 21412 31536 21418
rect 31484 21354 31536 21360
rect 31390 21176 31446 21185
rect 31390 21111 31446 21120
rect 31496 20806 31524 21354
rect 31208 20800 31260 20806
rect 31208 20742 31260 20748
rect 31484 20800 31536 20806
rect 31484 20742 31536 20748
rect 31116 20528 31168 20534
rect 31116 20470 31168 20476
rect 31024 20392 31076 20398
rect 31024 20334 31076 20340
rect 30932 20324 30984 20330
rect 30932 20266 30984 20272
rect 30840 20256 30892 20262
rect 30840 20198 30892 20204
rect 31116 20256 31168 20262
rect 31116 20198 31168 20204
rect 30748 18896 30800 18902
rect 30748 18838 30800 18844
rect 30656 18624 30708 18630
rect 30656 18566 30708 18572
rect 30564 17196 30616 17202
rect 30564 17138 30616 17144
rect 30564 16992 30616 16998
rect 30564 16934 30616 16940
rect 30576 16250 30604 16934
rect 30564 16244 30616 16250
rect 30564 16186 30616 16192
rect 30668 16182 30696 18566
rect 30748 17128 30800 17134
rect 30748 17070 30800 17076
rect 30656 16176 30708 16182
rect 30656 16118 30708 16124
rect 30760 15910 30788 17070
rect 30852 16182 30880 20198
rect 31128 19825 31156 20198
rect 31114 19816 31170 19825
rect 31114 19751 31170 19760
rect 31128 19718 31156 19751
rect 30932 19712 30984 19718
rect 30932 19654 30984 19660
rect 31116 19712 31168 19718
rect 31116 19654 31168 19660
rect 30944 18902 30972 19654
rect 30932 18896 30984 18902
rect 30932 18838 30984 18844
rect 30944 18737 30972 18838
rect 31024 18760 31076 18766
rect 30930 18728 30986 18737
rect 31024 18702 31076 18708
rect 31116 18760 31168 18766
rect 31116 18702 31168 18708
rect 30930 18663 30986 18672
rect 31036 18154 31064 18702
rect 31024 18148 31076 18154
rect 31024 18090 31076 18096
rect 30932 17876 30984 17882
rect 30932 17818 30984 17824
rect 30840 16176 30892 16182
rect 30840 16118 30892 16124
rect 30748 15904 30800 15910
rect 30748 15846 30800 15852
rect 30760 15434 30788 15846
rect 30748 15428 30800 15434
rect 30748 15370 30800 15376
rect 30562 15192 30618 15201
rect 30562 15127 30618 15136
rect 30576 15026 30604 15127
rect 30564 15020 30616 15026
rect 30564 14962 30616 14968
rect 30576 13841 30604 14962
rect 30656 14952 30708 14958
rect 30654 14920 30656 14929
rect 30708 14920 30710 14929
rect 30654 14855 30710 14864
rect 30760 14482 30788 15370
rect 30944 15094 30972 17818
rect 31128 16794 31156 18702
rect 31220 18426 31248 20742
rect 31484 20596 31536 20602
rect 31484 20538 31536 20544
rect 31300 20392 31352 20398
rect 31300 20334 31352 20340
rect 31312 19854 31340 20334
rect 31392 20324 31444 20330
rect 31392 20266 31444 20272
rect 31300 19848 31352 19854
rect 31300 19790 31352 19796
rect 31298 18864 31354 18873
rect 31298 18799 31354 18808
rect 31312 18698 31340 18799
rect 31300 18692 31352 18698
rect 31300 18634 31352 18640
rect 31208 18420 31260 18426
rect 31208 18362 31260 18368
rect 31404 17882 31432 20266
rect 31496 19446 31524 20538
rect 31588 19802 31616 21422
rect 31772 21049 31800 21626
rect 31758 21040 31814 21049
rect 31758 20975 31814 20984
rect 31588 19774 31708 19802
rect 31576 19712 31628 19718
rect 31576 19654 31628 19660
rect 31484 19440 31536 19446
rect 31484 19382 31536 19388
rect 31588 18630 31616 19654
rect 31680 19310 31708 19774
rect 31772 19446 31800 20975
rect 31864 20534 31892 22066
rect 32140 22030 32168 22986
rect 32312 22092 32364 22098
rect 32232 22052 32312 22080
rect 32128 22024 32180 22030
rect 32128 21966 32180 21972
rect 32140 21894 32168 21966
rect 32128 21888 32180 21894
rect 32128 21830 32180 21836
rect 31944 21344 31996 21350
rect 31944 21286 31996 21292
rect 31956 21078 31984 21286
rect 31944 21072 31996 21078
rect 31944 21014 31996 21020
rect 31852 20528 31904 20534
rect 31852 20470 31904 20476
rect 31956 20466 31984 21014
rect 32140 20874 32168 21830
rect 32128 20868 32180 20874
rect 32128 20810 32180 20816
rect 32140 20534 32168 20810
rect 32128 20528 32180 20534
rect 32128 20470 32180 20476
rect 31944 20460 31996 20466
rect 31944 20402 31996 20408
rect 32232 19786 32260 22052
rect 32312 22034 32364 22040
rect 32416 21894 32444 23734
rect 32508 23225 32536 26200
rect 33152 24682 33180 26200
rect 33324 24880 33376 24886
rect 33324 24822 33376 24828
rect 33140 24676 33192 24682
rect 33140 24618 33192 24624
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 32862 24304 32918 24313
rect 32862 24239 32918 24248
rect 32680 23724 32732 23730
rect 32680 23666 32732 23672
rect 32494 23216 32550 23225
rect 32494 23151 32550 23160
rect 32692 21894 32720 23666
rect 32772 22636 32824 22642
rect 32772 22578 32824 22584
rect 32784 22234 32812 22578
rect 32772 22228 32824 22234
rect 32772 22170 32824 22176
rect 32404 21888 32456 21894
rect 32404 21830 32456 21836
rect 32680 21888 32732 21894
rect 32680 21830 32732 21836
rect 32312 21004 32364 21010
rect 32312 20946 32364 20952
rect 32324 20398 32352 20946
rect 32416 20942 32444 21830
rect 32876 21457 32904 24239
rect 33336 24206 33364 24822
rect 33508 24336 33560 24342
rect 33508 24278 33560 24284
rect 33324 24200 33376 24206
rect 33324 24142 33376 24148
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 33336 23322 33364 24142
rect 33324 23316 33376 23322
rect 33324 23258 33376 23264
rect 33520 23186 33548 24278
rect 33782 23896 33838 23905
rect 33782 23831 33838 23840
rect 33796 23798 33824 23831
rect 33784 23792 33836 23798
rect 33690 23760 33746 23769
rect 33784 23734 33836 23740
rect 33690 23695 33746 23704
rect 33598 23352 33654 23361
rect 33598 23287 33654 23296
rect 33508 23180 33560 23186
rect 33508 23122 33560 23128
rect 33416 23044 33468 23050
rect 33416 22986 33468 22992
rect 33428 22642 33456 22986
rect 33416 22636 33468 22642
rect 33416 22578 33468 22584
rect 33520 22574 33548 23122
rect 33612 22710 33640 23287
rect 33600 22704 33652 22710
rect 33600 22646 33652 22652
rect 33508 22568 33560 22574
rect 33508 22510 33560 22516
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 33520 22094 33548 22510
rect 33336 22066 33548 22094
rect 32862 21448 32918 21457
rect 32862 21383 32918 21392
rect 32404 20936 32456 20942
rect 32404 20878 32456 20884
rect 32496 20936 32548 20942
rect 32496 20878 32548 20884
rect 32508 20602 32536 20878
rect 32496 20596 32548 20602
rect 32496 20538 32548 20544
rect 32312 20392 32364 20398
rect 32312 20334 32364 20340
rect 32588 20392 32640 20398
rect 32588 20334 32640 20340
rect 32770 20360 32826 20369
rect 32220 19780 32272 19786
rect 32220 19722 32272 19728
rect 32128 19712 32180 19718
rect 32128 19654 32180 19660
rect 31852 19508 31904 19514
rect 31852 19450 31904 19456
rect 31760 19440 31812 19446
rect 31760 19382 31812 19388
rect 31668 19304 31720 19310
rect 31668 19246 31720 19252
rect 31668 18760 31720 18766
rect 31668 18702 31720 18708
rect 31576 18624 31628 18630
rect 31576 18566 31628 18572
rect 31392 17876 31444 17882
rect 31392 17818 31444 17824
rect 31392 17740 31444 17746
rect 31392 17682 31444 17688
rect 31484 17740 31536 17746
rect 31536 17700 31616 17728
rect 31484 17682 31536 17688
rect 31404 17377 31432 17682
rect 31484 17604 31536 17610
rect 31484 17546 31536 17552
rect 31390 17368 31446 17377
rect 31390 17303 31446 17312
rect 31496 17202 31524 17546
rect 31392 17196 31444 17202
rect 31392 17138 31444 17144
rect 31484 17196 31536 17202
rect 31484 17138 31536 17144
rect 31116 16788 31168 16794
rect 31116 16730 31168 16736
rect 31208 16448 31260 16454
rect 31208 16390 31260 16396
rect 31300 16448 31352 16454
rect 31300 16390 31352 16396
rect 31220 16046 31248 16390
rect 31208 16040 31260 16046
rect 31208 15982 31260 15988
rect 31208 15904 31260 15910
rect 31208 15846 31260 15852
rect 31116 15564 31168 15570
rect 31116 15506 31168 15512
rect 31024 15360 31076 15366
rect 31024 15302 31076 15308
rect 30932 15088 30984 15094
rect 30932 15030 30984 15036
rect 30748 14476 30800 14482
rect 30748 14418 30800 14424
rect 31036 14278 31064 15302
rect 31024 14272 31076 14278
rect 31024 14214 31076 14220
rect 31128 14074 31156 15506
rect 31220 15434 31248 15846
rect 31208 15428 31260 15434
rect 31208 15370 31260 15376
rect 31220 15337 31248 15370
rect 31206 15328 31262 15337
rect 31206 15263 31262 15272
rect 31116 14068 31168 14074
rect 31116 14010 31168 14016
rect 31128 13938 31156 14010
rect 31220 14006 31248 15263
rect 31312 15162 31340 16390
rect 31300 15156 31352 15162
rect 31300 15098 31352 15104
rect 31208 14000 31260 14006
rect 31208 13942 31260 13948
rect 31116 13932 31168 13938
rect 31116 13874 31168 13880
rect 30562 13832 30618 13841
rect 30562 13767 30618 13776
rect 30840 13728 30892 13734
rect 30840 13670 30892 13676
rect 30472 13388 30524 13394
rect 30472 13330 30524 13336
rect 30196 13320 30248 13326
rect 30196 13262 30248 13268
rect 30562 13288 30618 13297
rect 30562 13223 30618 13232
rect 30196 12912 30248 12918
rect 30196 12854 30248 12860
rect 30208 10470 30236 12854
rect 30472 11620 30524 11626
rect 30472 11562 30524 11568
rect 30484 11286 30512 11562
rect 30472 11280 30524 11286
rect 30472 11222 30524 11228
rect 30472 10600 30524 10606
rect 30472 10542 30524 10548
rect 30196 10464 30248 10470
rect 30196 10406 30248 10412
rect 30024 9948 30144 9976
rect 30380 9988 30432 9994
rect 30024 9518 30052 9948
rect 30380 9930 30432 9936
rect 30104 9648 30156 9654
rect 30104 9590 30156 9596
rect 30116 9518 30144 9590
rect 30012 9512 30064 9518
rect 30012 9454 30064 9460
rect 30104 9512 30156 9518
rect 30104 9454 30156 9460
rect 30024 9110 30052 9454
rect 30012 9104 30064 9110
rect 30012 9046 30064 9052
rect 30392 8838 30420 9930
rect 30484 9382 30512 10542
rect 30472 9376 30524 9382
rect 30472 9318 30524 9324
rect 30380 8832 30432 8838
rect 30380 8774 30432 8780
rect 30472 8560 30524 8566
rect 30472 8502 30524 8508
rect 29920 7948 29972 7954
rect 29920 7890 29972 7896
rect 30484 7818 30512 8502
rect 30576 8090 30604 13223
rect 30852 11694 30880 13670
rect 31220 13326 31248 13942
rect 31404 13394 31432 17138
rect 31484 15904 31536 15910
rect 31484 15846 31536 15852
rect 31392 13388 31444 13394
rect 31392 13330 31444 13336
rect 31208 13320 31260 13326
rect 31260 13280 31340 13308
rect 31208 13262 31260 13268
rect 31312 12918 31340 13280
rect 31300 12912 31352 12918
rect 31300 12854 31352 12860
rect 31312 12306 31340 12854
rect 31300 12300 31352 12306
rect 31300 12242 31352 12248
rect 31496 12238 31524 15846
rect 31588 14482 31616 17700
rect 31680 16454 31708 18702
rect 31668 16448 31720 16454
rect 31668 16390 31720 16396
rect 31668 16176 31720 16182
rect 31668 16118 31720 16124
rect 31680 14550 31708 16118
rect 31864 15638 31892 19450
rect 32140 18358 32168 19654
rect 32496 19508 32548 19514
rect 32496 19450 32548 19456
rect 32404 19304 32456 19310
rect 32404 19246 32456 19252
rect 32128 18352 32180 18358
rect 32128 18294 32180 18300
rect 31944 18216 31996 18222
rect 31944 18158 31996 18164
rect 31956 16658 31984 18158
rect 32128 17536 32180 17542
rect 32128 17478 32180 17484
rect 32312 17536 32364 17542
rect 32312 17478 32364 17484
rect 31944 16652 31996 16658
rect 31944 16594 31996 16600
rect 31944 16516 31996 16522
rect 31944 16458 31996 16464
rect 31852 15632 31904 15638
rect 31852 15574 31904 15580
rect 31760 15020 31812 15026
rect 31760 14962 31812 14968
rect 31668 14544 31720 14550
rect 31668 14486 31720 14492
rect 31576 14476 31628 14482
rect 31576 14418 31628 14424
rect 31484 12232 31536 12238
rect 31484 12174 31536 12180
rect 31392 12096 31444 12102
rect 31392 12038 31444 12044
rect 31404 11830 31432 12038
rect 31588 11914 31616 14418
rect 31668 13184 31720 13190
rect 31668 13126 31720 13132
rect 31496 11886 31616 11914
rect 31392 11824 31444 11830
rect 31392 11766 31444 11772
rect 31116 11756 31168 11762
rect 31116 11698 31168 11704
rect 30840 11688 30892 11694
rect 30840 11630 30892 11636
rect 30748 11008 30800 11014
rect 30748 10950 30800 10956
rect 30840 11008 30892 11014
rect 30840 10950 30892 10956
rect 30656 10600 30708 10606
rect 30656 10542 30708 10548
rect 30668 10130 30696 10542
rect 30656 10124 30708 10130
rect 30656 10066 30708 10072
rect 30656 9648 30708 9654
rect 30656 9590 30708 9596
rect 30668 9382 30696 9590
rect 30656 9376 30708 9382
rect 30656 9318 30708 9324
rect 30668 8838 30696 9318
rect 30656 8832 30708 8838
rect 30656 8774 30708 8780
rect 30668 8498 30696 8774
rect 30656 8492 30708 8498
rect 30656 8434 30708 8440
rect 30564 8084 30616 8090
rect 30564 8026 30616 8032
rect 30576 7886 30604 8026
rect 30564 7880 30616 7886
rect 30564 7822 30616 7828
rect 30472 7812 30524 7818
rect 30472 7754 30524 7760
rect 30484 7002 30512 7754
rect 30668 7750 30696 8434
rect 30656 7744 30708 7750
rect 30656 7686 30708 7692
rect 30472 6996 30524 7002
rect 30472 6938 30524 6944
rect 29644 3664 29696 3670
rect 29644 3606 29696 3612
rect 29000 3596 29052 3602
rect 29000 3538 29052 3544
rect 28816 3052 28868 3058
rect 28816 2994 28868 3000
rect 29012 2650 29040 3538
rect 29656 3126 29684 3606
rect 29644 3120 29696 3126
rect 29644 3062 29696 3068
rect 29656 2990 29684 3062
rect 30668 2990 30696 7686
rect 30760 6390 30788 10950
rect 30852 10470 30880 10950
rect 31128 10810 31156 11698
rect 31496 11200 31524 11886
rect 31576 11824 31628 11830
rect 31576 11766 31628 11772
rect 31404 11172 31524 11200
rect 31404 11082 31432 11172
rect 31392 11076 31444 11082
rect 31392 11018 31444 11024
rect 31484 11076 31536 11082
rect 31588 11064 31616 11766
rect 31536 11036 31616 11064
rect 31484 11018 31536 11024
rect 31116 10804 31168 10810
rect 31116 10746 31168 10752
rect 30840 10464 30892 10470
rect 30840 10406 30892 10412
rect 31404 10266 31432 11018
rect 31392 10260 31444 10266
rect 31392 10202 31444 10208
rect 31496 9500 31524 11018
rect 31680 9586 31708 13126
rect 31772 12434 31800 14962
rect 31852 14952 31904 14958
rect 31850 14920 31852 14929
rect 31904 14920 31906 14929
rect 31850 14855 31906 14864
rect 31852 14408 31904 14414
rect 31852 14350 31904 14356
rect 31864 12986 31892 14350
rect 31956 13938 31984 16458
rect 32036 16244 32088 16250
rect 32036 16186 32088 16192
rect 32048 15978 32076 16186
rect 32036 15972 32088 15978
rect 32036 15914 32088 15920
rect 31944 13932 31996 13938
rect 31944 13874 31996 13880
rect 31852 12980 31904 12986
rect 31852 12922 31904 12928
rect 32036 12436 32088 12442
rect 31772 12406 31892 12434
rect 31760 12300 31812 12306
rect 31760 12242 31812 12248
rect 31772 12102 31800 12242
rect 31760 12096 31812 12102
rect 31760 12038 31812 12044
rect 31772 11830 31800 12038
rect 31864 11898 31892 12406
rect 32140 12434 32168 17478
rect 32324 17338 32352 17478
rect 32312 17332 32364 17338
rect 32312 17274 32364 17280
rect 32220 17196 32272 17202
rect 32220 17138 32272 17144
rect 32232 16658 32260 17138
rect 32312 17060 32364 17066
rect 32312 17002 32364 17008
rect 32220 16652 32272 16658
rect 32220 16594 32272 16600
rect 32324 15366 32352 17002
rect 32416 16046 32444 19246
rect 32404 16040 32456 16046
rect 32404 15982 32456 15988
rect 32312 15360 32364 15366
rect 32312 15302 32364 15308
rect 32312 14952 32364 14958
rect 32312 14894 32364 14900
rect 32324 13870 32352 14894
rect 32416 14362 32444 15982
rect 32508 14550 32536 19450
rect 32600 18086 32628 20334
rect 32770 20295 32772 20304
rect 32824 20295 32826 20304
rect 32772 20266 32824 20272
rect 32876 19446 32904 21383
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 33140 21004 33192 21010
rect 33140 20946 33192 20952
rect 33152 20890 33180 20946
rect 32968 20862 33180 20890
rect 32968 20806 32996 20862
rect 32956 20800 33008 20806
rect 32956 20742 33008 20748
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 33336 20074 33364 22066
rect 33416 21888 33468 21894
rect 33416 21830 33468 21836
rect 33428 21690 33456 21830
rect 33416 21684 33468 21690
rect 33416 21626 33468 21632
rect 33704 21622 33732 23695
rect 33796 23254 33824 23734
rect 33784 23248 33836 23254
rect 33784 23190 33836 23196
rect 33784 22976 33836 22982
rect 33784 22918 33836 22924
rect 33692 21616 33744 21622
rect 33506 21584 33562 21593
rect 33692 21558 33744 21564
rect 33506 21519 33508 21528
rect 33560 21519 33562 21528
rect 33508 21490 33560 21496
rect 33416 21480 33468 21486
rect 33416 21422 33468 21428
rect 33428 21128 33456 21422
rect 33428 21100 33640 21128
rect 33508 21004 33560 21010
rect 33508 20946 33560 20952
rect 33336 20046 33456 20074
rect 33324 19984 33376 19990
rect 33324 19926 33376 19932
rect 32864 19440 32916 19446
rect 32864 19382 32916 19388
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 33336 18970 33364 19926
rect 33428 19718 33456 20046
rect 33416 19712 33468 19718
rect 33416 19654 33468 19660
rect 33324 18964 33376 18970
rect 33324 18906 33376 18912
rect 33048 18896 33100 18902
rect 33048 18838 33100 18844
rect 33060 18578 33088 18838
rect 32692 18550 33088 18578
rect 33416 18624 33468 18630
rect 33416 18566 33468 18572
rect 32692 18290 32720 18550
rect 32680 18284 32732 18290
rect 32680 18226 32732 18232
rect 32588 18080 32640 18086
rect 32588 18022 32640 18028
rect 32692 17542 32720 18226
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 32864 17808 32916 17814
rect 32864 17750 32916 17756
rect 32680 17536 32732 17542
rect 32876 17524 32904 17750
rect 32956 17740 33008 17746
rect 32956 17682 33008 17688
rect 32968 17626 32996 17682
rect 33428 17626 33456 18566
rect 33520 17746 33548 20946
rect 33612 18358 33640 21100
rect 33796 19854 33824 22918
rect 33980 22273 34008 26302
rect 34426 26200 34482 27000
rect 35070 26200 35126 27000
rect 35714 26200 35770 27000
rect 36358 26330 36414 27000
rect 36358 26302 36492 26330
rect 36358 26200 36414 26302
rect 34152 24132 34204 24138
rect 34152 24074 34204 24080
rect 34060 24064 34112 24070
rect 34060 24006 34112 24012
rect 34072 23497 34100 24006
rect 34058 23488 34114 23497
rect 34058 23423 34114 23432
rect 34060 22568 34112 22574
rect 34060 22510 34112 22516
rect 33966 22264 34022 22273
rect 33966 22199 34022 22208
rect 33876 22092 33928 22098
rect 34072 22094 34100 22510
rect 34164 22438 34192 24074
rect 34336 23180 34388 23186
rect 34336 23122 34388 23128
rect 34348 22778 34376 23122
rect 34244 22772 34296 22778
rect 34244 22714 34296 22720
rect 34336 22772 34388 22778
rect 34336 22714 34388 22720
rect 34256 22545 34284 22714
rect 34242 22536 34298 22545
rect 34242 22471 34298 22480
rect 34152 22432 34204 22438
rect 34152 22374 34204 22380
rect 34256 22094 34284 22471
rect 33876 22034 33928 22040
rect 33980 22066 34100 22094
rect 34164 22066 34284 22094
rect 33784 19848 33836 19854
rect 33784 19790 33836 19796
rect 33888 19689 33916 22034
rect 33874 19680 33930 19689
rect 33874 19615 33930 19624
rect 33980 18970 34008 22066
rect 34060 19916 34112 19922
rect 34060 19858 34112 19864
rect 33968 18964 34020 18970
rect 33968 18906 34020 18912
rect 33600 18352 33652 18358
rect 33600 18294 33652 18300
rect 33600 18216 33652 18222
rect 33600 18158 33652 18164
rect 33508 17740 33560 17746
rect 33508 17682 33560 17688
rect 32968 17610 33272 17626
rect 32968 17604 33284 17610
rect 32968 17598 33232 17604
rect 33428 17598 33548 17626
rect 33232 17546 33284 17552
rect 33324 17536 33376 17542
rect 32876 17496 33088 17524
rect 32680 17478 32732 17484
rect 32588 17128 32640 17134
rect 32588 17070 32640 17076
rect 32600 16028 32628 17070
rect 32692 16454 32720 17478
rect 33060 17270 33088 17496
rect 33324 17478 33376 17484
rect 33048 17264 33100 17270
rect 33048 17206 33100 17212
rect 32956 17128 33008 17134
rect 32784 17088 32956 17116
rect 32784 16522 32812 17088
rect 32956 17070 33008 17076
rect 33060 16980 33088 17206
rect 32876 16952 33088 16980
rect 32772 16516 32824 16522
rect 32876 16504 32904 16952
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 32956 16516 33008 16522
rect 32876 16476 32956 16504
rect 32772 16458 32824 16464
rect 32956 16458 33008 16464
rect 32680 16448 32732 16454
rect 32680 16390 32732 16396
rect 32968 16250 32996 16458
rect 32956 16244 33008 16250
rect 32956 16186 33008 16192
rect 33336 16114 33364 17478
rect 33416 16448 33468 16454
rect 33416 16390 33468 16396
rect 33324 16108 33376 16114
rect 33324 16050 33376 16056
rect 32772 16040 32824 16046
rect 32600 16000 32772 16028
rect 32600 15706 32628 16000
rect 32772 15982 32824 15988
rect 32772 15904 32824 15910
rect 32772 15846 32824 15852
rect 32864 15904 32916 15910
rect 32864 15846 32916 15852
rect 32588 15700 32640 15706
rect 32588 15642 32640 15648
rect 32680 15360 32732 15366
rect 32680 15302 32732 15308
rect 32496 14544 32548 14550
rect 32496 14486 32548 14492
rect 32416 14334 32628 14362
rect 32496 13932 32548 13938
rect 32496 13874 32548 13880
rect 32312 13864 32364 13870
rect 32312 13806 32364 13812
rect 32404 12980 32456 12986
rect 32404 12922 32456 12928
rect 32140 12406 32260 12434
rect 32036 12378 32088 12384
rect 31852 11892 31904 11898
rect 31852 11834 31904 11840
rect 31760 11824 31812 11830
rect 31760 11766 31812 11772
rect 31852 11688 31904 11694
rect 31852 11630 31904 11636
rect 31864 10470 31892 11630
rect 32048 11218 32076 12378
rect 32128 12232 32180 12238
rect 32128 12174 32180 12180
rect 32036 11212 32088 11218
rect 32036 11154 32088 11160
rect 32048 11098 32076 11154
rect 31956 11070 32076 11098
rect 31760 10464 31812 10470
rect 31760 10406 31812 10412
rect 31852 10464 31904 10470
rect 31852 10406 31904 10412
rect 31772 9722 31800 10406
rect 31852 9988 31904 9994
rect 31852 9930 31904 9936
rect 31760 9716 31812 9722
rect 31760 9658 31812 9664
rect 31668 9580 31720 9586
rect 31668 9522 31720 9528
rect 31576 9512 31628 9518
rect 31496 9472 31576 9500
rect 31576 9454 31628 9460
rect 31760 9512 31812 9518
rect 31760 9454 31812 9460
rect 31864 9500 31892 9930
rect 31956 9654 31984 11070
rect 32140 11014 32168 12174
rect 32232 11898 32260 12406
rect 32416 12170 32444 12922
rect 32312 12164 32364 12170
rect 32312 12106 32364 12112
rect 32404 12164 32456 12170
rect 32404 12106 32456 12112
rect 32220 11892 32272 11898
rect 32220 11834 32272 11840
rect 32324 11830 32352 12106
rect 32312 11824 32364 11830
rect 32312 11766 32364 11772
rect 32036 11008 32088 11014
rect 32036 10950 32088 10956
rect 32128 11008 32180 11014
rect 32128 10950 32180 10956
rect 32048 10742 32076 10950
rect 32036 10736 32088 10742
rect 32036 10678 32088 10684
rect 32036 10464 32088 10470
rect 32036 10406 32088 10412
rect 31944 9648 31996 9654
rect 31944 9590 31996 9596
rect 31944 9512 31996 9518
rect 31864 9472 31944 9500
rect 31588 9382 31616 9454
rect 31772 9382 31800 9454
rect 31576 9376 31628 9382
rect 31576 9318 31628 9324
rect 31760 9376 31812 9382
rect 31760 9318 31812 9324
rect 30838 9072 30894 9081
rect 30838 9007 30894 9016
rect 31760 9036 31812 9042
rect 30852 8974 30880 9007
rect 31760 8978 31812 8984
rect 30840 8968 30892 8974
rect 30840 8910 30892 8916
rect 30932 8900 30984 8906
rect 30932 8842 30984 8848
rect 30944 8498 30972 8842
rect 31772 8498 31800 8978
rect 30932 8492 30984 8498
rect 30932 8434 30984 8440
rect 31116 8492 31168 8498
rect 31116 8434 31168 8440
rect 31760 8492 31812 8498
rect 31760 8434 31812 8440
rect 31128 7546 31156 8434
rect 31864 8362 31892 9472
rect 31944 9454 31996 9460
rect 32048 8566 32076 10406
rect 32140 10130 32168 10950
rect 32416 10606 32444 12106
rect 32404 10600 32456 10606
rect 32404 10542 32456 10548
rect 32128 10124 32180 10130
rect 32128 10066 32180 10072
rect 32140 9654 32168 10066
rect 32508 10062 32536 13874
rect 32600 11778 32628 14334
rect 32692 12782 32720 15302
rect 32784 14362 32812 15846
rect 32876 14498 32904 15846
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 33324 15360 33376 15366
rect 33428 15314 33456 16390
rect 33376 15308 33456 15314
rect 33324 15302 33456 15308
rect 33336 15286 33456 15302
rect 33324 14816 33376 14822
rect 33324 14758 33376 14764
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 32876 14470 32996 14498
rect 32968 14414 32996 14470
rect 32956 14408 33008 14414
rect 32784 14334 32904 14362
rect 32956 14350 33008 14356
rect 32772 14272 32824 14278
rect 32772 14214 32824 14220
rect 32680 12776 32732 12782
rect 32680 12718 32732 12724
rect 32784 11898 32812 14214
rect 32876 12434 32904 14334
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 33336 13444 33364 14758
rect 33428 14278 33456 15286
rect 33520 14822 33548 17598
rect 33612 17338 33640 18158
rect 33692 17876 33744 17882
rect 33692 17818 33744 17824
rect 33876 17876 33928 17882
rect 33876 17818 33928 17824
rect 33600 17332 33652 17338
rect 33600 17274 33652 17280
rect 33704 17066 33732 17818
rect 33888 17678 33916 17818
rect 33876 17672 33928 17678
rect 33876 17614 33928 17620
rect 33692 17060 33744 17066
rect 33692 17002 33744 17008
rect 33784 16992 33836 16998
rect 33784 16934 33836 16940
rect 33692 16652 33744 16658
rect 33692 16594 33744 16600
rect 33704 16250 33732 16594
rect 33796 16250 33824 16934
rect 34072 16726 34100 19858
rect 34164 19854 34192 22066
rect 34348 21894 34376 22714
rect 34336 21888 34388 21894
rect 34336 21830 34388 21836
rect 34242 21720 34298 21729
rect 34242 21655 34298 21664
rect 34256 21486 34284 21655
rect 34244 21480 34296 21486
rect 34244 21422 34296 21428
rect 34348 21010 34376 21830
rect 34440 21321 34468 26200
rect 34612 24744 34664 24750
rect 34612 24686 34664 24692
rect 34888 24744 34940 24750
rect 34888 24686 34940 24692
rect 34624 24138 34652 24686
rect 34702 24576 34758 24585
rect 34702 24511 34758 24520
rect 34612 24132 34664 24138
rect 34612 24074 34664 24080
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 34532 23050 34560 23462
rect 34612 23248 34664 23254
rect 34612 23190 34664 23196
rect 34520 23044 34572 23050
rect 34520 22986 34572 22992
rect 34624 22710 34652 23190
rect 34716 22817 34744 24511
rect 34796 24064 34848 24070
rect 34796 24006 34848 24012
rect 34702 22808 34758 22817
rect 34702 22743 34758 22752
rect 34612 22704 34664 22710
rect 34612 22646 34664 22652
rect 34612 21888 34664 21894
rect 34612 21830 34664 21836
rect 34426 21312 34482 21321
rect 34426 21247 34482 21256
rect 34336 21004 34388 21010
rect 34336 20946 34388 20952
rect 34336 20800 34388 20806
rect 34336 20742 34388 20748
rect 34152 19848 34204 19854
rect 34152 19790 34204 19796
rect 34152 19712 34204 19718
rect 34152 19654 34204 19660
rect 34060 16720 34112 16726
rect 34060 16662 34112 16668
rect 33968 16448 34020 16454
rect 33968 16390 34020 16396
rect 33692 16244 33744 16250
rect 33692 16186 33744 16192
rect 33784 16244 33836 16250
rect 33784 16186 33836 16192
rect 33704 15706 33732 16186
rect 33692 15700 33744 15706
rect 33692 15642 33744 15648
rect 33692 15360 33744 15366
rect 33692 15302 33744 15308
rect 33876 15360 33928 15366
rect 33876 15302 33928 15308
rect 33508 14816 33560 14822
rect 33508 14758 33560 14764
rect 33508 14340 33560 14346
rect 33508 14282 33560 14288
rect 33416 14272 33468 14278
rect 33416 14214 33468 14220
rect 33244 13416 33364 13444
rect 33244 12782 33272 13416
rect 33232 12776 33284 12782
rect 33232 12718 33284 12724
rect 33324 12640 33376 12646
rect 33324 12582 33376 12588
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 32876 12406 32996 12434
rect 32772 11892 32824 11898
rect 32772 11834 32824 11840
rect 32600 11750 32812 11778
rect 32588 11688 32640 11694
rect 32588 11630 32640 11636
rect 32600 11218 32628 11630
rect 32588 11212 32640 11218
rect 32588 11154 32640 11160
rect 32496 10056 32548 10062
rect 32496 9998 32548 10004
rect 32404 9920 32456 9926
rect 32404 9862 32456 9868
rect 32128 9648 32180 9654
rect 32128 9590 32180 9596
rect 32416 9178 32444 9862
rect 32496 9648 32548 9654
rect 32496 9590 32548 9596
rect 32404 9172 32456 9178
rect 32404 9114 32456 9120
rect 32508 9042 32536 9590
rect 32496 9036 32548 9042
rect 32324 8996 32496 9024
rect 32036 8560 32088 8566
rect 32036 8502 32088 8508
rect 32324 8498 32352 8996
rect 32496 8978 32548 8984
rect 32312 8492 32364 8498
rect 32312 8434 32364 8440
rect 32600 8430 32628 11154
rect 32784 10742 32812 11750
rect 32968 11642 32996 12406
rect 33336 12102 33364 12582
rect 33324 12096 33376 12102
rect 33324 12038 33376 12044
rect 32876 11614 32996 11642
rect 32772 10736 32824 10742
rect 32772 10678 32824 10684
rect 32876 10266 32904 11614
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 32956 11008 33008 11014
rect 32956 10950 33008 10956
rect 32968 10810 32996 10950
rect 32956 10804 33008 10810
rect 32956 10746 33008 10752
rect 33336 10674 33364 12038
rect 33324 10668 33376 10674
rect 33324 10610 33376 10616
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 32864 10260 32916 10266
rect 32864 10202 32916 10208
rect 32772 10124 32824 10130
rect 32772 10066 32824 10072
rect 32680 9988 32732 9994
rect 32680 9930 32732 9936
rect 31944 8424 31996 8430
rect 31944 8366 31996 8372
rect 32220 8424 32272 8430
rect 32220 8366 32272 8372
rect 32588 8424 32640 8430
rect 32588 8366 32640 8372
rect 31852 8356 31904 8362
rect 31852 8298 31904 8304
rect 31956 8294 31984 8366
rect 31944 8288 31996 8294
rect 31944 8230 31996 8236
rect 31392 7744 31444 7750
rect 31392 7686 31444 7692
rect 31404 7546 31432 7686
rect 31116 7540 31168 7546
rect 31116 7482 31168 7488
rect 31392 7540 31444 7546
rect 31392 7482 31444 7488
rect 31956 7478 31984 8230
rect 32232 7954 32260 8366
rect 32588 8016 32640 8022
rect 32588 7958 32640 7964
rect 32220 7948 32272 7954
rect 32220 7890 32272 7896
rect 32600 7750 32628 7958
rect 32692 7886 32720 9930
rect 32784 9450 32812 10066
rect 32772 9444 32824 9450
rect 32772 9386 32824 9392
rect 32864 9376 32916 9382
rect 32864 9318 32916 9324
rect 32772 8900 32824 8906
rect 32772 8842 32824 8848
rect 32784 8634 32812 8842
rect 32876 8838 32904 9318
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 33048 9036 33100 9042
rect 33048 8978 33100 8984
rect 32864 8832 32916 8838
rect 32864 8774 32916 8780
rect 32772 8628 32824 8634
rect 32772 8570 32824 8576
rect 32864 8560 32916 8566
rect 32916 8508 32996 8514
rect 32864 8502 32996 8508
rect 32876 8486 32996 8502
rect 32968 8430 32996 8486
rect 32956 8424 33008 8430
rect 32956 8366 33008 8372
rect 33060 8294 33088 8978
rect 33140 8832 33192 8838
rect 33140 8774 33192 8780
rect 33152 8566 33180 8774
rect 33140 8560 33192 8566
rect 33140 8502 33192 8508
rect 33048 8288 33100 8294
rect 33048 8230 33100 8236
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 32680 7880 32732 7886
rect 32680 7822 32732 7828
rect 32588 7744 32640 7750
rect 32588 7686 32640 7692
rect 31944 7472 31996 7478
rect 31944 7414 31996 7420
rect 32600 7206 32628 7686
rect 32588 7200 32640 7206
rect 32588 7142 32640 7148
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 30748 6384 30800 6390
rect 30748 6326 30800 6332
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 32772 4616 32824 4622
rect 32772 4558 32824 4564
rect 29644 2984 29696 2990
rect 29644 2926 29696 2932
rect 30656 2984 30708 2990
rect 30656 2926 30708 2932
rect 27620 2644 27672 2650
rect 27620 2586 27672 2592
rect 29000 2644 29052 2650
rect 29000 2586 29052 2592
rect 32784 2582 32812 4558
rect 32864 4072 32916 4078
rect 32864 4014 32916 4020
rect 32876 2650 32904 4014
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 33428 3670 33456 14214
rect 33520 12986 33548 14282
rect 33704 14006 33732 15302
rect 33888 15162 33916 15302
rect 33876 15156 33928 15162
rect 33876 15098 33928 15104
rect 33784 14952 33836 14958
rect 33784 14894 33836 14900
rect 33796 14618 33824 14894
rect 33980 14890 34008 16390
rect 34072 15502 34100 16662
rect 34060 15496 34112 15502
rect 34060 15438 34112 15444
rect 33968 14884 34020 14890
rect 33968 14826 34020 14832
rect 34072 14770 34100 15438
rect 33980 14742 34100 14770
rect 33784 14612 33836 14618
rect 33784 14554 33836 14560
rect 33692 14000 33744 14006
rect 33692 13942 33744 13948
rect 33784 13524 33836 13530
rect 33784 13466 33836 13472
rect 33600 13252 33652 13258
rect 33600 13194 33652 13200
rect 33692 13252 33744 13258
rect 33692 13194 33744 13200
rect 33508 12980 33560 12986
rect 33508 12922 33560 12928
rect 33520 11778 33548 12922
rect 33612 12306 33640 13194
rect 33704 12986 33732 13194
rect 33692 12980 33744 12986
rect 33692 12922 33744 12928
rect 33600 12300 33652 12306
rect 33600 12242 33652 12248
rect 33796 11898 33824 13466
rect 33876 13388 33928 13394
rect 33876 13330 33928 13336
rect 33888 12918 33916 13330
rect 33876 12912 33928 12918
rect 33876 12854 33928 12860
rect 33784 11892 33836 11898
rect 33784 11834 33836 11840
rect 33520 11750 33640 11778
rect 33508 11688 33560 11694
rect 33508 11630 33560 11636
rect 33520 11286 33548 11630
rect 33508 11280 33560 11286
rect 33508 11222 33560 11228
rect 33612 8838 33640 11750
rect 33876 11620 33928 11626
rect 33876 11562 33928 11568
rect 33888 10470 33916 11562
rect 33980 11150 34008 14742
rect 34164 13938 34192 19654
rect 34244 19372 34296 19378
rect 34244 19314 34296 19320
rect 34256 18630 34284 19314
rect 34348 18970 34376 20742
rect 34520 20392 34572 20398
rect 34520 20334 34572 20340
rect 34428 19236 34480 19242
rect 34428 19178 34480 19184
rect 34440 18970 34468 19178
rect 34336 18964 34388 18970
rect 34336 18906 34388 18912
rect 34428 18964 34480 18970
rect 34428 18906 34480 18912
rect 34334 18864 34390 18873
rect 34532 18834 34560 20334
rect 34334 18799 34336 18808
rect 34388 18799 34390 18808
rect 34520 18828 34572 18834
rect 34336 18770 34388 18776
rect 34520 18770 34572 18776
rect 34244 18624 34296 18630
rect 34244 18566 34296 18572
rect 34152 13932 34204 13938
rect 34152 13874 34204 13880
rect 34060 13864 34112 13870
rect 34060 13806 34112 13812
rect 34072 13326 34100 13806
rect 34060 13320 34112 13326
rect 34060 13262 34112 13268
rect 34072 12986 34100 13262
rect 34060 12980 34112 12986
rect 34060 12922 34112 12928
rect 34060 12844 34112 12850
rect 34060 12786 34112 12792
rect 34072 11354 34100 12786
rect 34256 12434 34284 18566
rect 34624 18465 34652 21830
rect 34716 21418 34744 22743
rect 34808 22098 34836 24006
rect 34900 22681 34928 24686
rect 34980 23792 35032 23798
rect 34980 23734 35032 23740
rect 34992 23662 35020 23734
rect 34980 23656 35032 23662
rect 34980 23598 35032 23604
rect 35084 23322 35112 26200
rect 35254 24440 35310 24449
rect 35254 24375 35310 24384
rect 35164 24132 35216 24138
rect 35164 24074 35216 24080
rect 35176 24041 35204 24074
rect 35268 24070 35296 24375
rect 35256 24064 35308 24070
rect 35162 24032 35218 24041
rect 35256 24006 35308 24012
rect 35624 24064 35676 24070
rect 35624 24006 35676 24012
rect 35162 23967 35218 23976
rect 35636 23798 35664 24006
rect 35624 23792 35676 23798
rect 35624 23734 35676 23740
rect 35348 23656 35400 23662
rect 35348 23598 35400 23604
rect 35438 23624 35494 23633
rect 35072 23316 35124 23322
rect 35072 23258 35124 23264
rect 35360 23186 35388 23598
rect 35438 23559 35440 23568
rect 35492 23559 35494 23568
rect 35440 23530 35492 23536
rect 35532 23520 35584 23526
rect 35532 23462 35584 23468
rect 35348 23180 35400 23186
rect 35348 23122 35400 23128
rect 35438 23080 35494 23089
rect 35438 23015 35494 23024
rect 35164 22976 35216 22982
rect 35164 22918 35216 22924
rect 34886 22672 34942 22681
rect 34886 22607 34942 22616
rect 34796 22092 34848 22098
rect 34796 22034 34848 22040
rect 34900 21622 34928 22607
rect 35176 22438 35204 22918
rect 35256 22636 35308 22642
rect 35256 22578 35308 22584
rect 35164 22432 35216 22438
rect 35164 22374 35216 22380
rect 34980 22094 35032 22098
rect 35176 22094 35204 22374
rect 34980 22092 35204 22094
rect 35032 22066 35204 22092
rect 34980 22034 35032 22040
rect 34888 21616 34940 21622
rect 34888 21558 34940 21564
rect 34888 21480 34940 21486
rect 34888 21422 34940 21428
rect 34704 21412 34756 21418
rect 34704 21354 34756 21360
rect 34900 21078 34928 21422
rect 35164 21344 35216 21350
rect 35164 21286 35216 21292
rect 34888 21072 34940 21078
rect 34888 21014 34940 21020
rect 34702 20496 34758 20505
rect 34702 20431 34758 20440
rect 34716 19446 34744 20431
rect 34796 20392 34848 20398
rect 34796 20334 34848 20340
rect 34808 19446 34836 20334
rect 34900 20330 34928 21014
rect 35072 20868 35124 20874
rect 35072 20810 35124 20816
rect 35084 20466 35112 20810
rect 35072 20460 35124 20466
rect 35072 20402 35124 20408
rect 34888 20324 34940 20330
rect 34888 20266 34940 20272
rect 34980 20324 35032 20330
rect 34980 20266 35032 20272
rect 34992 20058 35020 20266
rect 34980 20052 35032 20058
rect 34980 19994 35032 20000
rect 35072 19916 35124 19922
rect 35072 19858 35124 19864
rect 34886 19816 34942 19825
rect 34886 19751 34888 19760
rect 34940 19751 34942 19760
rect 34980 19780 35032 19786
rect 34888 19722 34940 19728
rect 34980 19722 35032 19728
rect 34992 19514 35020 19722
rect 34980 19508 35032 19514
rect 34980 19450 35032 19456
rect 34704 19440 34756 19446
rect 34704 19382 34756 19388
rect 34796 19440 34848 19446
rect 34796 19382 34848 19388
rect 34716 18630 34744 19382
rect 34888 19372 34940 19378
rect 34888 19314 34940 19320
rect 34980 19372 35032 19378
rect 34980 19314 35032 19320
rect 34900 18630 34928 19314
rect 34992 19281 35020 19314
rect 34978 19272 35034 19281
rect 34978 19207 35034 19216
rect 34704 18624 34756 18630
rect 34704 18566 34756 18572
rect 34888 18624 34940 18630
rect 34888 18566 34940 18572
rect 34610 18456 34666 18465
rect 34992 18442 35020 19207
rect 34610 18391 34666 18400
rect 34900 18414 35020 18442
rect 34336 18352 34388 18358
rect 34336 18294 34388 18300
rect 34348 17814 34376 18294
rect 34612 18216 34664 18222
rect 34612 18158 34664 18164
rect 34336 17808 34388 17814
rect 34336 17750 34388 17756
rect 34624 17746 34652 18158
rect 34612 17740 34664 17746
rect 34612 17682 34664 17688
rect 34520 17536 34572 17542
rect 34520 17478 34572 17484
rect 34428 16040 34480 16046
rect 34532 16028 34560 17478
rect 34624 16794 34652 17682
rect 34900 17490 34928 18414
rect 35084 17678 35112 19858
rect 35072 17672 35124 17678
rect 35072 17614 35124 17620
rect 35072 17536 35124 17542
rect 34900 17462 35020 17490
rect 35072 17478 35124 17484
rect 34796 17128 34848 17134
rect 34796 17070 34848 17076
rect 34612 16788 34664 16794
rect 34612 16730 34664 16736
rect 34612 16448 34664 16454
rect 34612 16390 34664 16396
rect 34480 16000 34560 16028
rect 34428 15982 34480 15988
rect 34334 13832 34390 13841
rect 34334 13767 34390 13776
rect 34348 12850 34376 13767
rect 34440 13190 34468 15982
rect 34624 15434 34652 16390
rect 34808 16250 34836 17070
rect 34796 16244 34848 16250
rect 34796 16186 34848 16192
rect 34808 15570 34836 16186
rect 34796 15564 34848 15570
rect 34796 15506 34848 15512
rect 34612 15428 34664 15434
rect 34612 15370 34664 15376
rect 34808 14482 34836 15506
rect 34888 14952 34940 14958
rect 34888 14894 34940 14900
rect 34796 14476 34848 14482
rect 34796 14418 34848 14424
rect 34612 14340 34664 14346
rect 34612 14282 34664 14288
rect 34428 13184 34480 13190
rect 34428 13126 34480 13132
rect 34336 12844 34388 12850
rect 34336 12786 34388 12792
rect 34440 12434 34468 13126
rect 34624 12442 34652 14282
rect 34900 14278 34928 14894
rect 34888 14272 34940 14278
rect 34888 14214 34940 14220
rect 34704 13796 34756 13802
rect 34704 13738 34756 13744
rect 34164 12406 34284 12434
rect 34348 12406 34468 12434
rect 34612 12436 34664 12442
rect 34060 11348 34112 11354
rect 34060 11290 34112 11296
rect 33968 11144 34020 11150
rect 33968 11086 34020 11092
rect 33876 10464 33928 10470
rect 33876 10406 33928 10412
rect 34164 9976 34192 12406
rect 34348 12102 34376 12406
rect 34612 12378 34664 12384
rect 34520 12368 34572 12374
rect 34520 12310 34572 12316
rect 34244 12096 34296 12102
rect 34244 12038 34296 12044
rect 34336 12096 34388 12102
rect 34336 12038 34388 12044
rect 34256 11898 34284 12038
rect 34244 11892 34296 11898
rect 34244 11834 34296 11840
rect 34256 10674 34284 11834
rect 34244 10668 34296 10674
rect 34244 10610 34296 10616
rect 34244 9988 34296 9994
rect 34164 9948 34244 9976
rect 34244 9930 34296 9936
rect 34152 9512 34204 9518
rect 34256 9489 34284 9930
rect 34152 9454 34204 9460
rect 34242 9480 34298 9489
rect 33876 9104 33928 9110
rect 33876 9046 33928 9052
rect 33600 8832 33652 8838
rect 33600 8774 33652 8780
rect 33612 8616 33640 8774
rect 33888 8634 33916 9046
rect 34164 9042 34192 9454
rect 34242 9415 34298 9424
rect 34256 9110 34284 9415
rect 34244 9104 34296 9110
rect 34244 9046 34296 9052
rect 34152 9036 34204 9042
rect 34152 8978 34204 8984
rect 34256 8838 34284 9046
rect 34244 8832 34296 8838
rect 34244 8774 34296 8780
rect 33876 8628 33928 8634
rect 33612 8588 33732 8616
rect 33704 8294 33732 8588
rect 33876 8570 33928 8576
rect 33692 8288 33744 8294
rect 33692 8230 33744 8236
rect 33416 3664 33468 3670
rect 33416 3606 33468 3612
rect 34348 2774 34376 12038
rect 34428 10192 34480 10198
rect 34428 10134 34480 10140
rect 34440 7478 34468 10134
rect 34532 7954 34560 12310
rect 34612 11552 34664 11558
rect 34612 11494 34664 11500
rect 34624 11354 34652 11494
rect 34612 11348 34664 11354
rect 34612 11290 34664 11296
rect 34716 10606 34744 13738
rect 34888 13320 34940 13326
rect 34888 13262 34940 13268
rect 34900 12918 34928 13262
rect 34888 12912 34940 12918
rect 34888 12854 34940 12860
rect 34796 12708 34848 12714
rect 34796 12650 34848 12656
rect 34808 11898 34836 12650
rect 34900 12238 34928 12854
rect 34992 12434 35020 17462
rect 35084 17338 35112 17478
rect 35072 17332 35124 17338
rect 35072 17274 35124 17280
rect 35176 17202 35204 21286
rect 35268 18766 35296 22578
rect 35452 22234 35480 23015
rect 35544 22778 35572 23462
rect 35728 23186 35756 26200
rect 36360 24200 36412 24206
rect 36360 24142 36412 24148
rect 36084 24064 36136 24070
rect 36084 24006 36136 24012
rect 35992 23724 36044 23730
rect 35992 23666 36044 23672
rect 35716 23180 35768 23186
rect 35716 23122 35768 23128
rect 35532 22772 35584 22778
rect 35532 22714 35584 22720
rect 35544 22234 35572 22714
rect 35440 22228 35492 22234
rect 35440 22170 35492 22176
rect 35532 22228 35584 22234
rect 35532 22170 35584 22176
rect 35452 22094 35480 22170
rect 35452 22066 35572 22094
rect 35348 20392 35400 20398
rect 35400 20340 35480 20346
rect 35348 20334 35480 20340
rect 35360 20318 35480 20334
rect 35346 20088 35402 20097
rect 35452 20058 35480 20318
rect 35346 20023 35402 20032
rect 35440 20052 35492 20058
rect 35360 19553 35388 20023
rect 35440 19994 35492 20000
rect 35346 19544 35402 19553
rect 35346 19479 35402 19488
rect 35348 19440 35400 19446
rect 35452 19428 35480 19994
rect 35544 19854 35572 22066
rect 35808 21956 35860 21962
rect 35808 21898 35860 21904
rect 35820 21350 35848 21898
rect 36004 21894 36032 23666
rect 36096 23361 36124 24006
rect 36082 23352 36138 23361
rect 36082 23287 36138 23296
rect 36372 23254 36400 24142
rect 36360 23248 36412 23254
rect 36360 23190 36412 23196
rect 36360 22500 36412 22506
rect 36360 22442 36412 22448
rect 35992 21888 36044 21894
rect 35992 21830 36044 21836
rect 36268 21888 36320 21894
rect 36268 21830 36320 21836
rect 35900 21684 35952 21690
rect 35900 21626 35952 21632
rect 35716 21344 35768 21350
rect 35716 21286 35768 21292
rect 35808 21344 35860 21350
rect 35808 21286 35860 21292
rect 35728 21146 35756 21286
rect 35716 21140 35768 21146
rect 35716 21082 35768 21088
rect 35716 20256 35768 20262
rect 35716 20198 35768 20204
rect 35728 19922 35756 20198
rect 35820 19922 35848 21286
rect 35716 19916 35768 19922
rect 35716 19858 35768 19864
rect 35808 19916 35860 19922
rect 35808 19858 35860 19864
rect 35532 19848 35584 19854
rect 35532 19790 35584 19796
rect 35400 19400 35480 19428
rect 35348 19382 35400 19388
rect 35256 18760 35308 18766
rect 35256 18702 35308 18708
rect 35256 17672 35308 17678
rect 35256 17614 35308 17620
rect 35164 17196 35216 17202
rect 35164 17138 35216 17144
rect 35164 16040 35216 16046
rect 35164 15982 35216 15988
rect 35176 14346 35204 15982
rect 35164 14340 35216 14346
rect 35164 14282 35216 14288
rect 35176 14006 35204 14282
rect 35164 14000 35216 14006
rect 35164 13942 35216 13948
rect 35162 13288 35218 13297
rect 35162 13223 35164 13232
rect 35216 13223 35218 13232
rect 35164 13194 35216 13200
rect 35176 12986 35204 13194
rect 35164 12980 35216 12986
rect 35164 12922 35216 12928
rect 35268 12782 35296 17614
rect 35346 17368 35402 17377
rect 35346 17303 35402 17312
rect 35360 16658 35388 17303
rect 35348 16652 35400 16658
rect 35348 16594 35400 16600
rect 35452 15473 35480 19400
rect 35532 19372 35584 19378
rect 35532 19314 35584 19320
rect 35544 18426 35572 19314
rect 35624 18692 35676 18698
rect 35624 18634 35676 18640
rect 35532 18420 35584 18426
rect 35532 18362 35584 18368
rect 35636 18086 35664 18634
rect 35716 18284 35768 18290
rect 35716 18226 35768 18232
rect 35624 18080 35676 18086
rect 35624 18022 35676 18028
rect 35532 17536 35584 17542
rect 35530 17504 35532 17513
rect 35584 17504 35586 17513
rect 35530 17439 35586 17448
rect 35544 17270 35572 17439
rect 35532 17264 35584 17270
rect 35532 17206 35584 17212
rect 35544 16590 35572 17206
rect 35624 16992 35676 16998
rect 35624 16934 35676 16940
rect 35532 16584 35584 16590
rect 35532 16526 35584 16532
rect 35532 16108 35584 16114
rect 35532 16050 35584 16056
rect 35544 15706 35572 16050
rect 35532 15700 35584 15706
rect 35532 15642 35584 15648
rect 35438 15464 35494 15473
rect 35438 15399 35494 15408
rect 35544 15416 35572 15642
rect 35636 15609 35664 16934
rect 35622 15600 35678 15609
rect 35622 15535 35678 15544
rect 35624 15428 35676 15434
rect 35544 15388 35624 15416
rect 35624 15370 35676 15376
rect 35636 14346 35664 15370
rect 35624 14340 35676 14346
rect 35624 14282 35676 14288
rect 35636 13705 35664 14282
rect 35622 13696 35678 13705
rect 35622 13631 35678 13640
rect 35636 13190 35664 13631
rect 35728 13530 35756 18226
rect 35820 16454 35848 19858
rect 35912 19446 35940 21626
rect 36176 21480 36228 21486
rect 36176 21422 36228 21428
rect 36082 20768 36138 20777
rect 36082 20703 36138 20712
rect 36096 20330 36124 20703
rect 36188 20602 36216 21422
rect 36176 20596 36228 20602
rect 36176 20538 36228 20544
rect 36084 20324 36136 20330
rect 36084 20266 36136 20272
rect 36280 19786 36308 21830
rect 36372 20874 36400 22442
rect 36464 21457 36492 26302
rect 37002 26200 37058 27000
rect 37646 26200 37702 27000
rect 38290 26200 38346 27000
rect 38934 26200 38990 27000
rect 39578 26200 39634 27000
rect 40222 26200 40278 27000
rect 42154 26330 42210 27000
rect 42154 26302 42748 26330
rect 42154 26200 42210 26302
rect 36728 24268 36780 24274
rect 36728 24210 36780 24216
rect 36634 21992 36690 22001
rect 36634 21927 36690 21936
rect 36544 21888 36596 21894
rect 36544 21830 36596 21836
rect 36450 21448 36506 21457
rect 36450 21383 36506 21392
rect 36360 20868 36412 20874
rect 36360 20810 36412 20816
rect 36372 20534 36400 20810
rect 36360 20528 36412 20534
rect 36360 20470 36412 20476
rect 36556 20330 36584 21830
rect 36648 21185 36676 21927
rect 36634 21176 36690 21185
rect 36740 21146 36768 24210
rect 36820 24132 36872 24138
rect 36820 24074 36872 24080
rect 36832 21894 36860 24074
rect 36912 23520 36964 23526
rect 36912 23462 36964 23468
rect 36924 23050 36952 23462
rect 36912 23044 36964 23050
rect 36912 22986 36964 22992
rect 37016 22001 37044 26200
rect 37280 24268 37332 24274
rect 37280 24210 37332 24216
rect 37188 23248 37240 23254
rect 37188 23190 37240 23196
rect 37096 22976 37148 22982
rect 37096 22918 37148 22924
rect 37108 22506 37136 22918
rect 37096 22500 37148 22506
rect 37096 22442 37148 22448
rect 37200 22137 37228 23190
rect 37186 22128 37242 22137
rect 37186 22063 37242 22072
rect 37002 21992 37058 22001
rect 37002 21927 37058 21936
rect 37188 21956 37240 21962
rect 37188 21898 37240 21904
rect 36820 21888 36872 21894
rect 36820 21830 36872 21836
rect 36910 21720 36966 21729
rect 36910 21655 36966 21664
rect 36924 21486 36952 21655
rect 37200 21486 37228 21898
rect 37292 21894 37320 24210
rect 37372 23520 37424 23526
rect 37372 23462 37424 23468
rect 37384 23322 37412 23462
rect 37554 23352 37610 23361
rect 37372 23316 37424 23322
rect 37372 23258 37424 23264
rect 37464 23316 37516 23322
rect 37554 23287 37610 23296
rect 37464 23258 37516 23264
rect 37476 22778 37504 23258
rect 37464 22772 37516 22778
rect 37464 22714 37516 22720
rect 37568 22438 37596 23287
rect 37660 22778 37688 26200
rect 37924 25288 37976 25294
rect 37924 25230 37976 25236
rect 37738 24440 37794 24449
rect 37738 24375 37794 24384
rect 37752 24206 37780 24375
rect 37832 24268 37884 24274
rect 37832 24210 37884 24216
rect 37740 24200 37792 24206
rect 37740 24142 37792 24148
rect 37740 24064 37792 24070
rect 37738 24032 37740 24041
rect 37844 24052 37872 24210
rect 37936 24206 37964 25230
rect 37924 24200 37976 24206
rect 37924 24142 37976 24148
rect 38108 24132 38160 24138
rect 38028 24092 38108 24120
rect 38028 24052 38056 24092
rect 38108 24074 38160 24080
rect 37792 24032 37794 24041
rect 37844 24024 38056 24052
rect 37738 23967 37794 23976
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 37648 22772 37700 22778
rect 37648 22714 37700 22720
rect 38304 22681 38332 26200
rect 38948 24818 38976 26200
rect 39592 24886 39620 26200
rect 39580 24880 39632 24886
rect 39580 24822 39632 24828
rect 38936 24812 38988 24818
rect 38936 24754 38988 24760
rect 40236 24682 40264 26200
rect 42064 24812 42116 24818
rect 42064 24754 42116 24760
rect 40316 24744 40368 24750
rect 40316 24686 40368 24692
rect 39948 24676 40000 24682
rect 39948 24618 40000 24624
rect 40224 24676 40276 24682
rect 40224 24618 40276 24624
rect 39488 24608 39540 24614
rect 39488 24550 39540 24556
rect 38660 24404 38712 24410
rect 38660 24346 38712 24352
rect 39304 24404 39356 24410
rect 39304 24346 39356 24352
rect 38672 24313 38700 24346
rect 38658 24304 38714 24313
rect 38658 24239 38714 24248
rect 38660 24064 38712 24070
rect 38712 24024 38792 24052
rect 38660 24006 38712 24012
rect 38568 23656 38620 23662
rect 38568 23598 38620 23604
rect 38580 23202 38608 23598
rect 38580 23186 38700 23202
rect 38384 23180 38436 23186
rect 38580 23180 38712 23186
rect 38580 23174 38660 23180
rect 38384 23122 38436 23128
rect 38660 23122 38712 23128
rect 38290 22672 38346 22681
rect 38290 22607 38346 22616
rect 37556 22432 37608 22438
rect 38396 22409 38424 23122
rect 38660 22976 38712 22982
rect 38660 22918 38712 22924
rect 38566 22808 38622 22817
rect 38566 22743 38568 22752
rect 38620 22743 38622 22752
rect 38568 22714 38620 22720
rect 38672 22710 38700 22918
rect 38764 22778 38792 24024
rect 39212 23724 39264 23730
rect 39212 23666 39264 23672
rect 39224 22953 39252 23666
rect 39316 23089 39344 24346
rect 39500 24206 39528 24550
rect 39854 24440 39910 24449
rect 39854 24375 39856 24384
rect 39908 24375 39910 24384
rect 39856 24346 39908 24352
rect 39764 24336 39816 24342
rect 39764 24278 39816 24284
rect 39488 24200 39540 24206
rect 39488 24142 39540 24148
rect 39672 24132 39724 24138
rect 39672 24074 39724 24080
rect 39684 23798 39712 24074
rect 39672 23792 39724 23798
rect 39672 23734 39724 23740
rect 39396 23656 39448 23662
rect 39396 23598 39448 23604
rect 39488 23656 39540 23662
rect 39488 23598 39540 23604
rect 39302 23080 39358 23089
rect 39302 23015 39358 23024
rect 39210 22944 39266 22953
rect 39210 22879 39266 22888
rect 38752 22772 38804 22778
rect 38752 22714 38804 22720
rect 38660 22704 38712 22710
rect 38660 22646 38712 22652
rect 38844 22704 38896 22710
rect 38844 22646 38896 22652
rect 38672 22488 38700 22646
rect 38580 22460 38700 22488
rect 37556 22374 37608 22380
rect 38382 22400 38438 22409
rect 38382 22335 38438 22344
rect 38580 22094 38608 22460
rect 38752 22432 38804 22438
rect 38672 22380 38752 22386
rect 38672 22374 38804 22380
rect 38672 22358 38792 22374
rect 38672 22234 38700 22358
rect 38856 22250 38884 22646
rect 39120 22432 39172 22438
rect 39120 22374 39172 22380
rect 38764 22234 38884 22250
rect 38660 22228 38712 22234
rect 38660 22170 38712 22176
rect 38764 22228 38896 22234
rect 38764 22222 38844 22228
rect 38764 22114 38792 22222
rect 38844 22170 38896 22176
rect 38488 22066 38608 22094
rect 38672 22086 38792 22114
rect 38842 22128 38898 22137
rect 37556 21956 37608 21962
rect 38384 21956 38436 21962
rect 37608 21916 37780 21944
rect 37556 21898 37608 21904
rect 37280 21888 37332 21894
rect 37280 21830 37332 21836
rect 37464 21888 37516 21894
rect 37464 21830 37516 21836
rect 37292 21622 37320 21830
rect 37476 21690 37504 21830
rect 37464 21684 37516 21690
rect 37464 21626 37516 21632
rect 37556 21684 37608 21690
rect 37752 21672 37780 21916
rect 38488 21944 38516 22066
rect 38436 21916 38516 21944
rect 38384 21898 38436 21904
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 37752 21644 38148 21672
rect 37556 21626 37608 21632
rect 37280 21616 37332 21622
rect 37280 21558 37332 21564
rect 36912 21480 36964 21486
rect 36912 21422 36964 21428
rect 37188 21480 37240 21486
rect 37188 21422 37240 21428
rect 36634 21111 36690 21120
rect 36728 21140 36780 21146
rect 36728 21082 36780 21088
rect 36636 20596 36688 20602
rect 36636 20538 36688 20544
rect 36648 20398 36676 20538
rect 36636 20392 36688 20398
rect 36636 20334 36688 20340
rect 36544 20324 36596 20330
rect 36544 20266 36596 20272
rect 36820 20256 36872 20262
rect 36820 20198 36872 20204
rect 36452 19916 36504 19922
rect 36452 19858 36504 19864
rect 36268 19780 36320 19786
rect 36268 19722 36320 19728
rect 35992 19712 36044 19718
rect 35992 19654 36044 19660
rect 35900 19440 35952 19446
rect 35900 19382 35952 19388
rect 35900 19304 35952 19310
rect 35900 19246 35952 19252
rect 35912 16522 35940 19246
rect 35900 16516 35952 16522
rect 35900 16458 35952 16464
rect 35808 16448 35860 16454
rect 35808 16390 35860 16396
rect 35806 16008 35862 16017
rect 35806 15943 35862 15952
rect 35820 14521 35848 15943
rect 35912 15570 35940 16458
rect 35900 15564 35952 15570
rect 35900 15506 35952 15512
rect 36004 15094 36032 19654
rect 36084 19304 36136 19310
rect 36084 19246 36136 19252
rect 36096 18601 36124 19246
rect 36082 18592 36138 18601
rect 36082 18527 36138 18536
rect 36360 18284 36412 18290
rect 36360 18226 36412 18232
rect 36372 18086 36400 18226
rect 36464 18222 36492 19858
rect 36544 19712 36596 19718
rect 36544 19654 36596 19660
rect 36556 19514 36584 19654
rect 36544 19508 36596 19514
rect 36544 19450 36596 19456
rect 36728 19372 36780 19378
rect 36728 19314 36780 19320
rect 36636 19168 36688 19174
rect 36636 19110 36688 19116
rect 36544 18828 36596 18834
rect 36544 18770 36596 18776
rect 36452 18216 36504 18222
rect 36452 18158 36504 18164
rect 36360 18080 36412 18086
rect 36360 18022 36412 18028
rect 36188 17326 36492 17354
rect 36188 17134 36216 17326
rect 36360 17196 36412 17202
rect 36360 17138 36412 17144
rect 36176 17128 36228 17134
rect 36176 17070 36228 17076
rect 36084 17060 36136 17066
rect 36084 17002 36136 17008
rect 36096 16674 36124 17002
rect 36372 16794 36400 17138
rect 36464 16794 36492 17326
rect 36360 16788 36412 16794
rect 36360 16730 36412 16736
rect 36452 16788 36504 16794
rect 36452 16730 36504 16736
rect 36096 16646 36308 16674
rect 36084 16516 36136 16522
rect 36084 16458 36136 16464
rect 36096 16046 36124 16458
rect 36084 16040 36136 16046
rect 36084 15982 36136 15988
rect 36280 15094 36308 16646
rect 36452 15360 36504 15366
rect 36452 15302 36504 15308
rect 35992 15088 36044 15094
rect 35992 15030 36044 15036
rect 36268 15088 36320 15094
rect 36268 15030 36320 15036
rect 35900 15020 35952 15026
rect 35900 14962 35952 14968
rect 35912 14929 35940 14962
rect 36084 14952 36136 14958
rect 35898 14920 35954 14929
rect 36268 14952 36320 14958
rect 36136 14912 36216 14940
rect 36084 14894 36136 14900
rect 35898 14855 35954 14864
rect 35806 14512 35862 14521
rect 35806 14447 35862 14456
rect 36084 13932 36136 13938
rect 36084 13874 36136 13880
rect 35992 13864 36044 13870
rect 35992 13806 36044 13812
rect 35716 13524 35768 13530
rect 35716 13466 35768 13472
rect 35624 13184 35676 13190
rect 35624 13126 35676 13132
rect 35256 12776 35308 12782
rect 35256 12718 35308 12724
rect 35624 12776 35676 12782
rect 35624 12718 35676 12724
rect 35636 12646 35664 12718
rect 35624 12640 35676 12646
rect 35624 12582 35676 12588
rect 35636 12442 35664 12582
rect 35624 12436 35676 12442
rect 34992 12406 35204 12434
rect 34888 12232 34940 12238
rect 34888 12174 34940 12180
rect 34796 11892 34848 11898
rect 34796 11834 34848 11840
rect 34900 11694 34928 12174
rect 34980 11892 35032 11898
rect 34980 11834 35032 11840
rect 34888 11688 34940 11694
rect 34888 11630 34940 11636
rect 34992 11234 35020 11834
rect 35072 11620 35124 11626
rect 35072 11562 35124 11568
rect 35084 11354 35112 11562
rect 35072 11348 35124 11354
rect 35072 11290 35124 11296
rect 34992 11206 35112 11234
rect 34704 10600 34756 10606
rect 34704 10542 34756 10548
rect 34716 10130 34744 10542
rect 34796 10464 34848 10470
rect 34796 10406 34848 10412
rect 34704 10124 34756 10130
rect 34704 10066 34756 10072
rect 34808 8974 34836 10406
rect 34888 10056 34940 10062
rect 34888 9998 34940 10004
rect 34900 9722 34928 9998
rect 34888 9716 34940 9722
rect 34888 9658 34940 9664
rect 35084 9042 35112 11206
rect 35176 10577 35204 12406
rect 35624 12378 35676 12384
rect 35440 12096 35492 12102
rect 35440 12038 35492 12044
rect 35452 11694 35480 12038
rect 35900 11824 35952 11830
rect 35900 11766 35952 11772
rect 35440 11688 35492 11694
rect 35440 11630 35492 11636
rect 35624 11552 35676 11558
rect 35624 11494 35676 11500
rect 35636 10674 35664 11494
rect 35912 11218 35940 11766
rect 36004 11286 36032 13806
rect 36096 11898 36124 13874
rect 36188 12102 36216 14912
rect 36268 14894 36320 14900
rect 36176 12096 36228 12102
rect 36176 12038 36228 12044
rect 36084 11892 36136 11898
rect 36084 11834 36136 11840
rect 35992 11280 36044 11286
rect 35992 11222 36044 11228
rect 35900 11212 35952 11218
rect 35900 11154 35952 11160
rect 35900 11076 35952 11082
rect 35900 11018 35952 11024
rect 35624 10668 35676 10674
rect 35624 10610 35676 10616
rect 35162 10568 35218 10577
rect 35162 10503 35218 10512
rect 35624 10532 35676 10538
rect 35624 10474 35676 10480
rect 35636 10282 35664 10474
rect 35544 10254 35664 10282
rect 35164 10124 35216 10130
rect 35164 10066 35216 10072
rect 35176 9722 35204 10066
rect 35440 9988 35492 9994
rect 35544 9976 35572 10254
rect 35492 9948 35572 9976
rect 35440 9930 35492 9936
rect 35808 9920 35860 9926
rect 35808 9862 35860 9868
rect 35164 9716 35216 9722
rect 35164 9658 35216 9664
rect 35532 9376 35584 9382
rect 35532 9318 35584 9324
rect 35544 9042 35572 9318
rect 34980 9036 35032 9042
rect 34980 8978 35032 8984
rect 35072 9036 35124 9042
rect 35072 8978 35124 8984
rect 35532 9036 35584 9042
rect 35532 8978 35584 8984
rect 34796 8968 34848 8974
rect 34796 8910 34848 8916
rect 34992 8634 35020 8978
rect 35256 8832 35308 8838
rect 35256 8774 35308 8780
rect 35624 8832 35676 8838
rect 35624 8774 35676 8780
rect 34980 8628 35032 8634
rect 34980 8570 35032 8576
rect 35268 8090 35296 8774
rect 35636 8566 35664 8774
rect 35624 8560 35676 8566
rect 35624 8502 35676 8508
rect 35820 8498 35848 9862
rect 35912 9518 35940 11018
rect 36084 9920 36136 9926
rect 36084 9862 36136 9868
rect 36096 9722 36124 9862
rect 36084 9716 36136 9722
rect 36084 9658 36136 9664
rect 35992 9648 36044 9654
rect 35992 9590 36044 9596
rect 35900 9512 35952 9518
rect 35900 9454 35952 9460
rect 36004 8634 36032 9590
rect 36280 9110 36308 14894
rect 36360 14544 36412 14550
rect 36360 14486 36412 14492
rect 36372 13734 36400 14486
rect 36360 13728 36412 13734
rect 36360 13670 36412 13676
rect 36464 13274 36492 15302
rect 36556 14890 36584 18770
rect 36648 17542 36676 19110
rect 36740 17746 36768 19314
rect 36832 19281 36860 20198
rect 36818 19272 36874 19281
rect 36818 19207 36874 19216
rect 36832 19174 36860 19207
rect 36820 19168 36872 19174
rect 36820 19110 36872 19116
rect 36832 18057 36860 19110
rect 36924 18426 36952 21422
rect 37004 20800 37056 20806
rect 37004 20742 37056 20748
rect 37016 20058 37044 20742
rect 37096 20528 37148 20534
rect 37096 20470 37148 20476
rect 37004 20052 37056 20058
rect 37004 19994 37056 20000
rect 37016 19514 37044 19994
rect 37004 19508 37056 19514
rect 37004 19450 37056 19456
rect 37108 19009 37136 20470
rect 37188 20460 37240 20466
rect 37188 20402 37240 20408
rect 37094 19000 37150 19009
rect 37094 18935 37150 18944
rect 36912 18420 36964 18426
rect 36912 18362 36964 18368
rect 36818 18048 36874 18057
rect 36818 17983 36874 17992
rect 36728 17740 36780 17746
rect 36728 17682 36780 17688
rect 36636 17536 36688 17542
rect 36636 17478 36688 17484
rect 36728 16992 36780 16998
rect 36728 16934 36780 16940
rect 36636 16788 36688 16794
rect 36636 16730 36688 16736
rect 36544 14884 36596 14890
rect 36544 14826 36596 14832
rect 36648 14618 36676 16730
rect 36636 14612 36688 14618
rect 36636 14554 36688 14560
rect 36648 13802 36676 14554
rect 36740 14006 36768 16934
rect 36924 16776 36952 18362
rect 37004 18352 37056 18358
rect 37004 18294 37056 18300
rect 37016 17610 37044 18294
rect 37096 18080 37148 18086
rect 37096 18022 37148 18028
rect 37004 17604 37056 17610
rect 37004 17546 37056 17552
rect 36832 16748 36952 16776
rect 36832 16658 36860 16748
rect 36820 16652 36872 16658
rect 36820 16594 36872 16600
rect 36832 16522 36860 16594
rect 36820 16516 36872 16522
rect 36820 16458 36872 16464
rect 37108 16250 37136 18022
rect 37200 17066 37228 20402
rect 37292 18630 37320 21558
rect 37568 21486 37596 21626
rect 37740 21548 37792 21554
rect 37740 21490 37792 21496
rect 37556 21480 37608 21486
rect 37556 21422 37608 21428
rect 37568 21350 37596 21422
rect 37752 21350 37780 21490
rect 38120 21350 38148 21644
rect 38292 21616 38344 21622
rect 38292 21558 38344 21564
rect 37556 21344 37608 21350
rect 37556 21286 37608 21292
rect 37740 21344 37792 21350
rect 37740 21286 37792 21292
rect 38108 21344 38160 21350
rect 38108 21286 38160 21292
rect 37568 20874 37596 21286
rect 37648 21140 37700 21146
rect 37648 21082 37700 21088
rect 37556 20868 37608 20874
rect 37556 20810 37608 20816
rect 37370 20632 37426 20641
rect 37370 20567 37426 20576
rect 37384 19854 37412 20567
rect 37464 20392 37516 20398
rect 37464 20334 37516 20340
rect 37372 19848 37424 19854
rect 37372 19790 37424 19796
rect 37372 19372 37424 19378
rect 37372 19314 37424 19320
rect 37384 18698 37412 19314
rect 37372 18692 37424 18698
rect 37372 18634 37424 18640
rect 37280 18624 37332 18630
rect 37280 18566 37332 18572
rect 37384 18426 37412 18634
rect 37372 18420 37424 18426
rect 37372 18362 37424 18368
rect 37476 18290 37504 20334
rect 37568 19718 37596 20810
rect 37660 20398 37688 21082
rect 38304 20806 38332 21558
rect 38396 21146 38424 21898
rect 38384 21140 38436 21146
rect 38384 21082 38436 21088
rect 38396 20890 38424 21082
rect 38672 21010 38700 22086
rect 38842 22063 38844 22072
rect 38896 22063 38898 22072
rect 38844 22034 38896 22040
rect 39132 21842 39160 22374
rect 39408 22098 39436 23598
rect 39500 23361 39528 23598
rect 39486 23352 39542 23361
rect 39486 23287 39542 23296
rect 39488 23180 39540 23186
rect 39488 23122 39540 23128
rect 39500 22642 39528 23122
rect 39672 22976 39724 22982
rect 39672 22918 39724 22924
rect 39488 22636 39540 22642
rect 39488 22578 39540 22584
rect 39500 22234 39528 22578
rect 39488 22228 39540 22234
rect 39488 22170 39540 22176
rect 39396 22092 39448 22098
rect 39500 22094 39528 22170
rect 39500 22066 39620 22094
rect 39396 22034 39448 22040
rect 39040 21814 39160 21842
rect 39040 21350 39068 21814
rect 39120 21684 39172 21690
rect 39120 21626 39172 21632
rect 39212 21684 39264 21690
rect 39212 21626 39264 21632
rect 38844 21344 38896 21350
rect 38844 21286 38896 21292
rect 39028 21344 39080 21350
rect 39028 21286 39080 21292
rect 38660 21004 38712 21010
rect 38660 20946 38712 20952
rect 38396 20874 38516 20890
rect 38384 20868 38516 20874
rect 38436 20862 38516 20868
rect 38384 20810 38436 20816
rect 38292 20800 38344 20806
rect 38292 20742 38344 20748
rect 38382 20768 38438 20777
rect 37950 20700 38258 20709
rect 38382 20703 38438 20712
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 37648 20392 37700 20398
rect 37648 20334 37700 20340
rect 37740 20256 37792 20262
rect 37740 20198 37792 20204
rect 37648 19916 37700 19922
rect 37648 19858 37700 19864
rect 37556 19712 37608 19718
rect 37556 19654 37608 19660
rect 37568 18630 37596 19654
rect 37556 18624 37608 18630
rect 37556 18566 37608 18572
rect 37464 18284 37516 18290
rect 37464 18226 37516 18232
rect 37280 18216 37332 18222
rect 37332 18164 37412 18170
rect 37280 18158 37412 18164
rect 37292 18142 37412 18158
rect 37384 18136 37412 18142
rect 37568 18136 37596 18566
rect 37384 18108 37596 18136
rect 37280 18080 37332 18086
rect 37280 18022 37332 18028
rect 37292 17864 37320 18022
rect 37292 17836 37504 17864
rect 37280 17740 37332 17746
rect 37280 17682 37332 17688
rect 37188 17060 37240 17066
rect 37188 17002 37240 17008
rect 37188 16788 37240 16794
rect 37188 16730 37240 16736
rect 37200 16454 37228 16730
rect 37188 16448 37240 16454
rect 37188 16390 37240 16396
rect 37096 16244 37148 16250
rect 37096 16186 37148 16192
rect 37004 16040 37056 16046
rect 37004 15982 37056 15988
rect 37016 15162 37044 15982
rect 37004 15156 37056 15162
rect 37004 15098 37056 15104
rect 37096 14952 37148 14958
rect 37096 14894 37148 14900
rect 37108 14618 37136 14894
rect 37096 14612 37148 14618
rect 37096 14554 37148 14560
rect 37096 14476 37148 14482
rect 37096 14418 37148 14424
rect 36820 14340 36872 14346
rect 36820 14282 36872 14288
rect 36728 14000 36780 14006
rect 36728 13942 36780 13948
rect 36636 13796 36688 13802
rect 36636 13738 36688 13744
rect 36372 13258 36492 13274
rect 36648 13258 36676 13738
rect 36728 13728 36780 13734
rect 36726 13696 36728 13705
rect 36832 13716 36860 14282
rect 36780 13696 36860 13716
rect 36782 13688 36860 13696
rect 36726 13631 36782 13640
rect 36360 13252 36492 13258
rect 36412 13246 36492 13252
rect 36636 13252 36688 13258
rect 36360 13194 36412 13200
rect 36636 13194 36688 13200
rect 37004 12912 37056 12918
rect 37004 12854 37056 12860
rect 36636 12436 36688 12442
rect 36636 12378 36688 12384
rect 36648 12102 36676 12378
rect 36636 12096 36688 12102
rect 36636 12038 36688 12044
rect 36820 11756 36872 11762
rect 36820 11698 36872 11704
rect 36636 11688 36688 11694
rect 36636 11630 36688 11636
rect 36648 10742 36676 11630
rect 36832 10810 36860 11698
rect 36912 11212 36964 11218
rect 36912 11154 36964 11160
rect 36924 10810 36952 11154
rect 36820 10804 36872 10810
rect 36820 10746 36872 10752
rect 36912 10804 36964 10810
rect 36912 10746 36964 10752
rect 36636 10736 36688 10742
rect 36636 10678 36688 10684
rect 36452 10668 36504 10674
rect 36452 10610 36504 10616
rect 36360 10600 36412 10606
rect 36360 10542 36412 10548
rect 36372 9178 36400 10542
rect 36360 9172 36412 9178
rect 36360 9114 36412 9120
rect 36268 9104 36320 9110
rect 36266 9072 36268 9081
rect 36320 9072 36322 9081
rect 36266 9007 36322 9016
rect 36464 8906 36492 10610
rect 36648 10266 36676 10678
rect 36924 10266 36952 10746
rect 36636 10260 36688 10266
rect 36636 10202 36688 10208
rect 36912 10260 36964 10266
rect 36912 10202 36964 10208
rect 36924 9994 36952 10202
rect 36912 9988 36964 9994
rect 36912 9930 36964 9936
rect 36452 8900 36504 8906
rect 36452 8842 36504 8848
rect 35992 8628 36044 8634
rect 35992 8570 36044 8576
rect 35808 8492 35860 8498
rect 35808 8434 35860 8440
rect 35256 8084 35308 8090
rect 35256 8026 35308 8032
rect 34520 7948 34572 7954
rect 34520 7890 34572 7896
rect 34428 7472 34480 7478
rect 34428 7414 34480 7420
rect 37016 4758 37044 12854
rect 37108 12238 37136 14418
rect 37200 12918 37228 16390
rect 37292 15978 37320 17682
rect 37372 17604 37424 17610
rect 37372 17546 37424 17552
rect 37384 16232 37412 17546
rect 37476 16794 37504 17836
rect 37568 17678 37596 18108
rect 37556 17672 37608 17678
rect 37556 17614 37608 17620
rect 37464 16788 37516 16794
rect 37464 16730 37516 16736
rect 37568 16726 37596 17614
rect 37556 16720 37608 16726
rect 37556 16662 37608 16668
rect 37464 16652 37516 16658
rect 37464 16594 37516 16600
rect 37476 16538 37504 16594
rect 37476 16510 37596 16538
rect 37384 16204 37504 16232
rect 37372 16108 37424 16114
rect 37372 16050 37424 16056
rect 37280 15972 37332 15978
rect 37280 15914 37332 15920
rect 37292 15706 37320 15914
rect 37280 15700 37332 15706
rect 37280 15642 37332 15648
rect 37384 15570 37412 16050
rect 37372 15564 37424 15570
rect 37372 15506 37424 15512
rect 37384 15026 37412 15506
rect 37372 15020 37424 15026
rect 37372 14962 37424 14968
rect 37384 14482 37412 14962
rect 37476 14822 37504 16204
rect 37464 14816 37516 14822
rect 37464 14758 37516 14764
rect 37372 14476 37424 14482
rect 37372 14418 37424 14424
rect 37568 14278 37596 16510
rect 37660 15162 37688 19858
rect 37752 19242 37780 20198
rect 38396 20058 38424 20703
rect 38488 20534 38516 20862
rect 38476 20528 38528 20534
rect 38476 20470 38528 20476
rect 38384 20052 38436 20058
rect 38384 19994 38436 20000
rect 38488 19990 38516 20470
rect 38856 20058 38884 21286
rect 39040 20874 39068 21286
rect 39132 21010 39160 21626
rect 39120 21004 39172 21010
rect 39120 20946 39172 20952
rect 39028 20868 39080 20874
rect 39028 20810 39080 20816
rect 38844 20052 38896 20058
rect 38844 19994 38896 20000
rect 38476 19984 38528 19990
rect 38476 19926 38528 19932
rect 38384 19712 38436 19718
rect 38384 19654 38436 19660
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 37740 19236 37792 19242
rect 37740 19178 37792 19184
rect 37752 18358 37780 19178
rect 37832 19168 37884 19174
rect 37832 19110 37884 19116
rect 37740 18352 37792 18358
rect 37740 18294 37792 18300
rect 37844 18222 37872 19110
rect 38290 19000 38346 19009
rect 38290 18935 38346 18944
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 38200 18420 38252 18426
rect 38304 18408 38332 18935
rect 38252 18380 38332 18408
rect 38200 18362 38252 18368
rect 38016 18284 38068 18290
rect 38016 18226 38068 18232
rect 37740 18216 37792 18222
rect 37740 18158 37792 18164
rect 37832 18216 37884 18222
rect 37832 18158 37884 18164
rect 37752 15706 37780 18158
rect 37844 17134 37872 18158
rect 38028 18154 38056 18226
rect 38016 18148 38068 18154
rect 38016 18090 38068 18096
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 37832 17128 37884 17134
rect 37832 17070 37884 17076
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 37740 15700 37792 15706
rect 37740 15642 37792 15648
rect 37648 15156 37700 15162
rect 37648 15098 37700 15104
rect 37660 14278 37688 15098
rect 37752 15094 37780 15642
rect 38396 15337 38424 19654
rect 38488 19514 38516 19926
rect 39224 19922 39252 21626
rect 39408 20097 39436 22034
rect 39592 22030 39620 22066
rect 39580 22024 39632 22030
rect 39580 21966 39632 21972
rect 39592 21010 39620 21966
rect 39684 21894 39712 22918
rect 39672 21888 39724 21894
rect 39672 21830 39724 21836
rect 39684 21622 39712 21830
rect 39672 21616 39724 21622
rect 39672 21558 39724 21564
rect 39776 21010 39804 24278
rect 39856 24064 39908 24070
rect 39856 24006 39908 24012
rect 39868 23610 39896 24006
rect 39960 23730 39988 24618
rect 40132 24200 40184 24206
rect 40132 24142 40184 24148
rect 40040 24064 40092 24070
rect 40040 24006 40092 24012
rect 40052 23866 40080 24006
rect 40144 23866 40172 24142
rect 40328 24070 40356 24686
rect 41144 24132 41196 24138
rect 41144 24074 41196 24080
rect 40316 24064 40368 24070
rect 40316 24006 40368 24012
rect 40040 23860 40092 23866
rect 40040 23802 40092 23808
rect 40132 23860 40184 23866
rect 40132 23802 40184 23808
rect 40222 23760 40278 23769
rect 39948 23724 40000 23730
rect 40222 23695 40278 23704
rect 40316 23724 40368 23730
rect 39948 23666 40000 23672
rect 39868 23582 40172 23610
rect 40236 23594 40264 23695
rect 40316 23666 40368 23672
rect 40038 23488 40094 23497
rect 40038 23423 40094 23432
rect 40052 23254 40080 23423
rect 40040 23248 40092 23254
rect 40040 23190 40092 23196
rect 40040 22432 40092 22438
rect 40040 22374 40092 22380
rect 40052 21962 40080 22374
rect 40040 21956 40092 21962
rect 40040 21898 40092 21904
rect 39948 21888 40000 21894
rect 39948 21830 40000 21836
rect 39960 21690 39988 21830
rect 39948 21684 40000 21690
rect 39948 21626 40000 21632
rect 40144 21146 40172 23582
rect 40224 23588 40276 23594
rect 40224 23530 40276 23536
rect 40224 23044 40276 23050
rect 40224 22986 40276 22992
rect 40236 22234 40264 22986
rect 40224 22228 40276 22234
rect 40224 22170 40276 22176
rect 40328 22094 40356 23666
rect 40592 23656 40644 23662
rect 40776 23656 40828 23662
rect 40644 23604 40776 23610
rect 40592 23598 40828 23604
rect 40604 23582 40816 23598
rect 40684 23520 40736 23526
rect 40684 23462 40736 23468
rect 40592 22704 40644 22710
rect 40592 22646 40644 22652
rect 40604 22094 40632 22646
rect 40696 22642 40724 23462
rect 40684 22636 40736 22642
rect 40684 22578 40736 22584
rect 40236 22066 40356 22094
rect 40512 22066 40632 22094
rect 40236 21298 40264 22066
rect 40314 21720 40370 21729
rect 40314 21655 40370 21664
rect 40328 21486 40356 21655
rect 40316 21480 40368 21486
rect 40316 21422 40368 21428
rect 40236 21270 40356 21298
rect 40222 21176 40278 21185
rect 40132 21140 40184 21146
rect 40222 21111 40278 21120
rect 40132 21082 40184 21088
rect 40236 21078 40264 21111
rect 40224 21072 40276 21078
rect 40224 21014 40276 21020
rect 39580 21004 39632 21010
rect 39580 20946 39632 20952
rect 39764 21004 39816 21010
rect 39764 20946 39816 20952
rect 39592 20466 39620 20946
rect 39580 20460 39632 20466
rect 39632 20420 39712 20448
rect 39580 20402 39632 20408
rect 39394 20088 39450 20097
rect 39394 20023 39450 20032
rect 39212 19916 39264 19922
rect 39212 19858 39264 19864
rect 39396 19916 39448 19922
rect 39396 19858 39448 19864
rect 38476 19508 38528 19514
rect 38476 19450 38528 19456
rect 38488 18952 38516 19450
rect 39408 19446 39436 19858
rect 39396 19440 39448 19446
rect 39396 19382 39448 19388
rect 39408 18970 39436 19382
rect 39684 19378 39712 20420
rect 40132 20392 40184 20398
rect 40132 20334 40184 20340
rect 40040 19780 40092 19786
rect 40040 19722 40092 19728
rect 40052 19514 40080 19722
rect 40040 19508 40092 19514
rect 40040 19450 40092 19456
rect 39672 19372 39724 19378
rect 39672 19314 39724 19320
rect 40038 19272 40094 19281
rect 40038 19207 40094 19216
rect 39396 18964 39448 18970
rect 38488 18924 38792 18952
rect 38568 18828 38620 18834
rect 38568 18770 38620 18776
rect 38476 18624 38528 18630
rect 38476 18566 38528 18572
rect 38488 17882 38516 18566
rect 38476 17876 38528 17882
rect 38476 17818 38528 17824
rect 38580 16454 38608 18770
rect 38764 18358 38792 18924
rect 39396 18906 39448 18912
rect 40052 18737 40080 19207
rect 40038 18728 40094 18737
rect 39764 18692 39816 18698
rect 40038 18663 40094 18672
rect 39764 18634 39816 18640
rect 38752 18352 38804 18358
rect 38752 18294 38804 18300
rect 39776 18290 39804 18634
rect 40144 18630 40172 20334
rect 40328 19310 40356 21270
rect 40512 21146 40540 22066
rect 40696 21672 40724 22578
rect 41052 22228 41104 22234
rect 41052 22170 41104 22176
rect 40868 21888 40920 21894
rect 40868 21830 40920 21836
rect 40960 21888 41012 21894
rect 40960 21830 41012 21836
rect 40604 21644 40724 21672
rect 40500 21140 40552 21146
rect 40500 21082 40552 21088
rect 40406 20904 40462 20913
rect 40406 20839 40462 20848
rect 40420 20602 40448 20839
rect 40408 20596 40460 20602
rect 40408 20538 40460 20544
rect 40420 19514 40448 20538
rect 40408 19508 40460 19514
rect 40408 19450 40460 19456
rect 40316 19304 40368 19310
rect 40316 19246 40368 19252
rect 40132 18624 40184 18630
rect 40132 18566 40184 18572
rect 40224 18624 40276 18630
rect 40224 18566 40276 18572
rect 40040 18352 40092 18358
rect 40040 18294 40092 18300
rect 39764 18284 39816 18290
rect 39764 18226 39816 18232
rect 40052 17542 40080 18294
rect 38936 17536 38988 17542
rect 38936 17478 38988 17484
rect 40040 17536 40092 17542
rect 40040 17478 40092 17484
rect 38948 17202 38976 17478
rect 40052 17354 40080 17478
rect 39960 17326 40080 17354
rect 39960 17270 39988 17326
rect 40144 17270 40172 18566
rect 40236 18086 40264 18566
rect 40512 18329 40540 21082
rect 40604 20534 40632 21644
rect 40880 21622 40908 21830
rect 40868 21616 40920 21622
rect 40868 21558 40920 21564
rect 40684 21548 40736 21554
rect 40684 21490 40736 21496
rect 40696 21457 40724 21490
rect 40682 21448 40738 21457
rect 40682 21383 40738 21392
rect 40868 21344 40920 21350
rect 40866 21312 40868 21321
rect 40920 21312 40922 21321
rect 40866 21247 40922 21256
rect 40684 21004 40736 21010
rect 40684 20946 40736 20952
rect 40696 20806 40724 20946
rect 40684 20800 40736 20806
rect 40684 20742 40736 20748
rect 40592 20528 40644 20534
rect 40592 20470 40644 20476
rect 40684 20256 40736 20262
rect 40684 20198 40736 20204
rect 40498 18320 40554 18329
rect 40498 18255 40554 18264
rect 40224 18080 40276 18086
rect 40224 18022 40276 18028
rect 40222 17912 40278 17921
rect 40222 17847 40278 17856
rect 39948 17264 40000 17270
rect 39948 17206 40000 17212
rect 40132 17264 40184 17270
rect 40132 17206 40184 17212
rect 38936 17196 38988 17202
rect 38936 17138 38988 17144
rect 38752 16992 38804 16998
rect 38752 16934 38804 16940
rect 38844 16992 38896 16998
rect 38844 16934 38896 16940
rect 38764 16522 38792 16934
rect 38856 16658 38884 16934
rect 38844 16652 38896 16658
rect 38844 16594 38896 16600
rect 38752 16516 38804 16522
rect 38752 16458 38804 16464
rect 38568 16448 38620 16454
rect 38568 16390 38620 16396
rect 38580 16182 38608 16390
rect 38568 16176 38620 16182
rect 38568 16118 38620 16124
rect 38568 15904 38620 15910
rect 38568 15846 38620 15852
rect 38382 15328 38438 15337
rect 37950 15260 38258 15269
rect 38382 15263 38438 15272
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 37740 15088 37792 15094
rect 37740 15030 37792 15036
rect 38580 14618 38608 15846
rect 38764 15434 38792 16458
rect 38752 15428 38804 15434
rect 38752 15370 38804 15376
rect 38764 15094 38792 15370
rect 38752 15088 38804 15094
rect 38752 15030 38804 15036
rect 38764 14940 38792 15030
rect 38672 14912 38792 14940
rect 38568 14612 38620 14618
rect 38568 14554 38620 14560
rect 37556 14272 37608 14278
rect 37556 14214 37608 14220
rect 37648 14272 37700 14278
rect 37648 14214 37700 14220
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 38672 14006 38700 14912
rect 38752 14816 38804 14822
rect 38752 14758 38804 14764
rect 38660 14000 38712 14006
rect 38660 13942 38712 13948
rect 38200 13796 38252 13802
rect 38200 13738 38252 13744
rect 38212 13530 38240 13738
rect 38672 13530 38700 13942
rect 38200 13524 38252 13530
rect 38200 13466 38252 13472
rect 38660 13524 38712 13530
rect 38660 13466 38712 13472
rect 38212 13274 38240 13466
rect 38212 13246 38332 13274
rect 37464 13184 37516 13190
rect 37464 13126 37516 13132
rect 37648 13184 37700 13190
rect 37648 13126 37700 13132
rect 37188 12912 37240 12918
rect 37188 12854 37240 12860
rect 37476 12850 37504 13126
rect 37660 12918 37688 13126
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 37648 12912 37700 12918
rect 37648 12854 37700 12860
rect 37464 12844 37516 12850
rect 37464 12786 37516 12792
rect 37280 12708 37332 12714
rect 37280 12650 37332 12656
rect 37096 12232 37148 12238
rect 37096 12174 37148 12180
rect 37292 11830 37320 12650
rect 37372 12096 37424 12102
rect 37372 12038 37424 12044
rect 37280 11824 37332 11830
rect 37280 11766 37332 11772
rect 37384 10742 37412 12038
rect 37476 11218 37504 12786
rect 38304 12782 38332 13246
rect 38292 12776 38344 12782
rect 38292 12718 38344 12724
rect 38764 12306 38792 14758
rect 38844 13524 38896 13530
rect 38844 13466 38896 13472
rect 38856 13258 38884 13466
rect 38844 13252 38896 13258
rect 38844 13194 38896 13200
rect 38856 12850 38884 13194
rect 38844 12844 38896 12850
rect 38844 12786 38896 12792
rect 38384 12300 38436 12306
rect 38384 12242 38436 12248
rect 38752 12300 38804 12306
rect 38752 12242 38804 12248
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 38396 11762 38424 12242
rect 38856 12170 38884 12786
rect 38844 12164 38896 12170
rect 38844 12106 38896 12112
rect 38660 12096 38712 12102
rect 38660 12038 38712 12044
rect 38672 11898 38700 12038
rect 38660 11892 38712 11898
rect 38660 11834 38712 11840
rect 38384 11756 38436 11762
rect 38384 11698 38436 11704
rect 38016 11620 38068 11626
rect 38016 11562 38068 11568
rect 37464 11212 37516 11218
rect 37464 11154 37516 11160
rect 38028 11121 38056 11562
rect 38014 11112 38070 11121
rect 38396 11082 38424 11698
rect 38856 11354 38884 12106
rect 38844 11348 38896 11354
rect 38844 11290 38896 11296
rect 38014 11047 38070 11056
rect 38384 11076 38436 11082
rect 38384 11018 38436 11024
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 38856 10810 38884 11290
rect 38948 11014 38976 17138
rect 39488 16584 39540 16590
rect 39488 16526 39540 16532
rect 39762 16552 39818 16561
rect 39212 16040 39264 16046
rect 39212 15982 39264 15988
rect 39224 15434 39252 15982
rect 39500 15570 39528 16526
rect 39960 16522 39988 17206
rect 40236 16794 40264 17847
rect 40696 17746 40724 20198
rect 40972 19990 41000 21830
rect 41064 21690 41092 22170
rect 41052 21684 41104 21690
rect 41052 21626 41104 21632
rect 41052 21072 41104 21078
rect 41052 21014 41104 21020
rect 41064 20058 41092 21014
rect 41156 20788 41184 24074
rect 41510 23352 41566 23361
rect 41510 23287 41566 23296
rect 41524 23050 41552 23287
rect 41512 23044 41564 23050
rect 41512 22986 41564 22992
rect 41236 22976 41288 22982
rect 41236 22918 41288 22924
rect 41248 22522 41276 22918
rect 41418 22808 41474 22817
rect 41418 22743 41474 22752
rect 41432 22642 41460 22743
rect 42076 22642 42104 24754
rect 42248 24404 42300 24410
rect 42248 24346 42300 24352
rect 42616 24404 42668 24410
rect 42616 24346 42668 24352
rect 42260 23866 42288 24346
rect 42524 24336 42576 24342
rect 42524 24278 42576 24284
rect 42248 23860 42300 23866
rect 42248 23802 42300 23808
rect 41420 22636 41472 22642
rect 41420 22578 41472 22584
rect 42064 22636 42116 22642
rect 42064 22578 42116 22584
rect 41248 22494 41368 22522
rect 41236 22432 41288 22438
rect 41236 22374 41288 22380
rect 41248 21049 41276 22374
rect 41340 21894 41368 22494
rect 41328 21888 41380 21894
rect 41328 21830 41380 21836
rect 41328 21344 41380 21350
rect 41328 21286 41380 21292
rect 41340 21146 41368 21286
rect 41432 21146 41460 22578
rect 41878 22536 41934 22545
rect 41878 22471 41880 22480
rect 41932 22471 41934 22480
rect 41880 22442 41932 22448
rect 41788 21888 41840 21894
rect 41788 21830 41840 21836
rect 41880 21888 41932 21894
rect 41880 21830 41932 21836
rect 41512 21480 41564 21486
rect 41512 21422 41564 21428
rect 41604 21480 41656 21486
rect 41604 21422 41656 21428
rect 41328 21140 41380 21146
rect 41328 21082 41380 21088
rect 41420 21140 41472 21146
rect 41420 21082 41472 21088
rect 41234 21040 41290 21049
rect 41234 20975 41290 20984
rect 41328 20800 41380 20806
rect 41156 20760 41328 20788
rect 41328 20742 41380 20748
rect 41052 20052 41104 20058
rect 41052 19994 41104 20000
rect 40960 19984 41012 19990
rect 40960 19926 41012 19932
rect 40868 19848 40920 19854
rect 40868 19790 40920 19796
rect 40776 19712 40828 19718
rect 40776 19654 40828 19660
rect 40788 18426 40816 19654
rect 40880 19242 40908 19790
rect 41064 19786 41092 19994
rect 41052 19780 41104 19786
rect 41052 19722 41104 19728
rect 41234 19272 41290 19281
rect 40868 19236 40920 19242
rect 41234 19207 41290 19216
rect 40868 19178 40920 19184
rect 41052 19168 41104 19174
rect 41052 19110 41104 19116
rect 41064 18698 41092 19110
rect 41052 18692 41104 18698
rect 41052 18634 41104 18640
rect 40776 18420 40828 18426
rect 40776 18362 40828 18368
rect 41064 18358 41092 18634
rect 41052 18352 41104 18358
rect 41052 18294 41104 18300
rect 41064 17864 41092 18294
rect 40972 17836 41092 17864
rect 40868 17808 40920 17814
rect 40868 17750 40920 17756
rect 40684 17740 40736 17746
rect 40684 17682 40736 17688
rect 40684 17128 40736 17134
rect 40684 17070 40736 17076
rect 40224 16788 40276 16794
rect 40224 16730 40276 16736
rect 40236 16522 40264 16730
rect 40316 16652 40368 16658
rect 40316 16594 40368 16600
rect 39762 16487 39818 16496
rect 39948 16516 40000 16522
rect 39488 15564 39540 15570
rect 39488 15506 39540 15512
rect 39212 15428 39264 15434
rect 39212 15370 39264 15376
rect 39224 13394 39252 15370
rect 39670 14920 39726 14929
rect 39776 14890 39804 16487
rect 39948 16458 40000 16464
rect 40224 16516 40276 16522
rect 40224 16458 40276 16464
rect 39960 16182 39988 16458
rect 39948 16176 40000 16182
rect 39948 16118 40000 16124
rect 39960 15434 39988 16118
rect 40328 15910 40356 16594
rect 40696 16590 40724 17070
rect 40684 16584 40736 16590
rect 40684 16526 40736 16532
rect 40316 15904 40368 15910
rect 40316 15846 40368 15852
rect 40328 15570 40356 15846
rect 40316 15564 40368 15570
rect 40316 15506 40368 15512
rect 39948 15428 40000 15434
rect 39948 15370 40000 15376
rect 39670 14855 39672 14864
rect 39724 14855 39726 14864
rect 39764 14884 39816 14890
rect 39672 14826 39724 14832
rect 39764 14826 39816 14832
rect 39960 14618 39988 15370
rect 40130 15328 40186 15337
rect 40130 15263 40186 15272
rect 40144 15162 40172 15263
rect 40132 15156 40184 15162
rect 40132 15098 40184 15104
rect 40880 15026 40908 17750
rect 40972 17270 41000 17836
rect 41052 17740 41104 17746
rect 41052 17682 41104 17688
rect 40960 17264 41012 17270
rect 40960 17206 41012 17212
rect 40972 16794 41000 17206
rect 41064 17066 41092 17682
rect 41052 17060 41104 17066
rect 41052 17002 41104 17008
rect 40960 16788 41012 16794
rect 40960 16730 41012 16736
rect 41248 16726 41276 19207
rect 41340 18193 41368 20742
rect 41524 19417 41552 21422
rect 41616 20942 41644 21422
rect 41800 21418 41828 21830
rect 41892 21729 41920 21830
rect 41878 21720 41934 21729
rect 42076 21690 42104 22578
rect 42432 22024 42484 22030
rect 42432 21966 42484 21972
rect 41878 21655 41934 21664
rect 42064 21684 42116 21690
rect 42064 21626 42116 21632
rect 41788 21412 41840 21418
rect 41788 21354 41840 21360
rect 42444 21010 42472 21966
rect 42536 21622 42564 24278
rect 42628 24070 42656 24346
rect 42720 24290 42748 26302
rect 42798 26200 42854 27000
rect 43442 26200 43498 27000
rect 44086 26200 44142 27000
rect 44730 26200 44786 27000
rect 45374 26200 45430 27000
rect 46018 26330 46074 27000
rect 46662 26330 46718 27000
rect 46018 26302 46336 26330
rect 46018 26200 46074 26302
rect 43902 24712 43958 24721
rect 43902 24647 43958 24656
rect 43996 24676 44048 24682
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 43916 24410 43944 24647
rect 43996 24618 44048 24624
rect 43904 24404 43956 24410
rect 43904 24346 43956 24352
rect 42720 24262 42840 24290
rect 42812 24206 42840 24262
rect 42800 24200 42852 24206
rect 42800 24142 42852 24148
rect 43812 24200 43864 24206
rect 43812 24142 43864 24148
rect 43904 24200 43956 24206
rect 43904 24142 43956 24148
rect 42616 24064 42668 24070
rect 42616 24006 42668 24012
rect 42708 24064 42760 24070
rect 42708 24006 42760 24012
rect 42720 23798 42748 24006
rect 42708 23792 42760 23798
rect 42708 23734 42760 23740
rect 42720 23594 42748 23734
rect 42800 23724 42852 23730
rect 42800 23666 42852 23672
rect 42708 23588 42760 23594
rect 42708 23530 42760 23536
rect 42812 23474 42840 23666
rect 42720 23446 42840 23474
rect 43536 23520 43588 23526
rect 43536 23462 43588 23468
rect 42720 23050 42748 23446
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 42800 23316 42852 23322
rect 42800 23258 42852 23264
rect 42708 23044 42760 23050
rect 42708 22986 42760 22992
rect 42616 22568 42668 22574
rect 42616 22510 42668 22516
rect 42628 22409 42656 22510
rect 42614 22400 42670 22409
rect 42614 22335 42670 22344
rect 42524 21616 42576 21622
rect 42524 21558 42576 21564
rect 42628 21146 42656 22335
rect 42720 22234 42748 22986
rect 42708 22228 42760 22234
rect 42708 22170 42760 22176
rect 42812 22094 42840 23258
rect 43350 23216 43406 23225
rect 43350 23151 43406 23160
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 42720 22066 42840 22094
rect 42892 22092 42944 22098
rect 42720 21962 42748 22066
rect 42892 22034 42944 22040
rect 42800 22024 42852 22030
rect 42798 21992 42800 22001
rect 42852 21992 42854 22001
rect 42708 21956 42760 21962
rect 42798 21927 42854 21936
rect 42708 21898 42760 21904
rect 42720 21622 42748 21898
rect 42812 21622 42840 21927
rect 42708 21616 42760 21622
rect 42708 21558 42760 21564
rect 42800 21616 42852 21622
rect 42800 21558 42852 21564
rect 42904 21332 42932 22034
rect 43260 22024 43312 22030
rect 43260 21966 43312 21972
rect 43272 21554 43300 21966
rect 43260 21548 43312 21554
rect 43260 21490 43312 21496
rect 42812 21304 42932 21332
rect 42616 21140 42668 21146
rect 42616 21082 42668 21088
rect 42432 21004 42484 21010
rect 42432 20946 42484 20952
rect 41604 20936 41656 20942
rect 41604 20878 41656 20884
rect 41510 19408 41566 19417
rect 41510 19343 41566 19352
rect 42064 19168 42116 19174
rect 42812 19145 42840 21304
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 43364 21010 43392 23151
rect 43548 23050 43576 23462
rect 43720 23248 43772 23254
rect 43720 23190 43772 23196
rect 43536 23044 43588 23050
rect 43536 22986 43588 22992
rect 43628 23044 43680 23050
rect 43628 22986 43680 22992
rect 43444 22568 43496 22574
rect 43444 22510 43496 22516
rect 43352 21004 43404 21010
rect 43352 20946 43404 20952
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 42064 19110 42116 19116
rect 42798 19136 42854 19145
rect 42076 18970 42104 19110
rect 42798 19071 42854 19080
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 42064 18964 42116 18970
rect 42064 18906 42116 18912
rect 41326 18184 41382 18193
rect 41326 18119 41382 18128
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 43456 17814 43484 22510
rect 43536 22228 43588 22234
rect 43536 22170 43588 22176
rect 43548 21690 43576 22170
rect 43536 21684 43588 21690
rect 43536 21626 43588 21632
rect 43536 21344 43588 21350
rect 43640 21332 43668 22986
rect 43732 22166 43760 23190
rect 43720 22160 43772 22166
rect 43720 22102 43772 22108
rect 43824 22098 43852 24142
rect 43916 23225 43944 24142
rect 43902 23216 43958 23225
rect 43902 23151 43958 23160
rect 44008 22642 44036 24618
rect 44100 23118 44128 26200
rect 44456 24200 44508 24206
rect 44456 24142 44508 24148
rect 44272 24132 44324 24138
rect 44272 24074 44324 24080
rect 44088 23112 44140 23118
rect 44088 23054 44140 23060
rect 43996 22636 44048 22642
rect 43996 22578 44048 22584
rect 43904 22432 43956 22438
rect 43904 22374 43956 22380
rect 43812 22092 43864 22098
rect 43812 22034 43864 22040
rect 43916 21593 43944 22374
rect 44008 21690 44036 22578
rect 44100 22234 44128 23054
rect 44088 22228 44140 22234
rect 44088 22170 44140 22176
rect 44284 22166 44312 24074
rect 44272 22160 44324 22166
rect 44468 22137 44496 24142
rect 44744 24138 44772 26200
rect 45284 24880 45336 24886
rect 45284 24822 45336 24828
rect 45190 24304 45246 24313
rect 45190 24239 45246 24248
rect 44732 24132 44784 24138
rect 44732 24074 44784 24080
rect 44824 23724 44876 23730
rect 44824 23666 44876 23672
rect 44836 23322 44864 23666
rect 44824 23316 44876 23322
rect 44824 23258 44876 23264
rect 44730 22672 44786 22681
rect 44730 22607 44732 22616
rect 44784 22607 44786 22616
rect 44732 22578 44784 22584
rect 44548 22432 44600 22438
rect 44548 22374 44600 22380
rect 44272 22102 44324 22108
rect 44454 22128 44510 22137
rect 44454 22063 44510 22072
rect 43996 21684 44048 21690
rect 43996 21626 44048 21632
rect 43902 21584 43958 21593
rect 43902 21519 43958 21528
rect 43588 21304 43668 21332
rect 43536 21286 43588 21292
rect 44560 19825 44588 22374
rect 44744 22098 44772 22578
rect 45204 22506 45232 24239
rect 45296 22642 45324 24822
rect 45388 24426 45416 26200
rect 45388 24398 45600 24426
rect 45376 24268 45428 24274
rect 45376 24210 45428 24216
rect 45388 23118 45416 24210
rect 45572 24206 45600 24398
rect 46308 24206 46336 26302
rect 46662 26302 46888 26330
rect 46662 26200 46718 26302
rect 46754 25120 46810 25129
rect 46754 25055 46810 25064
rect 45560 24200 45612 24206
rect 45560 24142 45612 24148
rect 46204 24200 46256 24206
rect 46204 24142 46256 24148
rect 46296 24200 46348 24206
rect 46296 24142 46348 24148
rect 46020 24064 46072 24070
rect 46020 24006 46072 24012
rect 46112 24064 46164 24070
rect 46112 24006 46164 24012
rect 45928 23724 45980 23730
rect 45928 23666 45980 23672
rect 45940 23594 45968 23666
rect 45928 23588 45980 23594
rect 45928 23530 45980 23536
rect 45376 23112 45428 23118
rect 45376 23054 45428 23060
rect 45284 22636 45336 22642
rect 45284 22578 45336 22584
rect 45192 22500 45244 22506
rect 45192 22442 45244 22448
rect 45376 22432 45428 22438
rect 45376 22374 45428 22380
rect 45388 22137 45416 22374
rect 45374 22128 45430 22137
rect 44732 22092 44784 22098
rect 45374 22063 45430 22072
rect 44732 22034 44784 22040
rect 44546 19816 44602 19825
rect 44546 19751 44602 19760
rect 43444 17808 43496 17814
rect 43444 17750 43496 17756
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 46032 16794 46060 24006
rect 46124 23254 46152 24006
rect 46216 23866 46244 24142
rect 46204 23860 46256 23866
rect 46204 23802 46256 23808
rect 46662 23760 46718 23769
rect 46662 23695 46718 23704
rect 46204 23520 46256 23526
rect 46204 23462 46256 23468
rect 46112 23248 46164 23254
rect 46112 23190 46164 23196
rect 46112 22976 46164 22982
rect 46112 22918 46164 22924
rect 46124 22710 46152 22918
rect 46112 22704 46164 22710
rect 46112 22646 46164 22652
rect 46216 21690 46244 23462
rect 46676 23322 46704 23695
rect 46664 23316 46716 23322
rect 46664 23258 46716 23264
rect 46676 23118 46704 23258
rect 46664 23112 46716 23118
rect 46664 23054 46716 23060
rect 46768 22710 46796 25055
rect 46860 24120 46888 26302
rect 47306 26200 47362 27000
rect 47950 26200 48006 27000
rect 48594 26200 48650 27000
rect 49238 26200 49294 27000
rect 46860 24092 46980 24120
rect 46952 23798 46980 24092
rect 46940 23792 46992 23798
rect 46940 23734 46992 23740
rect 47320 23662 47348 26200
rect 47582 24712 47638 24721
rect 47582 24647 47638 24656
rect 47492 24268 47544 24274
rect 47492 24210 47544 24216
rect 47400 24132 47452 24138
rect 47400 24074 47452 24080
rect 47412 23730 47440 24074
rect 47400 23724 47452 23730
rect 47400 23666 47452 23672
rect 47308 23656 47360 23662
rect 47308 23598 47360 23604
rect 46940 23588 46992 23594
rect 46940 23530 46992 23536
rect 47124 23588 47176 23594
rect 47124 23530 47176 23536
rect 46846 23488 46902 23497
rect 46846 23423 46902 23432
rect 46756 22704 46808 22710
rect 46756 22646 46808 22652
rect 46204 21684 46256 21690
rect 46204 21626 46256 21632
rect 46216 20806 46244 21626
rect 46860 21554 46888 23423
rect 46952 23322 46980 23530
rect 46940 23316 46992 23322
rect 46940 23258 46992 23264
rect 47136 23118 47164 23530
rect 47320 23118 47348 23598
rect 47124 23112 47176 23118
rect 47124 23054 47176 23060
rect 47308 23112 47360 23118
rect 47308 23054 47360 23060
rect 47504 22982 47532 24210
rect 47032 22976 47084 22982
rect 46938 22944 46994 22953
rect 47032 22918 47084 22924
rect 47492 22976 47544 22982
rect 47492 22918 47544 22924
rect 46938 22879 46994 22888
rect 46952 22438 46980 22879
rect 46940 22432 46992 22438
rect 46940 22374 46992 22380
rect 47044 22234 47072 22918
rect 47596 22506 47624 24647
rect 47766 24304 47822 24313
rect 47766 24239 47822 24248
rect 47676 22976 47728 22982
rect 47676 22918 47728 22924
rect 47584 22500 47636 22506
rect 47584 22442 47636 22448
rect 47032 22228 47084 22234
rect 47032 22170 47084 22176
rect 47596 22030 47624 22442
rect 47584 22024 47636 22030
rect 47584 21966 47636 21972
rect 46848 21548 46900 21554
rect 46848 21490 46900 21496
rect 46860 21146 46888 21490
rect 46848 21140 46900 21146
rect 46848 21082 46900 21088
rect 47688 20913 47716 22918
rect 47780 22642 47808 24239
rect 47964 24188 47992 26200
rect 48226 25528 48282 25537
rect 48226 25463 48282 25472
rect 48240 24274 48268 25463
rect 48228 24268 48280 24274
rect 48228 24210 48280 24216
rect 48044 24200 48096 24206
rect 47872 24160 48044 24188
rect 47872 23866 47900 24160
rect 48044 24142 48096 24148
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 47860 23860 47912 23866
rect 47860 23802 47912 23808
rect 48412 22976 48464 22982
rect 48412 22918 48464 22924
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 47768 22636 47820 22642
rect 47768 22578 47820 22584
rect 48320 22432 48372 22438
rect 48320 22374 48372 22380
rect 47860 21888 47912 21894
rect 47860 21830 47912 21836
rect 47872 21690 47900 21830
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 47860 21684 47912 21690
rect 47860 21626 47912 21632
rect 47674 20904 47730 20913
rect 47674 20839 47730 20848
rect 46204 20800 46256 20806
rect 46204 20742 46256 20748
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 48332 19961 48360 22374
rect 48424 20369 48452 22918
rect 48608 22094 48636 26200
rect 48780 24200 48832 24206
rect 48778 24168 48780 24177
rect 48832 24168 48834 24177
rect 48778 24103 48834 24112
rect 49252 23730 49280 26200
rect 49240 23724 49292 23730
rect 49240 23666 49292 23672
rect 48688 23112 48740 23118
rect 48686 23080 48688 23089
rect 48740 23080 48742 23089
rect 48686 23015 48742 23024
rect 48700 22778 48728 23015
rect 48688 22772 48740 22778
rect 48688 22714 48740 22720
rect 49252 22506 49280 23666
rect 49424 23112 49476 23118
rect 49424 23054 49476 23060
rect 49436 22681 49464 23054
rect 49422 22672 49478 22681
rect 49332 22636 49384 22642
rect 49422 22607 49478 22616
rect 49332 22578 49384 22584
rect 49240 22500 49292 22506
rect 49240 22442 49292 22448
rect 48688 22432 48740 22438
rect 48688 22374 48740 22380
rect 48516 22066 48636 22094
rect 48516 22030 48544 22066
rect 48504 22024 48556 22030
rect 48504 21966 48556 21972
rect 48594 21856 48650 21865
rect 48594 21791 48650 21800
rect 48608 21554 48636 21791
rect 48596 21548 48648 21554
rect 48596 21490 48648 21496
rect 48608 21146 48636 21490
rect 48596 21140 48648 21146
rect 48596 21082 48648 21088
rect 48410 20360 48466 20369
rect 48410 20295 48466 20304
rect 48412 20256 48464 20262
rect 48412 20198 48464 20204
rect 48318 19952 48374 19961
rect 48318 19887 48374 19896
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 48424 19446 48452 20198
rect 48412 19440 48464 19446
rect 48412 19382 48464 19388
rect 48700 18873 48728 22374
rect 49344 22273 49372 22578
rect 49330 22264 49386 22273
rect 49436 22234 49464 22607
rect 49330 22199 49386 22208
rect 49424 22228 49476 22234
rect 49424 22170 49476 22176
rect 49056 21956 49108 21962
rect 49056 21898 49108 21904
rect 49240 21956 49292 21962
rect 49240 21898 49292 21904
rect 49068 20505 49096 21898
rect 49252 21457 49280 21898
rect 49332 21548 49384 21554
rect 49332 21490 49384 21496
rect 49238 21448 49294 21457
rect 49238 21383 49294 21392
rect 49148 21344 49200 21350
rect 49148 21286 49200 21292
rect 49160 20602 49188 21286
rect 49344 21078 49372 21490
rect 49332 21072 49384 21078
rect 49330 21040 49332 21049
rect 49384 21040 49386 21049
rect 49330 20975 49386 20984
rect 49332 20936 49384 20942
rect 49332 20878 49384 20884
rect 49344 20641 49372 20878
rect 49424 20868 49476 20874
rect 49424 20810 49476 20816
rect 49330 20632 49386 20641
rect 49148 20596 49200 20602
rect 49330 20567 49386 20576
rect 49148 20538 49200 20544
rect 49054 20496 49110 20505
rect 48780 20460 48832 20466
rect 49436 20466 49464 20810
rect 49054 20431 49110 20440
rect 49424 20460 49476 20466
rect 48780 20402 48832 20408
rect 49424 20402 49476 20408
rect 48792 20233 48820 20402
rect 48778 20224 48834 20233
rect 48778 20159 48834 20168
rect 48792 20058 48820 20159
rect 48780 20052 48832 20058
rect 48780 19994 48832 20000
rect 49436 19825 49464 20402
rect 49422 19816 49478 19825
rect 49332 19780 49384 19786
rect 49422 19751 49478 19760
rect 49332 19722 49384 19728
rect 49148 19712 49200 19718
rect 49148 19654 49200 19660
rect 49160 19281 49188 19654
rect 49344 19417 49372 19722
rect 49330 19408 49386 19417
rect 49240 19372 49292 19378
rect 49330 19343 49386 19352
rect 49240 19314 49292 19320
rect 49146 19272 49202 19281
rect 49146 19207 49202 19216
rect 49252 19009 49280 19314
rect 49424 19168 49476 19174
rect 49424 19110 49476 19116
rect 49238 19000 49294 19009
rect 49238 18935 49294 18944
rect 48686 18864 48742 18873
rect 48686 18799 48742 18808
rect 49436 18766 49464 19110
rect 48780 18760 48832 18766
rect 48780 18702 48832 18708
rect 49424 18760 49476 18766
rect 49424 18702 49476 18708
rect 48412 18624 48464 18630
rect 48412 18566 48464 18572
rect 48504 18624 48556 18630
rect 48792 18601 48820 18702
rect 48504 18566 48556 18572
rect 48778 18592 48834 18601
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 48424 18290 48452 18566
rect 48412 18284 48464 18290
rect 48412 18226 48464 18232
rect 48320 18080 48372 18086
rect 48320 18022 48372 18028
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 48332 17338 48360 18022
rect 48412 17604 48464 17610
rect 48412 17546 48464 17552
rect 48424 17338 48452 17546
rect 48320 17332 48372 17338
rect 48320 17274 48372 17280
rect 48412 17332 48464 17338
rect 48412 17274 48464 17280
rect 48228 17264 48280 17270
rect 48516 17241 48544 18566
rect 48778 18527 48834 18536
rect 48792 18426 48820 18527
rect 48780 18420 48832 18426
rect 48780 18362 48832 18368
rect 49332 18284 49384 18290
rect 49332 18226 49384 18232
rect 49344 17785 49372 18226
rect 49436 18193 49464 18702
rect 49422 18184 49478 18193
rect 49422 18119 49478 18128
rect 49330 17776 49386 17785
rect 49330 17711 49386 17720
rect 49332 17672 49384 17678
rect 49332 17614 49384 17620
rect 48688 17536 48740 17542
rect 48688 17478 48740 17484
rect 49148 17536 49200 17542
rect 49148 17478 49200 17484
rect 48700 17270 48728 17478
rect 48688 17264 48740 17270
rect 48228 17206 48280 17212
rect 48502 17232 48558 17241
rect 41328 16788 41380 16794
rect 46020 16788 46072 16794
rect 41380 16748 41460 16776
rect 41328 16730 41380 16736
rect 41236 16720 41288 16726
rect 41236 16662 41288 16668
rect 41248 16522 41276 16662
rect 41236 16516 41288 16522
rect 41236 16458 41288 16464
rect 40960 16448 41012 16454
rect 40960 16390 41012 16396
rect 40972 16250 41000 16390
rect 41432 16250 41460 16748
rect 46020 16730 46072 16736
rect 48240 16561 48268 17206
rect 48688 17206 48740 17212
rect 48502 17167 48558 17176
rect 48780 17196 48832 17202
rect 48780 17138 48832 17144
rect 48792 16969 48820 17138
rect 49056 17128 49108 17134
rect 49054 17096 49056 17105
rect 49108 17096 49110 17105
rect 49054 17031 49110 17040
rect 48778 16960 48834 16969
rect 48778 16895 48834 16904
rect 48792 16794 48820 16895
rect 48780 16788 48832 16794
rect 48780 16730 48832 16736
rect 49160 16697 49188 17478
rect 49344 17377 49372 17614
rect 49330 17368 49386 17377
rect 49330 17303 49386 17312
rect 49146 16688 49202 16697
rect 49146 16623 49202 16632
rect 49424 16584 49476 16590
rect 48226 16552 48282 16561
rect 49424 16526 49476 16532
rect 48226 16487 48282 16496
rect 49148 16448 49200 16454
rect 49148 16390 49200 16396
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 40960 16244 41012 16250
rect 40960 16186 41012 16192
rect 41420 16244 41472 16250
rect 41420 16186 41472 16192
rect 41432 15706 41460 16186
rect 49160 16153 49188 16390
rect 49436 16153 49464 16526
rect 49146 16144 49202 16153
rect 48688 16108 48740 16114
rect 49422 16144 49478 16153
rect 49146 16079 49202 16088
rect 49332 16108 49384 16114
rect 48688 16050 48740 16056
rect 49422 16079 49478 16088
rect 49332 16050 49384 16056
rect 41788 16040 41840 16046
rect 41788 15982 41840 15988
rect 41420 15700 41472 15706
rect 41420 15642 41472 15648
rect 41800 15638 41828 15982
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 48700 15706 48728 16050
rect 49146 16008 49202 16017
rect 49146 15943 49148 15952
rect 49200 15943 49202 15952
rect 49148 15914 49200 15920
rect 49344 15745 49372 16050
rect 49330 15736 49386 15745
rect 48688 15700 48740 15706
rect 49330 15671 49386 15680
rect 48688 15642 48740 15648
rect 41788 15632 41840 15638
rect 41788 15574 41840 15580
rect 49332 15496 49384 15502
rect 49332 15438 49384 15444
rect 49344 15337 49372 15438
rect 49330 15328 49386 15337
rect 47950 15260 48258 15269
rect 49330 15263 49386 15272
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 48412 15088 48464 15094
rect 48412 15030 48464 15036
rect 49146 15056 49202 15065
rect 40868 15020 40920 15026
rect 40868 14962 40920 14968
rect 45652 14816 45704 14822
rect 45652 14758 45704 14764
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 39948 14612 40000 14618
rect 39948 14554 40000 14560
rect 39488 14272 39540 14278
rect 39488 14214 39540 14220
rect 39500 14006 39528 14214
rect 41328 14068 41380 14074
rect 41328 14010 41380 14016
rect 39488 14000 39540 14006
rect 39488 13942 39540 13948
rect 39212 13388 39264 13394
rect 39212 13330 39264 13336
rect 41340 13326 41368 14010
rect 45664 13938 45692 14758
rect 48320 14272 48372 14278
rect 48320 14214 48372 14220
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 47032 14068 47084 14074
rect 47032 14010 47084 14016
rect 45652 13932 45704 13938
rect 45652 13874 45704 13880
rect 46296 13864 46348 13870
rect 46296 13806 46348 13812
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 46308 13326 46336 13806
rect 41328 13320 41380 13326
rect 41328 13262 41380 13268
rect 46296 13320 46348 13326
rect 46296 13262 46348 13268
rect 39580 13184 39632 13190
rect 39580 13126 39632 13132
rect 45928 13184 45980 13190
rect 45928 13126 45980 13132
rect 39304 12776 39356 12782
rect 39304 12718 39356 12724
rect 39316 12646 39344 12718
rect 39304 12640 39356 12646
rect 39304 12582 39356 12588
rect 39316 12442 39344 12582
rect 39212 12436 39264 12442
rect 39212 12378 39264 12384
rect 39304 12436 39356 12442
rect 39304 12378 39356 12384
rect 39028 11756 39080 11762
rect 39028 11698 39080 11704
rect 38936 11008 38988 11014
rect 38936 10950 38988 10956
rect 38844 10804 38896 10810
rect 38844 10746 38896 10752
rect 37372 10736 37424 10742
rect 37372 10678 37424 10684
rect 38948 10062 38976 10950
rect 38936 10056 38988 10062
rect 38936 9998 38988 10004
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 38752 8424 38804 8430
rect 38752 8366 38804 8372
rect 38764 7886 38792 8366
rect 39040 8022 39068 11698
rect 39224 11694 39252 12378
rect 39212 11688 39264 11694
rect 39212 11630 39264 11636
rect 39592 11354 39620 13126
rect 40316 12980 40368 12986
rect 40316 12922 40368 12928
rect 40038 12880 40094 12889
rect 40038 12815 40040 12824
rect 40092 12815 40094 12824
rect 40040 12786 40092 12792
rect 40130 12200 40186 12209
rect 40130 12135 40132 12144
rect 40184 12135 40186 12144
rect 40132 12106 40184 12112
rect 40144 11898 40172 12106
rect 40132 11892 40184 11898
rect 40132 11834 40184 11840
rect 40224 11552 40276 11558
rect 40224 11494 40276 11500
rect 39580 11348 39632 11354
rect 39580 11290 39632 11296
rect 39592 11150 39620 11290
rect 40236 11150 40264 11494
rect 39580 11144 39632 11150
rect 39580 11086 39632 11092
rect 40224 11144 40276 11150
rect 40224 11086 40276 11092
rect 40040 8628 40092 8634
rect 40040 8570 40092 8576
rect 39028 8016 39080 8022
rect 39028 7958 39080 7964
rect 38752 7880 38804 7886
rect 38752 7822 38804 7828
rect 38660 7744 38712 7750
rect 38660 7686 38712 7692
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 38672 7478 38700 7686
rect 38660 7472 38712 7478
rect 38660 7414 38712 7420
rect 37280 7200 37332 7206
rect 37280 7142 37332 7148
rect 37924 7200 37976 7206
rect 37924 7142 37976 7148
rect 37292 5302 37320 7142
rect 37936 6934 37964 7142
rect 38476 6996 38528 7002
rect 38476 6938 38528 6944
rect 37924 6928 37976 6934
rect 37924 6870 37976 6876
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 37648 6112 37700 6118
rect 37648 6054 37700 6060
rect 37660 5914 37688 6054
rect 37648 5908 37700 5914
rect 37648 5850 37700 5856
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 38488 5302 38516 6938
rect 40052 6390 40080 8570
rect 40328 8566 40356 12922
rect 45940 12850 45968 13126
rect 47044 12850 47072 14010
rect 48332 13954 48360 14214
rect 48424 14074 48452 15030
rect 49146 14991 49202 15000
rect 49332 15020 49384 15026
rect 49056 14408 49108 14414
rect 49054 14376 49056 14385
rect 49108 14376 49110 14385
rect 49054 14311 49110 14320
rect 49160 14074 49188 14991
rect 49332 14962 49384 14968
rect 49344 14929 49372 14962
rect 49330 14920 49386 14929
rect 49330 14855 49386 14864
rect 49238 14512 49294 14521
rect 49238 14447 49294 14456
rect 49252 14414 49280 14447
rect 49240 14408 49292 14414
rect 49240 14350 49292 14356
rect 49238 14104 49294 14113
rect 48412 14068 48464 14074
rect 48412 14010 48464 14016
rect 49148 14068 49200 14074
rect 49238 14039 49294 14048
rect 49148 14010 49200 14016
rect 49252 14006 49280 14039
rect 48240 13938 48360 13954
rect 49240 14000 49292 14006
rect 49240 13942 49292 13948
rect 48228 13932 48360 13938
rect 48280 13926 48360 13932
rect 48228 13874 48280 13880
rect 48240 13705 48268 13874
rect 48226 13696 48282 13705
rect 48226 13631 48282 13640
rect 49148 13320 49200 13326
rect 49146 13288 49148 13297
rect 49200 13288 49202 13297
rect 49146 13223 49202 13232
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 49146 12880 49202 12889
rect 45928 12844 45980 12850
rect 45928 12786 45980 12792
rect 47032 12844 47084 12850
rect 49146 12815 49148 12824
rect 47032 12786 47084 12792
rect 49200 12815 49202 12824
rect 49148 12786 49200 12792
rect 42708 12708 42760 12714
rect 42708 12650 42760 12656
rect 40960 12096 41012 12102
rect 40960 12038 41012 12044
rect 40972 11830 41000 12038
rect 40960 11824 41012 11830
rect 40960 11766 41012 11772
rect 42720 11218 42748 12650
rect 47952 12640 48004 12646
rect 47952 12582 48004 12588
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 47124 12368 47176 12374
rect 47124 12310 47176 12316
rect 46112 12096 46164 12102
rect 46112 12038 46164 12044
rect 46124 11762 46152 12038
rect 46112 11756 46164 11762
rect 46112 11698 46164 11704
rect 46756 11620 46808 11626
rect 46756 11562 46808 11568
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 44088 11348 44140 11354
rect 44088 11290 44140 11296
rect 42708 11212 42760 11218
rect 42708 11154 42760 11160
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 44100 10062 44128 11290
rect 45744 11076 45796 11082
rect 45744 11018 45796 11024
rect 45756 10062 45784 11018
rect 46768 10062 46796 11562
rect 46940 11076 46992 11082
rect 46940 11018 46992 11024
rect 46952 10674 46980 11018
rect 46940 10668 46992 10674
rect 46940 10610 46992 10616
rect 46940 10532 46992 10538
rect 46940 10474 46992 10480
rect 44088 10056 44140 10062
rect 44088 9998 44140 10004
rect 45744 10056 45796 10062
rect 45744 9998 45796 10004
rect 46756 10056 46808 10062
rect 46756 9998 46808 10004
rect 42708 9988 42760 9994
rect 42708 9930 42760 9936
rect 46204 9988 46256 9994
rect 46204 9930 46256 9936
rect 42720 8634 42748 9930
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 43720 9172 43772 9178
rect 43720 9114 43772 9120
rect 42708 8628 42760 8634
rect 42708 8570 42760 8576
rect 40316 8560 40368 8566
rect 40316 8502 40368 8508
rect 40224 8424 40276 8430
rect 40224 8366 40276 8372
rect 40132 7812 40184 7818
rect 40132 7754 40184 7760
rect 40144 6798 40172 7754
rect 40132 6792 40184 6798
rect 40132 6734 40184 6740
rect 40040 6384 40092 6390
rect 40040 6326 40092 6332
rect 37280 5296 37332 5302
rect 37280 5238 37332 5244
rect 38476 5296 38528 5302
rect 38476 5238 38528 5244
rect 40040 5092 40092 5098
rect 40040 5034 40092 5040
rect 37832 5024 37884 5030
rect 37832 4966 37884 4972
rect 37844 4826 37872 4966
rect 37832 4820 37884 4826
rect 37832 4762 37884 4768
rect 37004 4752 37056 4758
rect 37004 4694 37056 4700
rect 37372 4480 37424 4486
rect 37372 4422 37424 4428
rect 39764 4480 39816 4486
rect 39764 4422 39816 4428
rect 37384 4282 37412 4422
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 37372 4276 37424 4282
rect 37372 4218 37424 4224
rect 39212 3528 39264 3534
rect 39212 3470 39264 3476
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 37740 3188 37792 3194
rect 37740 3130 37792 3136
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 34348 2746 34468 2774
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 32864 2644 32916 2650
rect 32864 2586 32916 2592
rect 34440 2582 34468 2746
rect 32772 2576 32824 2582
rect 32772 2518 32824 2524
rect 34428 2576 34480 2582
rect 34428 2518 34480 2524
rect 37752 2514 37780 3130
rect 38292 2916 38344 2922
rect 38292 2858 38344 2864
rect 37740 2508 37792 2514
rect 37740 2450 37792 2456
rect 38304 2446 38332 2858
rect 27160 2440 27212 2446
rect 29000 2440 29052 2446
rect 27160 2382 27212 2388
rect 28920 2388 29000 2394
rect 28920 2382 29052 2388
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 33140 2440 33192 2446
rect 33140 2382 33192 2388
rect 34980 2440 35032 2446
rect 34980 2382 35032 2388
rect 38292 2440 38344 2446
rect 38292 2382 38344 2388
rect 28920 2366 29040 2382
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 28644 870 28764 898
rect 28644 800 28672 870
rect 18156 734 18368 762
rect 20166 0 20222 800
rect 22282 0 22338 800
rect 24398 0 24454 800
rect 26514 0 26570 800
rect 28630 0 28686 800
rect 28736 762 28764 870
rect 28920 762 28948 2366
rect 30760 800 30788 2382
rect 33152 1578 33180 2382
rect 32876 1550 33180 1578
rect 32876 800 32904 1550
rect 34992 800 35020 2382
rect 37096 2304 37148 2310
rect 37096 2246 37148 2252
rect 37108 800 37136 2246
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 39224 800 39252 3470
rect 39776 3058 39804 4422
rect 40052 3602 40080 5034
rect 40236 4758 40264 8366
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 43732 5710 43760 9114
rect 44180 9036 44232 9042
rect 44180 8978 44232 8984
rect 44192 8566 44220 8978
rect 45468 8628 45520 8634
rect 45468 8570 45520 8576
rect 44180 8560 44232 8566
rect 44180 8502 44232 8508
rect 45480 8498 45508 8570
rect 46216 8498 46244 9930
rect 45468 8492 45520 8498
rect 45468 8434 45520 8440
rect 46204 8492 46256 8498
rect 46204 8434 46256 8440
rect 46848 8424 46900 8430
rect 46848 8366 46900 8372
rect 44916 8356 44968 8362
rect 44916 8298 44968 8304
rect 44928 7410 44956 8298
rect 46860 7993 46888 8366
rect 46846 7984 46902 7993
rect 46846 7919 46902 7928
rect 46952 7886 46980 10474
rect 47032 10124 47084 10130
rect 47032 10066 47084 10072
rect 46940 7880 46992 7886
rect 46940 7822 46992 7828
rect 47044 7410 47072 10066
rect 47136 9586 47164 12310
rect 47964 12238 47992 12582
rect 49146 12472 49202 12481
rect 49146 12407 49202 12416
rect 49160 12306 49188 12407
rect 49148 12300 49200 12306
rect 49148 12242 49200 12248
rect 47952 12232 48004 12238
rect 47952 12174 48004 12180
rect 49146 12064 49202 12073
rect 47950 11996 48258 12005
rect 49146 11999 49202 12008
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 49160 11830 49188 11999
rect 49148 11824 49200 11830
rect 49148 11766 49200 11772
rect 49146 11656 49202 11665
rect 49146 11591 49202 11600
rect 47768 11552 47820 11558
rect 47768 11494 47820 11500
rect 47308 9988 47360 9994
rect 47308 9930 47360 9936
rect 47320 9625 47348 9930
rect 47306 9616 47362 9625
rect 47124 9580 47176 9586
rect 47306 9551 47362 9560
rect 47124 9522 47176 9528
rect 47780 8974 47808 11494
rect 49160 11218 49188 11591
rect 49238 11248 49294 11257
rect 49148 11212 49200 11218
rect 49238 11183 49294 11192
rect 49148 11154 49200 11160
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 49146 10840 49202 10849
rect 49146 10775 49202 10784
rect 49160 10130 49188 10775
rect 49252 10742 49280 11183
rect 49240 10736 49292 10742
rect 49240 10678 49292 10684
rect 49238 10432 49294 10441
rect 49238 10367 49294 10376
rect 49148 10124 49200 10130
rect 49148 10066 49200 10072
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 49252 9654 49280 10367
rect 49330 10024 49386 10033
rect 49330 9959 49386 9968
rect 49240 9648 49292 9654
rect 49240 9590 49292 9596
rect 49146 9208 49202 9217
rect 49146 9143 49202 9152
rect 47676 8968 47728 8974
rect 47676 8910 47728 8916
rect 47768 8968 47820 8974
rect 47768 8910 47820 8916
rect 47584 8628 47636 8634
rect 47584 8570 47636 8576
rect 47308 7472 47360 7478
rect 47308 7414 47360 7420
rect 44916 7404 44968 7410
rect 44916 7346 44968 7352
rect 47032 7404 47084 7410
rect 47032 7346 47084 7352
rect 45836 7200 45888 7206
rect 45836 7142 45888 7148
rect 43720 5704 43772 5710
rect 43720 5646 43772 5652
rect 45744 5636 45796 5642
rect 45744 5578 45796 5584
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 40224 4752 40276 4758
rect 40224 4694 40276 4700
rect 45652 4276 45704 4282
rect 45652 4218 45704 4224
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 40040 3596 40092 3602
rect 40040 3538 40092 3544
rect 45560 3460 45612 3466
rect 45560 3402 45612 3408
rect 39764 3052 39816 3058
rect 39764 2994 39816 3000
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 41328 2508 41380 2514
rect 41328 2450 41380 2456
rect 41340 800 41368 2450
rect 43444 2304 43496 2310
rect 43444 2246 43496 2252
rect 43456 800 43484 2246
rect 45572 800 45600 3402
rect 45664 2446 45692 4218
rect 45756 3058 45784 5578
rect 45848 5234 45876 7142
rect 46940 6928 46992 6934
rect 46940 6870 46992 6876
rect 45836 5228 45888 5234
rect 45836 5170 45888 5176
rect 46952 4146 46980 6870
rect 47032 6180 47084 6186
rect 47032 6122 47084 6128
rect 45836 4140 45888 4146
rect 45836 4082 45888 4088
rect 46940 4140 46992 4146
rect 46940 4082 46992 4088
rect 45848 3534 45876 4082
rect 46664 4072 46716 4078
rect 46664 4014 46716 4020
rect 45836 3528 45888 3534
rect 45836 3470 45888 3476
rect 45744 3052 45796 3058
rect 45744 2994 45796 3000
rect 45652 2440 45704 2446
rect 45652 2382 45704 2388
rect 46676 1465 46704 4014
rect 47044 3534 47072 6122
rect 47216 5908 47268 5914
rect 47216 5850 47268 5856
rect 47124 4820 47176 4826
rect 47124 4762 47176 4768
rect 47032 3528 47084 3534
rect 47032 3470 47084 3476
rect 46756 2984 46808 2990
rect 46756 2926 46808 2932
rect 46848 2984 46900 2990
rect 46848 2926 46900 2932
rect 46768 1873 46796 2926
rect 46860 2689 46888 2926
rect 46846 2680 46902 2689
rect 46846 2615 46902 2624
rect 47136 2446 47164 4762
rect 47228 3058 47256 5850
rect 47320 4622 47348 7414
rect 47596 5710 47624 8570
rect 47688 6322 47716 8910
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 49160 8566 49188 9143
rect 49344 9042 49372 9959
rect 49332 9036 49384 9042
rect 49332 8978 49384 8984
rect 49238 8800 49294 8809
rect 49238 8735 49294 8744
rect 49148 8560 49200 8566
rect 49148 8502 49200 8508
rect 47768 8356 47820 8362
rect 47768 8298 47820 8304
rect 47780 6798 47808 8298
rect 49252 7954 49280 8735
rect 49330 8392 49386 8401
rect 49330 8327 49386 8336
rect 49240 7948 49292 7954
rect 49240 7890 49292 7896
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 49146 7576 49202 7585
rect 49146 7511 49202 7520
rect 47860 7268 47912 7274
rect 47860 7210 47912 7216
rect 47768 6792 47820 6798
rect 47768 6734 47820 6740
rect 47676 6316 47728 6322
rect 47676 6258 47728 6264
rect 47584 5704 47636 5710
rect 47584 5646 47636 5652
rect 47872 5234 47900 7210
rect 49160 6866 49188 7511
rect 49344 7478 49372 8327
rect 49332 7472 49384 7478
rect 49332 7414 49384 7420
rect 49330 7168 49386 7177
rect 49330 7103 49386 7112
rect 49148 6860 49200 6866
rect 49148 6802 49200 6808
rect 49238 6760 49294 6769
rect 48688 6724 48740 6730
rect 49238 6695 49294 6704
rect 48688 6666 48740 6672
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 48700 6361 48728 6666
rect 48686 6352 48742 6361
rect 48686 6287 48742 6296
rect 49146 5944 49202 5953
rect 49146 5879 49202 5888
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 49160 5302 49188 5879
rect 49252 5778 49280 6695
rect 49344 6390 49372 7103
rect 49332 6384 49384 6390
rect 49332 6326 49384 6332
rect 49240 5772 49292 5778
rect 49240 5714 49292 5720
rect 49422 5536 49478 5545
rect 49422 5471 49478 5480
rect 49148 5296 49200 5302
rect 49148 5238 49200 5244
rect 47860 5228 47912 5234
rect 47860 5170 47912 5176
rect 48320 5160 48372 5166
rect 48320 5102 48372 5108
rect 49330 5128 49386 5137
rect 48332 4729 48360 5102
rect 49330 5063 49386 5072
rect 48318 4720 48374 4729
rect 48318 4655 48374 4664
rect 47308 4616 47360 4622
rect 47308 4558 47360 4564
rect 47676 4548 47728 4554
rect 47676 4490 47728 4496
rect 47688 3942 47716 4490
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 49146 4312 49202 4321
rect 49146 4247 49202 4256
rect 47676 3936 47728 3942
rect 47676 3878 47728 3884
rect 47216 3052 47268 3058
rect 47216 2994 47268 3000
rect 47124 2440 47176 2446
rect 47124 2382 47176 2388
rect 46754 1864 46810 1873
rect 46754 1799 46810 1808
rect 46662 1456 46718 1465
rect 46662 1391 46718 1400
rect 47688 800 47716 3878
rect 49160 3602 49188 4247
rect 49344 4146 49372 5063
rect 49436 4690 49464 5471
rect 49424 4684 49476 4690
rect 49424 4626 49476 4632
rect 49792 4480 49844 4486
rect 49792 4422 49844 4428
rect 49332 4140 49384 4146
rect 49332 4082 49384 4088
rect 49238 3904 49294 3913
rect 49238 3839 49294 3848
rect 49148 3596 49200 3602
rect 49148 3538 49200 3544
rect 49146 3496 49202 3505
rect 48688 3460 48740 3466
rect 49146 3431 49202 3440
rect 48688 3402 48740 3408
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 48700 3097 48728 3402
rect 48686 3088 48742 3097
rect 48686 3023 48742 3032
rect 49160 2514 49188 3431
rect 49252 3126 49280 3839
rect 49240 3120 49292 3126
rect 49240 3062 49292 3068
rect 49148 2508 49200 2514
rect 49148 2450 49200 2456
rect 48504 2372 48556 2378
rect 48504 2314 48556 2320
rect 48516 2281 48544 2314
rect 48502 2272 48558 2281
rect 47950 2204 48258 2213
rect 48502 2207 48558 2216
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 49804 800 49832 4422
rect 28736 734 28948 762
rect 30746 0 30802 800
rect 32862 0 32918 800
rect 34978 0 35034 800
rect 37094 0 37150 800
rect 39210 0 39266 800
rect 41326 0 41382 800
rect 43442 0 43498 800
rect 45558 0 45614 800
rect 47674 0 47730 800
rect 49790 0 49846 800
<< via2 >>
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2778 24384 2834 24440
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 3054 23160 3110 23216
rect 2870 22752 2926 22808
rect 1766 21528 1822 21584
rect 1030 20712 1086 20768
rect 1306 20304 1362 20360
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 3238 21956 3294 21992
rect 3238 21936 3240 21956
rect 3240 21936 3292 21956
rect 3292 21936 3294 21956
rect 3422 25608 3478 25664
rect 3698 25200 3754 25256
rect 3606 24812 3662 24848
rect 3606 24792 3608 24812
rect 3608 24792 3660 24812
rect 3660 24792 3662 24812
rect 3514 23976 3570 24032
rect 3422 23588 3478 23624
rect 3422 23568 3424 23588
rect 3424 23568 3476 23588
rect 3476 23568 3478 23588
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2778 21120 2834 21176
rect 1766 19896 1822 19952
rect 1490 18672 1546 18728
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2870 19488 2926 19544
rect 2778 19080 2834 19136
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 3974 19352 4030 19408
rect 1766 18264 1822 18320
rect 4158 22480 4214 22536
rect 1398 17856 1454 17912
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 1766 17448 1822 17504
rect 938 17040 994 17096
rect 1030 16632 1086 16688
rect 1030 16224 1086 16280
rect 1030 15816 1086 15872
rect 938 15428 994 15464
rect 938 15408 940 15428
rect 940 15408 992 15428
rect 992 15408 994 15428
rect 938 15020 994 15056
rect 938 15000 940 15020
rect 940 15000 992 15020
rect 992 15000 994 15020
rect 938 14592 994 14648
rect 1030 14184 1086 14240
rect 1766 13776 1822 13832
rect 1306 12960 1362 13016
rect 1214 12552 1270 12608
rect 1214 12144 1270 12200
rect 1306 11736 1362 11792
rect 1306 11328 1362 11384
rect 1582 10920 1638 10976
rect 1306 10512 1362 10568
rect 1214 10104 1270 10160
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 5354 18808 5410 18864
rect 7930 24248 7986 24304
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 6550 21548 6606 21584
rect 6550 21528 6552 21548
rect 6552 21528 6604 21548
rect 6604 21528 6606 21548
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 9034 21548 9090 21584
rect 9034 21528 9036 21548
rect 9036 21528 9088 21548
rect 9088 21528 9090 21548
rect 8390 20884 8392 20904
rect 8392 20884 8444 20904
rect 8444 20884 8446 20904
rect 8390 20848 8446 20884
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 3514 13368 3570 13424
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2686 11736 2742 11792
rect 1306 9716 1362 9752
rect 1306 9696 1308 9716
rect 1308 9696 1360 9716
rect 1360 9696 1362 9716
rect 1766 9444 1822 9480
rect 1766 9424 1768 9444
rect 1768 9424 1820 9444
rect 1820 9424 1822 9444
rect 1306 9288 1362 9344
rect 1306 8900 1362 8936
rect 1306 8880 1308 8900
rect 1308 8880 1360 8900
rect 1360 8880 1362 8900
rect 1214 8472 1270 8528
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 9586 15952 9642 16008
rect 11334 23024 11390 23080
rect 10690 20576 10746 20632
rect 10598 19624 10654 19680
rect 10598 17720 10654 17776
rect 10506 16088 10562 16144
rect 11886 22092 11942 22128
rect 11886 22072 11888 22092
rect 11888 22072 11940 22092
rect 11940 22072 11942 22092
rect 11702 21428 11704 21448
rect 11704 21428 11756 21448
rect 11756 21428 11758 21448
rect 11702 21392 11758 21428
rect 12070 19760 12126 19816
rect 11242 18808 11298 18864
rect 11150 18128 11206 18184
rect 10414 14456 10470 14512
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 1306 8084 1362 8120
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 1306 8064 1308 8084
rect 1308 8064 1360 8084
rect 1360 8064 1362 8084
rect 1306 7656 1362 7712
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 1306 7248 1362 7304
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 11242 13776 11298 13832
rect 11150 13096 11206 13152
rect 1214 6840 1270 6896
rect 1306 6432 1362 6488
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 11886 17040 11942 17096
rect 12622 20984 12678 21040
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12898 20984 12954 21040
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12254 17176 12310 17232
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12346 14900 12348 14920
rect 12348 14900 12400 14920
rect 12400 14900 12402 14920
rect 12346 14864 12402 14900
rect 12162 12688 12218 12744
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 13542 16396 13544 16416
rect 13544 16396 13596 16416
rect 13596 16396 13598 16416
rect 13542 16360 13598 16396
rect 13542 15972 13598 16008
rect 13542 15952 13544 15972
rect 13544 15952 13596 15972
rect 13596 15952 13598 15972
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12438 12144 12494 12200
rect 1306 6024 1362 6080
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 1306 5652 1308 5672
rect 1308 5652 1360 5672
rect 1360 5652 1362 5672
rect 1306 5616 1362 5652
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 2778 5208 2834 5264
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 1306 4820 1362 4856
rect 1306 4800 1308 4820
rect 1308 4800 1360 4820
rect 1360 4800 1362 4820
rect 1306 4392 1362 4448
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 1398 3984 1454 4040
rect 5354 3984 5410 4040
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 1306 3576 1362 3632
rect 1122 3440 1178 3496
rect 1306 3188 1362 3224
rect 1306 3168 1308 3188
rect 1308 3168 1360 3188
rect 1360 3168 1362 3188
rect 1306 2760 1362 2816
rect 1306 2388 1308 2408
rect 1308 2388 1360 2408
rect 1360 2388 1362 2408
rect 1306 2352 1362 2388
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 1214 1944 1270 2000
rect 1306 1536 1362 1592
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 13358 12552 13414 12608
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 13358 12008 13414 12064
rect 14094 20596 14150 20632
rect 14094 20576 14096 20596
rect 14096 20576 14148 20596
rect 14148 20576 14150 20596
rect 14094 18264 14150 18320
rect 14830 18692 14886 18728
rect 14830 18672 14832 18692
rect 14832 18672 14884 18692
rect 14884 18672 14886 18692
rect 15014 18128 15070 18184
rect 15566 21528 15622 21584
rect 15474 19896 15530 19952
rect 14002 16360 14058 16416
rect 14830 16396 14832 16416
rect 14832 16396 14884 16416
rect 14884 16396 14886 16416
rect 13726 12552 13782 12608
rect 14830 16360 14886 16396
rect 14186 16088 14242 16144
rect 14554 16088 14610 16144
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 13450 10920 13506 10976
rect 13450 10548 13452 10568
rect 13452 10548 13504 10568
rect 13504 10548 13506 10568
rect 13450 10512 13506 10548
rect 15842 19624 15898 19680
rect 16210 20304 16266 20360
rect 15106 16632 15162 16688
rect 14554 13368 14610 13424
rect 14554 13096 14610 13152
rect 14830 15036 14832 15056
rect 14832 15036 14884 15056
rect 14884 15036 14886 15056
rect 14830 15000 14886 15036
rect 14830 12960 14886 13016
rect 14830 10920 14886 10976
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 15290 12980 15346 13016
rect 15290 12960 15292 12980
rect 15292 12960 15344 12980
rect 15344 12960 15346 12980
rect 16026 19252 16028 19272
rect 16028 19252 16080 19272
rect 16080 19252 16082 19272
rect 16026 19216 16082 19252
rect 16302 18692 16358 18728
rect 16302 18672 16304 18692
rect 16304 18672 16356 18692
rect 16356 18672 16358 18692
rect 15842 16088 15898 16144
rect 16026 15952 16082 16008
rect 15842 15408 15898 15464
rect 15842 12164 15898 12200
rect 15842 12144 15844 12164
rect 15844 12144 15896 12164
rect 15896 12144 15898 12164
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 16578 17992 16634 18048
rect 16302 16632 16358 16688
rect 16486 13640 16542 13696
rect 16302 12688 16358 12744
rect 16210 12416 16266 12472
rect 16026 10920 16082 10976
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 18602 21392 18658 21448
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17406 18692 17462 18728
rect 17406 18672 17408 18692
rect 17408 18672 17460 18692
rect 17460 18672 17462 18692
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17406 16940 17408 16960
rect 17408 16940 17460 16960
rect 17460 16940 17462 16960
rect 17406 16904 17462 16940
rect 17498 16632 17554 16688
rect 17222 15544 17278 15600
rect 16762 12144 16818 12200
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 19798 22616 19854 22672
rect 19614 22072 19670 22128
rect 19338 19352 19394 19408
rect 18970 17176 19026 17232
rect 18510 15020 18566 15056
rect 18510 15000 18512 15020
rect 18512 15000 18564 15020
rect 18564 15000 18566 15020
rect 18510 14864 18566 14920
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17406 12960 17462 13016
rect 17222 12280 17278 12336
rect 17222 12044 17224 12064
rect 17224 12044 17276 12064
rect 17276 12044 17278 12064
rect 17222 12008 17278 12044
rect 16946 11736 17002 11792
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18510 13232 18566 13288
rect 19338 18692 19394 18728
rect 19338 18672 19340 18692
rect 19340 18672 19392 18692
rect 19392 18672 19394 18692
rect 21270 23724 21326 23760
rect 21270 23704 21272 23724
rect 21272 23704 21324 23724
rect 21324 23704 21326 23724
rect 21270 22072 21326 22128
rect 19338 17992 19394 18048
rect 19154 15544 19210 15600
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 20350 18808 20406 18864
rect 20626 19216 20682 19272
rect 20350 17992 20406 18048
rect 21270 19508 21326 19544
rect 21270 19488 21272 19508
rect 21272 19488 21324 19508
rect 21324 19488 21326 19508
rect 19246 13232 19302 13288
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 20074 14320 20130 14376
rect 20074 13776 20130 13832
rect 20810 15700 20866 15736
rect 20810 15680 20812 15700
rect 20812 15680 20864 15700
rect 20864 15680 20866 15700
rect 20626 11756 20682 11792
rect 20626 11736 20628 11756
rect 20628 11736 20680 11756
rect 20680 11736 20682 11756
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 23294 23024 23350 23080
rect 22282 21800 22338 21856
rect 21914 20984 21970 21040
rect 21454 18572 21456 18592
rect 21456 18572 21508 18592
rect 21508 18572 21510 18592
rect 21454 18536 21510 18572
rect 21178 15544 21234 15600
rect 21822 16904 21878 16960
rect 21454 14456 21510 14512
rect 21638 14320 21694 14376
rect 21454 13096 21510 13152
rect 21362 10104 21418 10160
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 23110 21836 23112 21856
rect 23112 21836 23164 21856
rect 23164 21836 23166 21856
rect 23110 21800 23166 21836
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23754 22208 23810 22264
rect 22374 18400 22430 18456
rect 22098 17040 22154 17096
rect 23754 20848 23810 20904
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22558 17992 22614 18048
rect 22466 17312 22522 17368
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 23018 18536 23074 18592
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 23938 20032 23994 20088
rect 22466 16496 22522 16552
rect 22558 15700 22614 15736
rect 22558 15680 22560 15700
rect 22560 15680 22612 15700
rect 22612 15680 22614 15700
rect 22098 12960 22154 13016
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 23662 16768 23718 16824
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22742 12824 22798 12880
rect 22558 12280 22614 12336
rect 22926 12980 22982 13016
rect 22926 12960 22928 12980
rect 22928 12960 22980 12980
rect 22980 12960 22982 12980
rect 23018 12688 23074 12744
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 25778 24284 25780 24304
rect 25780 24284 25832 24304
rect 25832 24284 25834 24304
rect 25778 24248 25834 24284
rect 24766 22480 24822 22536
rect 25318 22924 25320 22944
rect 25320 22924 25372 22944
rect 25372 22924 25374 22944
rect 25318 22888 25374 22924
rect 25134 22344 25190 22400
rect 24490 22072 24546 22128
rect 24122 19488 24178 19544
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 24490 20168 24546 20224
rect 24950 21392 25006 21448
rect 25042 19624 25098 19680
rect 24582 16768 24638 16824
rect 25042 18284 25098 18320
rect 25042 18264 25044 18284
rect 25044 18264 25096 18284
rect 25096 18264 25098 18284
rect 24766 17176 24822 17232
rect 25226 20168 25282 20224
rect 25870 20848 25926 20904
rect 26054 21548 26110 21584
rect 26054 21528 26056 21548
rect 26056 21528 26108 21548
rect 26108 21528 26110 21548
rect 25594 18944 25650 19000
rect 25594 18400 25650 18456
rect 25410 17992 25466 18048
rect 25778 17212 25780 17232
rect 25780 17212 25832 17232
rect 25832 17212 25834 17232
rect 25778 17176 25834 17212
rect 24858 15952 24914 16008
rect 24674 13368 24730 13424
rect 24030 11056 24086 11112
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 24858 11736 24914 11792
rect 25778 16768 25834 16824
rect 26606 24132 26662 24168
rect 26606 24112 26608 24132
rect 26608 24112 26660 24132
rect 26660 24112 26662 24132
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 26146 19896 26202 19952
rect 26330 19896 26386 19952
rect 26054 19216 26110 19272
rect 25962 18264 26018 18320
rect 26330 18128 26386 18184
rect 25686 16088 25742 16144
rect 27618 21936 27674 21992
rect 28446 23704 28502 23760
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 28262 22228 28318 22264
rect 28262 22208 28264 22228
rect 28264 22208 28316 22228
rect 28316 22208 28318 22228
rect 27434 20984 27490 21040
rect 26698 19488 26754 19544
rect 26054 15272 26110 15328
rect 26054 13096 26110 13152
rect 26790 16768 26846 16824
rect 26238 12980 26294 13016
rect 26238 12960 26240 12980
rect 26240 12960 26292 12980
rect 26292 12960 26294 12980
rect 26422 12844 26478 12880
rect 26422 12824 26424 12844
rect 26424 12824 26476 12844
rect 26476 12824 26478 12844
rect 25962 12688 26018 12744
rect 26790 15544 26846 15600
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 27802 21120 27858 21176
rect 28814 21428 28816 21448
rect 28816 21428 28868 21448
rect 28868 21428 28870 21448
rect 28814 21392 28870 21428
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 27526 18944 27582 19000
rect 27710 19488 27766 19544
rect 27986 19932 27988 19952
rect 27988 19932 28040 19952
rect 28040 19932 28042 19952
rect 27986 19896 28042 19932
rect 28446 19896 28502 19952
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 27710 17332 27766 17368
rect 28354 19352 28410 19408
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 27710 17312 27712 17332
rect 27712 17312 27764 17332
rect 27764 17312 27766 17332
rect 28262 17176 28318 17232
rect 27710 17040 27766 17096
rect 27434 16768 27490 16824
rect 27066 15408 27122 15464
rect 27158 15308 27160 15328
rect 27160 15308 27212 15328
rect 27212 15308 27214 15328
rect 27158 15272 27214 15308
rect 27250 15020 27306 15056
rect 27250 15000 27252 15020
rect 27252 15000 27304 15020
rect 27304 15000 27306 15020
rect 26238 10104 26294 10160
rect 24858 4020 24860 4040
rect 24860 4020 24912 4040
rect 24912 4020 24914 4040
rect 24858 3984 24914 4020
rect 25778 3440 25834 3496
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 27802 16768 27858 16824
rect 27986 16652 28042 16688
rect 27986 16632 27988 16652
rect 27988 16632 28040 16652
rect 28040 16632 28042 16652
rect 28814 19624 28870 19680
rect 28722 18672 28778 18728
rect 28446 17992 28502 18048
rect 28722 18128 28778 18184
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 28998 18844 29000 18864
rect 29000 18844 29052 18864
rect 29052 18844 29054 18864
rect 28998 18808 29054 18844
rect 30194 23568 30250 23624
rect 29642 22616 29698 22672
rect 29734 22344 29790 22400
rect 29642 20984 29698 21040
rect 29182 15272 29238 15328
rect 28998 15136 29054 15192
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 27250 10104 27306 10160
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 28446 12824 28502 12880
rect 28630 11056 28686 11112
rect 30010 21140 30066 21176
rect 30010 21120 30012 21140
rect 30012 21120 30064 21140
rect 30064 21120 30066 21140
rect 29642 18400 29698 18456
rect 29826 19352 29882 19408
rect 30194 21936 30250 21992
rect 30746 22752 30802 22808
rect 30654 22652 30656 22672
rect 30656 22652 30708 22672
rect 30708 22652 30710 22672
rect 30654 22616 30710 22652
rect 30378 21392 30434 21448
rect 30378 20576 30434 20632
rect 30102 20304 30158 20360
rect 30194 18536 30250 18592
rect 29918 17448 29974 17504
rect 30746 21392 30802 21448
rect 30654 20712 30710 20768
rect 30378 17448 30434 17504
rect 29918 15680 29974 15736
rect 29734 12280 29790 12336
rect 29642 12144 29698 12200
rect 30010 11056 30066 11112
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 31942 24656 31998 24712
rect 31482 22480 31538 22536
rect 32126 23840 32182 23896
rect 31206 21548 31262 21584
rect 31206 21528 31208 21548
rect 31208 21528 31260 21548
rect 31260 21528 31262 21548
rect 31390 21120 31446 21176
rect 31114 19760 31170 19816
rect 30930 18672 30986 18728
rect 30562 15136 30618 15192
rect 30654 14900 30656 14920
rect 30656 14900 30708 14920
rect 30708 14900 30710 14920
rect 30654 14864 30710 14900
rect 31298 18808 31354 18864
rect 31758 20984 31814 21040
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32862 24248 32918 24304
rect 32494 23160 32550 23216
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 33782 23840 33838 23896
rect 33690 23704 33746 23760
rect 33598 23296 33654 23352
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 32862 21392 32918 21448
rect 31390 17312 31446 17368
rect 31206 15272 31262 15328
rect 30562 13776 30618 13832
rect 30562 13232 30618 13288
rect 31850 14900 31852 14920
rect 31852 14900 31904 14920
rect 31904 14900 31906 14920
rect 31850 14864 31906 14900
rect 32770 20324 32826 20360
rect 32770 20304 32772 20324
rect 32772 20304 32824 20324
rect 32824 20304 32826 20324
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 33506 21548 33562 21584
rect 33506 21528 33508 21548
rect 33508 21528 33560 21548
rect 33560 21528 33562 21548
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 34058 23432 34114 23488
rect 33966 22208 34022 22264
rect 34242 22480 34298 22536
rect 33874 19624 33930 19680
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 30838 9016 30894 9072
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 34242 21664 34298 21720
rect 34702 24520 34758 24576
rect 34702 22752 34758 22808
rect 34426 21256 34482 21312
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 34334 18828 34390 18864
rect 34334 18808 34336 18828
rect 34336 18808 34388 18828
rect 34388 18808 34390 18828
rect 35254 24384 35310 24440
rect 35162 23976 35218 24032
rect 35438 23588 35494 23624
rect 35438 23568 35440 23588
rect 35440 23568 35492 23588
rect 35492 23568 35494 23588
rect 35438 23024 35494 23080
rect 34886 22616 34942 22672
rect 34702 20440 34758 20496
rect 34886 19780 34942 19816
rect 34886 19760 34888 19780
rect 34888 19760 34940 19780
rect 34940 19760 34942 19780
rect 34978 19216 35034 19272
rect 34610 18400 34666 18456
rect 34334 13776 34390 13832
rect 34242 9424 34298 9480
rect 35346 20032 35402 20088
rect 35346 19488 35402 19544
rect 36082 23296 36138 23352
rect 35162 13252 35218 13288
rect 35162 13232 35164 13252
rect 35164 13232 35216 13252
rect 35216 13232 35218 13252
rect 35346 17312 35402 17368
rect 35530 17484 35532 17504
rect 35532 17484 35584 17504
rect 35584 17484 35586 17504
rect 35530 17448 35586 17484
rect 35438 15408 35494 15464
rect 35622 15544 35678 15600
rect 35622 13640 35678 13696
rect 36082 20712 36138 20768
rect 36634 21936 36690 21992
rect 36450 21392 36506 21448
rect 36634 21120 36690 21176
rect 37186 22072 37242 22128
rect 37002 21936 37058 21992
rect 36910 21664 36966 21720
rect 37554 23296 37610 23352
rect 37738 24384 37794 24440
rect 37738 24012 37740 24032
rect 37740 24012 37792 24032
rect 37792 24012 37794 24032
rect 37738 23976 37794 24012
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 38658 24248 38714 24304
rect 38290 22616 38346 22672
rect 38566 22772 38622 22808
rect 38566 22752 38568 22772
rect 38568 22752 38620 22772
rect 38620 22752 38622 22772
rect 39854 24404 39910 24440
rect 39854 24384 39856 24404
rect 39856 24384 39908 24404
rect 39908 24384 39910 24404
rect 39302 23024 39358 23080
rect 39210 22888 39266 22944
rect 38382 22344 38438 22400
rect 38842 22092 38898 22128
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 35806 15952 35862 16008
rect 36082 18536 36138 18592
rect 35898 14864 35954 14920
rect 35806 14456 35862 14512
rect 35162 10512 35218 10568
rect 36818 19216 36874 19272
rect 37094 18944 37150 19000
rect 36818 17992 36874 18048
rect 37370 20576 37426 20632
rect 38842 22072 38844 22092
rect 38844 22072 38896 22092
rect 38896 22072 38898 22092
rect 39486 23296 39542 23352
rect 38382 20712 38438 20768
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 36726 13676 36728 13696
rect 36728 13676 36780 13696
rect 36780 13676 36782 13696
rect 36726 13640 36782 13676
rect 36266 9052 36268 9072
rect 36268 9052 36320 9072
rect 36320 9052 36322 9072
rect 36266 9016 36322 9052
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 38290 18944 38346 19000
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 40222 23704 40278 23760
rect 40038 23432 40094 23488
rect 40314 21664 40370 21720
rect 40222 21120 40278 21176
rect 39394 20032 39450 20088
rect 40038 19216 40094 19272
rect 40038 18672 40094 18728
rect 40406 20848 40462 20904
rect 40682 21392 40738 21448
rect 40866 21292 40868 21312
rect 40868 21292 40920 21312
rect 40920 21292 40922 21312
rect 40866 21256 40922 21292
rect 40498 18264 40554 18320
rect 40222 17856 40278 17912
rect 38382 15272 38438 15328
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 38014 11056 38070 11112
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 39762 16496 39818 16552
rect 41510 23296 41566 23352
rect 41418 22752 41474 22808
rect 41878 22500 41934 22536
rect 41878 22480 41880 22500
rect 41880 22480 41932 22500
rect 41932 22480 41934 22500
rect 41234 20984 41290 21040
rect 41234 19216 41290 19272
rect 39670 14884 39726 14920
rect 39670 14864 39672 14884
rect 39672 14864 39724 14884
rect 39724 14864 39726 14884
rect 40130 15272 40186 15328
rect 41878 21664 41934 21720
rect 43902 24656 43958 24712
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 42614 22344 42670 22400
rect 43350 23160 43406 23216
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 42798 21972 42800 21992
rect 42800 21972 42852 21992
rect 42852 21972 42854 21992
rect 42798 21936 42854 21972
rect 41510 19352 41566 19408
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 42798 19080 42854 19136
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 41326 18128 41382 18184
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 43902 23160 43958 23216
rect 45190 24248 45246 24304
rect 44730 22636 44786 22672
rect 44730 22616 44732 22636
rect 44732 22616 44784 22636
rect 44784 22616 44786 22636
rect 44454 22072 44510 22128
rect 43902 21528 43958 21584
rect 46754 25064 46810 25120
rect 45374 22072 45430 22128
rect 44546 19760 44602 19816
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 46662 23704 46718 23760
rect 47582 24656 47638 24712
rect 46846 23432 46902 23488
rect 46938 22888 46994 22944
rect 47766 24248 47822 24304
rect 48226 25472 48282 25528
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 47674 20848 47730 20904
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 48778 24148 48780 24168
rect 48780 24148 48832 24168
rect 48832 24148 48834 24168
rect 48778 24112 48834 24148
rect 48686 23060 48688 23080
rect 48688 23060 48740 23080
rect 48740 23060 48742 23080
rect 48686 23024 48742 23060
rect 49422 22616 49478 22672
rect 48594 21800 48650 21856
rect 48410 20304 48466 20360
rect 48318 19896 48374 19952
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 49330 22208 49386 22264
rect 49238 21392 49294 21448
rect 49330 21020 49332 21040
rect 49332 21020 49384 21040
rect 49384 21020 49386 21040
rect 49330 20984 49386 21020
rect 49330 20576 49386 20632
rect 49054 20440 49110 20496
rect 48778 20168 48834 20224
rect 49422 19760 49478 19816
rect 49330 19352 49386 19408
rect 49146 19216 49202 19272
rect 49238 18944 49294 19000
rect 48686 18808 48742 18864
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 48778 18536 48834 18592
rect 49422 18128 49478 18184
rect 49330 17720 49386 17776
rect 48502 17176 48558 17232
rect 49054 17076 49056 17096
rect 49056 17076 49108 17096
rect 49108 17076 49110 17096
rect 49054 17040 49110 17076
rect 48778 16904 48834 16960
rect 49330 17312 49386 17368
rect 49146 16632 49202 16688
rect 48226 16496 48282 16552
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 49146 16088 49202 16144
rect 49422 16088 49478 16144
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 49146 15972 49202 16008
rect 49146 15952 49148 15972
rect 49148 15952 49200 15972
rect 49200 15952 49202 15972
rect 49330 15680 49386 15736
rect 49330 15272 49386 15328
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 40038 12844 40094 12880
rect 40038 12824 40040 12844
rect 40040 12824 40092 12844
rect 40092 12824 40094 12844
rect 40130 12164 40186 12200
rect 40130 12144 40132 12164
rect 40132 12144 40184 12164
rect 40184 12144 40186 12164
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 49146 15000 49202 15056
rect 49054 14356 49056 14376
rect 49056 14356 49108 14376
rect 49108 14356 49110 14376
rect 49054 14320 49110 14356
rect 49330 14864 49386 14920
rect 49238 14456 49294 14512
rect 49238 14048 49294 14104
rect 48226 13640 48282 13696
rect 49146 13268 49148 13288
rect 49148 13268 49200 13288
rect 49200 13268 49202 13288
rect 49146 13232 49202 13268
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 49146 12844 49202 12880
rect 49146 12824 49148 12844
rect 49148 12824 49200 12844
rect 49200 12824 49202 12844
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 46846 7928 46902 7984
rect 49146 12416 49202 12472
rect 49146 12008 49202 12064
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 49146 11600 49202 11656
rect 47306 9560 47362 9616
rect 49238 11192 49294 11248
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 49146 10784 49202 10840
rect 49238 10376 49294 10432
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 49330 9968 49386 10024
rect 49146 9152 49202 9208
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 46846 2624 46902 2680
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 49238 8744 49294 8800
rect 49330 8336 49386 8392
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 49146 7520 49202 7576
rect 49330 7112 49386 7168
rect 49238 6704 49294 6760
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 48686 6296 48742 6352
rect 49146 5888 49202 5944
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 49422 5480 49478 5536
rect 49330 5072 49386 5128
rect 48318 4664 48374 4720
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 49146 4256 49202 4312
rect 46754 1808 46810 1864
rect 46662 1400 46718 1456
rect 49238 3848 49294 3904
rect 49146 3440 49202 3496
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 48686 3032 48742 3088
rect 48502 2216 48558 2272
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
<< metal3 >>
rect 0 25666 800 25696
rect 3417 25666 3483 25669
rect 0 25664 3483 25666
rect 0 25608 3422 25664
rect 3478 25608 3483 25664
rect 0 25606 3483 25608
rect 0 25576 800 25606
rect 3417 25603 3483 25606
rect 48221 25530 48287 25533
rect 50200 25530 51000 25560
rect 48221 25528 51000 25530
rect 48221 25472 48226 25528
rect 48282 25472 51000 25528
rect 48221 25470 51000 25472
rect 48221 25467 48287 25470
rect 50200 25440 51000 25470
rect 0 25258 800 25288
rect 3693 25258 3759 25261
rect 0 25256 3759 25258
rect 0 25200 3698 25256
rect 3754 25200 3759 25256
rect 0 25198 3759 25200
rect 0 25168 800 25198
rect 3693 25195 3759 25198
rect 46749 25122 46815 25125
rect 50200 25122 51000 25152
rect 46749 25120 51000 25122
rect 46749 25064 46754 25120
rect 46810 25064 51000 25120
rect 46749 25062 51000 25064
rect 46749 25059 46815 25062
rect 50200 25032 51000 25062
rect 0 24850 800 24880
rect 3601 24850 3667 24853
rect 0 24848 3667 24850
rect 0 24792 3606 24848
rect 3662 24792 3667 24848
rect 0 24790 3667 24792
rect 0 24760 800 24790
rect 3601 24787 3667 24790
rect 31937 24714 32003 24717
rect 43897 24714 43963 24717
rect 31937 24712 43963 24714
rect 31937 24656 31942 24712
rect 31998 24656 43902 24712
rect 43958 24656 43963 24712
rect 31937 24654 43963 24656
rect 31937 24651 32003 24654
rect 43897 24651 43963 24654
rect 47577 24714 47643 24717
rect 50200 24714 51000 24744
rect 47577 24712 51000 24714
rect 47577 24656 47582 24712
rect 47638 24656 51000 24712
rect 47577 24654 51000 24656
rect 47577 24651 47643 24654
rect 50200 24624 51000 24654
rect 34697 24578 34763 24581
rect 34697 24576 41430 24578
rect 34697 24520 34702 24576
rect 34758 24520 41430 24576
rect 34697 24518 41430 24520
rect 34697 24515 34763 24518
rect 2946 24512 3262 24513
rect 0 24442 800 24472
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 2773 24442 2839 24445
rect 0 24440 2839 24442
rect 0 24384 2778 24440
rect 2834 24384 2839 24440
rect 0 24382 2839 24384
rect 0 24352 800 24382
rect 2773 24379 2839 24382
rect 35249 24442 35315 24445
rect 37733 24442 37799 24445
rect 39849 24442 39915 24445
rect 35249 24440 39915 24442
rect 35249 24384 35254 24440
rect 35310 24384 37738 24440
rect 37794 24384 39854 24440
rect 39910 24384 39915 24440
rect 35249 24382 39915 24384
rect 35249 24379 35315 24382
rect 37733 24379 37799 24382
rect 39849 24379 39915 24382
rect 7925 24306 7991 24309
rect 25773 24306 25839 24309
rect 7925 24304 25839 24306
rect 7925 24248 7930 24304
rect 7986 24248 25778 24304
rect 25834 24248 25839 24304
rect 7925 24246 25839 24248
rect 7925 24243 7991 24246
rect 25773 24243 25839 24246
rect 32857 24306 32923 24309
rect 38653 24306 38719 24309
rect 32857 24304 38719 24306
rect 32857 24248 32862 24304
rect 32918 24248 38658 24304
rect 38714 24248 38719 24304
rect 32857 24246 38719 24248
rect 41370 24306 41430 24518
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 45185 24306 45251 24309
rect 41370 24304 45251 24306
rect 41370 24248 45190 24304
rect 45246 24248 45251 24304
rect 41370 24246 45251 24248
rect 32857 24243 32923 24246
rect 38653 24243 38719 24246
rect 45185 24243 45251 24246
rect 47761 24306 47827 24309
rect 50200 24306 51000 24336
rect 47761 24304 51000 24306
rect 47761 24248 47766 24304
rect 47822 24248 51000 24304
rect 47761 24246 51000 24248
rect 47761 24243 47827 24246
rect 50200 24216 51000 24246
rect 26601 24170 26667 24173
rect 48773 24170 48839 24173
rect 26601 24168 48839 24170
rect 26601 24112 26606 24168
rect 26662 24112 48778 24168
rect 48834 24112 48839 24168
rect 26601 24110 48839 24112
rect 26601 24107 26667 24110
rect 48773 24107 48839 24110
rect 0 24034 800 24064
rect 3509 24034 3575 24037
rect 0 24032 3575 24034
rect 0 23976 3514 24032
rect 3570 23976 3575 24032
rect 0 23974 3575 23976
rect 0 23944 800 23974
rect 3509 23971 3575 23974
rect 35157 24034 35223 24037
rect 37733 24034 37799 24037
rect 35157 24032 37799 24034
rect 35157 23976 35162 24032
rect 35218 23976 37738 24032
rect 37794 23976 37799 24032
rect 35157 23974 37799 23976
rect 35157 23971 35223 23974
rect 37733 23971 37799 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 32121 23898 32187 23901
rect 33777 23898 33843 23901
rect 50200 23898 51000 23928
rect 32121 23896 33843 23898
rect 32121 23840 32126 23896
rect 32182 23840 33782 23896
rect 33838 23840 33843 23896
rect 32121 23838 33843 23840
rect 32121 23835 32187 23838
rect 33777 23835 33843 23838
rect 48454 23838 51000 23898
rect 21265 23762 21331 23765
rect 28441 23762 28507 23765
rect 21265 23760 28507 23762
rect 21265 23704 21270 23760
rect 21326 23704 28446 23760
rect 28502 23704 28507 23760
rect 21265 23702 28507 23704
rect 21265 23699 21331 23702
rect 28441 23699 28507 23702
rect 33685 23762 33751 23765
rect 40217 23762 40283 23765
rect 33685 23760 40283 23762
rect 33685 23704 33690 23760
rect 33746 23704 40222 23760
rect 40278 23704 40283 23760
rect 33685 23702 40283 23704
rect 33685 23699 33751 23702
rect 40217 23699 40283 23702
rect 46657 23762 46723 23765
rect 48454 23762 48514 23838
rect 50200 23808 51000 23838
rect 46657 23760 48514 23762
rect 46657 23704 46662 23760
rect 46718 23704 48514 23760
rect 46657 23702 48514 23704
rect 46657 23699 46723 23702
rect 0 23626 800 23656
rect 3417 23626 3483 23629
rect 0 23624 3483 23626
rect 0 23568 3422 23624
rect 3478 23568 3483 23624
rect 0 23566 3483 23568
rect 0 23536 800 23566
rect 3417 23563 3483 23566
rect 30189 23626 30255 23629
rect 35433 23626 35499 23629
rect 30189 23624 35499 23626
rect 30189 23568 30194 23624
rect 30250 23568 35438 23624
rect 35494 23568 35499 23624
rect 30189 23566 35499 23568
rect 30189 23563 30255 23566
rect 35433 23563 35499 23566
rect 34053 23490 34119 23493
rect 40033 23490 40099 23493
rect 34053 23488 40099 23490
rect 34053 23432 34058 23488
rect 34114 23432 40038 23488
rect 40094 23432 40099 23488
rect 34053 23430 40099 23432
rect 34053 23427 34119 23430
rect 40033 23427 40099 23430
rect 46841 23490 46907 23493
rect 50200 23490 51000 23520
rect 46841 23488 51000 23490
rect 46841 23432 46846 23488
rect 46902 23432 51000 23488
rect 46841 23430 51000 23432
rect 46841 23427 46907 23430
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 50200 23400 51000 23430
rect 42946 23359 43262 23360
rect 33593 23354 33659 23357
rect 36077 23354 36143 23357
rect 33593 23352 36143 23354
rect 33593 23296 33598 23352
rect 33654 23296 36082 23352
rect 36138 23296 36143 23352
rect 33593 23294 36143 23296
rect 33593 23291 33659 23294
rect 36077 23291 36143 23294
rect 37549 23354 37615 23357
rect 39481 23354 39547 23357
rect 41505 23354 41571 23357
rect 37549 23352 41571 23354
rect 37549 23296 37554 23352
rect 37610 23296 39486 23352
rect 39542 23296 41510 23352
rect 41566 23296 41571 23352
rect 37549 23294 41571 23296
rect 37549 23291 37615 23294
rect 39481 23291 39547 23294
rect 41505 23291 41571 23294
rect 0 23218 800 23248
rect 3049 23218 3115 23221
rect 0 23216 3115 23218
rect 0 23160 3054 23216
rect 3110 23160 3115 23216
rect 0 23158 3115 23160
rect 0 23128 800 23158
rect 3049 23155 3115 23158
rect 32489 23218 32555 23221
rect 43345 23218 43411 23221
rect 43897 23218 43963 23221
rect 32489 23216 43963 23218
rect 32489 23160 32494 23216
rect 32550 23160 43350 23216
rect 43406 23160 43902 23216
rect 43958 23160 43963 23216
rect 32489 23158 43963 23160
rect 32489 23155 32555 23158
rect 43345 23155 43411 23158
rect 43897 23155 43963 23158
rect 11329 23082 11395 23085
rect 23289 23082 23355 23085
rect 11329 23080 23355 23082
rect 11329 23024 11334 23080
rect 11390 23024 23294 23080
rect 23350 23024 23355 23080
rect 11329 23022 23355 23024
rect 11329 23019 11395 23022
rect 23289 23019 23355 23022
rect 35433 23082 35499 23085
rect 39297 23082 39363 23085
rect 35433 23080 39363 23082
rect 35433 23024 35438 23080
rect 35494 23024 39302 23080
rect 39358 23024 39363 23080
rect 35433 23022 39363 23024
rect 35433 23019 35499 23022
rect 39297 23019 39363 23022
rect 48681 23082 48747 23085
rect 50200 23082 51000 23112
rect 48681 23080 51000 23082
rect 48681 23024 48686 23080
rect 48742 23024 51000 23080
rect 48681 23022 51000 23024
rect 48681 23019 48747 23022
rect 50200 22992 51000 23022
rect 25313 22948 25379 22949
rect 25262 22884 25268 22948
rect 25332 22946 25379 22948
rect 39205 22946 39271 22949
rect 46933 22946 46999 22949
rect 25332 22944 25424 22946
rect 25374 22888 25424 22944
rect 25332 22886 25424 22888
rect 39205 22944 46999 22946
rect 39205 22888 39210 22944
rect 39266 22888 46938 22944
rect 46994 22888 46999 22944
rect 39205 22886 46999 22888
rect 25332 22884 25379 22886
rect 25313 22883 25379 22884
rect 39205 22883 39271 22886
rect 46933 22883 46999 22886
rect 7946 22880 8262 22881
rect 0 22810 800 22840
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 47946 22815 48262 22816
rect 2865 22810 2931 22813
rect 0 22808 2931 22810
rect 0 22752 2870 22808
rect 2926 22752 2931 22808
rect 0 22750 2931 22752
rect 0 22720 800 22750
rect 2865 22747 2931 22750
rect 30741 22810 30807 22813
rect 34697 22810 34763 22813
rect 30741 22808 34763 22810
rect 30741 22752 30746 22808
rect 30802 22752 34702 22808
rect 34758 22752 34763 22808
rect 30741 22750 34763 22752
rect 30741 22747 30807 22750
rect 34697 22747 34763 22750
rect 38561 22810 38627 22813
rect 41413 22810 41479 22813
rect 38561 22808 41479 22810
rect 38561 22752 38566 22808
rect 38622 22752 41418 22808
rect 41474 22752 41479 22808
rect 38561 22750 41479 22752
rect 38561 22747 38627 22750
rect 41413 22747 41479 22750
rect 19793 22674 19859 22677
rect 29637 22674 29703 22677
rect 19793 22672 29703 22674
rect 19793 22616 19798 22672
rect 19854 22616 29642 22672
rect 29698 22616 29703 22672
rect 19793 22614 29703 22616
rect 19793 22611 19859 22614
rect 29637 22611 29703 22614
rect 30649 22674 30715 22677
rect 34881 22674 34947 22677
rect 30649 22672 34947 22674
rect 30649 22616 30654 22672
rect 30710 22616 34886 22672
rect 34942 22616 34947 22672
rect 30649 22614 34947 22616
rect 30649 22611 30715 22614
rect 34881 22611 34947 22614
rect 38285 22674 38351 22677
rect 44725 22674 44791 22677
rect 38285 22672 44791 22674
rect 38285 22616 38290 22672
rect 38346 22616 44730 22672
rect 44786 22616 44791 22672
rect 38285 22614 44791 22616
rect 38285 22611 38351 22614
rect 44725 22611 44791 22614
rect 49417 22674 49483 22677
rect 50200 22674 51000 22704
rect 49417 22672 51000 22674
rect 49417 22616 49422 22672
rect 49478 22616 51000 22672
rect 49417 22614 51000 22616
rect 49417 22611 49483 22614
rect 50200 22584 51000 22614
rect 4153 22538 4219 22541
rect 2086 22536 4219 22538
rect 2086 22480 4158 22536
rect 4214 22480 4219 22536
rect 2086 22478 4219 22480
rect 0 22402 800 22432
rect 2086 22402 2146 22478
rect 4153 22475 4219 22478
rect 24761 22538 24827 22541
rect 31477 22538 31543 22541
rect 24761 22536 31543 22538
rect 24761 22480 24766 22536
rect 24822 22480 31482 22536
rect 31538 22480 31543 22536
rect 24761 22478 31543 22480
rect 24761 22475 24827 22478
rect 31477 22475 31543 22478
rect 34237 22538 34303 22541
rect 41873 22538 41939 22541
rect 34237 22536 41939 22538
rect 34237 22480 34242 22536
rect 34298 22480 41878 22536
rect 41934 22480 41939 22536
rect 34237 22478 41939 22480
rect 34237 22475 34303 22478
rect 41873 22475 41939 22478
rect 0 22342 2146 22402
rect 25129 22402 25195 22405
rect 29729 22402 29795 22405
rect 25129 22400 29795 22402
rect 25129 22344 25134 22400
rect 25190 22344 29734 22400
rect 29790 22344 29795 22400
rect 25129 22342 29795 22344
rect 0 22312 800 22342
rect 25129 22339 25195 22342
rect 29729 22339 29795 22342
rect 38377 22402 38443 22405
rect 42609 22402 42675 22405
rect 38377 22400 42675 22402
rect 38377 22344 38382 22400
rect 38438 22344 42614 22400
rect 42670 22344 42675 22400
rect 38377 22342 42675 22344
rect 38377 22339 38443 22342
rect 42609 22339 42675 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 23749 22266 23815 22269
rect 28257 22266 28323 22269
rect 23749 22264 28323 22266
rect 23749 22208 23754 22264
rect 23810 22208 28262 22264
rect 28318 22208 28323 22264
rect 23749 22206 28323 22208
rect 23749 22203 23815 22206
rect 28257 22203 28323 22206
rect 33961 22266 34027 22269
rect 49325 22266 49391 22269
rect 50200 22266 51000 22296
rect 33961 22264 41430 22266
rect 33961 22208 33966 22264
rect 34022 22208 41430 22264
rect 33961 22206 41430 22208
rect 33961 22203 34027 22206
rect 11881 22130 11947 22133
rect 19609 22130 19675 22133
rect 11881 22128 19675 22130
rect 11881 22072 11886 22128
rect 11942 22072 19614 22128
rect 19670 22072 19675 22128
rect 11881 22070 19675 22072
rect 11881 22067 11947 22070
rect 19609 22067 19675 22070
rect 21265 22130 21331 22133
rect 24485 22130 24551 22133
rect 21265 22128 24551 22130
rect 21265 22072 21270 22128
rect 21326 22072 24490 22128
rect 24546 22072 24551 22128
rect 21265 22070 24551 22072
rect 21265 22067 21331 22070
rect 24485 22067 24551 22070
rect 37181 22130 37247 22133
rect 38837 22130 38903 22133
rect 37181 22128 38903 22130
rect 37181 22072 37186 22128
rect 37242 22072 38842 22128
rect 38898 22072 38903 22128
rect 37181 22070 38903 22072
rect 41370 22130 41430 22206
rect 49325 22264 51000 22266
rect 49325 22208 49330 22264
rect 49386 22208 51000 22264
rect 49325 22206 51000 22208
rect 49325 22203 49391 22206
rect 50200 22176 51000 22206
rect 44449 22130 44515 22133
rect 45369 22130 45435 22133
rect 41370 22128 45435 22130
rect 41370 22072 44454 22128
rect 44510 22072 45374 22128
rect 45430 22072 45435 22128
rect 41370 22070 45435 22072
rect 37181 22067 37247 22070
rect 38837 22067 38903 22070
rect 44449 22067 44515 22070
rect 45369 22067 45435 22070
rect 0 21994 800 22024
rect 3233 21994 3299 21997
rect 0 21992 3299 21994
rect 0 21936 3238 21992
rect 3294 21936 3299 21992
rect 0 21934 3299 21936
rect 0 21904 800 21934
rect 3233 21931 3299 21934
rect 27613 21994 27679 21997
rect 30189 21994 30255 21997
rect 36629 21994 36695 21997
rect 27613 21992 30255 21994
rect 27613 21936 27618 21992
rect 27674 21936 30194 21992
rect 30250 21936 30255 21992
rect 27613 21934 30255 21936
rect 27613 21931 27679 21934
rect 30189 21931 30255 21934
rect 31710 21992 36695 21994
rect 31710 21936 36634 21992
rect 36690 21936 36695 21992
rect 31710 21934 36695 21936
rect 22277 21858 22343 21861
rect 23105 21858 23171 21861
rect 22277 21856 23171 21858
rect 22277 21800 22282 21856
rect 22338 21800 23110 21856
rect 23166 21800 23171 21856
rect 22277 21798 23171 21800
rect 22277 21795 22343 21798
rect 23105 21795 23171 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 31710 21722 31770 21934
rect 36629 21931 36695 21934
rect 36997 21994 37063 21997
rect 42793 21994 42859 21997
rect 36997 21992 42859 21994
rect 36997 21936 37002 21992
rect 37058 21936 42798 21992
rect 42854 21936 42859 21992
rect 36997 21934 42859 21936
rect 36997 21931 37063 21934
rect 42793 21931 42859 21934
rect 48589 21858 48655 21861
rect 50200 21858 51000 21888
rect 48589 21856 51000 21858
rect 48589 21800 48594 21856
rect 48650 21800 51000 21856
rect 48589 21798 51000 21800
rect 48589 21795 48655 21798
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 50200 21768 51000 21798
rect 47946 21727 48262 21728
rect 28398 21662 31770 21722
rect 34237 21722 34303 21725
rect 36905 21722 36971 21725
rect 34237 21720 36971 21722
rect 34237 21664 34242 21720
rect 34298 21664 36910 21720
rect 36966 21664 36971 21720
rect 34237 21662 36971 21664
rect 0 21586 800 21616
rect 1761 21586 1827 21589
rect 0 21584 1827 21586
rect 0 21528 1766 21584
rect 1822 21528 1827 21584
rect 0 21526 1827 21528
rect 0 21496 800 21526
rect 1761 21523 1827 21526
rect 6545 21586 6611 21589
rect 9029 21586 9095 21589
rect 6545 21584 9095 21586
rect 6545 21528 6550 21584
rect 6606 21528 9034 21584
rect 9090 21528 9095 21584
rect 6545 21526 9095 21528
rect 6545 21523 6611 21526
rect 9029 21523 9095 21526
rect 15561 21586 15627 21589
rect 26049 21586 26115 21589
rect 28398 21586 28458 21662
rect 34237 21659 34303 21662
rect 36905 21659 36971 21662
rect 40309 21722 40375 21725
rect 41873 21722 41939 21725
rect 40309 21720 41939 21722
rect 40309 21664 40314 21720
rect 40370 21664 41878 21720
rect 41934 21664 41939 21720
rect 40309 21662 41939 21664
rect 40309 21659 40375 21662
rect 41873 21659 41939 21662
rect 15561 21584 25882 21586
rect 15561 21528 15566 21584
rect 15622 21528 25882 21584
rect 15561 21526 25882 21528
rect 15561 21523 15627 21526
rect 11697 21450 11763 21453
rect 18597 21450 18663 21453
rect 24945 21450 25011 21453
rect 11697 21448 25011 21450
rect 11697 21392 11702 21448
rect 11758 21392 18602 21448
rect 18658 21392 24950 21448
rect 25006 21392 25011 21448
rect 11697 21390 25011 21392
rect 25822 21450 25882 21526
rect 26049 21584 28458 21586
rect 26049 21528 26054 21584
rect 26110 21528 28458 21584
rect 26049 21526 28458 21528
rect 31201 21586 31267 21589
rect 33501 21586 33567 21589
rect 43897 21586 43963 21589
rect 31201 21584 43963 21586
rect 31201 21528 31206 21584
rect 31262 21528 33506 21584
rect 33562 21528 43902 21584
rect 43958 21528 43963 21584
rect 31201 21526 43963 21528
rect 26049 21523 26115 21526
rect 31201 21523 31267 21526
rect 33501 21523 33567 21526
rect 43897 21523 43963 21526
rect 28809 21450 28875 21453
rect 30373 21450 30439 21453
rect 25822 21448 30439 21450
rect 25822 21392 28814 21448
rect 28870 21392 30378 21448
rect 30434 21392 30439 21448
rect 25822 21390 30439 21392
rect 11697 21387 11763 21390
rect 18597 21387 18663 21390
rect 24945 21387 25011 21390
rect 28809 21387 28875 21390
rect 30373 21387 30439 21390
rect 30741 21450 30807 21453
rect 32857 21450 32923 21453
rect 30741 21448 32923 21450
rect 30741 21392 30746 21448
rect 30802 21392 32862 21448
rect 32918 21392 32923 21448
rect 30741 21390 32923 21392
rect 30741 21387 30807 21390
rect 32857 21387 32923 21390
rect 36445 21450 36511 21453
rect 40677 21450 40743 21453
rect 36445 21448 40743 21450
rect 36445 21392 36450 21448
rect 36506 21392 40682 21448
rect 40738 21392 40743 21448
rect 36445 21390 40743 21392
rect 36445 21387 36511 21390
rect 40677 21387 40743 21390
rect 49233 21450 49299 21453
rect 50200 21450 51000 21480
rect 49233 21448 51000 21450
rect 49233 21392 49238 21448
rect 49294 21392 51000 21448
rect 49233 21390 51000 21392
rect 49233 21387 49299 21390
rect 50200 21360 51000 21390
rect 34421 21314 34487 21317
rect 40861 21314 40927 21317
rect 34421 21312 40927 21314
rect 34421 21256 34426 21312
rect 34482 21256 40866 21312
rect 40922 21256 40927 21312
rect 34421 21254 40927 21256
rect 34421 21251 34487 21254
rect 40861 21251 40927 21254
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 0 21088 800 21118
rect 2773 21115 2839 21118
rect 27797 21178 27863 21181
rect 30005 21178 30071 21181
rect 31385 21178 31451 21181
rect 27797 21176 31451 21178
rect 27797 21120 27802 21176
rect 27858 21120 30010 21176
rect 30066 21120 31390 21176
rect 31446 21120 31451 21176
rect 27797 21118 31451 21120
rect 27797 21115 27863 21118
rect 30005 21115 30071 21118
rect 31385 21115 31451 21118
rect 36629 21178 36695 21181
rect 40217 21178 40283 21181
rect 36629 21176 40283 21178
rect 36629 21120 36634 21176
rect 36690 21120 40222 21176
rect 40278 21120 40283 21176
rect 36629 21118 40283 21120
rect 36629 21115 36695 21118
rect 40217 21115 40283 21118
rect 12617 21042 12683 21045
rect 12893 21042 12959 21045
rect 21909 21042 21975 21045
rect 27429 21042 27495 21045
rect 29637 21042 29703 21045
rect 12617 21040 25882 21042
rect 12617 20984 12622 21040
rect 12678 20984 12898 21040
rect 12954 20984 21914 21040
rect 21970 20984 25882 21040
rect 12617 20982 25882 20984
rect 12617 20979 12683 20982
rect 12893 20979 12959 20982
rect 21909 20979 21975 20982
rect 25822 20909 25882 20982
rect 27429 21040 29703 21042
rect 27429 20984 27434 21040
rect 27490 20984 29642 21040
rect 29698 20984 29703 21040
rect 27429 20982 29703 20984
rect 27429 20979 27495 20982
rect 29637 20979 29703 20982
rect 31753 21042 31819 21045
rect 41229 21042 41295 21045
rect 31753 21040 41295 21042
rect 31753 20984 31758 21040
rect 31814 20984 41234 21040
rect 41290 20984 41295 21040
rect 31753 20982 41295 20984
rect 31753 20979 31819 20982
rect 41229 20979 41295 20982
rect 49325 21042 49391 21045
rect 50200 21042 51000 21072
rect 49325 21040 51000 21042
rect 49325 20984 49330 21040
rect 49386 20984 51000 21040
rect 49325 20982 51000 20984
rect 49325 20979 49391 20982
rect 50200 20952 51000 20982
rect 8385 20906 8451 20909
rect 23749 20906 23815 20909
rect 8385 20904 23815 20906
rect 8385 20848 8390 20904
rect 8446 20848 23754 20904
rect 23810 20848 23815 20904
rect 8385 20846 23815 20848
rect 25822 20906 25931 20909
rect 40401 20906 40467 20909
rect 47669 20906 47735 20909
rect 25822 20904 40467 20906
rect 25822 20848 25870 20904
rect 25926 20848 40406 20904
rect 40462 20848 40467 20904
rect 25822 20846 40467 20848
rect 8385 20843 8451 20846
rect 23749 20843 23815 20846
rect 25865 20843 25931 20846
rect 40401 20843 40467 20846
rect 41370 20904 47735 20906
rect 41370 20848 47674 20904
rect 47730 20848 47735 20904
rect 41370 20846 47735 20848
rect 0 20770 800 20800
rect 1025 20770 1091 20773
rect 0 20768 1091 20770
rect 0 20712 1030 20768
rect 1086 20712 1091 20768
rect 0 20710 1091 20712
rect 0 20680 800 20710
rect 1025 20707 1091 20710
rect 30649 20770 30715 20773
rect 36077 20770 36143 20773
rect 30649 20768 36143 20770
rect 30649 20712 30654 20768
rect 30710 20712 36082 20768
rect 36138 20712 36143 20768
rect 30649 20710 36143 20712
rect 30649 20707 30715 20710
rect 36077 20707 36143 20710
rect 38377 20770 38443 20773
rect 41370 20770 41430 20846
rect 47669 20843 47735 20846
rect 38377 20768 41430 20770
rect 38377 20712 38382 20768
rect 38438 20712 41430 20768
rect 38377 20710 41430 20712
rect 38377 20707 38443 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 10685 20634 10751 20637
rect 14089 20634 14155 20637
rect 10685 20632 14155 20634
rect 10685 20576 10690 20632
rect 10746 20576 14094 20632
rect 14150 20576 14155 20632
rect 10685 20574 14155 20576
rect 10685 20571 10751 20574
rect 14089 20571 14155 20574
rect 30373 20634 30439 20637
rect 37365 20634 37431 20637
rect 30373 20632 37431 20634
rect 30373 20576 30378 20632
rect 30434 20576 37370 20632
rect 37426 20576 37431 20632
rect 30373 20574 37431 20576
rect 30373 20571 30439 20574
rect 37365 20571 37431 20574
rect 49325 20634 49391 20637
rect 50200 20634 51000 20664
rect 49325 20632 51000 20634
rect 49325 20576 49330 20632
rect 49386 20576 51000 20632
rect 49325 20574 51000 20576
rect 49325 20571 49391 20574
rect 50200 20544 51000 20574
rect 34697 20498 34763 20501
rect 49049 20498 49115 20501
rect 34697 20496 49115 20498
rect 34697 20440 34702 20496
rect 34758 20440 49054 20496
rect 49110 20440 49115 20496
rect 34697 20438 49115 20440
rect 34697 20435 34763 20438
rect 49049 20435 49115 20438
rect 0 20362 800 20392
rect 1301 20362 1367 20365
rect 0 20360 1367 20362
rect 0 20304 1306 20360
rect 1362 20304 1367 20360
rect 0 20302 1367 20304
rect 0 20272 800 20302
rect 1301 20299 1367 20302
rect 16205 20362 16271 20365
rect 30097 20362 30163 20365
rect 16205 20360 30163 20362
rect 16205 20304 16210 20360
rect 16266 20304 30102 20360
rect 30158 20304 30163 20360
rect 16205 20302 30163 20304
rect 16205 20299 16271 20302
rect 30097 20299 30163 20302
rect 32765 20362 32831 20365
rect 48405 20362 48471 20365
rect 32765 20360 48471 20362
rect 32765 20304 32770 20360
rect 32826 20304 48410 20360
rect 48466 20304 48471 20360
rect 32765 20302 48471 20304
rect 32765 20299 32831 20302
rect 48405 20299 48471 20302
rect 24485 20226 24551 20229
rect 25221 20226 25287 20229
rect 24485 20224 25287 20226
rect 24485 20168 24490 20224
rect 24546 20168 25226 20224
rect 25282 20168 25287 20224
rect 24485 20166 25287 20168
rect 24485 20163 24551 20166
rect 25221 20163 25287 20166
rect 48773 20226 48839 20229
rect 50200 20226 51000 20256
rect 48773 20224 51000 20226
rect 48773 20168 48778 20224
rect 48834 20168 51000 20224
rect 48773 20166 51000 20168
rect 48773 20163 48839 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 50200 20136 51000 20166
rect 42946 20095 43262 20096
rect 23933 20090 23999 20093
rect 35341 20090 35407 20093
rect 39389 20090 39455 20093
rect 23933 20088 28504 20090
rect 23933 20032 23938 20088
rect 23994 20032 28504 20088
rect 23933 20030 28504 20032
rect 23933 20027 23999 20030
rect 0 19954 800 19984
rect 28444 19957 28504 20030
rect 35341 20088 39455 20090
rect 35341 20032 35346 20088
rect 35402 20032 39394 20088
rect 39450 20032 39455 20088
rect 35341 20030 39455 20032
rect 35341 20027 35407 20030
rect 39389 20027 39455 20030
rect 1761 19954 1827 19957
rect 0 19952 1827 19954
rect 0 19896 1766 19952
rect 1822 19896 1827 19952
rect 0 19894 1827 19896
rect 0 19864 800 19894
rect 1761 19891 1827 19894
rect 15469 19954 15535 19957
rect 26141 19954 26207 19957
rect 15469 19952 26207 19954
rect 15469 19896 15474 19952
rect 15530 19896 26146 19952
rect 26202 19896 26207 19952
rect 15469 19894 26207 19896
rect 15469 19891 15535 19894
rect 26141 19891 26207 19894
rect 26325 19954 26391 19957
rect 27981 19954 28047 19957
rect 26325 19952 28047 19954
rect 26325 19896 26330 19952
rect 26386 19896 27986 19952
rect 28042 19896 28047 19952
rect 26325 19894 28047 19896
rect 26325 19891 26391 19894
rect 27981 19891 28047 19894
rect 28441 19954 28507 19957
rect 48313 19954 48379 19957
rect 28441 19952 48379 19954
rect 28441 19896 28446 19952
rect 28502 19896 48318 19952
rect 48374 19896 48379 19952
rect 28441 19894 48379 19896
rect 28441 19891 28507 19894
rect 48313 19891 48379 19894
rect 12065 19818 12131 19821
rect 22134 19818 22140 19820
rect 12065 19816 22140 19818
rect 12065 19760 12070 19816
rect 12126 19760 22140 19816
rect 12065 19758 22140 19760
rect 12065 19755 12131 19758
rect 22134 19756 22140 19758
rect 22204 19756 22210 19820
rect 31109 19818 31175 19821
rect 26558 19816 31175 19818
rect 26558 19760 31114 19816
rect 31170 19760 31175 19816
rect 26558 19758 31175 19760
rect 10593 19682 10659 19685
rect 15837 19682 15903 19685
rect 10593 19680 15903 19682
rect 10593 19624 10598 19680
rect 10654 19624 15842 19680
rect 15898 19624 15903 19680
rect 10593 19622 15903 19624
rect 22142 19682 22202 19756
rect 25037 19682 25103 19685
rect 26558 19682 26618 19758
rect 31109 19755 31175 19758
rect 34881 19818 34947 19821
rect 44541 19818 44607 19821
rect 34881 19816 44607 19818
rect 34881 19760 34886 19816
rect 34942 19760 44546 19816
rect 44602 19760 44607 19816
rect 34881 19758 44607 19760
rect 34881 19755 34947 19758
rect 44541 19755 44607 19758
rect 49417 19818 49483 19821
rect 50200 19818 51000 19848
rect 49417 19816 51000 19818
rect 49417 19760 49422 19816
rect 49478 19760 51000 19816
rect 49417 19758 51000 19760
rect 49417 19755 49483 19758
rect 50200 19728 51000 19758
rect 22142 19680 26618 19682
rect 22142 19624 25042 19680
rect 25098 19624 26618 19680
rect 22142 19622 26618 19624
rect 28809 19682 28875 19685
rect 33869 19682 33935 19685
rect 28809 19680 33935 19682
rect 28809 19624 28814 19680
rect 28870 19624 33874 19680
rect 33930 19624 33935 19680
rect 28809 19622 33935 19624
rect 10593 19619 10659 19622
rect 15837 19619 15903 19622
rect 25037 19619 25103 19622
rect 28809 19619 28875 19622
rect 33869 19619 33935 19622
rect 7946 19616 8262 19617
rect 0 19546 800 19576
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 2865 19546 2931 19549
rect 0 19544 2931 19546
rect 0 19488 2870 19544
rect 2926 19488 2931 19544
rect 0 19486 2931 19488
rect 0 19456 800 19486
rect 2865 19483 2931 19486
rect 21265 19546 21331 19549
rect 24117 19546 24183 19549
rect 21265 19544 24183 19546
rect 21265 19488 21270 19544
rect 21326 19488 24122 19544
rect 24178 19488 24183 19544
rect 21265 19486 24183 19488
rect 21265 19483 21331 19486
rect 24117 19483 24183 19486
rect 26693 19546 26759 19549
rect 27705 19546 27771 19549
rect 35341 19546 35407 19549
rect 26693 19544 27771 19546
rect 26693 19488 26698 19544
rect 26754 19488 27710 19544
rect 27766 19488 27771 19544
rect 26693 19486 27771 19488
rect 26693 19483 26759 19486
rect 27705 19483 27771 19486
rect 28398 19544 35407 19546
rect 28398 19488 35346 19544
rect 35402 19488 35407 19544
rect 28398 19486 35407 19488
rect 28398 19413 28458 19486
rect 35341 19483 35407 19486
rect 3969 19410 4035 19413
rect 19333 19410 19399 19413
rect 28349 19410 28458 19413
rect 3969 19408 12450 19410
rect 3969 19352 3974 19408
rect 4030 19352 12450 19408
rect 3969 19350 12450 19352
rect 3969 19347 4035 19350
rect 12390 19274 12450 19350
rect 19333 19408 28458 19410
rect 19333 19352 19338 19408
rect 19394 19352 28354 19408
rect 28410 19352 28458 19408
rect 19333 19350 28458 19352
rect 29821 19410 29887 19413
rect 41505 19410 41571 19413
rect 29821 19408 41571 19410
rect 29821 19352 29826 19408
rect 29882 19352 41510 19408
rect 41566 19352 41571 19408
rect 29821 19350 41571 19352
rect 19333 19347 19399 19350
rect 28349 19347 28415 19350
rect 29821 19347 29887 19350
rect 41505 19347 41571 19350
rect 49325 19410 49391 19413
rect 50200 19410 51000 19440
rect 49325 19408 51000 19410
rect 49325 19352 49330 19408
rect 49386 19352 51000 19408
rect 49325 19350 51000 19352
rect 49325 19347 49391 19350
rect 50200 19320 51000 19350
rect 16021 19274 16087 19277
rect 12390 19272 16087 19274
rect 12390 19216 16026 19272
rect 16082 19216 16087 19272
rect 12390 19214 16087 19216
rect 16021 19211 16087 19214
rect 20621 19274 20687 19277
rect 26049 19274 26115 19277
rect 20621 19272 26115 19274
rect 20621 19216 20626 19272
rect 20682 19216 26054 19272
rect 26110 19216 26115 19272
rect 20621 19214 26115 19216
rect 20621 19211 20687 19214
rect 26049 19211 26115 19214
rect 34973 19274 35039 19277
rect 36813 19274 36879 19277
rect 34973 19272 36879 19274
rect 34973 19216 34978 19272
rect 35034 19216 36818 19272
rect 36874 19216 36879 19272
rect 34973 19214 36879 19216
rect 34973 19211 35039 19214
rect 36813 19211 36879 19214
rect 40033 19274 40099 19277
rect 41229 19274 41295 19277
rect 49141 19274 49207 19277
rect 40033 19272 49207 19274
rect 40033 19216 40038 19272
rect 40094 19216 41234 19272
rect 41290 19216 49146 19272
rect 49202 19216 49207 19272
rect 40033 19214 49207 19216
rect 40033 19211 40099 19214
rect 41229 19211 41295 19214
rect 49141 19211 49207 19214
rect 0 19138 800 19168
rect 2773 19138 2839 19141
rect 42793 19138 42859 19141
rect 0 19136 2839 19138
rect 0 19080 2778 19136
rect 2834 19080 2839 19136
rect 0 19078 2839 19080
rect 0 19048 800 19078
rect 2773 19075 2839 19078
rect 33366 19136 42859 19138
rect 33366 19080 42798 19136
rect 42854 19080 42859 19136
rect 33366 19078 42859 19080
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 25589 19002 25655 19005
rect 27521 19002 27587 19005
rect 25589 19000 27587 19002
rect 25589 18944 25594 19000
rect 25650 18944 27526 19000
rect 27582 18944 27587 19000
rect 25589 18942 27587 18944
rect 25589 18939 25655 18942
rect 27521 18939 27587 18942
rect 5349 18866 5415 18869
rect 11237 18866 11303 18869
rect 5349 18864 11303 18866
rect 5349 18808 5354 18864
rect 5410 18808 11242 18864
rect 11298 18808 11303 18864
rect 5349 18806 11303 18808
rect 5349 18803 5415 18806
rect 11237 18803 11303 18806
rect 20345 18866 20411 18869
rect 28993 18866 29059 18869
rect 20345 18864 29059 18866
rect 20345 18808 20350 18864
rect 20406 18808 28998 18864
rect 29054 18808 29059 18864
rect 20345 18806 29059 18808
rect 20345 18803 20411 18806
rect 28993 18803 29059 18806
rect 31293 18866 31359 18869
rect 33366 18866 33426 19078
rect 42793 19075 42859 19078
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 37089 19002 37155 19005
rect 38285 19002 38351 19005
rect 37089 19000 38351 19002
rect 37089 18944 37094 19000
rect 37150 18944 38290 19000
rect 38346 18944 38351 19000
rect 37089 18942 38351 18944
rect 37089 18939 37155 18942
rect 38285 18939 38351 18942
rect 49233 19002 49299 19005
rect 50200 19002 51000 19032
rect 49233 19000 51000 19002
rect 49233 18944 49238 19000
rect 49294 18944 51000 19000
rect 49233 18942 51000 18944
rect 49233 18939 49299 18942
rect 50200 18912 51000 18942
rect 31293 18864 33426 18866
rect 31293 18808 31298 18864
rect 31354 18808 33426 18864
rect 31293 18806 33426 18808
rect 34329 18866 34395 18869
rect 48681 18866 48747 18869
rect 34329 18864 48747 18866
rect 34329 18808 34334 18864
rect 34390 18808 48686 18864
rect 48742 18808 48747 18864
rect 34329 18806 48747 18808
rect 31293 18803 31359 18806
rect 34329 18803 34395 18806
rect 48681 18803 48747 18806
rect 0 18730 800 18760
rect 1485 18730 1551 18733
rect 0 18728 1551 18730
rect 0 18672 1490 18728
rect 1546 18672 1551 18728
rect 0 18670 1551 18672
rect 0 18640 800 18670
rect 1485 18667 1551 18670
rect 14825 18730 14891 18733
rect 16297 18730 16363 18733
rect 14825 18728 16363 18730
rect 14825 18672 14830 18728
rect 14886 18672 16302 18728
rect 16358 18672 16363 18728
rect 14825 18670 16363 18672
rect 14825 18667 14891 18670
rect 16297 18667 16363 18670
rect 17401 18730 17467 18733
rect 19333 18730 19399 18733
rect 28717 18730 28783 18733
rect 17401 18728 28783 18730
rect 17401 18672 17406 18728
rect 17462 18672 19338 18728
rect 19394 18672 28722 18728
rect 28778 18672 28783 18728
rect 17401 18670 28783 18672
rect 17401 18667 17467 18670
rect 19333 18667 19399 18670
rect 28717 18667 28783 18670
rect 30925 18730 30991 18733
rect 40033 18730 40099 18733
rect 30925 18728 40099 18730
rect 30925 18672 30930 18728
rect 30986 18672 40038 18728
rect 40094 18672 40099 18728
rect 30925 18670 40099 18672
rect 30925 18667 30991 18670
rect 40033 18667 40099 18670
rect 21449 18594 21515 18597
rect 23013 18594 23079 18597
rect 21449 18592 23079 18594
rect 21449 18536 21454 18592
rect 21510 18536 23018 18592
rect 23074 18536 23079 18592
rect 21449 18534 23079 18536
rect 21449 18531 21515 18534
rect 23013 18531 23079 18534
rect 30189 18594 30255 18597
rect 36077 18594 36143 18597
rect 30189 18592 36143 18594
rect 30189 18536 30194 18592
rect 30250 18536 36082 18592
rect 36138 18536 36143 18592
rect 30189 18534 36143 18536
rect 30189 18531 30255 18534
rect 36077 18531 36143 18534
rect 48773 18594 48839 18597
rect 50200 18594 51000 18624
rect 48773 18592 51000 18594
rect 48773 18536 48778 18592
rect 48834 18536 51000 18592
rect 48773 18534 51000 18536
rect 48773 18531 48839 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 50200 18504 51000 18534
rect 47946 18463 48262 18464
rect 22369 18458 22435 18461
rect 25589 18458 25655 18461
rect 22369 18456 25655 18458
rect 22369 18400 22374 18456
rect 22430 18400 25594 18456
rect 25650 18400 25655 18456
rect 22369 18398 25655 18400
rect 22369 18395 22435 18398
rect 25589 18395 25655 18398
rect 29637 18458 29703 18461
rect 34605 18458 34671 18461
rect 29637 18456 34671 18458
rect 29637 18400 29642 18456
rect 29698 18400 34610 18456
rect 34666 18400 34671 18456
rect 29637 18398 34671 18400
rect 29637 18395 29703 18398
rect 34605 18395 34671 18398
rect 0 18322 800 18352
rect 1761 18322 1827 18325
rect 0 18320 1827 18322
rect 0 18264 1766 18320
rect 1822 18264 1827 18320
rect 0 18262 1827 18264
rect 0 18232 800 18262
rect 1761 18259 1827 18262
rect 14089 18322 14155 18325
rect 25037 18322 25103 18325
rect 25957 18322 26023 18325
rect 40493 18322 40559 18325
rect 14089 18320 25882 18322
rect 14089 18264 14094 18320
rect 14150 18264 25042 18320
rect 25098 18264 25882 18320
rect 14089 18262 25882 18264
rect 14089 18259 14155 18262
rect 25037 18259 25103 18262
rect 11145 18186 11211 18189
rect 15009 18186 15075 18189
rect 11145 18184 15075 18186
rect 11145 18128 11150 18184
rect 11206 18128 15014 18184
rect 15070 18128 15075 18184
rect 11145 18126 15075 18128
rect 25822 18186 25882 18262
rect 25957 18320 40559 18322
rect 25957 18264 25962 18320
rect 26018 18264 40498 18320
rect 40554 18264 40559 18320
rect 25957 18262 40559 18264
rect 25957 18259 26023 18262
rect 40493 18259 40559 18262
rect 26325 18186 26391 18189
rect 25822 18184 26391 18186
rect 25822 18128 26330 18184
rect 26386 18128 26391 18184
rect 25822 18126 26391 18128
rect 11145 18123 11211 18126
rect 15009 18123 15075 18126
rect 26325 18123 26391 18126
rect 28717 18186 28783 18189
rect 41321 18186 41387 18189
rect 28717 18184 41387 18186
rect 28717 18128 28722 18184
rect 28778 18128 41326 18184
rect 41382 18128 41387 18184
rect 28717 18126 41387 18128
rect 28717 18123 28783 18126
rect 41321 18123 41387 18126
rect 49417 18186 49483 18189
rect 50200 18186 51000 18216
rect 49417 18184 51000 18186
rect 49417 18128 49422 18184
rect 49478 18128 51000 18184
rect 49417 18126 51000 18128
rect 49417 18123 49483 18126
rect 50200 18096 51000 18126
rect 16573 18050 16639 18053
rect 19333 18050 19399 18053
rect 16573 18048 19399 18050
rect 16573 17992 16578 18048
rect 16634 17992 19338 18048
rect 19394 17992 19399 18048
rect 16573 17990 19399 17992
rect 16573 17987 16639 17990
rect 19333 17987 19399 17990
rect 20345 18050 20411 18053
rect 22553 18050 22619 18053
rect 20345 18048 22619 18050
rect 20345 17992 20350 18048
rect 20406 17992 22558 18048
rect 22614 17992 22619 18048
rect 20345 17990 22619 17992
rect 20345 17987 20411 17990
rect 22553 17987 22619 17990
rect 25405 18050 25471 18053
rect 28441 18050 28507 18053
rect 25405 18048 28507 18050
rect 25405 17992 25410 18048
rect 25466 17992 28446 18048
rect 28502 17992 28507 18048
rect 25405 17990 28507 17992
rect 25405 17987 25471 17990
rect 28441 17987 28507 17990
rect 36813 18050 36879 18053
rect 36813 18048 38578 18050
rect 36813 17992 36818 18048
rect 36874 17992 38578 18048
rect 36813 17990 38578 17992
rect 36813 17987 36879 17990
rect 2946 17984 3262 17985
rect 0 17914 800 17944
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 1393 17914 1459 17917
rect 0 17912 1459 17914
rect 0 17856 1398 17912
rect 1454 17856 1459 17912
rect 0 17854 1459 17856
rect 38518 17914 38578 17990
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 40217 17914 40283 17917
rect 38518 17912 40283 17914
rect 38518 17856 40222 17912
rect 40278 17856 40283 17912
rect 38518 17854 40283 17856
rect 0 17824 800 17854
rect 1393 17851 1459 17854
rect 40217 17851 40283 17854
rect 10593 17778 10659 17781
rect 25262 17778 25268 17780
rect 10593 17776 25268 17778
rect 10593 17720 10598 17776
rect 10654 17720 25268 17776
rect 10593 17718 25268 17720
rect 10593 17715 10659 17718
rect 25262 17716 25268 17718
rect 25332 17716 25338 17780
rect 49325 17778 49391 17781
rect 50200 17778 51000 17808
rect 49325 17776 51000 17778
rect 49325 17720 49330 17776
rect 49386 17720 51000 17776
rect 49325 17718 51000 17720
rect 49325 17715 49391 17718
rect 50200 17688 51000 17718
rect 0 17506 800 17536
rect 1761 17506 1827 17509
rect 0 17504 1827 17506
rect 0 17448 1766 17504
rect 1822 17448 1827 17504
rect 0 17446 1827 17448
rect 0 17416 800 17446
rect 1761 17443 1827 17446
rect 29913 17506 29979 17509
rect 30373 17506 30439 17509
rect 35525 17506 35591 17509
rect 29913 17504 35591 17506
rect 29913 17448 29918 17504
rect 29974 17448 30378 17504
rect 30434 17448 35530 17504
rect 35586 17448 35591 17504
rect 29913 17446 35591 17448
rect 29913 17443 29979 17446
rect 30373 17443 30439 17446
rect 35525 17443 35591 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 22461 17370 22527 17373
rect 27705 17370 27771 17373
rect 22461 17368 27771 17370
rect 22461 17312 22466 17368
rect 22522 17312 27710 17368
rect 27766 17312 27771 17368
rect 22461 17310 27771 17312
rect 22461 17307 22527 17310
rect 27705 17307 27771 17310
rect 31385 17370 31451 17373
rect 35341 17370 35407 17373
rect 31385 17368 35407 17370
rect 31385 17312 31390 17368
rect 31446 17312 35346 17368
rect 35402 17312 35407 17368
rect 31385 17310 35407 17312
rect 31385 17307 31451 17310
rect 35341 17307 35407 17310
rect 49325 17370 49391 17373
rect 50200 17370 51000 17400
rect 49325 17368 51000 17370
rect 49325 17312 49330 17368
rect 49386 17312 51000 17368
rect 49325 17310 51000 17312
rect 49325 17307 49391 17310
rect 12249 17234 12315 17237
rect 18965 17234 19031 17237
rect 24761 17234 24827 17237
rect 25773 17234 25839 17237
rect 12249 17232 25839 17234
rect 12249 17176 12254 17232
rect 12310 17176 18970 17232
rect 19026 17176 24766 17232
rect 24822 17176 25778 17232
rect 25834 17176 25839 17232
rect 12249 17174 25839 17176
rect 27708 17234 27768 17307
rect 50200 17280 51000 17310
rect 28257 17234 28323 17237
rect 48497 17234 48563 17237
rect 27708 17232 48563 17234
rect 27708 17176 28262 17232
rect 28318 17176 48502 17232
rect 48558 17176 48563 17232
rect 27708 17174 48563 17176
rect 12249 17171 12315 17174
rect 18965 17171 19031 17174
rect 24761 17171 24827 17174
rect 25773 17171 25839 17174
rect 28257 17171 28323 17174
rect 48497 17171 48563 17174
rect 0 17098 800 17128
rect 933 17098 999 17101
rect 0 17096 999 17098
rect 0 17040 938 17096
rect 994 17040 999 17096
rect 0 17038 999 17040
rect 0 17008 800 17038
rect 933 17035 999 17038
rect 11881 17098 11947 17101
rect 22093 17100 22159 17101
rect 14222 17098 14228 17100
rect 11881 17096 14228 17098
rect 11881 17040 11886 17096
rect 11942 17040 14228 17096
rect 11881 17038 14228 17040
rect 11881 17035 11947 17038
rect 14222 17036 14228 17038
rect 14292 17036 14298 17100
rect 22093 17096 22140 17100
rect 22204 17098 22210 17100
rect 27705 17098 27771 17101
rect 49049 17098 49115 17101
rect 22093 17040 22098 17096
rect 22093 17036 22140 17040
rect 22204 17038 22250 17098
rect 27705 17096 49115 17098
rect 27705 17040 27710 17096
rect 27766 17040 49054 17096
rect 49110 17040 49115 17096
rect 27705 17038 49115 17040
rect 22204 17036 22210 17038
rect 22093 17035 22159 17036
rect 27705 17035 27771 17038
rect 49049 17035 49115 17038
rect 17401 16962 17467 16965
rect 21817 16962 21883 16965
rect 17401 16960 21883 16962
rect 17401 16904 17406 16960
rect 17462 16904 21822 16960
rect 21878 16904 21883 16960
rect 17401 16902 21883 16904
rect 17401 16899 17467 16902
rect 21817 16899 21883 16902
rect 48773 16962 48839 16965
rect 50200 16962 51000 16992
rect 48773 16960 51000 16962
rect 48773 16904 48778 16960
rect 48834 16904 51000 16960
rect 48773 16902 51000 16904
rect 48773 16899 48839 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 50200 16872 51000 16902
rect 42946 16831 43262 16832
rect 23657 16826 23723 16829
rect 24577 16826 24643 16829
rect 25773 16826 25839 16829
rect 26785 16826 26851 16829
rect 27429 16826 27495 16829
rect 27797 16826 27863 16829
rect 23657 16824 27863 16826
rect 23657 16768 23662 16824
rect 23718 16768 24582 16824
rect 24638 16768 25778 16824
rect 25834 16768 26790 16824
rect 26846 16768 27434 16824
rect 27490 16768 27802 16824
rect 27858 16768 27863 16824
rect 23657 16766 27863 16768
rect 23657 16763 23723 16766
rect 24577 16763 24643 16766
rect 25773 16763 25839 16766
rect 26785 16763 26851 16766
rect 27429 16763 27495 16766
rect 27797 16763 27863 16766
rect 0 16690 800 16720
rect 1025 16690 1091 16693
rect 0 16688 1091 16690
rect 0 16632 1030 16688
rect 1086 16632 1091 16688
rect 0 16630 1091 16632
rect 0 16600 800 16630
rect 1025 16627 1091 16630
rect 15101 16692 15167 16693
rect 15101 16688 15148 16692
rect 15212 16690 15218 16692
rect 16297 16690 16363 16693
rect 17493 16690 17559 16693
rect 15101 16632 15106 16688
rect 15101 16628 15148 16632
rect 15212 16630 15258 16690
rect 16297 16688 17559 16690
rect 16297 16632 16302 16688
rect 16358 16632 17498 16688
rect 17554 16632 17559 16688
rect 16297 16630 17559 16632
rect 15212 16628 15218 16630
rect 15101 16627 15167 16628
rect 16297 16627 16363 16630
rect 17493 16627 17559 16630
rect 27981 16690 28047 16693
rect 49141 16690 49207 16693
rect 27981 16688 49207 16690
rect 27981 16632 27986 16688
rect 28042 16632 49146 16688
rect 49202 16632 49207 16688
rect 27981 16630 49207 16632
rect 27981 16627 28047 16630
rect 49141 16627 49207 16630
rect 22461 16554 22527 16557
rect 39757 16554 39823 16557
rect 22461 16552 39823 16554
rect 22461 16496 22466 16552
rect 22522 16496 39762 16552
rect 39818 16496 39823 16552
rect 22461 16494 39823 16496
rect 22461 16491 22527 16494
rect 39757 16491 39823 16494
rect 48221 16554 48287 16557
rect 50200 16554 51000 16584
rect 48221 16552 51000 16554
rect 48221 16496 48226 16552
rect 48282 16496 51000 16552
rect 48221 16494 51000 16496
rect 48221 16491 48287 16494
rect 50200 16464 51000 16494
rect 13537 16418 13603 16421
rect 13997 16418 14063 16421
rect 14825 16418 14891 16421
rect 13537 16416 14891 16418
rect 13537 16360 13542 16416
rect 13598 16360 14002 16416
rect 14058 16360 14830 16416
rect 14886 16360 14891 16416
rect 13537 16358 14891 16360
rect 13537 16355 13603 16358
rect 13997 16355 14063 16358
rect 14825 16355 14891 16358
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 1025 16282 1091 16285
rect 0 16280 1091 16282
rect 0 16224 1030 16280
rect 1086 16224 1091 16280
rect 0 16222 1091 16224
rect 0 16192 800 16222
rect 1025 16219 1091 16222
rect 10501 16146 10567 16149
rect 14181 16146 14247 16149
rect 14549 16146 14615 16149
rect 15837 16146 15903 16149
rect 10501 16144 14106 16146
rect 10501 16088 10506 16144
rect 10562 16088 14106 16144
rect 10501 16086 14106 16088
rect 10501 16083 10567 16086
rect 9581 16010 9647 16013
rect 13537 16010 13603 16013
rect 9581 16008 13603 16010
rect 9581 15952 9586 16008
rect 9642 15952 13542 16008
rect 13598 15952 13603 16008
rect 9581 15950 13603 15952
rect 14046 16010 14106 16086
rect 14181 16144 15903 16146
rect 14181 16088 14186 16144
rect 14242 16088 14554 16144
rect 14610 16088 15842 16144
rect 15898 16088 15903 16144
rect 14181 16086 15903 16088
rect 14181 16083 14247 16086
rect 14549 16083 14615 16086
rect 15837 16083 15903 16086
rect 25681 16146 25747 16149
rect 49141 16146 49207 16149
rect 25681 16144 49207 16146
rect 25681 16088 25686 16144
rect 25742 16088 49146 16144
rect 49202 16088 49207 16144
rect 25681 16086 49207 16088
rect 25681 16083 25747 16086
rect 49141 16083 49207 16086
rect 49417 16146 49483 16149
rect 50200 16146 51000 16176
rect 49417 16144 51000 16146
rect 49417 16088 49422 16144
rect 49478 16088 51000 16144
rect 49417 16086 51000 16088
rect 49417 16083 49483 16086
rect 50200 16056 51000 16086
rect 16021 16010 16087 16013
rect 24853 16010 24919 16013
rect 14046 16008 24919 16010
rect 14046 15952 16026 16008
rect 16082 15952 24858 16008
rect 24914 15952 24919 16008
rect 14046 15950 24919 15952
rect 9581 15947 9647 15950
rect 13537 15947 13603 15950
rect 16021 15947 16087 15950
rect 24853 15947 24919 15950
rect 35801 16010 35867 16013
rect 49141 16010 49207 16013
rect 35801 16008 49207 16010
rect 35801 15952 35806 16008
rect 35862 15952 49146 16008
rect 49202 15952 49207 16008
rect 35801 15950 49207 15952
rect 35801 15947 35867 15950
rect 49141 15947 49207 15950
rect 0 15874 800 15904
rect 1025 15874 1091 15877
rect 0 15872 1091 15874
rect 0 15816 1030 15872
rect 1086 15816 1091 15872
rect 0 15814 1091 15816
rect 0 15784 800 15814
rect 1025 15811 1091 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 20805 15738 20871 15741
rect 22553 15738 22619 15741
rect 29913 15738 29979 15741
rect 20805 15736 22619 15738
rect 20805 15680 20810 15736
rect 20866 15680 22558 15736
rect 22614 15680 22619 15736
rect 20805 15678 22619 15680
rect 20805 15675 20871 15678
rect 22553 15675 22619 15678
rect 26558 15736 29979 15738
rect 26558 15680 29918 15736
rect 29974 15680 29979 15736
rect 26558 15678 29979 15680
rect 17217 15602 17283 15605
rect 19149 15602 19215 15605
rect 21173 15602 21239 15605
rect 17217 15600 21239 15602
rect 17217 15544 17222 15600
rect 17278 15544 19154 15600
rect 19210 15544 21178 15600
rect 21234 15544 21239 15600
rect 17217 15542 21239 15544
rect 17217 15539 17283 15542
rect 19149 15539 19215 15542
rect 21173 15539 21239 15542
rect 0 15466 800 15496
rect 933 15466 999 15469
rect 0 15464 999 15466
rect 0 15408 938 15464
rect 994 15408 999 15464
rect 0 15406 999 15408
rect 0 15376 800 15406
rect 933 15403 999 15406
rect 15837 15466 15903 15469
rect 26558 15466 26618 15678
rect 29913 15675 29979 15678
rect 49325 15738 49391 15741
rect 50200 15738 51000 15768
rect 49325 15736 51000 15738
rect 49325 15680 49330 15736
rect 49386 15680 51000 15736
rect 49325 15678 51000 15680
rect 49325 15675 49391 15678
rect 50200 15648 51000 15678
rect 26785 15602 26851 15605
rect 35617 15602 35683 15605
rect 26785 15600 35683 15602
rect 26785 15544 26790 15600
rect 26846 15544 35622 15600
rect 35678 15544 35683 15600
rect 26785 15542 35683 15544
rect 26785 15539 26851 15542
rect 35617 15539 35683 15542
rect 15837 15464 26618 15466
rect 15837 15408 15842 15464
rect 15898 15408 26618 15464
rect 15837 15406 26618 15408
rect 27061 15466 27127 15469
rect 35433 15466 35499 15469
rect 27061 15464 35499 15466
rect 27061 15408 27066 15464
rect 27122 15408 35438 15464
rect 35494 15408 35499 15464
rect 27061 15406 35499 15408
rect 15837 15403 15903 15406
rect 27061 15403 27127 15406
rect 35433 15403 35499 15406
rect 26049 15330 26115 15333
rect 27153 15330 27219 15333
rect 26049 15328 27219 15330
rect 26049 15272 26054 15328
rect 26110 15272 27158 15328
rect 27214 15272 27219 15328
rect 26049 15270 27219 15272
rect 26049 15267 26115 15270
rect 27153 15267 27219 15270
rect 29177 15330 29243 15333
rect 31201 15330 31267 15333
rect 29177 15328 31267 15330
rect 29177 15272 29182 15328
rect 29238 15272 31206 15328
rect 31262 15272 31267 15328
rect 29177 15270 31267 15272
rect 29177 15267 29243 15270
rect 31201 15267 31267 15270
rect 38377 15330 38443 15333
rect 40125 15330 40191 15333
rect 38377 15328 40191 15330
rect 38377 15272 38382 15328
rect 38438 15272 40130 15328
rect 40186 15272 40191 15328
rect 38377 15270 40191 15272
rect 38377 15267 38443 15270
rect 40125 15267 40191 15270
rect 49325 15330 49391 15333
rect 50200 15330 51000 15360
rect 49325 15328 51000 15330
rect 49325 15272 49330 15328
rect 49386 15272 51000 15328
rect 49325 15270 51000 15272
rect 49325 15267 49391 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 50200 15240 51000 15270
rect 47946 15199 48262 15200
rect 28993 15194 29059 15197
rect 30557 15194 30623 15197
rect 28993 15192 30623 15194
rect 28993 15136 28998 15192
rect 29054 15136 30562 15192
rect 30618 15136 30623 15192
rect 28993 15134 30623 15136
rect 28993 15131 29059 15134
rect 30557 15131 30623 15134
rect 0 15058 800 15088
rect 933 15058 999 15061
rect 0 15056 999 15058
rect 0 15000 938 15056
rect 994 15000 999 15056
rect 0 14998 999 15000
rect 0 14968 800 14998
rect 933 14995 999 14998
rect 14825 15058 14891 15061
rect 18505 15058 18571 15061
rect 14825 15056 18571 15058
rect 14825 15000 14830 15056
rect 14886 15000 18510 15056
rect 18566 15000 18571 15056
rect 14825 14998 18571 15000
rect 14825 14995 14891 14998
rect 18505 14995 18571 14998
rect 27245 15058 27311 15061
rect 49141 15058 49207 15061
rect 27245 15056 49207 15058
rect 27245 15000 27250 15056
rect 27306 15000 49146 15056
rect 49202 15000 49207 15056
rect 27245 14998 49207 15000
rect 27245 14995 27311 14998
rect 49141 14995 49207 14998
rect 12341 14922 12407 14925
rect 18505 14922 18571 14925
rect 12341 14920 18571 14922
rect 12341 14864 12346 14920
rect 12402 14864 18510 14920
rect 18566 14864 18571 14920
rect 12341 14862 18571 14864
rect 12341 14859 12407 14862
rect 18505 14859 18571 14862
rect 30649 14922 30715 14925
rect 31845 14922 31911 14925
rect 30649 14920 31911 14922
rect 30649 14864 30654 14920
rect 30710 14864 31850 14920
rect 31906 14864 31911 14920
rect 30649 14862 31911 14864
rect 30649 14859 30715 14862
rect 31845 14859 31911 14862
rect 35893 14922 35959 14925
rect 39665 14922 39731 14925
rect 35893 14920 39731 14922
rect 35893 14864 35898 14920
rect 35954 14864 39670 14920
rect 39726 14864 39731 14920
rect 35893 14862 39731 14864
rect 35893 14859 35959 14862
rect 39665 14859 39731 14862
rect 49325 14922 49391 14925
rect 50200 14922 51000 14952
rect 49325 14920 51000 14922
rect 49325 14864 49330 14920
rect 49386 14864 51000 14920
rect 49325 14862 51000 14864
rect 49325 14859 49391 14862
rect 50200 14832 51000 14862
rect 2946 14720 3262 14721
rect 0 14650 800 14680
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 933 14650 999 14653
rect 0 14648 999 14650
rect 0 14592 938 14648
rect 994 14592 999 14648
rect 0 14590 999 14592
rect 0 14560 800 14590
rect 933 14587 999 14590
rect 10409 14514 10475 14517
rect 21449 14514 21515 14517
rect 35801 14514 35867 14517
rect 10409 14512 35867 14514
rect 10409 14456 10414 14512
rect 10470 14456 21454 14512
rect 21510 14456 35806 14512
rect 35862 14456 35867 14512
rect 10409 14454 35867 14456
rect 10409 14451 10475 14454
rect 21449 14451 21515 14454
rect 35801 14451 35867 14454
rect 49233 14514 49299 14517
rect 50200 14514 51000 14544
rect 49233 14512 51000 14514
rect 49233 14456 49238 14512
rect 49294 14456 51000 14512
rect 49233 14454 51000 14456
rect 49233 14451 49299 14454
rect 50200 14424 51000 14454
rect 20069 14378 20135 14381
rect 21633 14378 21699 14381
rect 49049 14378 49115 14381
rect 20069 14376 49115 14378
rect 20069 14320 20074 14376
rect 20130 14320 21638 14376
rect 21694 14320 49054 14376
rect 49110 14320 49115 14376
rect 20069 14318 49115 14320
rect 20069 14315 20135 14318
rect 21633 14315 21699 14318
rect 49049 14315 49115 14318
rect 0 14242 800 14272
rect 1025 14242 1091 14245
rect 0 14240 1091 14242
rect 0 14184 1030 14240
rect 1086 14184 1091 14240
rect 0 14182 1091 14184
rect 0 14152 800 14182
rect 1025 14179 1091 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 49233 14106 49299 14109
rect 50200 14106 51000 14136
rect 49233 14104 51000 14106
rect 49233 14048 49238 14104
rect 49294 14048 51000 14104
rect 49233 14046 51000 14048
rect 49233 14043 49299 14046
rect 50200 14016 51000 14046
rect 0 13834 800 13864
rect 1761 13834 1827 13837
rect 0 13832 1827 13834
rect 0 13776 1766 13832
rect 1822 13776 1827 13832
rect 0 13774 1827 13776
rect 0 13744 800 13774
rect 1761 13771 1827 13774
rect 11237 13834 11303 13837
rect 20069 13834 20135 13837
rect 11237 13832 20135 13834
rect 11237 13776 11242 13832
rect 11298 13776 20074 13832
rect 20130 13776 20135 13832
rect 11237 13774 20135 13776
rect 11237 13771 11303 13774
rect 20069 13771 20135 13774
rect 30557 13834 30623 13837
rect 34329 13834 34395 13837
rect 30557 13832 34395 13834
rect 30557 13776 30562 13832
rect 30618 13776 34334 13832
rect 34390 13776 34395 13832
rect 30557 13774 34395 13776
rect 30557 13771 30623 13774
rect 34329 13771 34395 13774
rect 15142 13636 15148 13700
rect 15212 13698 15218 13700
rect 16481 13698 16547 13701
rect 15212 13696 16547 13698
rect 15212 13640 16486 13696
rect 16542 13640 16547 13696
rect 15212 13638 16547 13640
rect 15212 13636 15218 13638
rect 16481 13635 16547 13638
rect 35617 13698 35683 13701
rect 36721 13698 36787 13701
rect 35617 13696 36787 13698
rect 35617 13640 35622 13696
rect 35678 13640 36726 13696
rect 36782 13640 36787 13696
rect 35617 13638 36787 13640
rect 35617 13635 35683 13638
rect 36721 13635 36787 13638
rect 48221 13698 48287 13701
rect 50200 13698 51000 13728
rect 48221 13696 51000 13698
rect 48221 13640 48226 13696
rect 48282 13640 51000 13696
rect 48221 13638 51000 13640
rect 48221 13635 48287 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 50200 13608 51000 13638
rect 42946 13567 43262 13568
rect 0 13426 800 13456
rect 3509 13426 3575 13429
rect 0 13424 3575 13426
rect 0 13368 3514 13424
rect 3570 13368 3575 13424
rect 0 13366 3575 13368
rect 0 13336 800 13366
rect 3509 13363 3575 13366
rect 14549 13426 14615 13429
rect 24669 13426 24735 13429
rect 14549 13424 24735 13426
rect 14549 13368 14554 13424
rect 14610 13368 24674 13424
rect 24730 13368 24735 13424
rect 14549 13366 24735 13368
rect 14549 13363 14615 13366
rect 24669 13363 24735 13366
rect 18505 13290 18571 13293
rect 19241 13290 19307 13293
rect 30557 13290 30623 13293
rect 35157 13290 35223 13293
rect 18505 13288 35223 13290
rect 18505 13232 18510 13288
rect 18566 13232 19246 13288
rect 19302 13232 30562 13288
rect 30618 13232 35162 13288
rect 35218 13232 35223 13288
rect 18505 13230 35223 13232
rect 18505 13227 18571 13230
rect 19241 13227 19307 13230
rect 30557 13227 30623 13230
rect 35157 13227 35223 13230
rect 49141 13290 49207 13293
rect 50200 13290 51000 13320
rect 49141 13288 51000 13290
rect 49141 13232 49146 13288
rect 49202 13232 51000 13288
rect 49141 13230 51000 13232
rect 49141 13227 49207 13230
rect 50200 13200 51000 13230
rect 11145 13154 11211 13157
rect 14549 13154 14615 13157
rect 11145 13152 14615 13154
rect 11145 13096 11150 13152
rect 11206 13096 14554 13152
rect 14610 13096 14615 13152
rect 11145 13094 14615 13096
rect 11145 13091 11211 13094
rect 14549 13091 14615 13094
rect 21449 13154 21515 13157
rect 26049 13154 26115 13157
rect 21449 13152 26115 13154
rect 21449 13096 21454 13152
rect 21510 13096 26054 13152
rect 26110 13096 26115 13152
rect 21449 13094 26115 13096
rect 21449 13091 21515 13094
rect 26049 13091 26115 13094
rect 7946 13088 8262 13089
rect 0 13018 800 13048
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 1301 13018 1367 13021
rect 0 13016 1367 13018
rect 0 12960 1306 13016
rect 1362 12960 1367 13016
rect 0 12958 1367 12960
rect 0 12928 800 12958
rect 1301 12955 1367 12958
rect 14825 13018 14891 13021
rect 15285 13018 15351 13021
rect 17401 13018 17467 13021
rect 14825 13016 17467 13018
rect 14825 12960 14830 13016
rect 14886 12960 15290 13016
rect 15346 12960 17406 13016
rect 17462 12960 17467 13016
rect 14825 12958 17467 12960
rect 14825 12955 14891 12958
rect 15285 12955 15351 12958
rect 17401 12955 17467 12958
rect 22093 13018 22159 13021
rect 22921 13018 22987 13021
rect 26233 13018 26299 13021
rect 22093 13016 26299 13018
rect 22093 12960 22098 13016
rect 22154 12960 22926 13016
rect 22982 12960 26238 13016
rect 26294 12960 26299 13016
rect 22093 12958 26299 12960
rect 22093 12955 22159 12958
rect 22921 12955 22987 12958
rect 26233 12955 26299 12958
rect 22737 12882 22803 12885
rect 26417 12882 26483 12885
rect 22737 12880 26483 12882
rect 22737 12824 22742 12880
rect 22798 12824 26422 12880
rect 26478 12824 26483 12880
rect 22737 12822 26483 12824
rect 22737 12819 22803 12822
rect 26417 12819 26483 12822
rect 28441 12882 28507 12885
rect 40033 12882 40099 12885
rect 28441 12880 40099 12882
rect 28441 12824 28446 12880
rect 28502 12824 40038 12880
rect 40094 12824 40099 12880
rect 28441 12822 40099 12824
rect 28441 12819 28507 12822
rect 40033 12819 40099 12822
rect 49141 12882 49207 12885
rect 50200 12882 51000 12912
rect 49141 12880 51000 12882
rect 49141 12824 49146 12880
rect 49202 12824 51000 12880
rect 49141 12822 51000 12824
rect 49141 12819 49207 12822
rect 50200 12792 51000 12822
rect 12157 12746 12223 12749
rect 16297 12746 16363 12749
rect 12157 12744 16363 12746
rect 12157 12688 12162 12744
rect 12218 12688 16302 12744
rect 16358 12688 16363 12744
rect 12157 12686 16363 12688
rect 12157 12683 12223 12686
rect 16297 12683 16363 12686
rect 23013 12746 23079 12749
rect 25957 12746 26023 12749
rect 23013 12744 26023 12746
rect 23013 12688 23018 12744
rect 23074 12688 25962 12744
rect 26018 12688 26023 12744
rect 23013 12686 26023 12688
rect 23013 12683 23079 12686
rect 25957 12683 26023 12686
rect 0 12610 800 12640
rect 1209 12610 1275 12613
rect 0 12608 1275 12610
rect 0 12552 1214 12608
rect 1270 12552 1275 12608
rect 0 12550 1275 12552
rect 0 12520 800 12550
rect 1209 12547 1275 12550
rect 13353 12610 13419 12613
rect 13721 12610 13787 12613
rect 13353 12608 13787 12610
rect 13353 12552 13358 12608
rect 13414 12552 13726 12608
rect 13782 12552 13787 12608
rect 13353 12550 13787 12552
rect 13353 12547 13419 12550
rect 13721 12547 13787 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 14222 12412 14228 12476
rect 14292 12474 14298 12476
rect 16205 12474 16271 12477
rect 14292 12472 16271 12474
rect 14292 12416 16210 12472
rect 16266 12416 16271 12472
rect 14292 12414 16271 12416
rect 14292 12412 14298 12414
rect 16205 12411 16271 12414
rect 49141 12474 49207 12477
rect 50200 12474 51000 12504
rect 49141 12472 51000 12474
rect 49141 12416 49146 12472
rect 49202 12416 51000 12472
rect 49141 12414 51000 12416
rect 49141 12411 49207 12414
rect 50200 12384 51000 12414
rect 17217 12338 17283 12341
rect 22553 12338 22619 12341
rect 29729 12338 29795 12341
rect 17217 12336 29795 12338
rect 17217 12280 17222 12336
rect 17278 12280 22558 12336
rect 22614 12280 29734 12336
rect 29790 12280 29795 12336
rect 17217 12278 29795 12280
rect 17217 12275 17283 12278
rect 22553 12275 22619 12278
rect 29729 12275 29795 12278
rect 0 12202 800 12232
rect 1209 12202 1275 12205
rect 0 12200 1275 12202
rect 0 12144 1214 12200
rect 1270 12144 1275 12200
rect 0 12142 1275 12144
rect 0 12112 800 12142
rect 1209 12139 1275 12142
rect 12433 12202 12499 12205
rect 15837 12202 15903 12205
rect 16757 12202 16823 12205
rect 12433 12200 16823 12202
rect 12433 12144 12438 12200
rect 12494 12144 15842 12200
rect 15898 12144 16762 12200
rect 16818 12144 16823 12200
rect 12433 12142 16823 12144
rect 12433 12139 12499 12142
rect 15837 12139 15903 12142
rect 16757 12139 16823 12142
rect 29637 12202 29703 12205
rect 40125 12202 40191 12205
rect 29637 12200 40191 12202
rect 29637 12144 29642 12200
rect 29698 12144 40130 12200
rect 40186 12144 40191 12200
rect 29637 12142 40191 12144
rect 29637 12139 29703 12142
rect 40125 12139 40191 12142
rect 13353 12066 13419 12069
rect 17217 12066 17283 12069
rect 13353 12064 17283 12066
rect 13353 12008 13358 12064
rect 13414 12008 17222 12064
rect 17278 12008 17283 12064
rect 13353 12006 17283 12008
rect 13353 12003 13419 12006
rect 17217 12003 17283 12006
rect 49141 12066 49207 12069
rect 50200 12066 51000 12096
rect 49141 12064 51000 12066
rect 49141 12008 49146 12064
rect 49202 12008 51000 12064
rect 49141 12006 51000 12008
rect 49141 12003 49207 12006
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 50200 11976 51000 12006
rect 47946 11935 48262 11936
rect 0 11794 800 11824
rect 1301 11794 1367 11797
rect 0 11792 1367 11794
rect 0 11736 1306 11792
rect 1362 11736 1367 11792
rect 0 11734 1367 11736
rect 0 11704 800 11734
rect 1301 11731 1367 11734
rect 2681 11794 2747 11797
rect 16941 11794 17007 11797
rect 2681 11792 17007 11794
rect 2681 11736 2686 11792
rect 2742 11736 16946 11792
rect 17002 11736 17007 11792
rect 2681 11734 17007 11736
rect 2681 11731 2747 11734
rect 16941 11731 17007 11734
rect 20621 11794 20687 11797
rect 24853 11794 24919 11797
rect 20621 11792 24919 11794
rect 20621 11736 20626 11792
rect 20682 11736 24858 11792
rect 24914 11736 24919 11792
rect 20621 11734 24919 11736
rect 20621 11731 20687 11734
rect 24853 11731 24919 11734
rect 49141 11658 49207 11661
rect 50200 11658 51000 11688
rect 49141 11656 51000 11658
rect 49141 11600 49146 11656
rect 49202 11600 51000 11656
rect 49141 11598 51000 11600
rect 49141 11595 49207 11598
rect 50200 11568 51000 11598
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 1301 11386 1367 11389
rect 0 11384 1367 11386
rect 0 11328 1306 11384
rect 1362 11328 1367 11384
rect 0 11326 1367 11328
rect 0 11296 800 11326
rect 1301 11323 1367 11326
rect 49233 11250 49299 11253
rect 50200 11250 51000 11280
rect 49233 11248 51000 11250
rect 49233 11192 49238 11248
rect 49294 11192 51000 11248
rect 49233 11190 51000 11192
rect 49233 11187 49299 11190
rect 50200 11160 51000 11190
rect 24025 11114 24091 11117
rect 28625 11114 28691 11117
rect 24025 11112 28691 11114
rect 24025 11056 24030 11112
rect 24086 11056 28630 11112
rect 28686 11056 28691 11112
rect 24025 11054 28691 11056
rect 24025 11051 24091 11054
rect 28625 11051 28691 11054
rect 30005 11114 30071 11117
rect 38009 11114 38075 11117
rect 30005 11112 38075 11114
rect 30005 11056 30010 11112
rect 30066 11056 38014 11112
rect 38070 11056 38075 11112
rect 30005 11054 38075 11056
rect 30005 11051 30071 11054
rect 38009 11051 38075 11054
rect 0 10978 800 11008
rect 1577 10978 1643 10981
rect 0 10976 1643 10978
rect 0 10920 1582 10976
rect 1638 10920 1643 10976
rect 0 10918 1643 10920
rect 0 10888 800 10918
rect 1577 10915 1643 10918
rect 13445 10978 13511 10981
rect 14825 10978 14891 10981
rect 16021 10978 16087 10981
rect 13445 10976 16087 10978
rect 13445 10920 13450 10976
rect 13506 10920 14830 10976
rect 14886 10920 16026 10976
rect 16082 10920 16087 10976
rect 13445 10918 16087 10920
rect 13445 10915 13511 10918
rect 14825 10915 14891 10918
rect 16021 10915 16087 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 49141 10842 49207 10845
rect 50200 10842 51000 10872
rect 49141 10840 51000 10842
rect 49141 10784 49146 10840
rect 49202 10784 51000 10840
rect 49141 10782 51000 10784
rect 49141 10779 49207 10782
rect 50200 10752 51000 10782
rect 0 10570 800 10600
rect 1301 10570 1367 10573
rect 0 10568 1367 10570
rect 0 10512 1306 10568
rect 1362 10512 1367 10568
rect 0 10510 1367 10512
rect 0 10480 800 10510
rect 1301 10507 1367 10510
rect 13445 10570 13511 10573
rect 35157 10570 35223 10573
rect 13445 10568 35223 10570
rect 13445 10512 13450 10568
rect 13506 10512 35162 10568
rect 35218 10512 35223 10568
rect 13445 10510 35223 10512
rect 13445 10507 13511 10510
rect 35157 10507 35223 10510
rect 49233 10434 49299 10437
rect 50200 10434 51000 10464
rect 49233 10432 51000 10434
rect 49233 10376 49238 10432
rect 49294 10376 51000 10432
rect 49233 10374 51000 10376
rect 49233 10371 49299 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 50200 10344 51000 10374
rect 42946 10303 43262 10304
rect 0 10162 800 10192
rect 1209 10162 1275 10165
rect 0 10160 1275 10162
rect 0 10104 1214 10160
rect 1270 10104 1275 10160
rect 0 10102 1275 10104
rect 0 10072 800 10102
rect 1209 10099 1275 10102
rect 21357 10162 21423 10165
rect 26233 10162 26299 10165
rect 27245 10162 27311 10165
rect 21357 10160 27311 10162
rect 21357 10104 21362 10160
rect 21418 10104 26238 10160
rect 26294 10104 27250 10160
rect 27306 10104 27311 10160
rect 21357 10102 27311 10104
rect 21357 10099 21423 10102
rect 26233 10099 26299 10102
rect 27245 10099 27311 10102
rect 49325 10026 49391 10029
rect 50200 10026 51000 10056
rect 49325 10024 51000 10026
rect 49325 9968 49330 10024
rect 49386 9968 51000 10024
rect 49325 9966 51000 9968
rect 49325 9963 49391 9966
rect 50200 9936 51000 9966
rect 7946 9824 8262 9825
rect 0 9754 800 9784
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 1301 9754 1367 9757
rect 0 9752 1367 9754
rect 0 9696 1306 9752
rect 1362 9696 1367 9752
rect 0 9694 1367 9696
rect 0 9664 800 9694
rect 1301 9691 1367 9694
rect 47301 9618 47367 9621
rect 50200 9618 51000 9648
rect 47301 9616 51000 9618
rect 47301 9560 47306 9616
rect 47362 9560 51000 9616
rect 47301 9558 51000 9560
rect 47301 9555 47367 9558
rect 50200 9528 51000 9558
rect 1761 9482 1827 9485
rect 34237 9482 34303 9485
rect 1761 9480 34303 9482
rect 1761 9424 1766 9480
rect 1822 9424 34242 9480
rect 34298 9424 34303 9480
rect 1761 9422 34303 9424
rect 1761 9419 1827 9422
rect 34237 9419 34303 9422
rect 0 9346 800 9376
rect 1301 9346 1367 9349
rect 0 9344 1367 9346
rect 0 9288 1306 9344
rect 1362 9288 1367 9344
rect 0 9286 1367 9288
rect 0 9256 800 9286
rect 1301 9283 1367 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 49141 9210 49207 9213
rect 50200 9210 51000 9240
rect 49141 9208 51000 9210
rect 49141 9152 49146 9208
rect 49202 9152 51000 9208
rect 49141 9150 51000 9152
rect 49141 9147 49207 9150
rect 50200 9120 51000 9150
rect 30833 9074 30899 9077
rect 36261 9074 36327 9077
rect 30833 9072 36327 9074
rect 30833 9016 30838 9072
rect 30894 9016 36266 9072
rect 36322 9016 36327 9072
rect 30833 9014 36327 9016
rect 30833 9011 30899 9014
rect 36261 9011 36327 9014
rect 0 8938 800 8968
rect 1301 8938 1367 8941
rect 0 8936 1367 8938
rect 0 8880 1306 8936
rect 1362 8880 1367 8936
rect 0 8878 1367 8880
rect 0 8848 800 8878
rect 1301 8875 1367 8878
rect 49233 8802 49299 8805
rect 50200 8802 51000 8832
rect 49233 8800 51000 8802
rect 49233 8744 49238 8800
rect 49294 8744 51000 8800
rect 49233 8742 51000 8744
rect 49233 8739 49299 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 50200 8712 51000 8742
rect 47946 8671 48262 8672
rect 0 8530 800 8560
rect 1209 8530 1275 8533
rect 0 8528 1275 8530
rect 0 8472 1214 8528
rect 1270 8472 1275 8528
rect 0 8470 1275 8472
rect 0 8440 800 8470
rect 1209 8467 1275 8470
rect 49325 8394 49391 8397
rect 50200 8394 51000 8424
rect 49325 8392 51000 8394
rect 49325 8336 49330 8392
rect 49386 8336 51000 8392
rect 49325 8334 51000 8336
rect 49325 8331 49391 8334
rect 50200 8304 51000 8334
rect 2946 8192 3262 8193
rect 0 8122 800 8152
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 1301 8122 1367 8125
rect 0 8120 1367 8122
rect 0 8064 1306 8120
rect 1362 8064 1367 8120
rect 0 8062 1367 8064
rect 0 8032 800 8062
rect 1301 8059 1367 8062
rect 46841 7986 46907 7989
rect 50200 7986 51000 8016
rect 46841 7984 51000 7986
rect 46841 7928 46846 7984
rect 46902 7928 51000 7984
rect 46841 7926 51000 7928
rect 46841 7923 46907 7926
rect 50200 7896 51000 7926
rect 0 7714 800 7744
rect 1301 7714 1367 7717
rect 0 7712 1367 7714
rect 0 7656 1306 7712
rect 1362 7656 1367 7712
rect 0 7654 1367 7656
rect 0 7624 800 7654
rect 1301 7651 1367 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 49141 7578 49207 7581
rect 50200 7578 51000 7608
rect 49141 7576 51000 7578
rect 49141 7520 49146 7576
rect 49202 7520 51000 7576
rect 49141 7518 51000 7520
rect 49141 7515 49207 7518
rect 50200 7488 51000 7518
rect 0 7306 800 7336
rect 1301 7306 1367 7309
rect 0 7304 1367 7306
rect 0 7248 1306 7304
rect 1362 7248 1367 7304
rect 0 7246 1367 7248
rect 0 7216 800 7246
rect 1301 7243 1367 7246
rect 49325 7170 49391 7173
rect 50200 7170 51000 7200
rect 49325 7168 51000 7170
rect 49325 7112 49330 7168
rect 49386 7112 51000 7168
rect 49325 7110 51000 7112
rect 49325 7107 49391 7110
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 50200 7080 51000 7110
rect 42946 7039 43262 7040
rect 0 6898 800 6928
rect 1209 6898 1275 6901
rect 0 6896 1275 6898
rect 0 6840 1214 6896
rect 1270 6840 1275 6896
rect 0 6838 1275 6840
rect 0 6808 800 6838
rect 1209 6835 1275 6838
rect 49233 6762 49299 6765
rect 50200 6762 51000 6792
rect 49233 6760 51000 6762
rect 49233 6704 49238 6760
rect 49294 6704 51000 6760
rect 49233 6702 51000 6704
rect 49233 6699 49299 6702
rect 50200 6672 51000 6702
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 1301 6490 1367 6493
rect 0 6488 1367 6490
rect 0 6432 1306 6488
rect 1362 6432 1367 6488
rect 0 6430 1367 6432
rect 0 6400 800 6430
rect 1301 6427 1367 6430
rect 48681 6354 48747 6357
rect 50200 6354 51000 6384
rect 48681 6352 51000 6354
rect 48681 6296 48686 6352
rect 48742 6296 51000 6352
rect 48681 6294 51000 6296
rect 48681 6291 48747 6294
rect 50200 6264 51000 6294
rect 0 6082 800 6112
rect 1301 6082 1367 6085
rect 0 6080 1367 6082
rect 0 6024 1306 6080
rect 1362 6024 1367 6080
rect 0 6022 1367 6024
rect 0 5992 800 6022
rect 1301 6019 1367 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 49141 5946 49207 5949
rect 50200 5946 51000 5976
rect 49141 5944 51000 5946
rect 49141 5888 49146 5944
rect 49202 5888 51000 5944
rect 49141 5886 51000 5888
rect 49141 5883 49207 5886
rect 50200 5856 51000 5886
rect 0 5674 800 5704
rect 1301 5674 1367 5677
rect 0 5672 1367 5674
rect 0 5616 1306 5672
rect 1362 5616 1367 5672
rect 0 5614 1367 5616
rect 0 5584 800 5614
rect 1301 5611 1367 5614
rect 49417 5538 49483 5541
rect 50200 5538 51000 5568
rect 49417 5536 51000 5538
rect 49417 5480 49422 5536
rect 49478 5480 51000 5536
rect 49417 5478 51000 5480
rect 49417 5475 49483 5478
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 50200 5448 51000 5478
rect 47946 5407 48262 5408
rect 0 5266 800 5296
rect 2773 5266 2839 5269
rect 0 5264 2839 5266
rect 0 5208 2778 5264
rect 2834 5208 2839 5264
rect 0 5206 2839 5208
rect 0 5176 800 5206
rect 2773 5203 2839 5206
rect 49325 5130 49391 5133
rect 50200 5130 51000 5160
rect 49325 5128 51000 5130
rect 49325 5072 49330 5128
rect 49386 5072 51000 5128
rect 49325 5070 51000 5072
rect 49325 5067 49391 5070
rect 50200 5040 51000 5070
rect 2946 4928 3262 4929
rect 0 4858 800 4888
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 48313 4722 48379 4725
rect 50200 4722 51000 4752
rect 48313 4720 51000 4722
rect 48313 4664 48318 4720
rect 48374 4664 51000 4720
rect 48313 4662 51000 4664
rect 48313 4659 48379 4662
rect 50200 4632 51000 4662
rect 0 4450 800 4480
rect 1301 4450 1367 4453
rect 0 4448 1367 4450
rect 0 4392 1306 4448
rect 1362 4392 1367 4448
rect 0 4390 1367 4392
rect 0 4360 800 4390
rect 1301 4387 1367 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 49141 4314 49207 4317
rect 50200 4314 51000 4344
rect 49141 4312 51000 4314
rect 49141 4256 49146 4312
rect 49202 4256 51000 4312
rect 49141 4254 51000 4256
rect 49141 4251 49207 4254
rect 50200 4224 51000 4254
rect 0 4042 800 4072
rect 1393 4042 1459 4045
rect 0 4040 1459 4042
rect 0 3984 1398 4040
rect 1454 3984 1459 4040
rect 0 3982 1459 3984
rect 0 3952 800 3982
rect 1393 3979 1459 3982
rect 5349 4042 5415 4045
rect 24853 4042 24919 4045
rect 5349 4040 24919 4042
rect 5349 3984 5354 4040
rect 5410 3984 24858 4040
rect 24914 3984 24919 4040
rect 5349 3982 24919 3984
rect 5349 3979 5415 3982
rect 24853 3979 24919 3982
rect 49233 3906 49299 3909
rect 50200 3906 51000 3936
rect 49233 3904 51000 3906
rect 49233 3848 49238 3904
rect 49294 3848 51000 3904
rect 49233 3846 51000 3848
rect 49233 3843 49299 3846
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 50200 3816 51000 3846
rect 42946 3775 43262 3776
rect 0 3634 800 3664
rect 1301 3634 1367 3637
rect 0 3632 1367 3634
rect 0 3576 1306 3632
rect 1362 3576 1367 3632
rect 0 3574 1367 3576
rect 0 3544 800 3574
rect 1301 3571 1367 3574
rect 1117 3498 1183 3501
rect 25773 3498 25839 3501
rect 1117 3496 25839 3498
rect 1117 3440 1122 3496
rect 1178 3440 25778 3496
rect 25834 3440 25839 3496
rect 1117 3438 25839 3440
rect 1117 3435 1183 3438
rect 25773 3435 25839 3438
rect 49141 3498 49207 3501
rect 50200 3498 51000 3528
rect 49141 3496 51000 3498
rect 49141 3440 49146 3496
rect 49202 3440 51000 3496
rect 49141 3438 51000 3440
rect 49141 3435 49207 3438
rect 50200 3408 51000 3438
rect 7946 3296 8262 3297
rect 0 3226 800 3256
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 1301 3226 1367 3229
rect 0 3224 1367 3226
rect 0 3168 1306 3224
rect 1362 3168 1367 3224
rect 0 3166 1367 3168
rect 0 3136 800 3166
rect 1301 3163 1367 3166
rect 48681 3090 48747 3093
rect 50200 3090 51000 3120
rect 48681 3088 51000 3090
rect 48681 3032 48686 3088
rect 48742 3032 51000 3088
rect 48681 3030 51000 3032
rect 48681 3027 48747 3030
rect 50200 3000 51000 3030
rect 0 2818 800 2848
rect 1301 2818 1367 2821
rect 0 2816 1367 2818
rect 0 2760 1306 2816
rect 1362 2760 1367 2816
rect 0 2758 1367 2760
rect 0 2728 800 2758
rect 1301 2755 1367 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 46841 2682 46907 2685
rect 50200 2682 51000 2712
rect 46841 2680 51000 2682
rect 46841 2624 46846 2680
rect 46902 2624 51000 2680
rect 46841 2622 51000 2624
rect 46841 2619 46907 2622
rect 50200 2592 51000 2622
rect 0 2410 800 2440
rect 1301 2410 1367 2413
rect 0 2408 1367 2410
rect 0 2352 1306 2408
rect 1362 2352 1367 2408
rect 0 2350 1367 2352
rect 0 2320 800 2350
rect 1301 2347 1367 2350
rect 48497 2274 48563 2277
rect 50200 2274 51000 2304
rect 48497 2272 51000 2274
rect 48497 2216 48502 2272
rect 48558 2216 51000 2272
rect 48497 2214 51000 2216
rect 48497 2211 48563 2214
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 50200 2184 51000 2214
rect 47946 2143 48262 2144
rect 0 2002 800 2032
rect 1209 2002 1275 2005
rect 0 2000 1275 2002
rect 0 1944 1214 2000
rect 1270 1944 1275 2000
rect 0 1942 1275 1944
rect 0 1912 800 1942
rect 1209 1939 1275 1942
rect 46749 1866 46815 1869
rect 50200 1866 51000 1896
rect 46749 1864 51000 1866
rect 46749 1808 46754 1864
rect 46810 1808 51000 1864
rect 46749 1806 51000 1808
rect 46749 1803 46815 1806
rect 50200 1776 51000 1806
rect 0 1594 800 1624
rect 1301 1594 1367 1597
rect 0 1592 1367 1594
rect 0 1536 1306 1592
rect 1362 1536 1367 1592
rect 0 1534 1367 1536
rect 0 1504 800 1534
rect 1301 1531 1367 1534
rect 46657 1458 46723 1461
rect 50200 1458 51000 1488
rect 46657 1456 51000 1458
rect 46657 1400 46662 1456
rect 46718 1400 51000 1456
rect 46657 1398 51000 1400
rect 46657 1395 46723 1398
rect 50200 1368 51000 1398
<< via3 >>
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 25268 22944 25332 22948
rect 25268 22888 25318 22944
rect 25318 22888 25332 22944
rect 25268 22884 25332 22888
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 22140 19756 22204 19820
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 25268 17716 25332 17780
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 14228 17036 14292 17100
rect 22140 17096 22204 17100
rect 22140 17040 22154 17096
rect 22154 17040 22204 17096
rect 22140 17036 22204 17040
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 15148 16688 15212 16692
rect 15148 16632 15162 16688
rect 15162 16632 15212 16688
rect 15148 16628 15212 16632
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 15148 13636 15212 13700
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 14228 12412 14292 12476
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 17944 23968 18264 24528
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 27944 23968 28264 24528
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 25267 22948 25333 22949
rect 25267 22884 25268 22948
rect 25332 22884 25333 22948
rect 25267 22883 25333 22884
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22139 19820 22205 19821
rect 22139 19756 22140 19820
rect 22204 19756 22205 19820
rect 22139 19755 22205 19756
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 14227 17100 14293 17101
rect 14227 17036 14228 17100
rect 14292 17036 14293 17100
rect 14227 17035 14293 17036
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 14230 12477 14290 17035
rect 15147 16692 15213 16693
rect 15147 16628 15148 16692
rect 15212 16628 15213 16692
rect 15147 16627 15213 16628
rect 15150 13701 15210 16627
rect 17944 16352 18264 17376
rect 22142 17101 22202 19755
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22139 17100 22205 17101
rect 22139 17036 22140 17100
rect 22204 17036 22205 17100
rect 22139 17035 22205 17036
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 15147 13700 15213 13701
rect 15147 13636 15148 13700
rect 15212 13636 15213 13700
rect 15147 13635 15213 13636
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 14227 12476 14293 12477
rect 14227 12412 14228 12476
rect 14292 12412 14293 12476
rect 14227 12411 14293 12412
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 16896 23264 17920
rect 25270 17781 25330 22883
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27944 18528 28264 19552
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 25267 17780 25333 17781
rect 25267 17716 25268 17780
rect 25332 17716 25333 17780
rect 25267 17715 25333 17716
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 27944 17440 28264 18464
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27944 14176 28264 15200
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 24512 33264 24528
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 32944 19072 33264 20096
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32944 10368 33264 11392
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 23968 38264 24528
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 24512 43264 24528
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 23968 48264 24528
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_2  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14628 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1676037725
transform -1 0 11408 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1676037725
transform -1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1676037725
transform -1 0 6716 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1676037725
transform -1 0 10580 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1676037725
transform -1 0 11224 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform -1 0 14444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1676037725
transform -1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1676037725
transform -1 0 10672 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1676037725
transform -1 0 11224 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1676037725
transform -1 0 12052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform -1 0 9476 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1676037725
transform -1 0 15272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1676037725
transform -1 0 16376 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1676037725
transform -1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform -1 0 8004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform -1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform -1 0 12788 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform -1 0 15640 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform -1 0 8004 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1676037725
transform -1 0 12052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1676037725
transform -1 0 12512 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1676037725
transform -1 0 12144 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _127_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7820 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1676037725
transform -1 0 5520 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform -1 0 12052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1676037725
transform 1 0 7728 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1676037725
transform 1 0 3864 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1676037725
transform -1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1676037725
transform -1 0 6900 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1676037725
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1676037725
transform 1 0 37904 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform 1 0 37168 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1676037725
transform 1 0 43608 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 37628 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 37444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 43884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 38456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 37904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 44804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform 1 0 38640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 40204 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 39192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform 1 0 44068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1676037725
transform 1 0 40020 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1676037725
transform 1 0 38180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1676037725
transform 1 0 39652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1676037725
transform 1 0 44252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1676037725
transform 1 0 40020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1676037725
transform 1 0 39836 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 40020 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 44988 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 45540 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 39928 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1676037725
transform -1 0 46184 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1676037725
transform -1 0 46184 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1676037725
transform -1 0 45908 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform 1 0 44896 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1676037725
transform -1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1676037725
transform 1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1676037725
transform -1 0 5612 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _167_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1676037725
transform 1 0 6624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1676037725
transform 1 0 4692 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1676037725
transform -1 0 3680 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 1676037725
transform -1 0 2392 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1676037725
transform -1 0 6808 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp 1676037725
transform -1 0 4232 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1676037725
transform -1 0 26128 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1676037725
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1676037725
transform -1 0 13064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1676037725
transform 1 0 12328 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _179_
timestamp 1676037725
transform -1 0 13432 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1676037725
transform 1 0 14628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _181_
timestamp 1676037725
transform 1 0 13892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1676037725
transform -1 0 14812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1676037725
transform -1 0 7544 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1676037725
transform -1 0 23736 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1676037725
transform -1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1676037725
transform -1 0 19964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _187_
timestamp 1676037725
transform -1 0 22908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1676037725
transform -1 0 21528 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1676037725
transform -1 0 24932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1676037725
transform -1 0 27508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1676037725
transform -1 0 21528 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1676037725
transform 1 0 23184 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _194_
timestamp 1676037725
transform -1 0 16744 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1676037725
transform 1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1676037725
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 1676037725
transform -1 0 19688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1676037725
transform -1 0 20884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1676037725
transform -1 0 21528 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1676037725
transform -1 0 26680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1676037725
transform -1 0 10764 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1676037725
transform 1 0 9844 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1676037725
transform 1 0 10396 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1676037725
transform -1 0 10580 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1676037725
transform -1 0 13984 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1676037725
transform -1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1676037725
transform -1 0 10488 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1676037725
transform -1 0 10396 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1676037725
transform -1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1676037725
transform -1 0 15088 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1676037725
transform -1 0 11776 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1676037725
transform 1 0 11592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1676037725
transform -1 0 11960 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1676037725
transform -1 0 14904 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1676037725
transform -1 0 11408 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1676037725
transform 1 0 12236 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1676037725
transform -1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1676037725
transform -1 0 9384 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1676037725
transform 1 0 7452 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1676037725
transform -1 0 37076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1676037725
transform -1 0 38640 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A
timestamp 1676037725
transform 1 0 36800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A
timestamp 1676037725
transform -1 0 39100 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1676037725
transform -1 0 38180 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1676037725
transform -1 0 39192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1676037725
transform 1 0 37352 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1676037725
transform 1 0 37536 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1676037725
transform -1 0 39376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1676037725
transform -1 0 40940 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1676037725
transform -1 0 40020 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1676037725
transform -1 0 40756 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1676037725
transform -1 0 38916 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1676037725
transform -1 0 40388 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1676037725
transform 1 0 39560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1676037725
transform -1 0 40756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1676037725
transform -1 0 40572 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1676037725
transform -1 0 40664 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__A
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A
timestamp 1676037725
transform -1 0 26496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__A
timestamp 1676037725
transform -1 0 8464 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 19504 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20332 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 18216 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 18676 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18952 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 12696 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 16100 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 15640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 10856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10396 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 12420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11960 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14996 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 12880 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 11224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15088 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12328 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 15180 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A0
timestamp 1676037725
transform -1 0 21988 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 20516 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 15640 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 9476 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__S
timestamp 1676037725
transform -1 0 9844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 13616 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 9844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__S
timestamp 1676037725
transform -1 0 10212 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1676037725
transform -1 0 19504 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 19320 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 17940 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 17572 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__S
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 12328 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 16192 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 16744 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 16376 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 13340 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__S
timestamp 1676037725
transform 1 0 15180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 12788 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 10488 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 11592 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 16652 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 17940 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A0
timestamp 1676037725
transform -1 0 16008 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1676037725
transform -1 0 17204 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 24012 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23000 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform -1 0 23368 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 28244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 31004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1676037725
transform 1 0 28060 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1676037725
transform -1 0 24564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1676037725
transform 1 0 22172 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1676037725
transform 1 0 18768 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1676037725
transform 1 0 18952 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1676037725
transform -1 0 22724 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1676037725
transform 1 0 24656 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1676037725
transform 1 0 28428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1676037725
transform 1 0 28888 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1676037725
transform 1 0 34500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1676037725
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1676037725
transform 1 0 30360 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1676037725
transform -1 0 37168 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1676037725
transform 1 0 35328 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold3_A
timestamp 1676037725
transform -1 0 44528 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold4_A
timestamp 1676037725
transform -1 0 46644 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold6_A
timestamp 1676037725
transform -1 0 9476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform -1 0 3680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform -1 0 3220 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform -1 0 2484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform -1 0 2944 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform -1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform -1 0 2300 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1676037725
transform -1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1676037725
transform -1 0 2300 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1676037725
transform -1 0 3036 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1676037725
transform -1 0 3220 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1676037725
transform -1 0 2484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1676037725
transform -1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1676037725
transform -1 0 2300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1676037725
transform -1 0 3036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1676037725
transform -1 0 3220 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1676037725
transform -1 0 2484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1676037725
transform -1 0 2944 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1676037725
transform -1 0 2852 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1676037725
transform -1 0 2300 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1676037725
transform -1 0 3496 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1676037725
transform -1 0 2300 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1676037725
transform -1 0 4140 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1676037725
transform -1 0 2852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1676037725
transform -1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1676037725
transform -1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1676037725
transform -1 0 3036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1676037725
transform -1 0 3220 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1676037725
transform -1 0 2484 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1676037725
transform -1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1676037725
transform -1 0 3036 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1676037725
transform -1 0 48852 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1676037725
transform -1 0 48668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1676037725
transform -1 0 48852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1676037725
transform -1 0 48852 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1676037725
transform -1 0 48668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1676037725
transform -1 0 48668 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1676037725
transform -1 0 48852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1676037725
transform -1 0 48852 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1676037725
transform -1 0 48484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1676037725
transform -1 0 48024 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1676037725
transform -1 0 46920 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1676037725
transform -1 0 48208 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1676037725
transform -1 0 48668 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1676037725
transform -1 0 46828 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1676037725
transform -1 0 47288 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1676037725
transform -1 0 46460 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1676037725
transform -1 0 48208 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1676037725
transform 1 0 46552 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1676037725
transform -1 0 47932 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1676037725
transform 1 0 47932 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1676037725
transform -1 0 47748 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1676037725
transform -1 0 47104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1676037725
transform -1 0 48668 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1676037725
transform -1 0 48852 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1676037725
transform -1 0 48944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1676037725
transform -1 0 48852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1676037725
transform -1 0 48668 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1676037725
transform -1 0 48852 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1676037725
transform -1 0 48852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1676037725
transform -1 0 48668 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1676037725
transform -1 0 27048 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1676037725
transform -1 0 29716 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1676037725
transform -1 0 31832 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1676037725
transform -1 0 31188 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1676037725
transform -1 0 34316 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1676037725
transform -1 0 41952 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1676037725
transform -1 0 34868 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1676037725
transform -1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1676037725
transform -1 0 42964 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1676037725
transform -1 0 42780 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1676037725
transform -1 0 46000 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1676037725
transform -1 0 9568 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1676037725
transform -1 0 41032 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1676037725
transform -1 0 46552 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1676037725
transform -1 0 43148 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1676037725
transform -1 0 43332 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1676037725
transform -1 0 43148 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1676037725
transform -1 0 42596 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1676037725
transform -1 0 44712 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1676037725
transform -1 0 43516 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1676037725
transform -1 0 45816 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1676037725
transform -1 0 43976 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1676037725
transform -1 0 14260 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1676037725
transform -1 0 24656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1676037725
transform -1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1676037725
transform -1 0 31648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1676037725
transform -1 0 25300 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1676037725
transform -1 0 29164 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1676037725
transform -1 0 29072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1676037725
transform -1 0 29348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1676037725
transform -1 0 29716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1676037725
transform -1 0 31464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1676037725
transform -1 0 33580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1676037725
transform -1 0 35696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1676037725
transform -1 0 37168 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1676037725
transform -1 0 43332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1676037725
transform -1 0 45172 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1676037725
transform -1 0 46276 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1676037725
transform -1 0 47748 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1676037725
transform -1 0 47380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1676037725
transform -1 0 47932 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1676037725
transform -1 0 49312 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1676037725
transform -1 0 49496 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1676037725
transform -1 0 47472 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1676037725
transform -1 0 44896 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1676037725
transform -1 0 47472 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output174_A
timestamp 1676037725
transform -1 0 7268 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 27048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26588 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 24472 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22080 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1676037725
transform 1 0 19228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 19044 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 17020 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20608 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22080 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 20516 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23460 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 20700 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform -1 0 22172 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23184 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22724 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21160 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20792 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 19044 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20884 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25116 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 25300 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 27784 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 29072 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 27600 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 30176 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 30728 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 26680 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 29072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 27600 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21896 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 28152 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 31556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 34316 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 34224 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 36708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 38456 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform -1 0 37076 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 38456 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 38456 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform -1 0 39468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 39468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 37444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 38640 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 35880 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 36064 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 36892 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 33488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 34684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 33672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 34132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 31740 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 28980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 32752 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 33304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 34684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 32936 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 30176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 29072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform -1 0 45816 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 43608 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 33304 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 34040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 31832 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 34316 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 34224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 36892 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1676037725
transform 1 0 38456 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 39284 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 39468 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 39560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 37076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 37260 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 35512 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 39468 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 40388 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1676037725
transform 1 0 41032 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 40572 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 37628 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 39376 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 40204 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1676037725
transform 1 0 37444 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 40020 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 37260 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 39192 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 37444 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 37444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 37444 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 41124 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1676037725
transform 1 0 37628 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 40020 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 42044 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 40940 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 41032 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 41492 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 42044 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 40020 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 38916 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 35880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 27416 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26680 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26036 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26588 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25852 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23828 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13156 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 12328 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12972 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 14536 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 12696 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14352 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 19596 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_0__S
timestamp 1676037725
transform -1 0 31924 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 28336 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 28152 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 25852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 26220 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 26404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 19136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_3__S
timestamp 1676037725
transform -1 0 20700 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 30176 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 26404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 25208 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 25208 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 26220 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 25852 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 17756 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 27968 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 25484 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 25484 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 30176 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 26588 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 20332 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 27508 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 25760 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 24656 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__A0
timestamp 1676037725
transform -1 0 22356 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 22356 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 29440 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 25944 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 24104 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 22264 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 21896 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 28980 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 26680 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 25116 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_37.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 30912 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_37.mux_l2_in_1__A1
timestamp 1676037725
transform -1 0 24564 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_45.mux_l2_in_1__A1
timestamp 1676037725
transform -1 0 30544 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 25576 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_1__A1
timestamp 1676037725
transform -1 0 21252 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 30360 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 36064 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 34316 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__S
timestamp 1676037725
transform -1 0 34500 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 27600 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 27508 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__S
timestamp 1676037725
transform -1 0 27968 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1676037725
transform -1 0 34040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__A0
timestamp 1676037725
transform -1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 29532 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_0__S
timestamp 1676037725
transform -1 0 36892 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1676037725
transform -1 0 37812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 37444 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__S
timestamp 1676037725
transform -1 0 37076 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__A0
timestamp 1676037725
transform -1 0 30912 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__A1
timestamp 1676037725
transform -1 0 29440 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__S
timestamp 1676037725
transform -1 0 31924 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_0__S
timestamp 1676037725
transform -1 0 35880 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1676037725
transform -1 0 34592 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 33948 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 36616 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 36800 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 32752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_3__S
timestamp 1676037725
transform -1 0 33488 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 34316 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 34224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 34316 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 34500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 34316 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 30452 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_3__S
timestamp 1676037725
transform -1 0 32016 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 34684 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 34684 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 26220 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 26036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 31832 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 32292 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 29440 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 26036 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 30728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_1__A0
timestamp 1676037725
transform -1 0 29072 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 32016 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 25668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 33764 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 33304 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 30268 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 29072 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 27784 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 36892 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 35696 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 44712 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_1__S
timestamp 1676037725
transform -1 0 43976 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__A0
timestamp 1676037725
transform -1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 22908 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__S
timestamp 1676037725
transform -1 0 22908 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 28520 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 41216 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 39652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 46184 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 31096 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 36892 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 42780 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 29716 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 42596 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 42596 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_2__A0
timestamp 1676037725
transform -1 0 33856 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 34040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 42228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 34224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__A1
timestamp 1676037725
transform -1 0 34592 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 36892 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 41308 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 31740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 41032 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 41216 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l2_in_1__A1
timestamp 1676037725
transform -1 0 39192 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 41584 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 41952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 36892 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 41216 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 41400 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 36432 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 38824 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 39008 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 28520 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 28888 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 24656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 27140 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 27968 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 28336 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 21988 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 28612 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 24012 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_28.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21620 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_30.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21804 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 23184 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_32.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16008 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 19136 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_34.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 16928 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 27140 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 27508 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 23000 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_40.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 12236 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_40.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 12788 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_42.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_42.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17756 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_44.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 15088 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_46.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 10488 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_48.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 16836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_50.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 16744 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_58.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 25484 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_58.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 26680 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 20148 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16376 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18216 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 18952 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 16192 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 16100 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 13616 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 15456 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10764 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9476 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform -1 0 12788 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 15180 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 12604 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform -1 0 11040 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15272 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform -1 0 16376 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 20700 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform -1 0 16376 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform -1 0 16008 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 17112 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 16928 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 18308 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__254 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform -1 0 16376 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform -1 0 17480 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform -1 0 18676 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 19872 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform -1 0 11224 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform -1 0 13524 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 19504 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 17940 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform -1 0 13800 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform -1 0 13524 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__255
timestamp 1676037725
transform -1 0 13800 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 17112 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform -1 0 14720 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform -1 0 16008 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform -1 0 8556 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform -1 0 8740 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 18124 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 14444 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 16744 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform -1 0 10212 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__256
timestamp 1676037725
transform -1 0 11224 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform -1 0 12512 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform -1 0 12512 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 12328 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform -1 0 12972 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 15824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform -1 0 13800 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14352 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 15640 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 18308 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 15088 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13156 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 14352 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__257
timestamp 1676037725
transform -1 0 16008 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 16376 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 11960 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform -1 0 11868 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 14536 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 29072 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23552 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 22724 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21896 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform -1 0 27048 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform -1 0 23828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 20424 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20976 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform -1 0 26128 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 23000 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform -1 0 24104 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24196 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform -1 0 26496 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22264 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform -1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 18032 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28888 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 28980 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18952 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 17848 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 22448 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 22540 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform -1 0 18768 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 17940 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform -1 0 23000 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 23276 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 28796 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform -1 0 29256 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 33304 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 34040 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 29900 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 30728 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform -1 0 35604 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform -1 0 35880 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17
timestamp 1676037725
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24
timestamp 1676037725
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1676037725
transform 1 0 9476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10396 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132
timestamp 1676037725
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_159
timestamp 1676037725
transform 1 0 15732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1676037725
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1676037725
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_225 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_247
timestamp 1676037725
transform 1 0 23828 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1676037725
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_271
timestamp 1676037725
transform 1 0 26036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1676037725
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1676037725
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_299
timestamp 1676037725
transform 1 0 28612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1676037725
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_311
timestamp 1676037725
transform 1 0 29716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_326
timestamp 1676037725
transform 1 0 31096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1676037725
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_345
timestamp 1676037725
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_349
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_353
timestamp 1676037725
transform 1 0 33580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1676037725
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_372
timestamp 1676037725
transform 1 0 35328 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_376
timestamp 1676037725
transform 1 0 35696 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_388
timestamp 1676037725
transform 1 0 36800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1676037725
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_429
timestamp 1676037725
transform 1 0 40572 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1676037725
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_459
timestamp 1676037725
transform 1 0 43332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_471
timestamp 1676037725
transform 1 0 44436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1676037725
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_485
timestamp 1676037725
transform 1 0 45724 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1676037725
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1676037725
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_9
timestamp 1676037725
transform 1 0 1932 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_19
timestamp 1676037725
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_31
timestamp 1676037725
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_43
timestamp 1676037725
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_96
timestamp 1676037725
transform 1 0 9936 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1676037725
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1676037725
transform 1 0 12236 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_130
timestamp 1676037725
transform 1 0 13064 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_142
timestamp 1676037725
transform 1 0 14168 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1676037725
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_171
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1676037725
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_184
timestamp 1676037725
transform 1 0 18032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_201
timestamp 1676037725
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_208
timestamp 1676037725
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1676037725
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_235
timestamp 1676037725
transform 1 0 22724 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_239
timestamp 1676037725
transform 1 0 23092 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_247
timestamp 1676037725
transform 1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_271
timestamp 1676037725
transform 1 0 26036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1676037725
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_297
timestamp 1676037725
transform 1 0 28428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_301
timestamp 1676037725
transform 1 0 28796 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_323
timestamp 1676037725
transform 1 0 30820 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_327
timestamp 1676037725
transform 1 0 31188 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_465
timestamp 1676037725
transform 1 0 43884 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_482
timestamp 1676037725
transform 1 0 45448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1676037725
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1676037725
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_170
timestamp 1676037725
transform 1 0 16744 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_182
timestamp 1676037725
transform 1 0 17848 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1676037725
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_215
timestamp 1676037725
transform 1 0 20884 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_236
timestamp 1676037725
transform 1 0 22816 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_242
timestamp 1676037725
transform 1 0 23368 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_276
timestamp 1676037725
transform 1 0 26496 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_288
timestamp 1676037725
transform 1 0 27600 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_300
timestamp 1676037725
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_387
timestamp 1676037725
transform 1 0 36708 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_391
timestamp 1676037725
transform 1 0 37076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_403
timestamp 1676037725
transform 1 0 38180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_415
timestamp 1676037725
transform 1 0 39284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1676037725
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_479
timestamp 1676037725
transform 1 0 45172 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_485
timestamp 1676037725
transform 1 0 45724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_505
timestamp 1676037725
transform 1 0 47564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_9
timestamp 1676037725
transform 1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_17
timestamp 1676037725
transform 1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_23
timestamp 1676037725
transform 1 0 3220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_35
timestamp 1676037725
transform 1 0 4324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1676037725
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_229
timestamp 1676037725
transform 1 0 22172 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_233
timestamp 1676037725
transform 1 0 22540 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_240
timestamp 1676037725
transform 1 0 23184 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_247
timestamp 1676037725
transform 1 0 23828 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_272
timestamp 1676037725
transform 1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_304
timestamp 1676037725
transform 1 0 29072 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_316
timestamp 1676037725
transform 1 0 30176 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_328
timestamp 1676037725
transform 1 0 31280 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1676037725
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_507
timestamp 1676037725
transform 1 0 47748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1676037725
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_9
timestamp 1676037725
transform 1 0 1932 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_218
timestamp 1676037725
transform 1 0 21160 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_234
timestamp 1676037725
transform 1 0 22632 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_241
timestamp 1676037725
transform 1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1676037725
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_282
timestamp 1676037725
transform 1 0 27048 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_294
timestamp 1676037725
transform 1 0 28152 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1676037725
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_385
timestamp 1676037725
transform 1 0 36524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_390
timestamp 1676037725
transform 1 0 36984 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_396
timestamp 1676037725
transform 1 0 37536 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_404
timestamp 1676037725
transform 1 0 38272 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_408
timestamp 1676037725
transform 1 0 38640 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_491
timestamp 1676037725
transform 1 0 46276 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_497
timestamp 1676037725
transform 1 0 46828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_505
timestamp 1676037725
transform 1 0 47564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_201
timestamp 1676037725
transform 1 0 19596 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_213
timestamp 1676037725
transform 1 0 20700 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp 1676037725
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_395
timestamp 1676037725
transform 1 0 37444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_401
timestamp 1676037725
transform 1 0 37996 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_409
timestamp 1676037725
transform 1 0 38732 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_413
timestamp 1676037725
transform 1 0 39100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_425
timestamp 1676037725
transform 1 0 40204 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_437
timestamp 1676037725
transform 1 0 41308 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_445
timestamp 1676037725
transform 1 0 42044 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1676037725
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1676037725
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1676037725
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_17
timestamp 1676037725
transform 1 0 2668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1676037725
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_461
timestamp 1676037725
transform 1 0 43516 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_466
timestamp 1676037725
transform 1 0 43976 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_474
timestamp 1676037725
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_9
timestamp 1676037725
transform 1 0 1932 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_192
timestamp 1676037725
transform 1 0 18768 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_204
timestamp 1676037725
transform 1 0 19872 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_216
timestamp 1676037725
transform 1 0 20976 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_399
timestamp 1676037725
transform 1 0 37812 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_403
timestamp 1676037725
transform 1 0 38180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_415
timestamp 1676037725
transform 1 0 39284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_427
timestamp 1676037725
transform 1 0 40388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_439
timestamp 1676037725
transform 1 0 41492 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_469
timestamp 1676037725
transform 1 0 44252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_481
timestamp 1676037725
transform 1 0 45356 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_493
timestamp 1676037725
transform 1 0 46460 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_501
timestamp 1676037725
transform 1 0 47196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1676037725
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_9
timestamp 1676037725
transform 1 0 1932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_16
timestamp 1676037725
transform 1 0 2576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1676037725
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_183
timestamp 1676037725
transform 1 0 17940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_204
timestamp 1676037725
transform 1 0 19872 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_216
timestamp 1676037725
transform 1 0 20976 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_224
timestamp 1676037725
transform 1 0 21712 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_227
timestamp 1676037725
transform 1 0 21988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_239
timestamp 1676037725
transform 1 0 23092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_505
timestamp 1676037725
transform 1 0 47564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_9
timestamp 1676037725
transform 1 0 1932 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_13
timestamp 1676037725
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_25
timestamp 1676037725
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_37
timestamp 1676037725
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1676037725
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_185
timestamp 1676037725
transform 1 0 18124 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_188
timestamp 1676037725
transform 1 0 18400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_196
timestamp 1676037725
transform 1 0 19136 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_208
timestamp 1676037725
transform 1 0 20240 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_216
timestamp 1676037725
transform 1 0 20976 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_221
timestamp 1676037725
transform 1 0 21436 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_236
timestamp 1676037725
transform 1 0 22816 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_240
timestamp 1676037725
transform 1 0 23184 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_252
timestamp 1676037725
transform 1 0 24288 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_264
timestamp 1676037725
transform 1 0 25392 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1676037725
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_323
timestamp 1676037725
transform 1 0 30820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_327
timestamp 1676037725
transform 1 0 31188 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_333
timestamp 1676037725
transform 1 0 31740 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_342
timestamp 1676037725
transform 1 0 32568 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_346
timestamp 1676037725
transform 1 0 32936 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_358
timestamp 1676037725
transform 1 0 34040 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_370
timestamp 1676037725
transform 1 0 35144 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_382
timestamp 1676037725
transform 1 0 36248 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1676037725
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_396
timestamp 1676037725
transform 1 0 37536 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_402
timestamp 1676037725
transform 1 0 38088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_410
timestamp 1676037725
transform 1 0 38824 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_414
timestamp 1676037725
transform 1 0 39192 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_426
timestamp 1676037725
transform 1 0 40296 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_438
timestamp 1676037725
transform 1 0 41400 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_446
timestamp 1676037725
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_479
timestamp 1676037725
transform 1 0 45172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_491
timestamp 1676037725
transform 1 0 46276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1676037725
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_9
timestamp 1676037725
transform 1 0 1932 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_160
timestamp 1676037725
transform 1 0 15824 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_168
timestamp 1676037725
transform 1 0 16560 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 1676037725
transform 1 0 17480 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_191
timestamp 1676037725
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_219
timestamp 1676037725
transform 1 0 21252 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_225
timestamp 1676037725
transform 1 0 21804 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_236
timestamp 1676037725
transform 1 0 22816 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_240
timestamp 1676037725
transform 1 0 23184 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_314
timestamp 1676037725
transform 1 0 29992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_323
timestamp 1676037725
transform 1 0 30820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_334
timestamp 1676037725
transform 1 0 31832 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_338
timestamp 1676037725
transform 1 0 32200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_348
timestamp 1676037725
transform 1 0 33120 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_352
timestamp 1676037725
transform 1 0 33488 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_395
timestamp 1676037725
transform 1 0 37444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_398
timestamp 1676037725
transform 1 0 37720 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_404
timestamp 1676037725
transform 1 0 38272 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_412
timestamp 1676037725
transform 1 0 39008 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_416
timestamp 1676037725
transform 1 0 39376 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1676037725
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1676037725
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_133
timestamp 1676037725
transform 1 0 13340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_156
timestamp 1676037725
transform 1 0 15456 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_160
timestamp 1676037725
transform 1 0 15824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 1676037725
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp 1676037725
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_198
timestamp 1676037725
transform 1 0 19320 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_247
timestamp 1676037725
transform 1 0 23828 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_251
timestamp 1676037725
transform 1 0 24196 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_263
timestamp 1676037725
transform 1 0 25300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_275
timestamp 1676037725
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_321
timestamp 1676037725
transform 1 0 30636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1676037725
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_359
timestamp 1676037725
transform 1 0 34132 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_367
timestamp 1676037725
transform 1 0 34868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_379
timestamp 1676037725
transform 1 0 35972 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1676037725
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_398
timestamp 1676037725
transform 1 0 37720 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_410
timestamp 1676037725
transform 1 0 38824 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_414
timestamp 1676037725
transform 1 0 39192 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_422
timestamp 1676037725
transform 1 0 39928 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_429
timestamp 1676037725
transform 1 0 40572 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_433
timestamp 1676037725
transform 1 0 40940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_445
timestamp 1676037725
transform 1 0 42044 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_471
timestamp 1676037725
transform 1 0 44436 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_483
timestamp 1676037725
transform 1 0 45540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_502
timestamp 1676037725
transform 1 0 47288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1676037725
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_9
timestamp 1676037725
transform 1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_17
timestamp 1676037725
transform 1 0 2668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1676037725
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_146
timestamp 1676037725
transform 1 0 14536 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1676037725
transform 1 0 14996 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_162
timestamp 1676037725
transform 1 0 16008 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1676037725
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_190
timestamp 1676037725
transform 1 0 18584 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1676037725
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_226
timestamp 1676037725
transform 1 0 21896 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_259
timestamp 1676037725
transform 1 0 24932 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_269
timestamp 1676037725
transform 1 0 25852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_281
timestamp 1676037725
transform 1 0 26956 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_292
timestamp 1676037725
transform 1 0 27968 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_303
timestamp 1676037725
transform 1 0 28980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_314
timestamp 1676037725
transform 1 0 29992 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_318
timestamp 1676037725
transform 1 0 30360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_342
timestamp 1676037725
transform 1 0 32568 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_348
timestamp 1676037725
transform 1 0 33120 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_359
timestamp 1676037725
transform 1 0 34132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_376
timestamp 1676037725
transform 1 0 35696 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_384
timestamp 1676037725
transform 1 0 36432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_388
timestamp 1676037725
transform 1 0 36800 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_396
timestamp 1676037725
transform 1 0 37536 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_400
timestamp 1676037725
transform 1 0 37904 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_412
timestamp 1676037725
transform 1 0 39008 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_418
timestamp 1676037725
transform 1 0 39560 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_423
timestamp 1676037725
transform 1 0 40020 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_435
timestamp 1676037725
transform 1 0 41124 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_447
timestamp 1676037725
transform 1 0 42228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_459
timestamp 1676037725
transform 1 0 43332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_471
timestamp 1676037725
transform 1 0 44436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1676037725
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_501
timestamp 1676037725
transform 1 0 47196 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1676037725
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_9
timestamp 1676037725
transform 1 0 1932 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1676037725
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_129
timestamp 1676037725
transform 1 0 12972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1676037725
transform 1 0 15456 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1676037725
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_218
timestamp 1676037725
transform 1 0 21160 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_227
timestamp 1676037725
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_239
timestamp 1676037725
transform 1 0 23092 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_263
timestamp 1676037725
transform 1 0 25300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1676037725
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_307
timestamp 1676037725
transform 1 0 29348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_331
timestamp 1676037725
transform 1 0 31556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1676037725
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_339
timestamp 1676037725
transform 1 0 32292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_351
timestamp 1676037725
transform 1 0 33396 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_355
timestamp 1676037725
transform 1 0 33764 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_376
timestamp 1676037725
transform 1 0 35696 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_382
timestamp 1676037725
transform 1 0 36248 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1676037725
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1676037725
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1676037725
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1676037725
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1676037725
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1676037725
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1676037725
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1676037725
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_124
timestamp 1676037725
transform 1 0 12512 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_135
timestamp 1676037725
transform 1 0 13524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_163
timestamp 1676037725
transform 1 0 16100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1676037725
transform 1 0 16744 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_181
timestamp 1676037725
transform 1 0 17756 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_203
timestamp 1676037725
transform 1 0 19780 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_207
timestamp 1676037725
transform 1 0 20148 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_228
timestamp 1676037725
transform 1 0 22080 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_243
timestamp 1676037725
transform 1 0 23460 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_275
timestamp 1676037725
transform 1 0 26404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_279
timestamp 1676037725
transform 1 0 26772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_301
timestamp 1676037725
transform 1 0 28796 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_305
timestamp 1676037725
transform 1 0 29164 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_314
timestamp 1676037725
transform 1 0 29992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_338
timestamp 1676037725
transform 1 0 32200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_351
timestamp 1676037725
transform 1 0 33396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_358
timestamp 1676037725
transform 1 0 34040 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_387
timestamp 1676037725
transform 1 0 36708 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_391
timestamp 1676037725
transform 1 0 37076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_407
timestamp 1676037725
transform 1 0 38548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_411
timestamp 1676037725
transform 1 0 38916 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1676037725
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_427
timestamp 1676037725
transform 1 0 40388 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_431
timestamp 1676037725
transform 1 0 40756 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_443
timestamp 1676037725
transform 1 0 41860 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_455
timestamp 1676037725
transform 1 0 42964 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_467
timestamp 1676037725
transform 1 0 44068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_473
timestamp 1676037725
transform 1 0 44620 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_505
timestamp 1676037725
transform 1 0 47564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1676037725
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_9
timestamp 1676037725
transform 1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_17
timestamp 1676037725
transform 1 0 2668 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 1676037725
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1676037725
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_129
timestamp 1676037725
transform 1 0 12972 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_140
timestamp 1676037725
transform 1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1676037725
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_172
timestamp 1676037725
transform 1 0 16928 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_183
timestamp 1676037725
transform 1 0 17940 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1676037725
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1676037725
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_247
timestamp 1676037725
transform 1 0 23828 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_260
timestamp 1676037725
transform 1 0 25024 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_267
timestamp 1676037725
transform 1 0 25668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_277
timestamp 1676037725
transform 1 0 26588 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_292
timestamp 1676037725
transform 1 0 27968 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_296
timestamp 1676037725
transform 1 0 28336 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_299
timestamp 1676037725
transform 1 0 28612 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_312
timestamp 1676037725
transform 1 0 29808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_325
timestamp 1676037725
transform 1 0 31004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_332
timestamp 1676037725
transform 1 0 31648 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_348
timestamp 1676037725
transform 1 0 33120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_352
timestamp 1676037725
transform 1 0 33488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_376
timestamp 1676037725
transform 1 0 35696 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_389
timestamp 1676037725
transform 1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_397
timestamp 1676037725
transform 1 0 37628 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_409
timestamp 1676037725
transform 1 0 38732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_417
timestamp 1676037725
transform 1 0 39468 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_423
timestamp 1676037725
transform 1 0 40020 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_427
timestamp 1676037725
transform 1 0 40388 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_439
timestamp 1676037725
transform 1 0 41492 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1676037725
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1676037725
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1676037725
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1676037725
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1676037725
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1676037725
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1676037725
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_9
timestamp 1676037725
transform 1 0 1932 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_105
timestamp 1676037725
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_127
timestamp 1676037725
transform 1 0 12788 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1676037725
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_179
timestamp 1676037725
transform 1 0 17572 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_192
timestamp 1676037725
transform 1 0 18768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_201
timestamp 1676037725
transform 1 0 19596 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_206
timestamp 1676037725
transform 1 0 20056 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_230
timestamp 1676037725
transform 1 0 22264 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_237
timestamp 1676037725
transform 1 0 22908 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_275
timestamp 1676037725
transform 1 0 26404 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_279
timestamp 1676037725
transform 1 0 26772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_300
timestamp 1676037725
transform 1 0 28704 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_320
timestamp 1676037725
transform 1 0 30544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_324
timestamp 1676037725
transform 1 0 30912 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_346
timestamp 1676037725
transform 1 0 32936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_361
timestamp 1676037725
transform 1 0 34316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_367
timestamp 1676037725
transform 1 0 34868 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_375
timestamp 1676037725
transform 1 0 35604 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_399
timestamp 1676037725
transform 1 0 37812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_406
timestamp 1676037725
transform 1 0 38456 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_410
timestamp 1676037725
transform 1 0 38824 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_427
timestamp 1676037725
transform 1 0 40388 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_434
timestamp 1676037725
transform 1 0 41032 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_446
timestamp 1676037725
transform 1 0 42136 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_458
timestamp 1676037725
transform 1 0 43240 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_470
timestamp 1676037725
transform 1 0 44344 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_487
timestamp 1676037725
transform 1 0 45908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_499
timestamp 1676037725
transform 1 0 47012 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_507
timestamp 1676037725
transform 1 0 47748 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1676037725
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1676037725
transform 1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_16
timestamp 1676037725
transform 1 0 2576 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_20
timestamp 1676037725
transform 1 0 2944 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_32
timestamp 1676037725
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_44
timestamp 1676037725
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_115
timestamp 1676037725
transform 1 0 11684 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1676037725
transform 1 0 12144 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_131
timestamp 1676037725
transform 1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_148
timestamp 1676037725
transform 1 0 14720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_191
timestamp 1676037725
transform 1 0 18676 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_198
timestamp 1676037725
transform 1 0 19320 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1676037725
transform 1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_231
timestamp 1676037725
transform 1 0 22356 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1676037725
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_268
timestamp 1676037725
transform 1 0 25760 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_273
timestamp 1676037725
transform 1 0 26220 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1676037725
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_292
timestamp 1676037725
transform 1 0 27968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_296
timestamp 1676037725
transform 1 0 28336 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_318
timestamp 1676037725
transform 1 0 30360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_331
timestamp 1676037725
transform 1 0 31556 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_348
timestamp 1676037725
transform 1 0 33120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_361
timestamp 1676037725
transform 1 0 34316 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_367
timestamp 1676037725
transform 1 0 34868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1676037725
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_404
timestamp 1676037725
transform 1 0 38272 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_417
timestamp 1676037725
transform 1 0 39468 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_425
timestamp 1676037725
transform 1 0 40204 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_431
timestamp 1676037725
transform 1 0 40756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_443
timestamp 1676037725
transform 1 0 41860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1676037725
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1676037725
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_473
timestamp 1676037725
transform 1 0 44620 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_481
timestamp 1676037725
transform 1 0 45356 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_493
timestamp 1676037725
transform 1 0 46460 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_501
timestamp 1676037725
transform 1 0 47196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1676037725
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_19
timestamp 1676037725
transform 1 0 2852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_111
timestamp 1676037725
transform 1 0 11316 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_164
timestamp 1676037725
transform 1 0 16192 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_168
timestamp 1676037725
transform 1 0 16560 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1676037725
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_208
timestamp 1676037725
transform 1 0 20240 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_213
timestamp 1676037725
transform 1 0 20700 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_224
timestamp 1676037725
transform 1 0 21712 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_237
timestamp 1676037725
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_275
timestamp 1676037725
transform 1 0 26404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_279
timestamp 1676037725
transform 1 0 26772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_290
timestamp 1676037725
transform 1 0 27784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_294
timestamp 1676037725
transform 1 0 28152 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1676037725
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_331
timestamp 1676037725
transform 1 0 31556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_335
timestamp 1676037725
transform 1 0 31924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_387
timestamp 1676037725
transform 1 0 36708 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_400
timestamp 1676037725
transform 1 0 37904 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_413
timestamp 1676037725
transform 1 0 39100 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1676037725
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_427
timestamp 1676037725
transform 1 0 40388 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_434
timestamp 1676037725
transform 1 0 41032 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_441
timestamp 1676037725
transform 1 0 41676 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_453
timestamp 1676037725
transform 1 0 42780 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_465
timestamp 1676037725
transform 1 0 43884 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_473
timestamp 1676037725
transform 1 0 44620 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_485
timestamp 1676037725
transform 1 0 45724 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_490
timestamp 1676037725
transform 1 0 46184 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_502
timestamp 1676037725
transform 1 0 47288 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_508
timestamp 1676037725
transform 1 0 47840 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_9
timestamp 1676037725
transform 1 0 1932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_13
timestamp 1676037725
transform 1 0 2300 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_22
timestamp 1676037725
transform 1 0 3128 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_26
timestamp 1676037725
transform 1 0 3496 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_38
timestamp 1676037725
transform 1 0 4600 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1676037725
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_124
timestamp 1676037725
transform 1 0 12512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_128
timestamp 1676037725
transform 1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_150
timestamp 1676037725
transform 1 0 14904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1676037725
transform 1 0 15364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1676037725
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_173
timestamp 1676037725
transform 1 0 17020 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1676037725
transform 1 0 17480 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_193
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_206
timestamp 1676037725
transform 1 0 20056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_211
timestamp 1676037725
transform 1 0 20516 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_230
timestamp 1676037725
transform 1 0 22264 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_243
timestamp 1676037725
transform 1 0 23460 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_267
timestamp 1676037725
transform 1 0 25668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_277
timestamp 1676037725
transform 1 0 26588 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_306
timestamp 1676037725
transform 1 0 29256 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_311
timestamp 1676037725
transform 1 0 29716 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1676037725
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_348
timestamp 1676037725
transform 1 0 33120 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_356
timestamp 1676037725
transform 1 0 33856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_369
timestamp 1676037725
transform 1 0 35052 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_382
timestamp 1676037725
transform 1 0 36248 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_418
timestamp 1676037725
transform 1 0 39560 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_426
timestamp 1676037725
transform 1 0 40296 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_430
timestamp 1676037725
transform 1 0 40664 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_442
timestamp 1676037725
transform 1 0 41768 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1676037725
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1676037725
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_485
timestamp 1676037725
transform 1 0 45724 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_490
timestamp 1676037725
transform 1 0 46184 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_502
timestamp 1676037725
transform 1 0 47288 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1676037725
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1676037725
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_103
timestamp 1676037725
transform 1 0 10580 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_126
timestamp 1676037725
transform 1 0 12696 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_147
timestamp 1676037725
transform 1 0 14628 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1676037725
transform 1 0 14996 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1676037725
transform 1 0 16008 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1676037725
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_200
timestamp 1676037725
transform 1 0 19504 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_211
timestamp 1676037725
transform 1 0 20516 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_224
timestamp 1676037725
transform 1 0 21712 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_237
timestamp 1676037725
transform 1 0 22908 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_256
timestamp 1676037725
transform 1 0 24656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_267
timestamp 1676037725
transform 1 0 25668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_274
timestamp 1676037725
transform 1 0 26312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_280
timestamp 1676037725
transform 1 0 26864 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_292
timestamp 1676037725
transform 1 0 27968 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_295
timestamp 1676037725
transform 1 0 28244 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1676037725
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_320
timestamp 1676037725
transform 1 0 30544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_324
timestamp 1676037725
transform 1 0 30912 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_346
timestamp 1676037725
transform 1 0 32936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_359
timestamp 1676037725
transform 1 0 34132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1676037725
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_376
timestamp 1676037725
transform 1 0 35696 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_382
timestamp 1676037725
transform 1 0 36248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_404
timestamp 1676037725
transform 1 0 38272 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_408
timestamp 1676037725
transform 1 0 38640 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_416
timestamp 1676037725
transform 1 0 39376 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_433
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_440
timestamp 1676037725
transform 1 0 41584 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_452
timestamp 1676037725
transform 1 0 42688 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_464
timestamp 1676037725
transform 1 0 43792 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1676037725
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_29
timestamp 1676037725
transform 1 0 3772 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1676037725
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1676037725
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1676037725
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_97
timestamp 1676037725
transform 1 0 10028 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_124
timestamp 1676037725
transform 1 0 12512 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_128
timestamp 1676037725
transform 1 0 12880 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_155
timestamp 1676037725
transform 1 0 15364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_172
timestamp 1676037725
transform 1 0 16928 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_183
timestamp 1676037725
transform 1 0 17940 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_196
timestamp 1676037725
transform 1 0 19136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 1676037725
transform 1 0 19504 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_247
timestamp 1676037725
transform 1 0 23828 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_254
timestamp 1676037725
transform 1 0 24472 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1676037725
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_303
timestamp 1676037725
transform 1 0 28980 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_327
timestamp 1676037725
transform 1 0 31188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1676037725
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_359
timestamp 1676037725
transform 1 0 34132 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_372
timestamp 1676037725
transform 1 0 35328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_385
timestamp 1676037725
transform 1 0 36524 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1676037725
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_404
timestamp 1676037725
transform 1 0 38272 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_408
timestamp 1676037725
transform 1 0 38640 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_413
timestamp 1676037725
transform 1 0 39100 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_425
timestamp 1676037725
transform 1 0 40204 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_437
timestamp 1676037725
transform 1 0 41308 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_445
timestamp 1676037725
transform 1 0 42044 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1676037725
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_473
timestamp 1676037725
transform 1 0 44620 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_480
timestamp 1676037725
transform 1 0 45264 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_487
timestamp 1676037725
transform 1 0 45908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_499
timestamp 1676037725
transform 1 0 47012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1676037725
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_509
timestamp 1676037725
transform 1 0 47932 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_512
timestamp 1676037725
transform 1 0 48208 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_517
timestamp 1676037725
transform 1 0 48668 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1676037725
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1676037725
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_95
timestamp 1676037725
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_103
timestamp 1676037725
transform 1 0 10580 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_107
timestamp 1676037725
transform 1 0 10948 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_112
timestamp 1676037725
transform 1 0 11408 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_125
timestamp 1676037725
transform 1 0 12604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1676037725
transform 1 0 15272 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_158
timestamp 1676037725
transform 1 0 15640 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_162
timestamp 1676037725
transform 1 0 16008 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_175
timestamp 1676037725
transform 1 0 17204 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_183
timestamp 1676037725
transform 1 0 17940 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1676037725
transform 1 0 20884 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_238
timestamp 1676037725
transform 1 0 23000 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_242
timestamp 1676037725
transform 1 0 23368 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_245
timestamp 1676037725
transform 1 0 23644 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_257
timestamp 1676037725
transform 1 0 24748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_262
timestamp 1676037725
transform 1 0 25208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_286
timestamp 1676037725
transform 1 0 27416 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_299
timestamp 1676037725
transform 1 0 28612 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1676037725
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_320
timestamp 1676037725
transform 1 0 30544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_333
timestamp 1676037725
transform 1 0 31740 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_346
timestamp 1676037725
transform 1 0 32936 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_359
timestamp 1676037725
transform 1 0 34132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1676037725
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_387
timestamp 1676037725
transform 1 0 36708 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_411
timestamp 1676037725
transform 1 0 38916 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1676037725
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_425
timestamp 1676037725
transform 1 0 40204 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_437
timestamp 1676037725
transform 1 0 41308 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_449
timestamp 1676037725
transform 1 0 42412 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_461
timestamp 1676037725
transform 1 0 43516 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_473
timestamp 1676037725
transform 1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1676037725
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1676037725
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_513
timestamp 1676037725
transform 1 0 48300 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_519
timestamp 1676037725
transform 1 0 48852 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1676037725
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_21
timestamp 1676037725
transform 1 0 3036 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_33
timestamp 1676037725
transform 1 0 4140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_45
timestamp 1676037725
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1676037725
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_89
timestamp 1676037725
transform 1 0 9292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_99
timestamp 1676037725
transform 1 0 10212 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_104
timestamp 1676037725
transform 1 0 10672 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_115
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_126
timestamp 1676037725
transform 1 0 12696 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_130
timestamp 1676037725
transform 1 0 13064 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_153
timestamp 1676037725
transform 1 0 15180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_180
timestamp 1676037725
transform 1 0 17664 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_185
timestamp 1676037725
transform 1 0 18124 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_196
timestamp 1676037725
transform 1 0 19136 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_209
timestamp 1676037725
transform 1 0 20332 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_229
timestamp 1676037725
transform 1 0 22172 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_246
timestamp 1676037725
transform 1 0 23736 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_259
timestamp 1676037725
transform 1 0 24932 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_267
timestamp 1676037725
transform 1 0 25668 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1676037725
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_289
timestamp 1676037725
transform 1 0 27692 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_312
timestamp 1676037725
transform 1 0 29808 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_325
timestamp 1676037725
transform 1 0 31004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_332
timestamp 1676037725
transform 1 0 31648 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_348
timestamp 1676037725
transform 1 0 33120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_361
timestamp 1676037725
transform 1 0 34316 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_374
timestamp 1676037725
transform 1 0 35512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_387
timestamp 1676037725
transform 1 0 36708 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1676037725
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_415
timestamp 1676037725
transform 1 0 39284 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_428
timestamp 1676037725
transform 1 0 40480 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_435
timestamp 1676037725
transform 1 0 41124 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1676037725
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1676037725
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1676037725
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1676037725
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1676037725
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_519
timestamp 1676037725
transform 1 0 48852 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1676037725
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1676037725
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_61
timestamp 1676037725
transform 1 0 6716 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_73
timestamp 1676037725
transform 1 0 7820 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1676037725
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_87
timestamp 1676037725
transform 1 0 9108 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_99
timestamp 1676037725
transform 1 0 10212 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_103
timestamp 1676037725
transform 1 0 10580 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_125
timestamp 1676037725
transform 1 0 12604 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_152
timestamp 1676037725
transform 1 0 15088 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_156
timestamp 1676037725
transform 1 0 15456 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_166
timestamp 1676037725
transform 1 0 16376 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_179
timestamp 1676037725
transform 1 0 17572 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_185
timestamp 1676037725
transform 1 0 18124 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_191
timestamp 1676037725
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_201
timestamp 1676037725
transform 1 0 19596 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_213
timestamp 1676037725
transform 1 0 20700 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_217
timestamp 1676037725
transform 1 0 21068 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_227
timestamp 1676037725
transform 1 0 21988 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_233
timestamp 1676037725
transform 1 0 22540 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1676037725
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_265
timestamp 1676037725
transform 1 0 25484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_278
timestamp 1676037725
transform 1 0 26680 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_284
timestamp 1676037725
transform 1 0 27232 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_295
timestamp 1676037725
transform 1 0 28244 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_301
timestamp 1676037725
transform 1 0 28796 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_315
timestamp 1676037725
transform 1 0 30084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_339
timestamp 1676037725
transform 1 0 32292 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_352
timestamp 1676037725
transform 1 0 33488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_359
timestamp 1676037725
transform 1 0 34132 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1676037725
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_387
timestamp 1676037725
transform 1 0 36708 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_394
timestamp 1676037725
transform 1 0 37352 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_418
timestamp 1676037725
transform 1 0 39560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_443
timestamp 1676037725
transform 1 0 41860 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_447
timestamp 1676037725
transform 1 0 42228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_459
timestamp 1676037725
transform 1 0 43332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_471
timestamp 1676037725
transform 1 0 44436 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1676037725
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1676037725
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1676037725
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_513
timestamp 1676037725
transform 1 0 48300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_517
timestamp 1676037725
transform 1 0 48668 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_520
timestamp 1676037725
transform 1 0 48944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1676037725
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1676037725
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1676037725
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1676037725
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1676037725
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_73
timestamp 1676037725
transform 1 0 7820 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1676037725
transform 1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_91
timestamp 1676037725
transform 1 0 9476 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_99
timestamp 1676037725
transform 1 0 10212 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_104
timestamp 1676037725
transform 1 0 10672 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_116
timestamp 1676037725
transform 1 0 11776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_127
timestamp 1676037725
transform 1 0 12788 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_140
timestamp 1676037725
transform 1 0 13984 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1676037725
transform 1 0 15180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1676037725
transform 1 0 17204 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_186
timestamp 1676037725
transform 1 0 18216 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_194
timestamp 1676037725
transform 1 0 18952 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1676037725
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_233
timestamp 1676037725
transform 1 0 22540 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_237
timestamp 1676037725
transform 1 0 22908 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_248
timestamp 1676037725
transform 1 0 23920 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_254
timestamp 1676037725
transform 1 0 24472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_275
timestamp 1676037725
transform 1 0 26404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1676037725
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_292
timestamp 1676037725
transform 1 0 27968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_316
timestamp 1676037725
transform 1 0 30176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_329
timestamp 1676037725
transform 1 0 31372 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1676037725
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_348
timestamp 1676037725
transform 1 0 33120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_361
timestamp 1676037725
transform 1 0 34316 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_367
timestamp 1676037725
transform 1 0 34868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1676037725
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_398
timestamp 1676037725
transform 1 0 37720 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_402
timestamp 1676037725
transform 1 0 38088 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_423
timestamp 1676037725
transform 1 0 40020 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_427
timestamp 1676037725
transform 1 0 40388 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_437
timestamp 1676037725
transform 1 0 41308 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1676037725
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1676037725
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1676037725
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1676037725
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1676037725
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1676037725
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1676037725
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_519
timestamp 1676037725
transform 1 0 48852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1676037725
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_71
timestamp 1676037725
transform 1 0 7636 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1676037725
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_87
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_95
timestamp 1676037725
transform 1 0 9844 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_98
timestamp 1676037725
transform 1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_104
timestamp 1676037725
transform 1 0 10672 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_117
timestamp 1676037725
transform 1 0 11868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_125
timestamp 1676037725
transform 1 0 12604 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_143
timestamp 1676037725
transform 1 0 14260 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1676037725
transform 1 0 15272 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_167
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_171
timestamp 1676037725
transform 1 0 16836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_202
timestamp 1676037725
transform 1 0 19688 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_213
timestamp 1676037725
transform 1 0 20700 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_236
timestamp 1676037725
transform 1 0 22816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_240
timestamp 1676037725
transform 1 0 23184 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_258
timestamp 1676037725
transform 1 0 24840 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_286
timestamp 1676037725
transform 1 0 27416 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_290
timestamp 1676037725
transform 1 0 27784 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_302
timestamp 1676037725
transform 1 0 28888 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_320
timestamp 1676037725
transform 1 0 30544 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_337
timestamp 1676037725
transform 1 0 32108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_358
timestamp 1676037725
transform 1 0 34040 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_378
timestamp 1676037725
transform 1 0 35880 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_391
timestamp 1676037725
transform 1 0 37076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_395
timestamp 1676037725
transform 1 0 37444 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1676037725
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_432
timestamp 1676037725
transform 1 0 40848 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_440
timestamp 1676037725
transform 1 0 41584 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_452
timestamp 1676037725
transform 1 0 42688 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_464
timestamp 1676037725
transform 1 0 43792 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1676037725
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1676037725
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_513
timestamp 1676037725
transform 1 0 48300 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_519
timestamp 1676037725
transform 1 0 48852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1676037725
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_21
timestamp 1676037725
transform 1 0 3036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_33
timestamp 1676037725
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_45
timestamp 1676037725
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1676037725
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_89
timestamp 1676037725
transform 1 0 9292 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_99
timestamp 1676037725
transform 1 0 10212 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_119
timestamp 1676037725
transform 1 0 12052 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_124
timestamp 1676037725
transform 1 0 12512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_135
timestamp 1676037725
transform 1 0 13524 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_139
timestamp 1676037725
transform 1 0 13892 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_145
timestamp 1676037725
transform 1 0 14444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_153
timestamp 1676037725
transform 1 0 15180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1676037725
transform 1 0 17204 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1676037725
transform 1 0 17572 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_192
timestamp 1676037725
transform 1 0 18768 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_216
timestamp 1676037725
transform 1 0 20976 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_220
timestamp 1676037725
transform 1 0 21344 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_230
timestamp 1676037725
transform 1 0 22264 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_254
timestamp 1676037725
transform 1 0 24472 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_267
timestamp 1676037725
transform 1 0 25668 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_271
timestamp 1676037725
transform 1 0 26036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1676037725
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_294
timestamp 1676037725
transform 1 0 28152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_298
timestamp 1676037725
transform 1 0 28520 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_308
timestamp 1676037725
transform 1 0 29440 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_321
timestamp 1676037725
transform 1 0 30636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_360
timestamp 1676037725
transform 1 0 34224 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_375
timestamp 1676037725
transform 1 0 35604 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_388
timestamp 1676037725
transform 1 0 36800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_404
timestamp 1676037725
transform 1 0 38272 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_408
timestamp 1676037725
transform 1 0 38640 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_431
timestamp 1676037725
transform 1 0 40756 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_435
timestamp 1676037725
transform 1 0 41124 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1676037725
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1676037725
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1676037725
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1676037725
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1676037725
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_513
timestamp 1676037725
transform 1 0 48300 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_517
timestamp 1676037725
transform 1 0 48668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1676037725
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1676037725
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_101
timestamp 1676037725
transform 1 0 10396 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_123
timestamp 1676037725
transform 1 0 12420 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_127
timestamp 1676037725
transform 1 0 12788 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_131
timestamp 1676037725
transform 1 0 13156 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_163
timestamp 1676037725
transform 1 0 16100 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_168
timestamp 1676037725
transform 1 0 16560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_179
timestamp 1676037725
transform 1 0 17572 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_202
timestamp 1676037725
transform 1 0 19688 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_228
timestamp 1676037725
transform 1 0 22080 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_232
timestamp 1676037725
transform 1 0 22448 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_237
timestamp 1676037725
transform 1 0 22908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_264
timestamp 1676037725
transform 1 0 25392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_271
timestamp 1676037725
transform 1 0 26036 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_277
timestamp 1676037725
transform 1 0 26588 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_281
timestamp 1676037725
transform 1 0 26956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_302
timestamp 1676037725
transform 1 0 28888 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_311
timestamp 1676037725
transform 1 0 29716 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_324
timestamp 1676037725
transform 1 0 30912 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_337
timestamp 1676037725
transform 1 0 32108 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_341
timestamp 1676037725
transform 1 0 32476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_353
timestamp 1676037725
transform 1 0 33580 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_359
timestamp 1676037725
transform 1 0 34132 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_370
timestamp 1676037725
transform 1 0 35144 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_374
timestamp 1676037725
transform 1 0 35512 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_397
timestamp 1676037725
transform 1 0 37628 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_410
timestamp 1676037725
transform 1 0 38824 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_416
timestamp 1676037725
transform 1 0 39376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_427
timestamp 1676037725
transform 1 0 40388 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_437
timestamp 1676037725
transform 1 0 41308 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_449
timestamp 1676037725
transform 1 0 42412 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_461
timestamp 1676037725
transform 1 0 43516 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_473
timestamp 1676037725
transform 1 0 44620 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1676037725
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1676037725
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_513
timestamp 1676037725
transform 1 0 48300 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_519
timestamp 1676037725
transform 1 0 48852 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1676037725
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_21
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_28
timestamp 1676037725
transform 1 0 3680 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_32
timestamp 1676037725
transform 1 0 4048 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1676037725
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_75
timestamp 1676037725
transform 1 0 8004 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_87
timestamp 1676037725
transform 1 0 9108 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_97
timestamp 1676037725
transform 1 0 10028 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_135
timestamp 1676037725
transform 1 0 13524 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_148
timestamp 1676037725
transform 1 0 14720 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_154
timestamp 1676037725
transform 1 0 15272 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_159
timestamp 1676037725
transform 1 0 15732 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_173
timestamp 1676037725
transform 1 0 17020 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_179
timestamp 1676037725
transform 1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_192
timestamp 1676037725
transform 1 0 18768 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_196
timestamp 1676037725
transform 1 0 19136 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_199
timestamp 1676037725
transform 1 0 19412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_252
timestamp 1676037725
transform 1 0 24288 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_265
timestamp 1676037725
transform 1 0 25484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1676037725
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_292
timestamp 1676037725
transform 1 0 27968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_305
timestamp 1676037725
transform 1 0 29164 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_313
timestamp 1676037725
transform 1 0 29900 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_324
timestamp 1676037725
transform 1 0 30912 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_331
timestamp 1676037725
transform 1 0 31556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1676037725
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_348
timestamp 1676037725
transform 1 0 33120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_352
timestamp 1676037725
transform 1 0 33488 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_373
timestamp 1676037725
transform 1 0 35420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_377
timestamp 1676037725
transform 1 0 35788 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_387
timestamp 1676037725
transform 1 0 36708 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1676037725
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_399
timestamp 1676037725
transform 1 0 37812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_421
timestamp 1676037725
transform 1 0 39836 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_425
timestamp 1676037725
transform 1 0 40204 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_436
timestamp 1676037725
transform 1 0 41216 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1676037725
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1676037725
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1676037725
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1676037725
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1676037725
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_513
timestamp 1676037725
transform 1 0 48300 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_519
timestamp 1676037725
transform 1 0 48852 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1676037725
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1676037725
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_47
timestamp 1676037725
transform 1 0 5428 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_59
timestamp 1676037725
transform 1 0 6532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_71
timestamp 1676037725
transform 1 0 7636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_75
timestamp 1676037725
transform 1 0 8004 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1676037725
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_108
timestamp 1676037725
transform 1 0 11040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_112
timestamp 1676037725
transform 1 0 11408 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_115
timestamp 1676037725
transform 1 0 11684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_120
timestamp 1676037725
transform 1 0 12144 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_163
timestamp 1676037725
transform 1 0 16100 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_167
timestamp 1676037725
transform 1 0 16468 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_170
timestamp 1676037725
transform 1 0 16744 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1676037725
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_199
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_202
timestamp 1676037725
transform 1 0 19688 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_213
timestamp 1676037725
transform 1 0 20700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_226
timestamp 1676037725
transform 1 0 21896 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_264
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_288
timestamp 1676037725
transform 1 0 27600 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_300
timestamp 1676037725
transform 1 0 28704 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1676037725
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_320
timestamp 1676037725
transform 1 0 30544 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_328
timestamp 1676037725
transform 1 0 31280 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_339
timestamp 1676037725
transform 1 0 32292 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_352
timestamp 1676037725
transform 1 0 33488 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_371
timestamp 1676037725
transform 1 0 35236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_395
timestamp 1676037725
transform 1 0 37444 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_399
timestamp 1676037725
transform 1 0 37812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_410
timestamp 1676037725
transform 1 0 38824 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_443
timestamp 1676037725
transform 1 0 41860 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_447
timestamp 1676037725
transform 1 0 42228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_459
timestamp 1676037725
transform 1 0 43332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_471
timestamp 1676037725
transform 1 0 44436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1676037725
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1676037725
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1676037725
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_513
timestamp 1676037725
transform 1 0 48300 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_517
timestamp 1676037725
transform 1 0 48668 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1676037725
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1676037725
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1676037725
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_49
timestamp 1676037725
transform 1 0 5612 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1676037725
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_96
timestamp 1676037725
transform 1 0 9936 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_103
timestamp 1676037725
transform 1 0 10580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_116
timestamp 1676037725
transform 1 0 11776 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1676037725
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_146
timestamp 1676037725
transform 1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_152
timestamp 1676037725
transform 1 0 15088 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_158
timestamp 1676037725
transform 1 0 15640 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_180
timestamp 1676037725
transform 1 0 17664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_207
timestamp 1676037725
transform 1 0 20148 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_211
timestamp 1676037725
transform 1 0 20516 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1676037725
transform 1 0 23000 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_242
timestamp 1676037725
transform 1 0 23368 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_263
timestamp 1676037725
transform 1 0 25300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_267
timestamp 1676037725
transform 1 0 25668 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1676037725
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_293
timestamp 1676037725
transform 1 0 28060 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_306
timestamp 1676037725
transform 1 0 29256 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_310
timestamp 1676037725
transform 1 0 29624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_314
timestamp 1676037725
transform 1 0 29992 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_320
timestamp 1676037725
transform 1 0 30544 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1676037725
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_348
timestamp 1676037725
transform 1 0 33120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_361
timestamp 1676037725
transform 1 0 34316 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_374
timestamp 1676037725
transform 1 0 35512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_387
timestamp 1676037725
transform 1 0 36708 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1676037725
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_397
timestamp 1676037725
transform 1 0 37628 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_420
timestamp 1676037725
transform 1 0 39744 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_433
timestamp 1676037725
transform 1 0 40940 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_439
timestamp 1676037725
transform 1 0 41492 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1676037725
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1676037725
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1676037725
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1676037725
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1676037725
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1676037725
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_513
timestamp 1676037725
transform 1 0 48300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_519
timestamp 1676037725
transform 1 0 48852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1676037725
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1676037725
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_47
timestamp 1676037725
transform 1 0 5428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_67
timestamp 1676037725
transform 1 0 7268 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_71
timestamp 1676037725
transform 1 0 7636 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_75
timestamp 1676037725
transform 1 0 8004 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_93
timestamp 1676037725
transform 1 0 9660 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_99
timestamp 1676037725
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_106
timestamp 1676037725
transform 1 0 10856 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1676037725
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1676037725
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_154
timestamp 1676037725
transform 1 0 15272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_167
timestamp 1676037725
transform 1 0 16468 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1676037725
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_184
timestamp 1676037725
transform 1 0 18032 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_199
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_205
timestamp 1676037725
transform 1 0 19964 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1676037725
transform 1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_231
timestamp 1676037725
transform 1 0 22356 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_239
timestamp 1676037725
transform 1 0 23092 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_258
timestamp 1676037725
transform 1 0 24840 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_264
timestamp 1676037725
transform 1 0 25392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_275
timestamp 1676037725
transform 1 0 26404 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_288
timestamp 1676037725
transform 1 0 27600 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_301
timestamp 1676037725
transform 1 0 28796 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_305
timestamp 1676037725
transform 1 0 29164 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_320
timestamp 1676037725
transform 1 0 30544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_333
timestamp 1676037725
transform 1 0 31740 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_346
timestamp 1676037725
transform 1 0 32936 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_350
timestamp 1676037725
transform 1 0 33304 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_360
timestamp 1676037725
transform 1 0 34224 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_376
timestamp 1676037725
transform 1 0 35696 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_389
timestamp 1676037725
transform 1 0 36892 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_397
timestamp 1676037725
transform 1 0 37628 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_408
timestamp 1676037725
transform 1 0 38640 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_414
timestamp 1676037725
transform 1 0 39192 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_432
timestamp 1676037725
transform 1 0 40848 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_438
timestamp 1676037725
transform 1 0 41400 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_450
timestamp 1676037725
transform 1 0 42504 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_462
timestamp 1676037725
transform 1 0 43608 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_474
timestamp 1676037725
transform 1 0 44712 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1676037725
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1676037725
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_513
timestamp 1676037725
transform 1 0 48300 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_519
timestamp 1676037725
transform 1 0 48852 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1676037725
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_21
timestamp 1676037725
transform 1 0 3036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_41
timestamp 1676037725
transform 1 0 4876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_48
timestamp 1676037725
transform 1 0 5520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_75
timestamp 1676037725
transform 1 0 8004 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_83
timestamp 1676037725
transform 1 0 8740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_89
timestamp 1676037725
transform 1 0 9292 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_96
timestamp 1676037725
transform 1 0 9936 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_103
timestamp 1676037725
transform 1 0 10580 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_119
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_127
timestamp 1676037725
transform 1 0 12788 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_135
timestamp 1676037725
transform 1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_146
timestamp 1676037725
transform 1 0 14536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_153
timestamp 1676037725
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1676037725
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_171
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_193
timestamp 1676037725
transform 1 0 18860 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_199
timestamp 1676037725
transform 1 0 19412 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_236
timestamp 1676037725
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_243
timestamp 1676037725
transform 1 0 23460 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_267
timestamp 1676037725
transform 1 0 25668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_274
timestamp 1676037725
transform 1 0 26312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1676037725
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_304
timestamp 1676037725
transform 1 0 29072 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_317
timestamp 1676037725
transform 1 0 30268 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_330
timestamp 1676037725
transform 1 0 31464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_359
timestamp 1676037725
transform 1 0 34132 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_372
timestamp 1676037725
transform 1 0 35328 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_378
timestamp 1676037725
transform 1 0 35880 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1676037725
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_395
timestamp 1676037725
transform 1 0 37444 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_418
timestamp 1676037725
transform 1 0 39560 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_431
timestamp 1676037725
transform 1 0 40756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_438
timestamp 1676037725
transform 1 0 41400 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_444
timestamp 1676037725
transform 1 0 41952 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1676037725
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1676037725
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1676037725
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1676037725
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1676037725
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_513
timestamp 1676037725
transform 1 0 48300 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_517
timestamp 1676037725
transform 1 0 48668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1676037725
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1676037725
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1676037725
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_67
timestamp 1676037725
transform 1 0 7268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_71
timestamp 1676037725
transform 1 0 7636 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_76
timestamp 1676037725
transform 1 0 8096 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1676037725
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_91
timestamp 1676037725
transform 1 0 9476 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_98
timestamp 1676037725
transform 1 0 10120 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_105
timestamp 1676037725
transform 1 0 10764 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_112
timestamp 1676037725
transform 1 0 11408 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_120
timestamp 1676037725
transform 1 0 12144 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_124
timestamp 1676037725
transform 1 0 12512 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_130
timestamp 1676037725
transform 1 0 13064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_134
timestamp 1676037725
transform 1 0 13432 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_163
timestamp 1676037725
transform 1 0 16100 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_170
timestamp 1676037725
transform 1 0 16744 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_203
timestamp 1676037725
transform 1 0 19780 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_214
timestamp 1676037725
transform 1 0 20792 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_238
timestamp 1676037725
transform 1 0 23000 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_246
timestamp 1676037725
transform 1 0 23736 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_258
timestamp 1676037725
transform 1 0 24840 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_276
timestamp 1676037725
transform 1 0 26496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_282
timestamp 1676037725
transform 1 0 27048 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_287
timestamp 1676037725
transform 1 0 27508 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_292
timestamp 1676037725
transform 1 0 27968 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1676037725
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_314
timestamp 1676037725
transform 1 0 29992 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_320
timestamp 1676037725
transform 1 0 30544 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_332
timestamp 1676037725
transform 1 0 31648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_336
timestamp 1676037725
transform 1 0 32016 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_340
timestamp 1676037725
transform 1 0 32384 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1676037725
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_387
timestamp 1676037725
transform 1 0 36708 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_395
timestamp 1676037725
transform 1 0 37444 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_417
timestamp 1676037725
transform 1 0 39468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_432
timestamp 1676037725
transform 1 0 40848 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_445
timestamp 1676037725
transform 1 0 42044 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1676037725
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1676037725
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1676037725
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1676037725
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_501
timestamp 1676037725
transform 1 0 47196 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_507
timestamp 1676037725
transform 1 0 47748 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_512
timestamp 1676037725
transform 1 0 48208 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_519
timestamp 1676037725
transform 1 0 48852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_525
timestamp 1676037725
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1676037725
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_41
timestamp 1676037725
transform 1 0 4876 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_49
timestamp 1676037725
transform 1 0 5612 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1676037725
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_75
timestamp 1676037725
transform 1 0 8004 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_95
timestamp 1676037725
transform 1 0 9844 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_101
timestamp 1676037725
transform 1 0 10396 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1676037725
transform 1 0 11960 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_124
timestamp 1676037725
transform 1 0 12512 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_128
timestamp 1676037725
transform 1 0 12880 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_134
timestamp 1676037725
transform 1 0 13432 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_138
timestamp 1676037725
transform 1 0 13800 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_142
timestamp 1676037725
transform 1 0 14168 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_175
timestamp 1676037725
transform 1 0 17204 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_186
timestamp 1676037725
transform 1 0 18216 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_210
timestamp 1676037725
transform 1 0 20424 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_216
timestamp 1676037725
transform 1 0 20976 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_230
timestamp 1676037725
transform 1 0 22264 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_253
timestamp 1676037725
transform 1 0 24380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_266
timestamp 1676037725
transform 1 0 25576 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_272
timestamp 1676037725
transform 1 0 26128 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_292
timestamp 1676037725
transform 1 0 27968 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_305
timestamp 1676037725
transform 1 0 29164 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_318
timestamp 1676037725
transform 1 0 30360 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_331
timestamp 1676037725
transform 1 0 31556 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1676037725
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_341
timestamp 1676037725
transform 1 0 32476 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_345
timestamp 1676037725
transform 1 0 32844 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_358
timestamp 1676037725
transform 1 0 34040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_371
timestamp 1676037725
transform 1 0 35236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_375
timestamp 1676037725
transform 1 0 35604 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_385
timestamp 1676037725
transform 1 0 36524 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1676037725
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_399
timestamp 1676037725
transform 1 0 37812 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_421
timestamp 1676037725
transform 1 0 39836 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_431
timestamp 1676037725
transform 1 0 40756 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_434
timestamp 1676037725
transform 1 0 41032 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1676037725
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_461
timestamp 1676037725
transform 1 0 43516 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_466
timestamp 1676037725
transform 1 0 43976 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_478
timestamp 1676037725
transform 1 0 45080 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_490
timestamp 1676037725
transform 1 0 46184 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_502
timestamp 1676037725
transform 1 0 47288 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_505
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_510
timestamp 1676037725
transform 1 0 48024 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_517
timestamp 1676037725
transform 1 0 48668 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1676037725
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1676037725
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_47
timestamp 1676037725
transform 1 0 5428 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_67
timestamp 1676037725
transform 1 0 7268 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_75
timestamp 1676037725
transform 1 0 8004 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1676037725
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_103
timestamp 1676037725
transform 1 0 10580 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_107
timestamp 1676037725
transform 1 0 10948 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1676037725
transform 1 0 11960 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_125
timestamp 1676037725
transform 1 0 12604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_143
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_149
timestamp 1676037725
transform 1 0 14812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_173
timestamp 1676037725
transform 1 0 17020 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1676037725
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_215
timestamp 1676037725
transform 1 0 20884 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_219
timestamp 1676037725
transform 1 0 21252 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_230
timestamp 1676037725
transform 1 0 22264 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_243
timestamp 1676037725
transform 1 0 23460 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1676037725
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_268
timestamp 1676037725
transform 1 0 25760 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_279
timestamp 1676037725
transform 1 0 26772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_292
timestamp 1676037725
transform 1 0 27968 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_305
timestamp 1676037725
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_314
timestamp 1676037725
transform 1 0 29992 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_320
timestamp 1676037725
transform 1 0 30544 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_343
timestamp 1676037725
transform 1 0 32660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_356
timestamp 1676037725
transform 1 0 33856 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_376
timestamp 1676037725
transform 1 0 35696 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_389
timestamp 1676037725
transform 1 0 36892 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_414
timestamp 1676037725
transform 1 0 39192 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_423
timestamp 1676037725
transform 1 0 40020 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_434
timestamp 1676037725
transform 1 0 41032 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_447
timestamp 1676037725
transform 1 0 42228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_454
timestamp 1676037725
transform 1 0 42872 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_468
timestamp 1676037725
transform 1 0 44160 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_489
timestamp 1676037725
transform 1 0 46092 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_495
timestamp 1676037725
transform 1 0 46644 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_504
timestamp 1676037725
transform 1 0 47472 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_509
timestamp 1676037725
transform 1 0 47932 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_517
timestamp 1676037725
transform 1 0 48668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_21
timestamp 1676037725
transform 1 0 3036 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_29
timestamp 1676037725
transform 1 0 3772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1676037725
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_63
timestamp 1676037725
transform 1 0 6900 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_67
timestamp 1676037725
transform 1 0 7268 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_85
timestamp 1676037725
transform 1 0 8924 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_92
timestamp 1676037725
transform 1 0 9568 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_119
timestamp 1676037725
transform 1 0 12052 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_123
timestamp 1676037725
transform 1 0 12420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_141
timestamp 1676037725
transform 1 0 14076 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_148
timestamp 1676037725
transform 1 0 14720 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_191
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_197
timestamp 1676037725
transform 1 0 19228 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_220
timestamp 1676037725
transform 1 0 21344 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_248
timestamp 1676037725
transform 1 0 23920 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_256
timestamp 1676037725
transform 1 0 24656 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1676037725
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_286
timestamp 1676037725
transform 1 0 27416 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_290
timestamp 1676037725
transform 1 0 27784 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_313
timestamp 1676037725
transform 1 0 29900 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_326
timestamp 1676037725
transform 1 0 31096 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_333
timestamp 1676037725
transform 1 0 31740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_348
timestamp 1676037725
transform 1 0 33120 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_352
timestamp 1676037725
transform 1 0 33488 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_374
timestamp 1676037725
transform 1 0 35512 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_378
timestamp 1676037725
transform 1 0 35880 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_389
timestamp 1676037725
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_415
timestamp 1676037725
transform 1 0 39284 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_421
timestamp 1676037725
transform 1 0 39836 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_432
timestamp 1676037725
transform 1 0 40848 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_439
timestamp 1676037725
transform 1 0 41492 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_446
timestamp 1676037725
transform 1 0 42136 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_461
timestamp 1676037725
transform 1 0 43516 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_468
timestamp 1676037725
transform 1 0 44160 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_475
timestamp 1676037725
transform 1 0 44804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_482
timestamp 1676037725
transform 1 0 45448 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_488
timestamp 1676037725
transform 1 0 46000 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_497
timestamp 1676037725
transform 1 0 46828 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_502
timestamp 1676037725
transform 1 0 47288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_511
timestamp 1676037725
transform 1 0 48116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_517
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1676037725
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1676037725
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_35
timestamp 1676037725
transform 1 0 4324 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1676037725
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1676037725
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1676037725
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_91
timestamp 1676037725
transform 1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_98
timestamp 1676037725
transform 1 0 10120 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_118
timestamp 1676037725
transform 1 0 11960 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_145
timestamp 1676037725
transform 1 0 14444 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_150
timestamp 1676037725
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1676037725
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_199
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_205
timestamp 1676037725
transform 1 0 19964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_229
timestamp 1676037725
transform 1 0 22172 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_237
timestamp 1676037725
transform 1 0 22908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_259
timestamp 1676037725
transform 1 0 24932 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_265
timestamp 1676037725
transform 1 0 25484 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_287
timestamp 1676037725
transform 1 0 27508 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_300
timestamp 1676037725
transform 1 0 28704 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_320
timestamp 1676037725
transform 1 0 30544 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_324
timestamp 1676037725
transform 1 0 30912 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_327
timestamp 1676037725
transform 1 0 31188 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_350
timestamp 1676037725
transform 1 0 33304 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_357
timestamp 1676037725
transform 1 0 33948 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1676037725
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_367
timestamp 1676037725
transform 1 0 34868 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_389
timestamp 1676037725
transform 1 0 36892 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_413
timestamp 1676037725
transform 1 0 39100 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1676037725
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_432
timestamp 1676037725
transform 1 0 40848 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_436
timestamp 1676037725
transform 1 0 41216 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_462
timestamp 1676037725
transform 1 0 43608 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_466
timestamp 1676037725
transform 1 0 43976 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_472
timestamp 1676037725
transform 1 0 44528 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_477
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_482
timestamp 1676037725
transform 1 0 45448 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_486
timestamp 1676037725
transform 1 0 45816 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_492
timestamp 1676037725
transform 1 0 46368 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_496
timestamp 1676037725
transform 1 0 46736 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_501
timestamp 1676037725
transform 1 0 47196 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_509
timestamp 1676037725
transform 1 0 47932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_517
timestamp 1676037725
transform 1 0 48668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1676037725
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1676037725
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1676037725
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_63
timestamp 1676037725
transform 1 0 6900 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1676037725
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1676037725
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1676037725
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_126
timestamp 1676037725
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1676037725
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_188
timestamp 1676037725
transform 1 0 18400 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_212
timestamp 1676037725
transform 1 0 20608 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_217
timestamp 1676037725
transform 1 0 21068 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_237
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_250
timestamp 1676037725
transform 1 0 24104 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_256
timestamp 1676037725
transform 1 0 24656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1676037725
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_286
timestamp 1676037725
transform 1 0 27416 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_300
timestamp 1676037725
transform 1 0 28704 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_307
timestamp 1676037725
transform 1 0 29348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_311
timestamp 1676037725
transform 1 0 29716 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1676037725
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_348
timestamp 1676037725
transform 1 0 33120 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_352
timestamp 1676037725
transform 1 0 33488 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_373
timestamp 1676037725
transform 1 0 35420 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_377
timestamp 1676037725
transform 1 0 35788 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_387
timestamp 1676037725
transform 1 0 36708 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1676037725
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_404
timestamp 1676037725
transform 1 0 38272 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_408
timestamp 1676037725
transform 1 0 38640 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_419
timestamp 1676037725
transform 1 0 39652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_426
timestamp 1676037725
transform 1 0 40296 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_440
timestamp 1676037725
transform 1 0 41584 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_453
timestamp 1676037725
transform 1 0 42780 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_476
timestamp 1676037725
transform 1 0 44896 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_488
timestamp 1676037725
transform 1 0 46000 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_494
timestamp 1676037725
transform 1 0 46552 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_500
timestamp 1676037725
transform 1 0 47104 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_509
timestamp 1676037725
transform 1 0 47932 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_520
timestamp 1676037725
transform 1 0 48944 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_526
timestamp 1676037725
transform 1 0 49496 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1676037725
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1676037725
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1676037725
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1676037725
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1676037725
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1676037725
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1676037725
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1676037725
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1676037725
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1676037725
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_174
timestamp 1676037725
transform 1 0 17112 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1676037725
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1676037725
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_225
timestamp 1676037725
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_243
timestamp 1676037725
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_272
timestamp 1676037725
transform 1 0 26128 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_281
timestamp 1676037725
transform 1 0 26956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_287
timestamp 1676037725
transform 1 0 27508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_294
timestamp 1676037725
transform 1 0 28152 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_301
timestamp 1676037725
transform 1 0 28796 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1676037725
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_314
timestamp 1676037725
transform 1 0 29992 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_321
timestamp 1676037725
transform 1 0 30636 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_328
timestamp 1676037725
transform 1 0 31280 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1676037725
transform 1 0 32108 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_342
timestamp 1676037725
transform 1 0 32568 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_349
timestamp 1676037725
transform 1 0 33212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1676037725
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_376
timestamp 1676037725
transform 1 0 35696 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_389
timestamp 1676037725
transform 1 0 36892 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_393
timestamp 1676037725
transform 1 0 37260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_404
timestamp 1676037725
transform 1 0 38272 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_411
timestamp 1676037725
transform 1 0 38916 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_418
timestamp 1676037725
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_432
timestamp 1676037725
transform 1 0 40848 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_436
timestamp 1676037725
transform 1 0 41216 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_446
timestamp 1676037725
transform 1 0 42136 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_449
timestamp 1676037725
transform 1 0 42412 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_459
timestamp 1676037725
transform 1 0 43332 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_466
timestamp 1676037725
transform 1 0 43976 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_473
timestamp 1676037725
transform 1 0 44620 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_483
timestamp 1676037725
transform 1 0 45540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_491
timestamp 1676037725
transform 1 0 46276 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_499
timestamp 1676037725
transform 1 0 47012 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_503
timestamp 1676037725
transform 1 0 47380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_505
timestamp 1676037725
transform 1 0 47564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_511
timestamp 1676037725
transform 1 0 48116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_525
timestamp 1676037725
transform 1 0 49404 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 42136 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  hold2
timestamp 1676037725
transform -1 0 44896 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1676037725
transform -1 0 43332 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1676037725
transform -1 0 48944 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1676037725
transform -1 0 46000 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1676037725
transform 1 0 12328 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform -1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 46920 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform -1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input4 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1676037725
transform 1 0 1564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform -1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1676037725
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1676037725
transform -1 0 2484 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1676037725
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1676037725
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1676037725
transform -1 0 2484 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1676037725
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1676037725
transform 1 0 1564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform -1 0 2576 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1676037725
transform -1 0 2484 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1676037725
transform 1 0 1564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform -1 0 3128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1676037725
transform 1 0 1564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1676037725
transform 1 0 3404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1676037725
transform -1 0 2484 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input28
timestamp 1676037725
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 1676037725
transform 1 0 1564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1676037725
transform -1 0 2484 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1676037725
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 48392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1676037725
transform -1 0 49404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1676037725
transform -1 0 49404 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 48392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1676037725
transform -1 0 49404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1676037725
transform -1 0 49404 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1676037725
transform -1 0 49404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1676037725
transform 1 0 48392 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1676037725
transform -1 0 49404 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1676037725
transform -1 0 49404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1676037725
transform -1 0 49404 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1676037725
transform -1 0 49404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1676037725
transform 1 0 48392 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1676037725
transform -1 0 49404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1676037725
transform -1 0 49404 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1676037725
transform -1 0 48668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 47748 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1676037725
transform 1 0 46092 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1676037725
transform -1 0 48668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1676037725
transform 1 0 47656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 47012 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1676037725
transform 1 0 48484 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1676037725
transform -1 0 49404 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1676037725
transform -1 0 49404 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1676037725
transform 1 0 49128 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1676037725
transform -1 0 49404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1676037725
transform -1 0 49404 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1676037725
transform -1 0 49404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1676037725
transform 1 0 48392 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1676037725
transform -1 0 49404 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform -1 0 26312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1676037725
transform -1 0 29348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1676037725
transform -1 0 31280 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 32292 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1676037725
transform 1 0 32936 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1676037725
transform 1 0 38640 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1676037725
transform 1 0 33672 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1676037725
transform 1 0 39284 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1676037725
transform 1 0 43700 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1676037725
transform 1 0 40020 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1676037725
transform 1 0 44344 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1676037725
transform -1 0 11960 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1676037725
transform 1 0 41216 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1676037725
transform 1 0 40664 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1676037725
transform 1 0 42596 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input78
timestamp 1676037725
transform 1 0 43240 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1676037725
transform 1 0 42596 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1676037725
transform 1 0 41216 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1676037725
transform 1 0 44528 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1676037725
transform 1 0 41860 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1676037725
transform 1 0 45172 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1676037725
transform 1 0 43884 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input85
timestamp 1676037725
transform -1 0 12696 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input86
timestamp 1676037725
transform -1 0 22908 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1676037725
transform -1 0 24840 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1676037725
transform -1 0 30636 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1676037725
transform -1 0 24104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1676037725
transform -1 0 28152 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1676037725
transform -1 0 28060 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1676037725
transform -1 0 28796 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1676037725
transform 1 0 28980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1676037725
transform 1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1676037725
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1676037725
transform 1 0 35052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input97
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1676037725
transform 1 0 45172 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input99
timestamp 1676037725
transform 1 0 43516 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input100
timestamp 1676037725
transform -1 0 45724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1676037725
transform -1 0 47564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input102
timestamp 1676037725
transform -1 0 46828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1676037725
transform -1 0 46276 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input104
timestamp 1676037725
transform -1 0 47012 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input105
timestamp 1676037725
transform -1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input106
timestamp 1676037725
transform -1 0 47932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input107
timestamp 1676037725
transform -1 0 48116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input108
timestamp 1676037725
transform -1 0 48668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input109
timestamp 1676037725
transform -1 0 44528 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1676037725
transform -1 0 45540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output111 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40664 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform -1 0 4876 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform -1 0 3036 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform -1 0 3036 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform -1 0 3036 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform -1 0 3036 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform -1 0 3036 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform -1 0 3036 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform -1 0 3036 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform -1 0 4876 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform -1 0 3036 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform -1 0 3036 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform -1 0 3036 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform -1 0 3036 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform -1 0 5428 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform -1 0 5428 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform -1 0 7268 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform -1 0 7268 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform -1 0 5428 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform -1 0 7268 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 6532 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 8372 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 9108 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform -1 0 3036 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform -1 0 3036 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform -1 0 3036 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform -1 0 3036 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform -1 0 3036 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform -1 0 3036 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform -1 0 3036 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform -1 0 3036 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 45816 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 47932 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 47932 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 47932 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 47932 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 47932 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 45816 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1676037725
transform 1 0 47932 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1676037725
transform 1 0 47932 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1676037725
transform 1 0 47932 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1676037725
transform 1 0 43976 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1676037725
transform 1 0 46092 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1676037725
transform 1 0 47932 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1676037725
transform 1 0 47932 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1676037725
transform 1 0 47932 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1676037725
transform 1 0 47932 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1676037725
transform 1 0 47932 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1676037725
transform 1 0 47932 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1676037725
transform 1 0 47932 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1676037725
transform 1 0 47932 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1676037725
transform 1 0 47932 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1676037725
transform 1 0 45816 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1676037725
transform 1 0 45816 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1676037725
transform 1 0 47932 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1676037725
transform 1 0 47932 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1676037725
transform 1 0 47932 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1676037725
transform 1 0 45816 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1676037725
transform 1 0 47932 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1676037725
transform -1 0 5428 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1676037725
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1676037725
transform -1 0 9384 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1676037725
transform -1 0 11224 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1676037725
transform -1 0 11224 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1676037725
transform -1 0 11960 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1676037725
transform -1 0 11224 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1676037725
transform -1 0 14076 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1676037725
transform -1 0 13800 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1676037725
transform -1 0 13800 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1676037725
transform 1 0 13064 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1676037725
transform -1 0 4876 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1676037725
transform -1 0 16376 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1676037725
transform -1 0 16744 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1676037725
transform -1 0 16376 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1676037725
transform -1 0 18860 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1676037725
transform -1 0 16376 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1676037725
transform -1 0 18400 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1676037725
transform -1 0 18952 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1676037725
transform 1 0 21988 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1676037725
transform -1 0 21528 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1676037725
transform -1 0 3496 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1676037725
transform -1 0 4232 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1676037725
transform -1 0 6072 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1676037725
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1676037725
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1676037725
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output202
timestamp 1676037725
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output203
timestamp 1676037725
transform -1 0 13248 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output204
timestamp 1676037725
transform -1 0 15732 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output205
timestamp 1676037725
transform -1 0 18308 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output206
timestamp 1676037725
transform -1 0 19596 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output207
timestamp 1676037725
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output208
timestamp 1676037725
transform 1 0 22356 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output209
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output210
timestamp 1676037725
transform 1 0 27140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 29256 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 26404 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 24472 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 24104 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 22356 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17020 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18584 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 22080 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 18952 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19136 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 23828 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21068 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 22816 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 20976 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19596 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 21528 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 18952 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 22172 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 20608 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23828 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 25300 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25760 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 28888 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 27416 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27232 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 29900 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 26680 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25668 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 26680 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 23000 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22448 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28336 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 30452 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32200 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34868 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 36984 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34868 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 36432 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37444 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34868 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 35144 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 37812 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 33856 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34868 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 35696 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29992 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32108 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 32936 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27968 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29716 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 30360 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 26956 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 28796 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 32200 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 31096 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32292 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 32568 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29716 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 29348 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 26864 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 43608 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 30820 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 31832 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 31372 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 33672 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 35420 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35052 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 36708 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 34132 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32476 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 39284 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 39100 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 39192 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 37996 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 39468 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 39560 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 37628 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 33580 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35604 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 39744 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 39836 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 41860 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 40756 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 39560 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 38180 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 40020 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 39560 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37444 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 38916 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 34132 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 31188 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 27416 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 26680 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 25668 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23920 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 26404 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 25300 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 24104 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 23828 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 21528 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 21252 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 21252 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19320 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 22080 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 22264 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 18676 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 14904 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12972 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 16100 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 14536 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 13524 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 12420 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 16100 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 17020 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 18952 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30728 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27232 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_2_
timestamp 1676037725
transform -1 0 23460 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_1.mux_l1_in_3__258
timestamp 1676037725
transform 1 0 26036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_3_
timestamp 1676037725
transform -1 0 21712 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25852 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l2_in_1_
timestamp 1676037725
transform -1 0 23920 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19872 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_3.mux_l2_in_1__211
timestamp 1676037725
transform -1 0 15732 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l2_in_1_
timestamp 1676037725
transform -1 0 17572 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 16836 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9936 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25576 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24656 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_5.mux_l2_in_1__214
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18308 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l3_in_0_
timestamp 1676037725
transform 1 0 17388 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24656 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_2_
timestamp 1676037725
transform -1 0 20332 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23092 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l2_in_1_
timestamp 1676037725
transform -1 0 20516 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_7.mux_l2_in_1__216
timestamp 1676037725
transform -1 0 18952 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19872 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 17204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27968 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25760 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_2_
timestamp 1676037725
transform 1 0 20884 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_11.mux_l1_in_3__259
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_3_
timestamp 1676037725
transform 1 0 20700 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22080 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19504 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l3_in_0_
timestamp 1676037725
transform 1 0 17940 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24748 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_2_
timestamp 1676037725
transform 1 0 21160 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_13.mux_l2_in_1__260
timestamp 1676037725
transform -1 0 16744 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18124 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15640 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10580 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27876 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_2_
timestamp 1676037725
transform 1 0 21068 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_21.mux_l2_in_1__261
timestamp 1676037725
transform -1 0 17112 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18124 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l3_in_0_
timestamp 1676037725
transform 1 0 17388 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29532 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_1_
timestamp 1676037725
transform 1 0 26772 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_2_
timestamp 1676037725
transform 1 0 24104 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25668 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l2_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_29.mux_l2_in_1__262
timestamp 1676037725
transform -1 0 22908 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32108 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l1_in_1_
timestamp 1676037725
transform 1 0 29716 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l2_in_0_
timestamp 1676037725
transform 1 0 28336 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_37.mux_l2_in_1__212
timestamp 1676037725
transform 1 0 23828 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l2_in_1_
timestamp 1676037725
transform -1 0 24104 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18400 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 28336 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28336 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_45.mux_l2_in_1__213
timestamp 1676037725
transform -1 0 27968 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30268 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25944 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l2_in_1_
timestamp 1676037725
transform 1 0 22632 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_53.mux_l2_in_1__215
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19964 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_0_
timestamp 1676037725
transform -1 0 30268 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 33304 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_2_
timestamp 1676037725
transform -1 0 28612 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform -1 0 31832 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_0.mux_l2_in_1__217
timestamp 1676037725
transform -1 0 30084 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l2_in_1_
timestamp 1676037725
transform -1 0 31740 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l3_in_0_
timestamp 1676037725
transform -1 0 34316 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 39560 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform -1 0 34040 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_1_
timestamp 1676037725
transform -1 0 33120 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_2_
timestamp 1676037725
transform -1 0 30544 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform -1 0 36708 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_2.mux_l2_in_1__220
timestamp 1676037725
transform 1 0 33856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l2_in_1_
timestamp 1676037725
transform -1 0 34316 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l3_in_0_
timestamp 1676037725
transform -1 0 38824 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 41124 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform -1 0 35236 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 36248 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_2_
timestamp 1676037725
transform -1 0 30544 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform -1 0 36800 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l2_in_1_
timestamp 1676037725
transform -1 0 36524 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_4.mux_l2_in_1__224
timestamp 1676037725
transform -1 0 31832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l3_in_0_
timestamp 1676037725
transform -1 0 38272 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 41584 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform -1 0 35696 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform -1 0 33580 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_2_
timestamp 1676037725
transform -1 0 36248 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_6.mux_l1_in_3__227
timestamp 1676037725
transform 1 0 33764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_3_
timestamp 1676037725
transform -1 0 33120 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform -1 0 36708 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 38640 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l3_in_0_
timestamp 1676037725
transform -1 0 39100 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 41676 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform -1 0 34224 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_1_
timestamp 1676037725
transform -1 0 33488 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_2_
timestamp 1676037725
transform -1 0 34132 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_3_
timestamp 1676037725
transform -1 0 31832 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_10.mux_l1_in_3__218
timestamp 1676037725
transform -1 0 31188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform -1 0 35328 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l2_in_1_
timestamp 1676037725
transform -1 0 36892 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l3_in_0_
timestamp 1676037725
transform -1 0 38272 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 41032 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform -1 0 33120 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_1_
timestamp 1676037725
transform -1 0 33120 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_2_
timestamp 1676037725
transform -1 0 27968 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform -1 0 34132 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l2_in_1_
timestamp 1676037725
transform -1 0 33120 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_12.mux_l2_in_1__219
timestamp 1676037725
transform -1 0 29992 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l3_in_0_
timestamp 1676037725
transform -1 0 37904 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 41032 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30636 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_1_
timestamp 1676037725
transform -1 0 30636 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_2_
timestamp 1676037725
transform -1 0 27968 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l2_in_0_
timestamp 1676037725
transform -1 0 31372 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_20.mux_l2_in_1__221
timestamp 1676037725
transform 1 0 28980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l2_in_1_
timestamp 1676037725
transform -1 0 29256 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l3_in_0_
timestamp 1676037725
transform -1 0 34316 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 38456 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform -1 0 30544 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 30176 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_2_
timestamp 1676037725
transform -1 0 26496 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform -1 0 30544 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l2_in_1_
timestamp 1676037725
transform -1 0 31004 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_28.mux_l2_in_1__222
timestamp 1676037725
transform -1 0 29992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l3_in_0_
timestamp 1676037725
transform -1 0 33396 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 37904 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l1_in_0_
timestamp 1676037725
transform -1 0 32108 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l1_in_1_
timestamp 1676037725
transform -1 0 32936 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l2_in_0_
timestamp 1676037725
transform -1 0 33120 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l2_in_1_
timestamp 1676037725
transform -1 0 31832 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_36.mux_l2_in_1__223
timestamp 1676037725
transform 1 0 32292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l3_in_0_
timestamp 1676037725
transform -1 0 35696 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 39192 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform -1 0 30544 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_44.mux_l1_in_1__225
timestamp 1676037725
transform 1 0 29716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l1_in_1_
timestamp 1676037725
transform -1 0 28980 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform -1 0 33396 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 37720 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l1_in_0_
timestamp 1676037725
transform -1 0 29440 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l1_in_1_
timestamp 1676037725
transform -1 0 27784 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_52.mux_l1_in_1__226
timestamp 1676037725
transform -1 0 26680 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l2_in_0_
timestamp 1676037725
transform -1 0 33120 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 36800 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform -1 0 35696 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38824 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_2_
timestamp 1676037725
transform -1 0 24104 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_0.mux_l1_in_3__228
timestamp 1676037725
transform 1 0 29716 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 28428 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35880 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l2_in_1_
timestamp 1676037725
transform -1 0 29164 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 27140 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform -1 0 35696 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40020 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_2_
timestamp 1676037725
transform -1 0 31740 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 33028 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_2.mux_l2_in_1__234
timestamp 1676037725
transform -1 0 32844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 28428 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform -1 0 35328 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40020 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35696 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_4.mux_l2_in_1__244
timestamp 1676037725
transform 1 0 31280 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l2_in_1_
timestamp 1676037725
transform -1 0 30912 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 30820 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 27416 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 40204 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 41400 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_2_
timestamp 1676037725
transform -1 0 33488 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 36064 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_6.mux_l2_in_1__252
timestamp 1676037725
transform -1 0 35236 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33580 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29716 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1676037725
transform -1 0 38272 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 41216 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_2_
timestamp 1676037725
transform -1 0 34316 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l2_in_1_
timestamp 1676037725
transform -1 0 36892 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_8.mux_l2_in_1__253
timestamp 1676037725
transform 1 0 41124 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 36064 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 31464 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform -1 0 35512 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40112 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 36064 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l2_in_1_
timestamp 1676037725
transform -1 0 31740 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_10.mux_l2_in_1__229
timestamp 1676037725
transform 1 0 31372 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 31464 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 26404 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform -1 0 40848 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40388 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_12.mux_l2_in_1__230
timestamp 1676037725
transform -1 0 35144 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 37444 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 36064 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29716 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1676037725
transform -1 0 40756 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40480 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_14.mux_l2_in_1__231
timestamp 1676037725
transform 1 0 37444 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l2_in_1_
timestamp 1676037725
transform -1 0 35512 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37996 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1676037725
transform -1 0 40848 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40480 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_16.mux_l2_in_1__232
timestamp 1676037725
transform 1 0 37076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l2_in_1_
timestamp 1676037725
transform -1 0 35696 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l3_in_0_
timestamp 1676037725
transform 1 0 35880 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 28980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1676037725
transform -1 0 38640 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 39652 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l2_in_1_
timestamp 1676037725
transform -1 0 31556 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_18.mux_l2_in_1__233
timestamp 1676037725
transform 1 0 31372 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 25760 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27324 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_20.mux_l1_in_1__235
timestamp 1676037725
transform -1 0 25208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l1_in_1_
timestamp 1676037725
transform -1 0 25668 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24840 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25852 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_22.mux_l1_in_1__236
timestamp 1676037725
transform 1 0 24196 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22908 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20056 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l1_in_1_
timestamp 1676037725
transform -1 0 22908 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_24.mux_l1_in_1__237
timestamp 1676037725
transform -1 0 20056 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27416 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_26.mux_l1_in_1__238
timestamp 1676037725
transform 1 0 25392 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24196 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22080 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22264 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_28.mux_l2_in_0__239
timestamp 1676037725
transform 1 0 22632 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14904 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_30.mux_l2_in_0__240
timestamp 1676037725
transform -1 0 17480 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_32.mux_l2_in_0__241
timestamp 1676037725
transform 1 0 19044 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 12604 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19504 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19228 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_34.mux_l2_in_0__242
timestamp 1676037725
transform -1 0 19780 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14904 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25852 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_36.mux_l1_in_1__243
timestamp 1676037725
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21988 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 14536 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 13156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_40.mux_l2_in_0__245
timestamp 1676037725
transform 1 0 13064 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9752 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_42.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16744 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_42.mux_l2_in_0__246
timestamp 1676037725
transform -1 0 11224 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_42.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13892 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10488 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_44.mux_l2_in_0__247
timestamp 1676037725
transform -1 0 10580 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12512 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10304 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11868 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_46.mux_l2_in_0__248
timestamp 1676037725
transform -1 0 9936 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9016 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_48.mux_l2_in_0__249
timestamp 1676037725
transform -1 0 10764 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9200 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_50.mux_l2_in_0__250
timestamp 1676037725
transform -1 0 10120 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_58.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_58.mux_l2_in_0__251
timestamp 1676037725
transform -1 0 10120 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_58.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 26864 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 32016 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 37168 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 42320 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 47472 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 49238 26200 49294 27000 0 FreeSans 224 90 0 0 ccff_head_1
port 3 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1582 26200 1638 27000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[20]
port 18 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[21]
port 19 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[22]
port 20 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[23]
port 21 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[24]
port 22 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[25]
port 23 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[26]
port 24 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[27]
port 25 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[28]
port 26 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[29]
port 27 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 28 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 29 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 30 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 31 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 32 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 33 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 34 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 35 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 36 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 37 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 38 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 39 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 40 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 41 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 42 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 43 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 44 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 45 nsew signal tristate
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 46 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 47 nsew signal tristate
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 chanx_left_out[20]
port 48 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 chanx_left_out[21]
port 49 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 chanx_left_out[22]
port 50 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_out[23]
port 51 nsew signal tristate
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 chanx_left_out[24]
port 52 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 chanx_left_out[25]
port 53 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 chanx_left_out[26]
port 54 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 chanx_left_out[27]
port 55 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_out[28]
port 56 nsew signal tristate
flabel metal3 s 0 25576 800 25696 0 FreeSans 480 0 0 0 chanx_left_out[29]
port 57 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal3 s 50200 13608 51000 13728 0 FreeSans 480 0 0 0 chanx_right_in_0[0]
port 66 nsew signal input
flabel metal3 s 50200 17688 51000 17808 0 FreeSans 480 0 0 0 chanx_right_in_0[10]
port 67 nsew signal input
flabel metal3 s 50200 18096 51000 18216 0 FreeSans 480 0 0 0 chanx_right_in_0[11]
port 68 nsew signal input
flabel metal3 s 50200 18504 51000 18624 0 FreeSans 480 0 0 0 chanx_right_in_0[12]
port 69 nsew signal input
flabel metal3 s 50200 18912 51000 19032 0 FreeSans 480 0 0 0 chanx_right_in_0[13]
port 70 nsew signal input
flabel metal3 s 50200 19320 51000 19440 0 FreeSans 480 0 0 0 chanx_right_in_0[14]
port 71 nsew signal input
flabel metal3 s 50200 19728 51000 19848 0 FreeSans 480 0 0 0 chanx_right_in_0[15]
port 72 nsew signal input
flabel metal3 s 50200 20136 51000 20256 0 FreeSans 480 0 0 0 chanx_right_in_0[16]
port 73 nsew signal input
flabel metal3 s 50200 20544 51000 20664 0 FreeSans 480 0 0 0 chanx_right_in_0[17]
port 74 nsew signal input
flabel metal3 s 50200 20952 51000 21072 0 FreeSans 480 0 0 0 chanx_right_in_0[18]
port 75 nsew signal input
flabel metal3 s 50200 21360 51000 21480 0 FreeSans 480 0 0 0 chanx_right_in_0[19]
port 76 nsew signal input
flabel metal3 s 50200 14016 51000 14136 0 FreeSans 480 0 0 0 chanx_right_in_0[1]
port 77 nsew signal input
flabel metal3 s 50200 21768 51000 21888 0 FreeSans 480 0 0 0 chanx_right_in_0[20]
port 78 nsew signal input
flabel metal3 s 50200 22176 51000 22296 0 FreeSans 480 0 0 0 chanx_right_in_0[21]
port 79 nsew signal input
flabel metal3 s 50200 22584 51000 22704 0 FreeSans 480 0 0 0 chanx_right_in_0[22]
port 80 nsew signal input
flabel metal3 s 50200 22992 51000 23112 0 FreeSans 480 0 0 0 chanx_right_in_0[23]
port 81 nsew signal input
flabel metal3 s 50200 23400 51000 23520 0 FreeSans 480 0 0 0 chanx_right_in_0[24]
port 82 nsew signal input
flabel metal3 s 50200 23808 51000 23928 0 FreeSans 480 0 0 0 chanx_right_in_0[25]
port 83 nsew signal input
flabel metal3 s 50200 24216 51000 24336 0 FreeSans 480 0 0 0 chanx_right_in_0[26]
port 84 nsew signal input
flabel metal3 s 50200 24624 51000 24744 0 FreeSans 480 0 0 0 chanx_right_in_0[27]
port 85 nsew signal input
flabel metal3 s 50200 25032 51000 25152 0 FreeSans 480 0 0 0 chanx_right_in_0[28]
port 86 nsew signal input
flabel metal3 s 50200 25440 51000 25560 0 FreeSans 480 0 0 0 chanx_right_in_0[29]
port 87 nsew signal input
flabel metal3 s 50200 14424 51000 14544 0 FreeSans 480 0 0 0 chanx_right_in_0[2]
port 88 nsew signal input
flabel metal3 s 50200 14832 51000 14952 0 FreeSans 480 0 0 0 chanx_right_in_0[3]
port 89 nsew signal input
flabel metal3 s 50200 15240 51000 15360 0 FreeSans 480 0 0 0 chanx_right_in_0[4]
port 90 nsew signal input
flabel metal3 s 50200 15648 51000 15768 0 FreeSans 480 0 0 0 chanx_right_in_0[5]
port 91 nsew signal input
flabel metal3 s 50200 16056 51000 16176 0 FreeSans 480 0 0 0 chanx_right_in_0[6]
port 92 nsew signal input
flabel metal3 s 50200 16464 51000 16584 0 FreeSans 480 0 0 0 chanx_right_in_0[7]
port 93 nsew signal input
flabel metal3 s 50200 16872 51000 16992 0 FreeSans 480 0 0 0 chanx_right_in_0[8]
port 94 nsew signal input
flabel metal3 s 50200 17280 51000 17400 0 FreeSans 480 0 0 0 chanx_right_in_0[9]
port 95 nsew signal input
flabel metal3 s 50200 1368 51000 1488 0 FreeSans 480 0 0 0 chanx_right_out_0[0]
port 96 nsew signal tristate
flabel metal3 s 50200 5448 51000 5568 0 FreeSans 480 0 0 0 chanx_right_out_0[10]
port 97 nsew signal tristate
flabel metal3 s 50200 5856 51000 5976 0 FreeSans 480 0 0 0 chanx_right_out_0[11]
port 98 nsew signal tristate
flabel metal3 s 50200 6264 51000 6384 0 FreeSans 480 0 0 0 chanx_right_out_0[12]
port 99 nsew signal tristate
flabel metal3 s 50200 6672 51000 6792 0 FreeSans 480 0 0 0 chanx_right_out_0[13]
port 100 nsew signal tristate
flabel metal3 s 50200 7080 51000 7200 0 FreeSans 480 0 0 0 chanx_right_out_0[14]
port 101 nsew signal tristate
flabel metal3 s 50200 7488 51000 7608 0 FreeSans 480 0 0 0 chanx_right_out_0[15]
port 102 nsew signal tristate
flabel metal3 s 50200 7896 51000 8016 0 FreeSans 480 0 0 0 chanx_right_out_0[16]
port 103 nsew signal tristate
flabel metal3 s 50200 8304 51000 8424 0 FreeSans 480 0 0 0 chanx_right_out_0[17]
port 104 nsew signal tristate
flabel metal3 s 50200 8712 51000 8832 0 FreeSans 480 0 0 0 chanx_right_out_0[18]
port 105 nsew signal tristate
flabel metal3 s 50200 9120 51000 9240 0 FreeSans 480 0 0 0 chanx_right_out_0[19]
port 106 nsew signal tristate
flabel metal3 s 50200 1776 51000 1896 0 FreeSans 480 0 0 0 chanx_right_out_0[1]
port 107 nsew signal tristate
flabel metal3 s 50200 9528 51000 9648 0 FreeSans 480 0 0 0 chanx_right_out_0[20]
port 108 nsew signal tristate
flabel metal3 s 50200 9936 51000 10056 0 FreeSans 480 0 0 0 chanx_right_out_0[21]
port 109 nsew signal tristate
flabel metal3 s 50200 10344 51000 10464 0 FreeSans 480 0 0 0 chanx_right_out_0[22]
port 110 nsew signal tristate
flabel metal3 s 50200 10752 51000 10872 0 FreeSans 480 0 0 0 chanx_right_out_0[23]
port 111 nsew signal tristate
flabel metal3 s 50200 11160 51000 11280 0 FreeSans 480 0 0 0 chanx_right_out_0[24]
port 112 nsew signal tristate
flabel metal3 s 50200 11568 51000 11688 0 FreeSans 480 0 0 0 chanx_right_out_0[25]
port 113 nsew signal tristate
flabel metal3 s 50200 11976 51000 12096 0 FreeSans 480 0 0 0 chanx_right_out_0[26]
port 114 nsew signal tristate
flabel metal3 s 50200 12384 51000 12504 0 FreeSans 480 0 0 0 chanx_right_out_0[27]
port 115 nsew signal tristate
flabel metal3 s 50200 12792 51000 12912 0 FreeSans 480 0 0 0 chanx_right_out_0[28]
port 116 nsew signal tristate
flabel metal3 s 50200 13200 51000 13320 0 FreeSans 480 0 0 0 chanx_right_out_0[29]
port 117 nsew signal tristate
flabel metal3 s 50200 2184 51000 2304 0 FreeSans 480 0 0 0 chanx_right_out_0[2]
port 118 nsew signal tristate
flabel metal3 s 50200 2592 51000 2712 0 FreeSans 480 0 0 0 chanx_right_out_0[3]
port 119 nsew signal tristate
flabel metal3 s 50200 3000 51000 3120 0 FreeSans 480 0 0 0 chanx_right_out_0[4]
port 120 nsew signal tristate
flabel metal3 s 50200 3408 51000 3528 0 FreeSans 480 0 0 0 chanx_right_out_0[5]
port 121 nsew signal tristate
flabel metal3 s 50200 3816 51000 3936 0 FreeSans 480 0 0 0 chanx_right_out_0[6]
port 122 nsew signal tristate
flabel metal3 s 50200 4224 51000 4344 0 FreeSans 480 0 0 0 chanx_right_out_0[7]
port 123 nsew signal tristate
flabel metal3 s 50200 4632 51000 4752 0 FreeSans 480 0 0 0 chanx_right_out_0[8]
port 124 nsew signal tristate
flabel metal3 s 50200 5040 51000 5160 0 FreeSans 480 0 0 0 chanx_right_out_0[9]
port 125 nsew signal tristate
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 126 nsew signal input
flabel metal2 s 27986 26200 28042 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 127 nsew signal input
flabel metal2 s 28630 26200 28686 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 128 nsew signal input
flabel metal2 s 29274 26200 29330 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 129 nsew signal input
flabel metal2 s 29918 26200 29974 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 130 nsew signal input
flabel metal2 s 30562 26200 30618 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 131 nsew signal input
flabel metal2 s 31206 26200 31262 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 132 nsew signal input
flabel metal2 s 31850 26200 31906 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 133 nsew signal input
flabel metal2 s 32494 26200 32550 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 134 nsew signal input
flabel metal2 s 33138 26200 33194 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 135 nsew signal input
flabel metal2 s 33782 26200 33838 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 136 nsew signal input
flabel metal2 s 22190 26200 22246 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 137 nsew signal input
flabel metal2 s 34426 26200 34482 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 138 nsew signal input
flabel metal2 s 35070 26200 35126 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 139 nsew signal input
flabel metal2 s 35714 26200 35770 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 140 nsew signal input
flabel metal2 s 36358 26200 36414 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 141 nsew signal input
flabel metal2 s 37002 26200 37058 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 142 nsew signal input
flabel metal2 s 37646 26200 37702 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 143 nsew signal input
flabel metal2 s 38290 26200 38346 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 144 nsew signal input
flabel metal2 s 38934 26200 38990 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 145 nsew signal input
flabel metal2 s 39578 26200 39634 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 146 nsew signal input
flabel metal2 s 40222 26200 40278 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 147 nsew signal input
flabel metal2 s 22834 26200 22890 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 148 nsew signal input
flabel metal2 s 23478 26200 23534 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 149 nsew signal input
flabel metal2 s 24122 26200 24178 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 150 nsew signal input
flabel metal2 s 24766 26200 24822 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 151 nsew signal input
flabel metal2 s 25410 26200 25466 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 152 nsew signal input
flabel metal2 s 26054 26200 26110 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 153 nsew signal input
flabel metal2 s 26698 26200 26754 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 154 nsew signal input
flabel metal2 s 27342 26200 27398 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 155 nsew signal input
flabel metal2 s 2226 26200 2282 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 156 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 157 nsew signal tristate
flabel metal2 s 9310 26200 9366 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 158 nsew signal tristate
flabel metal2 s 9954 26200 10010 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 159 nsew signal tristate
flabel metal2 s 10598 26200 10654 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 160 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 161 nsew signal tristate
flabel metal2 s 11886 26200 11942 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 162 nsew signal tristate
flabel metal2 s 12530 26200 12586 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 163 nsew signal tristate
flabel metal2 s 13174 26200 13230 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 164 nsew signal tristate
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 165 nsew signal tristate
flabel metal2 s 14462 26200 14518 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 166 nsew signal tristate
flabel metal2 s 2870 26200 2926 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 167 nsew signal tristate
flabel metal2 s 15106 26200 15162 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 168 nsew signal tristate
flabel metal2 s 15750 26200 15806 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 169 nsew signal tristate
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 170 nsew signal tristate
flabel metal2 s 17038 26200 17094 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 171 nsew signal tristate
flabel metal2 s 17682 26200 17738 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 172 nsew signal tristate
flabel metal2 s 18326 26200 18382 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 173 nsew signal tristate
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 174 nsew signal tristate
flabel metal2 s 19614 26200 19670 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 175 nsew signal tristate
flabel metal2 s 20258 26200 20314 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 176 nsew signal tristate
flabel metal2 s 20902 26200 20958 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 177 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 178 nsew signal tristate
flabel metal2 s 4158 26200 4214 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 179 nsew signal tristate
flabel metal2 s 4802 26200 4858 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 180 nsew signal tristate
flabel metal2 s 5446 26200 5502 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 181 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 182 nsew signal tristate
flabel metal2 s 6734 26200 6790 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 183 nsew signal tristate
flabel metal2 s 7378 26200 7434 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 184 nsew signal tristate
flabel metal2 s 8022 26200 8078 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 185 nsew signal tristate
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 42154 26200 42210 27000 0 FreeSans 224 90 0 0 prog_reset
port 200 nsew signal input
flabel metal2 s 42798 26200 42854 27000 0 FreeSans 224 90 0 0 reset
port 201 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 202 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 203 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 204 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 205 nsew signal input
flabel metal2 s 43442 26200 43498 27000 0 FreeSans 224 90 0 0 test_enable
port 206 nsew signal input
flabel metal2 s 45374 26200 45430 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 207 nsew signal input
flabel metal2 s 46018 26200 46074 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 208 nsew signal input
flabel metal2 s 46662 26200 46718 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 209 nsew signal input
flabel metal2 s 47306 26200 47362 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 210 nsew signal input
flabel metal2 s 47950 26200 48006 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 211 nsew signal input
flabel metal2 s 48594 26200 48650 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 212 nsew signal input
flabel metal2 s 44086 26200 44142 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 213 nsew signal input
flabel metal2 s 44730 26200 44786 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 214 nsew signal input
flabel metal2 s 1122 0 1178 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_inpad_0_
port 215 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_1__pin_inpad_0_
port 216 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_2__pin_inpad_0_
port 217 nsew signal tristate
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_3__pin_inpad_0_
port 218 nsew signal tristate
rlabel metal1 25484 23936 25484 23936 0 VGND
rlabel metal1 25484 24480 25484 24480 0 VPWR
rlabel metal1 21850 4658 21850 4658 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 19872 4658 19872 4658 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal2 18906 6596 18906 6596 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 17480 6290 17480 6290 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 20424 20978 20424 20978 0 cbx_1__0_.cbx_8__0_.ccff_head
rlabel metal2 18630 9044 18630 9044 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
rlabel metal1 15778 16048 15778 16048 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
rlabel metal1 16790 13498 16790 13498 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
rlabel metal2 16422 9962 16422 9962 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
rlabel metal1 15226 9010 15226 9010 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
rlabel metal1 19734 14450 19734 14450 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
rlabel metal1 13662 15538 13662 15538 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
rlabel metal1 14122 9894 14122 9894 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
rlabel metal1 11040 11186 11040 11186 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
rlabel metal1 13570 9622 13570 9622 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
rlabel metal2 14950 13056 14950 13056 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
rlabel metal1 11546 12410 11546 12410 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
rlabel metal2 14950 16286 14950 16286 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
rlabel metal1 15778 14926 15778 14926 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
rlabel metal1 13156 16014 13156 16014 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
rlabel metal2 15502 14892 15502 14892 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17848 7786 17848 7786 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 19642 7276 19642 7276 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 15594 14246 15594 14246 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17618 14994 17618 14994 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 17526 14144 17526 14144 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16836 12682 16836 12682 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15916 11186 15916 11186 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16882 14042 16882 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 16974 8908 16974 8908 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 17066 9146 17066 9146 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 17710 7854 17710 7854 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 13018 15470 13018 15470 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15594 9860 15594 9860 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 16836 6766 16836 6766 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13432 15470 13432 15470 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17802 13974 17802 13974 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 15962 14416 15962 14416 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 14076 10098 14076 10098 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13662 15334 13662 15334 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 14950 14042 14950 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 14766 10234 14766 10234 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 16560 10778 16560 10778 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 15502 10268 15502 10268 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 9706 15810 9706 15810 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12374 10540 12374 10540 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 14858 7854 14858 7854 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 9798 15538 9798 15538 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18308 14586 18308 14586 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14582 14586 14582 14586 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 15824 10642 15824 10642 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11684 12954 11684 12954 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 13938 14042 13938 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 14398 11254 14398 11254 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 12558 11730 12558 11730 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 12512 12614 12512 12614 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 13662 16320 13662 16320 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12834 14586 12834 14586 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 13156 8942 13156 8942 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 14398 16184 14398 16184 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15870 15062 15870 15062 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17158 15130 17158 15130 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 14858 11356 14858 11356 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12834 16218 12834 16218 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 15042 14790 15042 14790 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 13754 14246 13754 14246 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 14214 14314 14214 14314 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 11684 16218 11684 16218 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 20332 3434 20332 3434 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal2 22218 2958 22218 2958 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 26312 3026 26312 3026 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 28842 4012 28842 4012 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 23506 2856 23506 2856 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 19113 2414 19113 2414 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal2 21298 3740 21298 3740 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 23161 4114 23161 4114 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 27600 2958 27600 2958 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal2 19090 4080 19090 4080 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 20654 4012 20654 4012 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal2 25898 4318 25898 4318 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 17296 3502 17296 3502 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 19090 6086 19090 6086 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 24564 3570 24564 3570 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 9522 2278 9522 2278 0 ccff_head
rlabel metal1 49082 23698 49082 23698 0 ccff_head_1
rlabel metal2 41354 1622 41354 1622 0 ccff_tail
rlabel metal2 1610 24524 1610 24524 0 ccff_tail_0
rlabel metal1 2990 2414 2990 2414 0 chanx_left_in[0]
rlabel metal1 1472 5678 1472 5678 0 chanx_left_in[10]
rlabel metal1 1472 6290 1472 6290 0 chanx_left_in[11]
rlabel metal1 1840 6766 1840 6766 0 chanx_left_in[12]
rlabel metal1 1472 6698 1472 6698 0 chanx_left_in[13]
rlabel metal1 1472 7378 1472 7378 0 chanx_left_in[14]
rlabel metal1 1472 7854 1472 7854 0 chanx_left_in[15]
rlabel metal1 1748 8058 1748 8058 0 chanx_left_in[16]
rlabel metal1 1794 8942 1794 8942 0 chanx_left_in[17]
rlabel metal1 1518 8874 1518 8874 0 chanx_left_in[18]
rlabel metal1 1472 9554 1472 9554 0 chanx_left_in[19]
rlabel metal1 1840 2346 1840 2346 0 chanx_left_in[1]
rlabel metal1 1748 9690 1748 9690 0 chanx_left_in[20]
rlabel metal1 2346 10676 2346 10676 0 chanx_left_in[21]
rlabel metal1 1472 10642 1472 10642 0 chanx_left_in[22]
rlabel metal2 1610 11033 1610 11033 0 chanx_left_in[23]
rlabel metal1 2346 11696 2346 11696 0 chanx_left_in[24]
rlabel metal1 1886 12274 1886 12274 0 chanx_left_in[25]
rlabel metal1 1426 11730 1426 11730 0 chanx_left_in[26]
rlabel metal2 1242 12699 1242 12699 0 chanx_left_in[27]
rlabel metal1 1518 12886 1518 12886 0 chanx_left_in[28]
rlabel metal2 3542 13651 3542 13651 0 chanx_left_in[29]
rlabel metal1 2208 2414 2208 2414 0 chanx_left_in[2]
rlabel metal1 1472 3026 1472 3026 0 chanx_left_in[3]
rlabel metal1 1748 3162 1748 3162 0 chanx_left_in[4]
rlabel metal1 2070 4114 2070 4114 0 chanx_left_in[5]
rlabel metal1 1564 4182 1564 4182 0 chanx_left_in[6]
rlabel metal1 1472 4590 1472 4590 0 chanx_left_in[7]
rlabel metal1 1748 4794 1748 4794 0 chanx_left_in[8]
rlabel metal1 2576 5678 2576 5678 0 chanx_left_in[9]
rlabel metal3 1234 13804 1234 13804 0 chanx_left_out[0]
rlabel metal3 1050 17884 1050 17884 0 chanx_left_out[10]
rlabel metal3 1234 18292 1234 18292 0 chanx_left_out[11]
rlabel metal3 1096 18700 1096 18700 0 chanx_left_out[12]
rlabel metal1 2645 20366 2645 20366 0 chanx_left_out[13]
rlabel metal2 2898 20247 2898 20247 0 chanx_left_out[14]
rlabel metal3 1234 19924 1234 19924 0 chanx_left_out[15]
rlabel metal3 1004 20332 1004 20332 0 chanx_left_out[16]
rlabel metal3 866 20740 866 20740 0 chanx_left_out[17]
rlabel metal1 2668 22542 2668 22542 0 chanx_left_out[18]
rlabel metal3 1234 21556 1234 21556 0 chanx_left_out[19]
rlabel metal3 866 14212 866 14212 0 chanx_left_out[1]
rlabel via2 3266 21947 3266 21947 0 chanx_left_out[20]
rlabel metal3 1395 22372 1395 22372 0 chanx_left_out[21]
rlabel metal3 1786 22780 1786 22780 0 chanx_left_out[22]
rlabel metal3 1878 23188 1878 23188 0 chanx_left_out[23]
rlabel metal3 2062 23596 2062 23596 0 chanx_left_out[24]
rlabel metal3 2108 24004 2108 24004 0 chanx_left_out[25]
rlabel metal3 1740 24412 1740 24412 0 chanx_left_out[26]
rlabel metal3 2154 24820 2154 24820 0 chanx_left_out[27]
rlabel metal3 2200 25228 2200 25228 0 chanx_left_out[28]
rlabel metal3 2062 25636 2062 25636 0 chanx_left_out[29]
rlabel metal3 820 14620 820 14620 0 chanx_left_out[2]
rlabel metal3 820 15028 820 15028 0 chanx_left_out[3]
rlabel metal3 820 15436 820 15436 0 chanx_left_out[4]
rlabel metal3 866 15844 866 15844 0 chanx_left_out[5]
rlabel metal3 866 16252 866 16252 0 chanx_left_out[6]
rlabel metal3 866 16660 866 16660 0 chanx_left_out[7]
rlabel metal3 820 17068 820 17068 0 chanx_left_out[8]
rlabel metal3 1234 17476 1234 17476 0 chanx_left_out[9]
rlabel metal1 48438 13906 48438 13906 0 chanx_right_in_0[0]
rlabel metal2 49358 18003 49358 18003 0 chanx_right_in_0[10]
rlabel metal1 49404 18734 49404 18734 0 chanx_right_in_0[11]
rlabel metal2 48806 18479 48806 18479 0 chanx_right_in_0[12]
rlabel metal2 49266 19159 49266 19159 0 chanx_right_in_0[13]
rlabel metal1 49312 19754 49312 19754 0 chanx_right_in_0[14]
rlabel metal1 49404 20434 49404 20434 0 chanx_right_in_0[15]
rlabel metal2 48806 20111 48806 20111 0 chanx_right_in_0[16]
rlabel metal2 49358 20757 49358 20757 0 chanx_right_in_0[17]
rlabel metal2 49358 21267 49358 21267 0 chanx_right_in_0[18]
rlabel metal2 49266 21675 49266 21675 0 chanx_right_in_0[19]
rlabel metal2 49266 14025 49266 14025 0 chanx_right_in_0[1]
rlabel metal2 48622 21675 48622 21675 0 chanx_right_in_0[20]
rlabel metal2 49358 22423 49358 22423 0 chanx_right_in_0[21]
rlabel metal1 49404 23086 49404 23086 0 chanx_right_in_0[22]
rlabel metal1 48668 23086 48668 23086 0 chanx_right_in_0[23]
rlabel metal1 47426 21522 47426 21522 0 chanx_right_in_0[24]
rlabel metal2 46690 23511 46690 23511 0 chanx_right_in_0[25]
rlabel metal2 47794 23443 47794 23443 0 chanx_right_in_0[26]
rlabel metal1 47748 21998 47748 21998 0 chanx_right_in_0[27]
rlabel metal1 47196 22678 47196 22678 0 chanx_right_in_0[28]
rlabel metal2 47518 23596 47518 23596 0 chanx_right_in_0[29]
rlabel metal2 49266 14433 49266 14433 0 chanx_right_in_0[2]
rlabel metal2 49358 14943 49358 14943 0 chanx_right_in_0[3]
rlabel metal2 49358 15385 49358 15385 0 chanx_right_in_0[4]
rlabel metal2 49358 15895 49358 15895 0 chanx_right_in_0[5]
rlabel metal1 49404 16558 49404 16558 0 chanx_right_in_0[6]
rlabel metal1 48760 17238 48760 17238 0 chanx_right_in_0[7]
rlabel metal2 48806 16847 48806 16847 0 chanx_right_in_0[8]
rlabel metal2 49358 17493 49358 17493 0 chanx_right_in_0[9]
rlabel metal2 46690 2737 46690 2737 0 chanx_right_out_0[0]
rlabel metal1 49312 4658 49312 4658 0 chanx_right_out_0[10]
rlabel metal2 49174 5593 49174 5593 0 chanx_right_out_0[11]
rlabel metal3 49504 6324 49504 6324 0 chanx_right_out_0[12]
rlabel metal1 49220 5746 49220 5746 0 chanx_right_out_0[13]
rlabel metal1 49266 6358 49266 6358 0 chanx_right_out_0[14]
rlabel metal3 49734 7548 49734 7548 0 chanx_right_out_0[15]
rlabel metal2 46874 8177 46874 8177 0 chanx_right_out_0[16]
rlabel metal1 49266 7446 49266 7446 0 chanx_right_out_0[17]
rlabel metal1 49220 7922 49220 7922 0 chanx_right_out_0[18]
rlabel metal2 49174 8857 49174 8857 0 chanx_right_out_0[19]
rlabel metal2 46782 2397 46782 2397 0 chanx_right_out_0[1]
rlabel metal3 48814 9588 48814 9588 0 chanx_right_out_0[20]
rlabel metal1 49266 9010 49266 9010 0 chanx_right_out_0[21]
rlabel metal1 49220 9622 49220 9622 0 chanx_right_out_0[22]
rlabel metal2 49174 10455 49174 10455 0 chanx_right_out_0[23]
rlabel metal1 49220 10710 49220 10710 0 chanx_right_out_0[24]
rlabel metal2 49174 11407 49174 11407 0 chanx_right_out_0[25]
rlabel metal2 49174 11917 49174 11917 0 chanx_right_out_0[26]
rlabel metal2 49174 12359 49174 12359 0 chanx_right_out_0[27]
rlabel via2 49174 12835 49174 12835 0 chanx_right_out_0[28]
rlabel metal3 49734 13260 49734 13260 0 chanx_right_out_0[29]
rlabel metal3 49412 2244 49412 2244 0 chanx_right_out_0[2]
rlabel metal2 46874 2805 46874 2805 0 chanx_right_out_0[3]
rlabel metal3 49504 3060 49504 3060 0 chanx_right_out_0[4]
rlabel metal2 49174 2975 49174 2975 0 chanx_right_out_0[5]
rlabel metal1 49220 3094 49220 3094 0 chanx_right_out_0[6]
rlabel metal2 49174 3927 49174 3927 0 chanx_right_out_0[7]
rlabel metal1 47610 5134 47610 5134 0 chanx_right_out_0[8]
rlabel metal1 49266 4114 49266 4114 0 chanx_right_out_0[9]
rlabel metal2 21574 24626 21574 24626 0 chany_top_in[0]
rlabel metal1 29118 23664 29118 23664 0 chany_top_in[10]
rlabel metal2 28658 25306 28658 25306 0 chany_top_in[11]
rlabel metal2 31602 24378 31602 24378 0 chany_top_in[12]
rlabel metal1 33258 24174 33258 24174 0 chany_top_in[13]
rlabel metal2 39698 23936 39698 23936 0 chany_top_in[14]
rlabel metal1 33488 23086 33488 23086 0 chany_top_in[15]
rlabel metal2 39514 24378 39514 24378 0 chany_top_in[16]
rlabel metal1 43148 20978 43148 20978 0 chany_top_in[17]
rlabel metal1 40112 23698 40112 23698 0 chany_top_in[18]
rlabel metal2 33994 24276 33994 24276 0 chany_top_in[19]
rlabel metal1 10672 22542 10672 22542 0 chany_top_in[1]
rlabel metal2 34454 23793 34454 23793 0 chany_top_in[20]
rlabel metal1 40710 23596 40710 23596 0 chany_top_in[21]
rlabel metal1 42826 21114 42826 21114 0 chany_top_in[22]
rlabel metal2 43286 21760 43286 21760 0 chany_top_in[23]
rlabel via2 42826 21981 42826 21981 0 chany_top_in[24]
rlabel via2 38594 22763 38594 22763 0 chany_top_in[25]
rlabel metal1 44712 22066 44712 22066 0 chany_top_in[26]
rlabel metal2 42090 23698 42090 23698 0 chany_top_in[27]
rlabel metal1 45356 22610 45356 22610 0 chany_top_in[28]
rlabel metal1 44068 22610 44068 22610 0 chany_top_in[29]
rlabel metal1 15226 23222 15226 23222 0 chany_top_in[2]
rlabel metal1 23184 23698 23184 23698 0 chany_top_in[3]
rlabel metal1 24104 21114 24104 21114 0 chany_top_in[4]
rlabel metal2 24794 25544 24794 25544 0 chany_top_in[5]
rlabel metal1 25346 23290 25346 23290 0 chany_top_in[6]
rlabel metal1 27094 24174 27094 24174 0 chany_top_in[7]
rlabel metal2 27830 23868 27830 23868 0 chany_top_in[8]
rlabel metal1 28566 24208 28566 24208 0 chany_top_in[9]
rlabel metal1 3266 22202 3266 22202 0 chany_top_out[0]
rlabel metal1 8464 24242 8464 24242 0 chany_top_out[10]
rlabel metal1 9062 23630 9062 23630 0 chany_top_out[11]
rlabel metal2 9982 24490 9982 24490 0 chany_top_out[12]
rlabel metal2 10626 24966 10626 24966 0 chany_top_out[13]
rlabel metal2 11270 24728 11270 24728 0 chany_top_out[14]
rlabel metal1 10718 24276 10718 24276 0 chany_top_out[15]
rlabel metal2 12703 26316 12703 26316 0 chany_top_out[16]
rlabel metal1 13340 23154 13340 23154 0 chany_top_out[17]
rlabel metal1 13570 24242 13570 24242 0 chany_top_out[18]
rlabel metal1 14352 23766 14352 23766 0 chany_top_out[19]
rlabel metal2 3135 26316 3135 26316 0 chany_top_out[1]
rlabel metal2 15134 24490 15134 24490 0 chany_top_out[20]
rlabel metal2 15778 24728 15778 24728 0 chany_top_out[21]
rlabel metal1 16146 23630 16146 23630 0 chany_top_out[22]
rlabel metal1 17342 22134 17342 22134 0 chany_top_out[23]
rlabel metal1 16790 24242 16790 24242 0 chany_top_out[24]
rlabel metal1 18124 23630 18124 23630 0 chany_top_out[25]
rlabel metal1 19458 22066 19458 22066 0 chany_top_out[26]
rlabel metal1 18446 24276 18446 24276 0 chany_top_out[27]
rlabel metal2 20286 25306 20286 25306 0 chany_top_out[28]
rlabel metal2 20930 25272 20930 25272 0 chany_top_out[29]
rlabel metal1 3266 24242 3266 24242 0 chany_top_out[2]
rlabel metal1 3956 23630 3956 23630 0 chany_top_out[3]
rlabel metal2 4830 24490 4830 24490 0 chany_top_out[4]
rlabel metal2 5474 24966 5474 24966 0 chany_top_out[5]
rlabel metal2 6118 24728 6118 24728 0 chany_top_out[6]
rlabel metal1 6302 24242 6302 24242 0 chany_top_out[7]
rlabel metal1 7682 22542 7682 22542 0 chany_top_out[8]
rlabel metal2 7866 23919 7866 23919 0 chany_top_out[9]
rlabel metal2 18722 17816 18722 17816 0 clknet_0_prog_clk
rlabel metal2 13662 5712 13662 5712 0 clknet_4_0_0_prog_clk
rlabel metal2 32154 11152 32154 11152 0 clknet_4_10_0_prog_clk
rlabel metal2 34086 13566 34086 13566 0 clknet_4_11_0_prog_clk
rlabel metal1 32338 17204 32338 17204 0 clknet_4_12_0_prog_clk
rlabel metal1 34316 20366 34316 20366 0 clknet_4_13_0_prog_clk
rlabel metal1 34868 15538 34868 15538 0 clknet_4_14_0_prog_clk
rlabel metal2 37582 17170 37582 17170 0 clknet_4_15_0_prog_clk
rlabel metal1 10626 12274 10626 12274 0 clknet_4_1_0_prog_clk
rlabel metal2 21022 3230 21022 3230 0 clknet_4_2_0_prog_clk
rlabel metal1 25622 12886 25622 12886 0 clknet_4_3_0_prog_clk
rlabel metal1 14950 19346 14950 19346 0 clknet_4_4_0_prog_clk
rlabel metal1 21252 14450 21252 14450 0 clknet_4_5_0_prog_clk
rlabel metal2 21758 23392 21758 23392 0 clknet_4_6_0_prog_clk
rlabel metal1 25484 19346 25484 19346 0 clknet_4_7_0_prog_clk
rlabel metal2 28842 5712 28842 5712 0 clknet_4_8_0_prog_clk
rlabel metal1 27002 13838 27002 13838 0 clknet_4_9_0_prog_clk
rlabel metal2 11730 1554 11730 1554 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 13846 1554 13846 1554 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 15962 1554 15962 1554 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 18078 823 18078 823 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 29118 2414 29118 2414 0 gfpga_pad_io_soc_in[0]
rlabel metal1 30912 2414 30912 2414 0 gfpga_pad_io_soc_in[1]
rlabel metal2 33166 1989 33166 1989 0 gfpga_pad_io_soc_in[2]
rlabel metal1 35144 2414 35144 2414 0 gfpga_pad_io_soc_in[3]
rlabel metal2 20194 1622 20194 1622 0 gfpga_pad_io_soc_out[0]
rlabel metal2 22310 1622 22310 1622 0 gfpga_pad_io_soc_out[1]
rlabel metal2 24426 1622 24426 1622 0 gfpga_pad_io_soc_out[2]
rlabel metal2 26542 1622 26542 1622 0 gfpga_pad_io_soc_out[3]
rlabel metal2 37122 1520 37122 1520 0 isol_n
rlabel metal1 11132 3026 11132 3026 0 net1
rlabel metal2 2714 10115 2714 10115 0 net10
rlabel metal1 33902 14246 33902 14246 0 net100
rlabel metal1 36938 16422 36938 16422 0 net101
rlabel metal1 34086 13226 34086 13226 0 net102
rlabel metal1 41538 16728 41538 16728 0 net103
rlabel metal1 17296 15334 17296 15334 0 net104
rlabel metal1 16054 17068 16054 17068 0 net105
rlabel metal3 44551 20876 44551 20876 0 net106
rlabel metal2 19366 19533 19366 19533 0 net107
rlabel metal1 41998 20774 41998 20774 0 net108
rlabel metal1 26910 15130 26910 15130 0 net109
rlabel metal1 2530 8840 2530 8840 0 net11
rlabel metal2 26450 24514 26450 24514 0 net110
rlabel metal1 39514 2414 39514 2414 0 net111
rlabel metal1 8050 18938 8050 18938 0 net112
rlabel metal1 2990 13362 2990 13362 0 net113
rlabel metal1 11316 17170 11316 17170 0 net114
rlabel metal2 9246 17816 9246 17816 0 net115
rlabel metal1 3174 19822 3174 19822 0 net116
rlabel via2 16054 19261 16054 19261 0 net117
rlabel metal1 11546 19278 11546 19278 0 net118
rlabel metal1 6670 18326 6670 18326 0 net119
rlabel metal1 4393 9078 4393 9078 0 net12
rlabel metal1 8096 20026 8096 20026 0 net120
rlabel metal2 12466 21539 12466 21539 0 net121
rlabel metal1 2990 22576 2990 22576 0 net122
rlabel metal1 2990 23120 2990 23120 0 net123
rlabel metal1 2990 13940 2990 13940 0 net124
rlabel metal1 11316 20434 11316 20434 0 net125
rlabel metal1 5382 20978 5382 20978 0 net126
rlabel metal1 9522 20944 9522 20944 0 net127
rlabel metal1 7544 20910 7544 20910 0 net128
rlabel metal1 6072 20570 6072 20570 0 net129
rlabel via2 1794 9435 1794 9435 0 net13
rlabel metal1 11408 22474 11408 22474 0 net130
rlabel metal1 7222 19754 7222 19754 0 net131
rlabel metal1 4830 22474 4830 22474 0 net132
rlabel metal1 7222 21386 7222 21386 0 net133
rlabel metal1 8004 22474 8004 22474 0 net134
rlabel metal1 6256 14382 6256 14382 0 net135
rlabel metal1 3588 14994 3588 14994 0 net136
rlabel metal2 10258 14994 10258 14994 0 net137
rlabel metal2 10902 15606 10902 15606 0 net138
rlabel metal2 14214 16864 14214 16864 0 net139
rlabel metal1 19527 2550 19527 2550 0 net14
rlabel metal1 3680 17170 3680 17170 0 net140
rlabel metal1 10304 16694 10304 16694 0 net141
rlabel metal1 10396 16218 10396 16218 0 net142
rlabel metal2 45862 3808 45862 3808 0 net143
rlabel metal1 47656 4590 47656 4590 0 net144
rlabel metal1 47932 5202 47932 5202 0 net145
rlabel metal2 40158 7276 40158 7276 0 net146
rlabel metal2 45494 8534 45494 8534 0 net147
rlabel metal1 47840 6290 47840 6290 0 net148
rlabel metal1 47886 6766 47886 6766 0 net149
rlabel metal2 2162 13566 2162 13566 0 net15
rlabel metal1 45402 8568 45402 8568 0 net150
rlabel metal2 47058 8738 47058 8738 0 net151
rlabel metal2 46966 9180 46966 9180 0 net152
rlabel metal2 46230 9214 46230 9214 0 net153
rlabel metal2 39790 3740 39790 3740 0 net154
rlabel metal2 45770 10540 45770 10540 0 net155
rlabel metal1 42826 11560 42826 11560 0 net156
rlabel metal2 47150 10948 47150 10948 0 net157
rlabel metal2 46782 10812 46782 10812 0 net158
rlabel metal1 47472 10642 47472 10642 0 net159
rlabel metal2 2530 11288 2530 11288 0 net16
rlabel metal2 42734 11934 42734 11934 0 net160
rlabel metal1 47058 11730 47058 11730 0 net161
rlabel metal2 47978 12410 47978 12410 0 net162
rlabel metal1 47518 12818 47518 12818 0 net163
rlabel metal2 46322 13566 46322 13566 0 net164
rlabel metal2 45678 3332 45678 3332 0 net165
rlabel metal2 45770 4318 45770 4318 0 net166
rlabel metal1 46138 3536 46138 3536 0 net167
rlabel metal2 47150 3604 47150 3604 0 net168
rlabel metal2 47242 4454 47242 4454 0 net169
rlabel metal1 4347 10506 4347 10506 0 net17
rlabel metal2 47058 4828 47058 4828 0 net170
rlabel metal1 42090 7208 42090 7208 0 net171
rlabel metal1 47472 4114 47472 4114 0 net172
rlabel metal1 7222 23222 7222 23222 0 net173
rlabel metal1 7682 24174 7682 24174 0 net174
rlabel metal1 9338 23732 9338 23732 0 net175
rlabel metal2 11178 23324 11178 23324 0 net176
rlabel metal1 11178 23664 11178 23664 0 net177
rlabel metal1 12144 22202 12144 22202 0 net178
rlabel metal1 11178 24140 11178 24140 0 net179
rlabel metal1 4347 11254 4347 11254 0 net18
rlabel metal1 14352 22610 14352 22610 0 net180
rlabel metal1 13892 21658 13892 21658 0 net181
rlabel metal1 14398 22066 14398 22066 0 net182
rlabel metal1 13110 23630 13110 23630 0 net183
rlabel metal1 4370 22950 4370 22950 0 net184
rlabel metal1 16514 22610 16514 22610 0 net185
rlabel metal1 19596 19958 19596 19958 0 net186
rlabel metal2 19642 23528 19642 23528 0 net187
rlabel metal1 18814 21964 18814 21964 0 net188
rlabel metal1 20930 21590 20930 21590 0 net189
rlabel metal1 3358 11526 3358 11526 0 net19
rlabel metal1 18676 23698 18676 23698 0 net190
rlabel metal2 19458 23018 19458 23018 0 net191
rlabel metal2 18906 24446 18906 24446 0 net192
rlabel metal2 21482 24004 21482 24004 0 net193
rlabel metal1 21390 24208 21390 24208 0 net194
rlabel metal1 3680 24174 3680 24174 0 net195
rlabel metal1 4278 18258 4278 18258 0 net196
rlabel metal2 6026 23052 6026 23052 0 net197
rlabel metal2 4738 23494 4738 23494 0 net198
rlabel metal1 4508 22746 4508 22746 0 net199
rlabel metal2 46966 23426 46966 23426 0 net2
rlabel metal1 4048 12206 4048 12206 0 net20
rlabel metal1 3496 23834 3496 23834 0 net200
rlabel metal2 7498 23324 7498 23324 0 net201
rlabel metal2 5566 23562 5566 23562 0 net202
rlabel metal1 13570 2414 13570 2414 0 net203
rlabel metal1 16560 2414 16560 2414 0 net204
rlabel metal1 18492 2414 18492 2414 0 net205
rlabel metal1 19550 3094 19550 3094 0 net206
rlabel metal1 19872 2414 19872 2414 0 net207
rlabel metal1 22264 2414 22264 2414 0 net208
rlabel metal1 24610 2380 24610 2380 0 net209
rlabel metal1 6670 11594 6670 11594 0 net21
rlabel metal1 26910 2822 26910 2822 0 net210
rlabel metal1 16836 17646 16836 17646 0 net211
rlabel metal2 23690 13209 23690 13209 0 net212
rlabel metal2 27922 21250 27922 21250 0 net213
rlabel metal1 18768 14042 18768 14042 0 net214
rlabel metal2 24610 20910 24610 20910 0 net215
rlabel metal1 19504 13226 19504 13226 0 net216
rlabel metal1 31188 14246 31188 14246 0 net217
rlabel metal2 31142 7990 31142 7990 0 net218
rlabel metal1 31878 10608 31878 10608 0 net219
rlabel metal1 4370 23086 4370 23086 0 net22
rlabel metal2 33902 15232 33902 15232 0 net220
rlabel metal1 28934 13294 28934 13294 0 net221
rlabel metal2 29946 9282 29946 9282 0 net222
rlabel metal2 31418 7616 31418 7616 0 net223
rlabel metal1 33948 14042 33948 14042 0 net224
rlabel metal1 29164 8874 29164 8874 0 net225
rlabel metal1 27002 11866 27002 11866 0 net226
rlabel metal2 32706 8908 32706 8908 0 net227
rlabel metal1 29302 19346 29302 19346 0 net228
rlabel metal1 31372 15130 31372 15130 0 net229
rlabel metal2 9522 14858 9522 14858 0 net23
rlabel metal1 36478 17306 36478 17306 0 net230
rlabel metal1 36064 15130 36064 15130 0 net231
rlabel metal1 35834 13226 35834 13226 0 net232
rlabel metal1 31280 10778 31280 10778 0 net233
rlabel metal1 33120 21658 33120 21658 0 net234
rlabel metal1 25208 13294 25208 13294 0 net235
rlabel metal1 24104 13838 24104 13838 0 net236
rlabel metal1 20102 11186 20102 11186 0 net237
rlabel metal1 25024 10642 25024 10642 0 net238
rlabel metal2 22678 10880 22678 10880 0 net239
rlabel metal2 20286 19550 20286 19550 0 net24
rlabel metal1 18377 12750 18377 12750 0 net240
rlabel metal1 18124 8398 18124 8398 0 net241
rlabel metal1 19688 10098 19688 10098 0 net242
rlabel metal1 22310 7854 22310 7854 0 net243
rlabel metal1 30912 18258 30912 18258 0 net244
rlabel metal1 13018 13362 13018 13362 0 net245
rlabel metal1 14122 18326 14122 18326 0 net246
rlabel metal1 12880 18734 12880 18734 0 net247
rlabel metal1 10350 18394 10350 18394 0 net248
rlabel via2 14122 20587 14122 20587 0 net249
rlabel metal1 4370 2414 4370 2414 0 net25
rlabel metal1 10166 20978 10166 20978 0 net250
rlabel metal1 10074 23222 10074 23222 0 net251
rlabel metal1 35236 18734 35236 18734 0 net252
rlabel metal1 40710 20366 40710 20366 0 net253
rlabel metal2 18722 9792 18722 9792 0 net254
rlabel metal1 16698 10710 16698 10710 0 net255
rlabel metal1 11638 13906 11638 13906 0 net256
rlabel metal1 16376 14314 16376 14314 0 net257
rlabel metal1 21390 12206 21390 12206 0 net258
rlabel metal1 21436 11798 21436 11798 0 net259
rlabel metal1 12788 10438 12788 10438 0 net26
rlabel metal2 18538 19754 18538 19754 0 net260
rlabel metal1 18492 19686 18492 19686 0 net261
rlabel metal1 23276 17578 23276 17578 0 net262
rlabel metal2 45402 23664 45402 23664 0 net263
rlabel metal2 42090 19040 42090 19040 0 net264
rlabel metal1 42366 24174 42366 24174 0 net265
rlabel metal2 47150 23324 47150 23324 0 net266
rlabel metal1 43424 23018 43424 23018 0 net267
rlabel metal1 10028 2550 10028 2550 0 net268
rlabel metal1 13938 2958 13938 2958 0 net269
rlabel metal2 17158 14552 17158 14552 0 net27
rlabel metal1 2530 4182 2530 4182 0 net28
rlabel metal1 4393 3978 4393 3978 0 net29
rlabel metal1 5083 2550 5083 2550 0 net3
rlabel metal1 37812 6358 37812 6358 0 net30
rlabel metal1 15870 17238 15870 17238 0 net31
rlabel metal2 13386 8670 13386 8670 0 net32
rlabel metal2 48438 14552 48438 14552 0 net33
rlabel metal2 48346 17680 48346 17680 0 net34
rlabel metal2 48530 17901 48530 17901 0 net35
rlabel metal2 48438 18428 48438 18428 0 net36
rlabel metal1 15364 19822 15364 19822 0 net37
rlabel metal2 49174 19465 49174 19465 0 net38
rlabel metal1 41630 20366 41630 20366 0 net39
rlabel metal1 1794 5576 1794 5576 0 net4
rlabel metal2 48438 19822 48438 19822 0 net40
rlabel metal2 40250 21097 40250 21097 0 net41
rlabel metal2 49174 20944 49174 20944 0 net42
rlabel metal2 49082 21199 49082 21199 0 net43
rlabel metal2 49174 14535 49174 14535 0 net44
rlabel metal2 41630 21182 41630 21182 0 net45
rlabel metal1 16238 16422 16238 16422 0 net46
rlabel metal2 43608 21318 43608 21318 0 net47
rlabel metal1 20194 14382 20194 14382 0 net48
rlabel metal2 41814 21624 41814 21624 0 net49
rlabel metal1 6532 6154 6532 6154 0 net5
rlabel metal1 41170 22746 41170 22746 0 net50
rlabel metal1 11500 22678 11500 22678 0 net51
rlabel metal1 46000 22134 46000 22134 0 net52
rlabel metal1 47012 22406 47012 22406 0 net53
rlabel via2 26634 24123 26634 24123 0 net54
rlabel via2 49082 14365 49082 14365 0 net55
rlabel metal2 39790 15691 39790 15691 0 net56
rlabel metal1 48944 15674 48944 15674 0 net57
rlabel via2 49174 15963 49174 15963 0 net58
rlabel metal2 49174 16269 49174 16269 0 net59
rlabel metal1 2530 6664 2530 6664 0 net6
rlabel via2 49082 17085 49082 17085 0 net60
rlabel metal2 48438 17442 48438 17442 0 net61
rlabel metal2 49174 17085 49174 17085 0 net62
rlabel metal1 26818 19482 26818 19482 0 net63
rlabel metal1 28336 18258 28336 18258 0 net64
rlabel metal1 28520 19686 28520 19686 0 net65
rlabel metal2 32338 23800 32338 23800 0 net66
rlabel metal1 32982 24276 32982 24276 0 net67
rlabel metal1 32798 19414 32798 19414 0 net68
rlabel metal1 33166 19822 33166 19822 0 net69
rlabel metal2 1794 6494 1794 6494 0 net7
rlabel metal1 35420 19822 35420 19822 0 net70
rlabel metal2 40342 24378 40342 24378 0 net71
rlabel metal1 33672 21590 33672 21590 0 net72
rlabel metal1 31832 20502 31832 20502 0 net73
rlabel metal1 14582 21896 14582 21896 0 net74
rlabel metal2 41538 20417 41538 20417 0 net75
rlabel metal2 36110 18921 36110 18921 0 net76
rlabel metal1 42435 17782 42435 17782 0 net77
rlabel metal2 42826 20213 42826 20213 0 net78
rlabel metal2 40342 21573 40342 21573 0 net79
rlabel metal2 18078 14586 18078 14586 0 net8
rlabel metal2 31786 21335 31786 21335 0 net80
rlabel metal1 34316 19754 34316 19754 0 net81
rlabel metal1 34684 19822 34684 19822 0 net82
rlabel metal1 34730 21454 34730 21454 0 net83
rlabel via2 33534 21539 33534 21539 0 net84
rlabel metal2 12374 24038 12374 24038 0 net85
rlabel metal1 32614 15980 32614 15980 0 net86
rlabel metal1 32982 15572 32982 15572 0 net87
rlabel metal1 33304 17714 33304 17714 0 net88
rlabel metal1 25162 22202 25162 22202 0 net89
rlabel metal1 1794 7752 1794 7752 0 net9
rlabel metal1 27738 19244 27738 19244 0 net90
rlabel metal1 28704 21998 28704 21998 0 net91
rlabel metal1 28428 17306 28428 17306 0 net92
rlabel metal1 27738 3570 27738 3570 0 net93
rlabel metal1 29256 2550 29256 2550 0 net94
rlabel metal1 32890 2550 32890 2550 0 net95
rlabel metal1 33994 2618 33994 2618 0 net96
rlabel metal2 37766 2822 37766 2822 0 net97
rlabel metal1 45034 23290 45034 23290 0 net98
rlabel metal1 43838 2516 43838 2516 0 net99
rlabel metal2 39238 2132 39238 2132 0 prog_clk
rlabel metal1 44114 22066 44114 22066 0 prog_reset
rlabel metal1 43378 2278 43378 2278 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 45586 2098 45586 2098 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 47702 2336 47702 2336 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 46690 4488 46690 4488 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 28796 11254 28796 11254 0 sb_1__0_.mem_left_track_1.ccff_head
rlabel metal1 23644 18666 23644 18666 0 sb_1__0_.mem_left_track_1.ccff_tail
rlabel metal2 29302 19040 29302 19040 0 sb_1__0_.mem_left_track_1.mem_out\[0\]
rlabel metal1 24334 17102 24334 17102 0 sb_1__0_.mem_left_track_1.mem_out\[1\]
rlabel metal1 21344 14314 21344 14314 0 sb_1__0_.mem_left_track_11.ccff_head
rlabel metal2 19182 17816 19182 17816 0 sb_1__0_.mem_left_track_11.ccff_tail
rlabel metal1 21436 13362 21436 13362 0 sb_1__0_.mem_left_track_11.mem_out\[0\]
rlabel metal1 21068 17238 21068 17238 0 sb_1__0_.mem_left_track_11.mem_out\[1\]
rlabel metal1 18446 21114 18446 21114 0 sb_1__0_.mem_left_track_13.ccff_tail
rlabel metal1 21344 18054 21344 18054 0 sb_1__0_.mem_left_track_13.mem_out\[0\]
rlabel metal1 19274 18802 19274 18802 0 sb_1__0_.mem_left_track_13.mem_out\[1\]
rlabel metal1 18262 21454 18262 21454 0 sb_1__0_.mem_left_track_21.ccff_tail
rlabel metal1 21528 18802 21528 18802 0 sb_1__0_.mem_left_track_21.mem_out\[0\]
rlabel metal1 19366 19890 19366 19890 0 sb_1__0_.mem_left_track_21.mem_out\[1\]
rlabel metal1 21390 19244 21390 19244 0 sb_1__0_.mem_left_track_29.ccff_tail
rlabel metal1 24196 20366 24196 20366 0 sb_1__0_.mem_left_track_29.mem_out\[0\]
rlabel metal2 24978 18496 24978 18496 0 sb_1__0_.mem_left_track_29.mem_out\[1\]
rlabel metal1 18860 20570 18860 20570 0 sb_1__0_.mem_left_track_3.ccff_tail
rlabel metal2 27646 21862 27646 21862 0 sb_1__0_.mem_left_track_3.mem_out\[0\]
rlabel metal1 17112 20366 17112 20366 0 sb_1__0_.mem_left_track_3.mem_out\[1\]
rlabel metal1 25760 16626 25760 16626 0 sb_1__0_.mem_left_track_37.ccff_tail
rlabel metal1 28244 18870 28244 18870 0 sb_1__0_.mem_left_track_37.mem_out\[0\]
rlabel metal1 26772 16626 26772 16626 0 sb_1__0_.mem_left_track_37.mem_out\[1\]
rlabel metal2 24886 23324 24886 23324 0 sb_1__0_.mem_left_track_45.ccff_tail
rlabel metal1 32890 22508 32890 22508 0 sb_1__0_.mem_left_track_45.mem_out\[0\]
rlabel metal1 28520 22066 28520 22066 0 sb_1__0_.mem_left_track_45.mem_out\[1\]
rlabel metal1 17986 16082 17986 16082 0 sb_1__0_.mem_left_track_5.ccff_tail
rlabel metal2 21114 20978 21114 20978 0 sb_1__0_.mem_left_track_5.mem_out\[0\]
rlabel metal1 18777 16762 18777 16762 0 sb_1__0_.mem_left_track_5.mem_out\[1\]
rlabel metal1 27462 22984 27462 22984 0 sb_1__0_.mem_left_track_53.mem_out\[0\]
rlabel metal1 23000 22066 23000 22066 0 sb_1__0_.mem_left_track_53.mem_out\[1\]
rlabel metal2 21942 14892 21942 14892 0 sb_1__0_.mem_left_track_7.mem_out\[0\]
rlabel metal2 22034 14688 22034 14688 0 sb_1__0_.mem_left_track_7.mem_out\[1\]
rlabel metal1 17480 21998 17480 21998 0 sb_1__0_.mem_right_track_0.ccff_head
rlabel metal2 32614 16388 32614 16388 0 sb_1__0_.mem_right_track_0.ccff_tail
rlabel metal1 29532 20366 29532 20366 0 sb_1__0_.mem_right_track_0.mem_out\[0\]
rlabel metal1 30452 15878 30452 15878 0 sb_1__0_.mem_right_track_0.mem_out\[1\]
rlabel metal1 37950 11050 37950 11050 0 sb_1__0_.mem_right_track_10.ccff_head
rlabel metal2 36662 10948 36662 10948 0 sb_1__0_.mem_right_track_10.ccff_tail
rlabel metal1 32890 15504 32890 15504 0 sb_1__0_.mem_right_track_10.mem_out\[0\]
rlabel metal1 34638 13804 34638 13804 0 sb_1__0_.mem_right_track_10.mem_out\[1\]
rlabel metal1 33120 13226 33120 13226 0 sb_1__0_.mem_right_track_12.ccff_tail
rlabel metal2 32430 15181 32430 15181 0 sb_1__0_.mem_right_track_12.mem_out\[0\]
rlabel metal1 31832 12954 31832 12954 0 sb_1__0_.mem_right_track_12.mem_out\[1\]
rlabel metal1 36800 16014 36800 16014 0 sb_1__0_.mem_right_track_2.ccff_tail
rlabel metal2 33534 21114 33534 21114 0 sb_1__0_.mem_right_track_2.mem_out\[0\]
rlabel metal1 35558 15538 35558 15538 0 sb_1__0_.mem_right_track_2.mem_out\[1\]
rlabel metal1 33626 11696 33626 11696 0 sb_1__0_.mem_right_track_20.ccff_tail
rlabel metal1 30038 17136 30038 17136 0 sb_1__0_.mem_right_track_20.mem_out\[0\]
rlabel metal1 29808 14926 29808 14926 0 sb_1__0_.mem_right_track_20.mem_out\[1\]
rlabel metal2 31878 9146 31878 9146 0 sb_1__0_.mem_right_track_28.ccff_tail
rlabel metal1 27324 9962 27324 9962 0 sb_1__0_.mem_right_track_28.mem_out\[0\]
rlabel metal1 30130 10574 30130 10574 0 sb_1__0_.mem_right_track_28.mem_out\[1\]
rlabel metal1 33994 8602 33994 8602 0 sb_1__0_.mem_right_track_36.ccff_tail
rlabel metal1 31924 14450 31924 14450 0 sb_1__0_.mem_right_track_36.mem_out\[0\]
rlabel metal1 32430 8398 32430 8398 0 sb_1__0_.mem_right_track_36.mem_out\[1\]
rlabel metal2 38226 13634 38226 13634 0 sb_1__0_.mem_right_track_4.ccff_tail
rlabel metal2 36846 16694 36846 16694 0 sb_1__0_.mem_right_track_4.mem_out\[0\]
rlabel metal2 36662 15674 36662 15674 0 sb_1__0_.mem_right_track_4.mem_out\[1\]
rlabel metal2 32798 9758 32798 9758 0 sb_1__0_.mem_right_track_44.ccff_tail
rlabel metal1 30038 16626 30038 16626 0 sb_1__0_.mem_right_track_44.mem_out\[0\]
rlabel metal1 28842 17068 28842 17068 0 sb_1__0_.mem_right_track_52.mem_out\[0\]
rlabel metal1 39422 12750 39422 12750 0 sb_1__0_.mem_right_track_6.mem_out\[0\]
rlabel metal2 36156 14926 36156 14926 0 sb_1__0_.mem_right_track_6.mem_out\[1\]
rlabel metal2 30314 23324 30314 23324 0 sb_1__0_.mem_top_track_0.ccff_tail
rlabel via1 35006 22073 35006 22073 0 sb_1__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 32522 21862 32522 21862 0 sb_1__0_.mem_top_track_0.mem_out\[1\]
rlabel metal1 37214 21114 37214 21114 0 sb_1__0_.mem_top_track_10.ccff_head
rlabel metal1 34040 18666 34040 18666 0 sb_1__0_.mem_top_track_10.ccff_tail
rlabel metal2 37766 19720 37766 19720 0 sb_1__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 34270 18190 34270 18190 0 sb_1__0_.mem_top_track_10.mem_out\[1\]
rlabel metal1 41538 18632 41538 18632 0 sb_1__0_.mem_top_track_12.ccff_tail
rlabel metal2 39422 19176 39422 19176 0 sb_1__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 37950 17102 37950 17102 0 sb_1__0_.mem_top_track_12.mem_out\[1\]
rlabel metal1 38548 16150 38548 16150 0 sb_1__0_.mem_top_track_14.ccff_tail
rlabel metal1 40112 18598 40112 18598 0 sb_1__0_.mem_top_track_14.mem_out\[0\]
rlabel metal1 38364 16626 38364 16626 0 sb_1__0_.mem_top_track_14.mem_out\[1\]
rlabel metal2 37766 16932 37766 16932 0 sb_1__0_.mem_top_track_16.ccff_tail
rlabel metal1 40158 15878 40158 15878 0 sb_1__0_.mem_top_track_16.mem_out\[0\]
rlabel metal2 41814 15810 41814 15810 0 sb_1__0_.mem_top_track_16.mem_out\[1\]
rlabel metal2 32338 14382 32338 14382 0 sb_1__0_.mem_top_track_18.ccff_tail
rlabel metal1 38594 14280 38594 14280 0 sb_1__0_.mem_top_track_18.mem_out\[0\]
rlabel metal2 37122 14756 37122 14756 0 sb_1__0_.mem_top_track_18.mem_out\[1\]
rlabel metal1 34086 23494 34086 23494 0 sb_1__0_.mem_top_track_2.ccff_tail
rlabel metal1 32437 19788 32437 19788 0 sb_1__0_.mem_top_track_2.mem_out\[0\]
rlabel metal1 35190 23630 35190 23630 0 sb_1__0_.mem_top_track_2.mem_out\[1\]
rlabel metal1 25576 14586 25576 14586 0 sb_1__0_.mem_top_track_20.ccff_tail
rlabel metal2 27094 13838 27094 13838 0 sb_1__0_.mem_top_track_20.mem_out\[0\]
rlabel metal1 23736 12750 23736 12750 0 sb_1__0_.mem_top_track_22.ccff_tail
rlabel metal1 25116 14042 25116 14042 0 sb_1__0_.mem_top_track_22.mem_out\[0\]
rlabel metal1 24656 11186 24656 11186 0 sb_1__0_.mem_top_track_24.ccff_tail
rlabel metal1 26634 12342 26634 12342 0 sb_1__0_.mem_top_track_24.mem_out\[0\]
rlabel metal1 22770 13396 22770 13396 0 sb_1__0_.mem_top_track_26.ccff_tail
rlabel metal1 27324 15538 27324 15538 0 sb_1__0_.mem_top_track_26.mem_out\[0\]
rlabel metal1 21390 10506 21390 10506 0 sb_1__0_.mem_top_track_28.ccff_tail
rlabel metal1 23644 9350 23644 9350 0 sb_1__0_.mem_top_track_28.mem_out\[0\]
rlabel metal1 19826 8602 19826 8602 0 sb_1__0_.mem_top_track_30.ccff_tail
rlabel metal1 21620 8602 21620 8602 0 sb_1__0_.mem_top_track_30.mem_out\[0\]
rlabel metal1 19596 9622 19596 9622 0 sb_1__0_.mem_top_track_32.ccff_tail
rlabel metal2 19458 9078 19458 9078 0 sb_1__0_.mem_top_track_32.mem_out\[0\]
rlabel metal1 20102 12750 20102 12750 0 sb_1__0_.mem_top_track_34.ccff_tail
rlabel metal2 21114 10132 21114 10132 0 sb_1__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 20884 11186 20884 11186 0 sb_1__0_.mem_top_track_36.ccff_tail
rlabel metal1 25622 14926 25622 14926 0 sb_1__0_.mem_top_track_36.mem_out\[0\]
rlabel metal2 32338 20672 32338 20672 0 sb_1__0_.mem_top_track_4.ccff_tail
rlabel metal2 36386 20672 36386 20672 0 sb_1__0_.mem_top_track_4.mem_out\[0\]
rlabel metal1 33212 20366 33212 20366 0 sb_1__0_.mem_top_track_4.mem_out\[1\]
rlabel metal2 13294 14212 13294 14212 0 sb_1__0_.mem_top_track_40.ccff_tail
rlabel metal1 14582 12376 14582 12376 0 sb_1__0_.mem_top_track_40.mem_out\[0\]
rlabel metal2 14582 18428 14582 18428 0 sb_1__0_.mem_top_track_42.ccff_tail
rlabel metal1 16928 15538 16928 15538 0 sb_1__0_.mem_top_track_42.mem_out\[0\]
rlabel metal1 12926 18802 12926 18802 0 sb_1__0_.mem_top_track_44.ccff_tail
rlabel metal1 15640 18938 15640 18938 0 sb_1__0_.mem_top_track_44.mem_out\[0\]
rlabel metal2 10994 19006 10994 19006 0 sb_1__0_.mem_top_track_46.ccff_tail
rlabel metal1 12466 14892 12466 14892 0 sb_1__0_.mem_top_track_46.mem_out\[0\]
rlabel metal2 14306 21352 14306 21352 0 sb_1__0_.mem_top_track_48.ccff_tail
rlabel metal1 15962 20842 15962 20842 0 sb_1__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 16192 22678 16192 22678 0 sb_1__0_.mem_top_track_50.ccff_tail
rlabel metal1 16928 21454 16928 21454 0 sb_1__0_.mem_top_track_50.mem_out\[0\]
rlabel metal2 18630 23698 18630 23698 0 sb_1__0_.mem_top_track_58.mem_out\[0\]
rlabel metal1 36846 23222 36846 23222 0 sb_1__0_.mem_top_track_6.ccff_tail
rlabel metal1 35374 20774 35374 20774 0 sb_1__0_.mem_top_track_6.mem_out\[0\]
rlabel metal2 37490 23018 37490 23018 0 sb_1__0_.mem_top_track_6.mem_out\[1\]
rlabel metal1 37352 21862 37352 21862 0 sb_1__0_.mem_top_track_8.mem_out\[0\]
rlabel metal1 39100 20842 39100 20842 0 sb_1__0_.mem_top_track_8.mem_out\[1\]
rlabel metal2 7268 22100 7268 22100 0 sb_1__0_.mux_left_track_1.out
rlabel metal2 26358 18428 26358 18428 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 26772 18394 26772 18394 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 23414 14484 23414 14484 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22494 12376 22494 12376 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 25070 17884 25070 17884 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24288 16218 24288 16218 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 21574 18020 21574 18020 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 8326 18360 8326 18360 0 sb_1__0_.mux_left_track_11.out
rlabel metal1 22862 18258 22862 18258 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24150 18394 24150 18394 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20930 14246 20930 14246 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20792 13668 20792 13668 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20930 18088 20930 18088 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 19504 15130 19504 15130 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 15226 18394 15226 18394 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 15916 16218 15916 16218 0 sb_1__0_.mux_left_track_13.out
rlabel metal2 21942 21760 21942 21760 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23874 21658 23874 21658 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21160 15334 21160 15334 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21482 21046 21482 21046 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18032 18938 18032 18938 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10810 19754 10810 19754 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 9706 21318 9706 21318 0 sb_1__0_.mux_left_track_21.out
rlabel metal2 27922 23562 27922 23562 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24150 22066 24150 22066 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20930 18938 20930 18938 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19458 21658 19458 21658 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18262 19686 18262 19686 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12558 21624 12558 21624 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 13616 17510 13616 17510 0 sb_1__0_.mux_left_track_29.out
rlabel metal2 26174 20910 26174 20910 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 26818 20434 26818 20434 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23966 15130 23966 15130 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21252 19482 21252 19482 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22816 17782 22816 17782 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13754 17578 13754 17578 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 9982 20740 9982 20740 0 sb_1__0_.mux_left_track_3.out
rlabel metal1 26680 21862 26680 21862 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22494 18632 22494 18632 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19734 18938 19734 18938 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17388 17850 17388 17850 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13570 19924 13570 19924 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18446 15368 18446 15368 0 sb_1__0_.mux_left_track_37.out
rlabel metal2 32154 19006 32154 19006 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 29256 18394 29256 18394 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23782 16660 23782 16660 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23874 13498 23874 13498 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 20930 15810 20930 15810 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8326 18768 8326 18768 0 sb_1__0_.mux_left_track_45.out
rlabel metal1 29670 21930 29670 21930 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 28336 22202 28336 22202 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 27324 21318 27324 21318 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23322 23001 23322 23001 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 5658 22644 5658 22644 0 sb_1__0_.mux_left_track_5.out
rlabel metal1 24058 20026 24058 20026 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24242 18122 24242 18122 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17894 15980 17894 15980 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 18354 15130 18354 15130 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16744 16218 16744 16218 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 12834 15946 12834 15946 0 sb_1__0_.mux_left_track_53.out
rlabel metal1 26542 21998 26542 21998 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21298 20808 21298 20808 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20792 20910 20792 20910 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13754 20944 13754 20944 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 14766 16014 14766 16014 0 sb_1__0_.mux_left_track_7.out
rlabel metal1 25484 15470 25484 15470 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24104 15402 24104 15402 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20148 11866 20148 11866 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20378 15572 20378 15572 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20378 13498 20378 13498 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 19642 15606 19642 15606 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 39514 14110 39514 14110 0 sb_1__0_.mux_right_track_0.out
rlabel metal1 30820 17238 30820 17238 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33350 13396 33350 13396 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 29900 14314 29900 14314 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 33810 16592 33810 16592 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 31694 15334 31694 15334 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 39146 14382 39146 14382 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 43539 11118 43539 11118 0 sb_1__0_.mux_right_track_10.out
rlabel metal1 34500 13906 34500 13906 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34316 13974 34316 13974 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35236 9146 35236 9146 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32292 8602 32292 8602 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 35696 13906 35696 13906 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 36846 11254 36846 11254 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 40526 11118 40526 11118 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 40986 11934 40986 11934 0 sb_1__0_.mux_right_track_12.out
rlabel metal1 33626 14484 33626 14484 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33350 14382 33350 14382 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32154 10472 32154 10472 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 36064 14450 36064 14450 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 34914 10778 34914 10778 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 39330 12206 39330 12206 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 45678 14348 45678 14348 0 sb_1__0_.mux_right_track_2.out
rlabel metal1 36064 19414 36064 19414 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34316 18394 34316 18394 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 33810 14756 33810 14756 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37490 17510 37490 17510 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 35880 14790 35880 14790 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 40894 16388 40894 16388 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 44252 10030 44252 10030 0 sb_1__0_.mux_right_track_20.out
rlabel metal2 30866 18190 30866 18190 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 30774 16218 30774 16218 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28336 11866 28336 11866 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33810 11764 33810 11764 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 33856 11866 33856 11866 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 38226 11220 38226 11220 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 44206 8772 44206 8772 0 sb_1__0_.mux_right_track_28.out
rlabel metal1 30268 13362 30268 13362 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 30176 13294 30176 13294 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 26450 9452 26450 9452 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 31510 13158 31510 13158 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32384 9690 32384 9690 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 37674 8976 37674 8976 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 44942 7854 44942 7854 0 sb_1__0_.mux_right_track_36.out
rlabel metal1 32108 17510 32108 17510 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 32844 14246 32844 14246 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35006 8942 35006 8942 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33534 8058 33534 8058 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 38962 8500 38962 8500 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 45954 12988 45954 12988 0 sb_1__0_.mux_right_track_4.out
rlabel metal1 35742 17170 35742 17170 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36340 16762 36340 16762 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32982 11628 32982 11628 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37260 13974 37260 13974 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 37168 14042 37168 14042 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 41354 13668 41354 13668 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 40066 7480 40066 7480 0 sb_1__0_.mux_right_track_44.out
rlabel metal2 31970 15198 31970 15198 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 32430 9520 32430 9520 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36662 8466 36662 8466 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 43746 7412 43746 7412 0 sb_1__0_.mux_right_track_52.out
rlabel metal1 32660 12750 32660 12750 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 29762 12954 29762 12954 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33948 12682 33948 12682 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 43585 12070 43585 12070 0 sb_1__0_.mux_right_track_6.out
rlabel metal1 36110 15062 36110 15062 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 36294 15861 36294 15861 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36754 12682 36754 12682 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 36064 7990 36064 7990 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 38180 14790 38180 14790 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 38686 11968 38686 11968 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 41446 12240 41446 12240 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 23460 21998 23460 21998 0 sb_1__0_.mux_top_track_0.out
rlabel metal1 35834 21862 35834 21862 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38502 23562 38502 23562 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 25852 19958 25852 19958 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 28612 19482 28612 19482 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel via2 35466 23579 35466 23579 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 29624 20774 29624 20774 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 27485 23698 27485 23698 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 21390 21454 21390 21454 0 sb_1__0_.mux_top_track_10.out
rlabel metal1 36018 19482 36018 19482 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40112 19482 40112 19482 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 31970 18870 31970 18870 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 31694 17578 31694 17578 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 31004 18938 31004 18938 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal3 27462 22372 27462 22372 0 sb_1__0_.mux_top_track_12.out
rlabel metal1 40848 18394 40848 18394 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36846 20502 36846 20502 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37352 17034 37352 17034 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 36110 20519 36110 20519 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19826 22831 19826 22831 0 sb_1__0_.mux_top_track_14.out
rlabel metal1 40848 17714 40848 17714 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39514 17850 39514 17850 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36018 14858 36018 14858 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37490 18870 37490 18870 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 20378 19295 20378 19295 0 sb_1__0_.mux_top_track_16.out
rlabel metal2 40986 16320 40986 16320 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38824 16218 38824 16218 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35696 13498 35696 13498 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33718 18088 33718 18088 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24702 17782 24702 17782 0 sb_1__0_.mux_top_track_18.out
rlabel metal2 40158 15215 40158 15215 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 39698 14875 39698 14875 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32246 14994 32246 14994 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 31510 15096 31510 15096 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel via2 21298 23715 21298 23715 0 sb_1__0_.mux_top_track_2.out
rlabel metal1 36800 23766 36800 23766 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38962 23834 38962 23834 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 31694 19720 31694 19720 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 35144 23834 35144 23834 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32890 21862 32890 21862 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 28658 23766 28658 23766 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 7912 23698 7912 23698 0 sb_1__0_.mux_top_track_20.out
rlabel metal1 26358 17306 26358 17306 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 25622 15334 25622 15334 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24472 17306 24472 17306 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20102 16456 20102 16456 0 sb_1__0_.mux_top_track_22.out
rlabel metal1 24656 15062 24656 15062 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 23322 13158 23322 13158 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21206 16456 21206 16456 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15732 18122 15732 18122 0 sb_1__0_.mux_top_track_24.out
rlabel metal1 26956 15878 26956 15878 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23276 12138 23276 12138 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17894 15844 17894 15844 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19412 17850 19412 17850 0 sb_1__0_.mux_top_track_26.out
rlabel metal1 23092 13158 23092 13158 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22678 13226 22678 13226 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22172 13498 22172 13498 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14490 17306 14490 17306 0 sb_1__0_.mux_top_track_28.out
rlabel metal2 22310 10200 22310 10200 0 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 15847 13668 15847 13668 0 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12788 17850 12788 17850 0 sb_1__0_.mux_top_track_30.out
rlabel metal1 20930 7514 20930 7514 0 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13432 12716 13432 12716 0 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12788 20774 12788 20774 0 sb_1__0_.mux_top_track_32.out
rlabel metal1 18262 10234 18262 10234 0 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12742 16524 12742 16524 0 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13662 24140 13662 24140 0 sb_1__0_.mux_top_track_34.out
rlabel metal1 19642 10778 19642 10778 0 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19182 12954 19182 12954 0 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14490 22100 14490 22100 0 sb_1__0_.mux_top_track_36.out
rlabel metal1 21206 12716 21206 12716 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21988 8058 21988 8058 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19274 12682 19274 12682 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 27370 23290 27370 23290 0 sb_1__0_.mux_top_track_4.out
rlabel metal1 35742 20570 35742 20570 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36800 21658 36800 21658 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 35742 21216 35742 21216 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 31050 18394 31050 18394 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 30866 20808 30866 20808 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 4002 24140 4002 24140 0 sb_1__0_.mux_top_track_40.out
rlabel metal1 13018 10778 13018 10778 0 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11546 14586 11546 14586 0 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6739 24174 6739 24174 0 sb_1__0_.mux_top_track_42.out
rlabel metal2 16790 17000 16790 17000 0 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13846 18122 13846 18122 0 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2162 23732 2162 23732 0 sb_1__0_.mux_top_track_44.out
rlabel metal2 15594 17952 15594 17952 0 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12466 19584 12466 19584 0 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3450 18292 3450 18292 0 sb_1__0_.mux_top_track_46.out
rlabel metal1 11868 15130 11868 15130 0 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10074 18054 10074 18054 0 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4922 23018 4922 23018 0 sb_1__0_.mux_top_track_48.out
rlabel metal1 15962 19482 15962 19482 0 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9430 20876 9430 20876 0 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6854 23664 6854 23664 0 sb_1__0_.mux_top_track_50.out
rlabel metal1 16974 18904 16974 18904 0 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9062 21930 9062 21930 0 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9246 23086 9246 23086 0 sb_1__0_.mux_top_track_58.out
rlabel metal1 16928 24310 16928 24310 0 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11086 24208 11086 24208 0 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20562 24378 20562 24378 0 sb_1__0_.mux_top_track_6.out
rlabel metal2 40250 22610 40250 22610 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 41400 21862 41400 21862 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33718 18938 33718 18938 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 40066 23341 40066 23341 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 35604 22474 35604 22474 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 33626 24072 33626 24072 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 31510 22457 31510 22457 0 sb_1__0_.mux_top_track_8.out
rlabel metal1 40158 20978 40158 20978 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40848 20842 40848 20842 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34638 19482 34638 19482 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 40112 21114 40112 21114 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 36662 24106 36662 24106 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 33626 23001 33626 23001 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 45908 24174 45908 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
rlabel metal1 46598 24174 46598 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
rlabel metal2 46966 23936 46966 23936 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
rlabel metal1 47610 23086 47610 23086 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
rlabel metal2 48024 24174 48024 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
rlabel metal1 47978 21930 47978 21930 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
rlabel metal1 44252 23086 44252 23086 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
rlabel metal1 45080 24106 45080 24106 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
rlabel metal2 1150 2115 1150 2115 0 top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 3266 1299 3266 1299 0 top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 5382 2387 5382 2387 0 top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 7498 2234 7498 2234 0 top_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 27000
<< end >>
