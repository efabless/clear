magic
tech sky130A
magscale 1 2
timestamp 1682557524
<< viali >>
rect 1777 24361 1811 24395
rect 6561 24361 6595 24395
rect 27353 24361 27387 24395
rect 34161 24361 34195 24395
rect 36093 24361 36127 24395
rect 37473 24361 37507 24395
rect 44649 24361 44683 24395
rect 45845 24361 45879 24395
rect 47225 24361 47259 24395
rect 21189 24293 21223 24327
rect 27905 24293 27939 24327
rect 34897 24293 34931 24327
rect 48053 24293 48087 24327
rect 3249 24225 3283 24259
rect 5825 24225 5859 24259
rect 8217 24225 8251 24259
rect 10977 24225 11011 24259
rect 13553 24225 13587 24259
rect 18705 24225 18739 24259
rect 22477 24225 22511 24259
rect 28457 24225 28491 24259
rect 32965 24225 32999 24259
rect 35541 24225 35575 24259
rect 36737 24225 36771 24259
rect 38117 24225 38151 24259
rect 39129 24225 39163 24259
rect 39313 24225 39347 24259
rect 40693 24225 40727 24259
rect 42165 24225 42199 24259
rect 46949 24225 46983 24259
rect 48789 24225 48823 24259
rect 2145 24157 2179 24191
rect 4169 24157 4203 24191
rect 4629 24157 4663 24191
rect 6745 24157 6779 24191
rect 7389 24157 7423 24191
rect 9229 24157 9263 24191
rect 9781 24157 9815 24191
rect 12541 24157 12575 24191
rect 15117 24157 15151 24191
rect 17049 24157 17083 24191
rect 17693 24157 17727 24191
rect 19441 24157 19475 24191
rect 22109 24157 22143 24191
rect 24041 24157 24075 24191
rect 24869 24157 24903 24191
rect 25973 24157 26007 24191
rect 26617 24157 26651 24191
rect 28273 24157 28307 24191
rect 29193 24157 29227 24191
rect 29745 24157 29779 24191
rect 30849 24157 30883 24191
rect 33517 24157 33551 24191
rect 35357 24157 35391 24191
rect 36553 24157 36587 24191
rect 37933 24157 37967 24191
rect 41261 24157 41295 24191
rect 42625 24157 42659 24191
rect 43729 24157 43763 24191
rect 45201 24157 45235 24191
rect 46305 24157 46339 24191
rect 48513 24157 48547 24191
rect 1593 24089 1627 24123
rect 11713 24089 11747 24123
rect 11897 24089 11931 24123
rect 16129 24089 16163 24123
rect 19717 24089 19751 24123
rect 27261 24089 27295 24123
rect 28365 24089 28399 24123
rect 31769 24089 31803 24123
rect 32781 24089 32815 24123
rect 39037 24089 39071 24123
rect 40509 24089 40543 24123
rect 44373 24089 44407 24123
rect 47869 24089 47903 24123
rect 3985 24021 4019 24055
rect 9137 24021 9171 24055
rect 9413 24021 9447 24055
rect 12081 24021 12115 24055
rect 14289 24021 14323 24055
rect 16865 24021 16899 24055
rect 21557 24021 21591 24055
rect 23857 24021 23891 24055
rect 24501 24021 24535 24055
rect 25513 24021 25547 24055
rect 29009 24021 29043 24055
rect 29377 24021 29411 24055
rect 30389 24021 30423 24055
rect 31493 24021 31527 24055
rect 32321 24021 32355 24055
rect 32689 24021 32723 24055
rect 34437 24021 34471 24055
rect 35265 24021 35299 24055
rect 36461 24021 36495 24055
rect 37841 24021 37875 24055
rect 38669 24021 38703 24055
rect 40049 24021 40083 24055
rect 40417 24021 40451 24055
rect 41889 24021 41923 24055
rect 43269 24021 43303 24055
rect 48329 24021 48363 24055
rect 2329 23817 2363 23851
rect 27629 23817 27663 23851
rect 30297 23817 30331 23851
rect 30665 23817 30699 23851
rect 35357 23817 35391 23851
rect 36001 23817 36035 23851
rect 40049 23817 40083 23851
rect 41889 23817 41923 23851
rect 42257 23817 42291 23851
rect 45201 23817 45235 23851
rect 48053 23817 48087 23851
rect 3985 23749 4019 23783
rect 9137 23749 9171 23783
rect 10701 23749 10735 23783
rect 14289 23749 14323 23783
rect 16129 23749 16163 23783
rect 18981 23749 19015 23783
rect 19901 23749 19935 23783
rect 25145 23749 25179 23783
rect 29469 23749 29503 23783
rect 31769 23749 31803 23783
rect 33609 23749 33643 23783
rect 37749 23749 37783 23783
rect 46949 23749 46983 23783
rect 1685 23681 1719 23715
rect 2973 23681 3007 23715
rect 4813 23681 4847 23715
rect 6469 23681 6503 23715
rect 6561 23681 6595 23715
rect 8125 23681 8159 23715
rect 9965 23681 9999 23715
rect 11805 23681 11839 23715
rect 12081 23681 12115 23715
rect 13277 23681 13311 23715
rect 15025 23681 15059 23715
rect 16865 23681 16899 23715
rect 17325 23681 17359 23715
rect 17877 23681 17911 23715
rect 22201 23681 22235 23715
rect 24225 23681 24259 23715
rect 27997 23681 28031 23715
rect 28825 23681 28859 23715
rect 31585 23681 31619 23715
rect 32505 23681 32539 23715
rect 33333 23681 33367 23715
rect 35909 23681 35943 23715
rect 36369 23681 36403 23715
rect 40417 23681 40451 23715
rect 41245 23681 41279 23715
rect 42625 23681 42659 23715
rect 43729 23681 43763 23715
rect 44373 23681 44407 23715
rect 44649 23681 44683 23715
rect 45109 23681 45143 23715
rect 46029 23681 46063 23715
rect 47225 23681 47259 23715
rect 47869 23681 47903 23715
rect 48697 23681 48731 23715
rect 5457 23613 5491 23647
rect 6837 23613 6871 23647
rect 19625 23613 19659 23647
rect 22477 23613 22511 23647
rect 23765 23613 23799 23647
rect 24869 23613 24903 23647
rect 28089 23613 28123 23647
rect 28273 23613 28307 23647
rect 30757 23613 30791 23647
rect 30941 23613 30975 23647
rect 35541 23613 35575 23647
rect 36461 23613 36495 23647
rect 36645 23613 36679 23647
rect 37473 23613 37507 23647
rect 39497 23613 39531 23647
rect 40509 23613 40543 23647
rect 40693 23613 40727 23647
rect 43269 23613 43303 23647
rect 45753 23613 45787 23647
rect 48973 23613 49007 23647
rect 26617 23545 26651 23579
rect 44833 23545 44867 23579
rect 47133 23545 47167 23579
rect 17141 23477 17175 23511
rect 21373 23477 21407 23511
rect 24317 23477 24351 23511
rect 26985 23477 27019 23511
rect 27169 23477 27203 23511
rect 29745 23477 29779 23511
rect 30021 23477 30055 23511
rect 32781 23477 32815 23511
rect 35081 23477 35115 23511
rect 37013 23477 37047 23511
rect 47685 23477 47719 23511
rect 3617 23273 3651 23307
rect 14657 23273 14691 23307
rect 24777 23273 24811 23307
rect 37013 23273 37047 23307
rect 37368 23273 37402 23307
rect 39037 23273 39071 23307
rect 44373 23273 44407 23307
rect 45845 23273 45879 23307
rect 3433 23205 3467 23239
rect 3985 23205 4019 23239
rect 31677 23205 31711 23239
rect 34253 23205 34287 23239
rect 36645 23205 36679 23239
rect 38853 23205 38887 23239
rect 46949 23205 46983 23239
rect 47225 23205 47259 23239
rect 6101 23137 6135 23171
rect 7849 23137 7883 23171
rect 11253 23137 11287 23171
rect 13369 23137 13403 23171
rect 14197 23137 14231 23171
rect 16405 23137 16439 23171
rect 20821 23137 20855 23171
rect 23673 23137 23707 23171
rect 25697 23137 25731 23171
rect 28273 23137 28307 23171
rect 29101 23137 29135 23171
rect 32137 23137 32171 23171
rect 34529 23137 34563 23171
rect 34897 23137 34931 23171
rect 37105 23137 37139 23171
rect 41705 23137 41739 23171
rect 41981 23137 42015 23171
rect 48053 23137 48087 23171
rect 1777 23069 1811 23103
rect 4261 23069 4295 23103
rect 5365 23069 5399 23103
rect 7389 23069 7423 23103
rect 9413 23069 9447 23103
rect 10517 23069 10551 23103
rect 12541 23069 12575 23103
rect 14841 23069 14875 23103
rect 15485 23069 15519 23103
rect 17141 23069 17175 23103
rect 20177 23069 20211 23103
rect 23397 23069 23431 23103
rect 25421 23069 25455 23103
rect 28089 23069 28123 23103
rect 29929 23069 29963 23103
rect 39497 23069 39531 23103
rect 40049 23069 40083 23103
rect 40325 23069 40359 23103
rect 44281 23069 44315 23103
rect 45201 23069 45235 23103
rect 46305 23069 46339 23103
rect 47409 23069 47443 23103
rect 48513 23069 48547 23103
rect 2789 23001 2823 23035
rect 9137 23001 9171 23035
rect 17417 23001 17451 23035
rect 19441 23001 19475 23035
rect 21097 23001 21131 23035
rect 22845 23001 22879 23035
rect 24685 23001 24719 23035
rect 27997 23001 28031 23035
rect 28917 23001 28951 23035
rect 30205 23001 30239 23035
rect 32413 23001 32447 23035
rect 35173 23001 35207 23035
rect 43729 23001 43763 23035
rect 49157 23001 49191 23035
rect 4905 22933 4939 22967
rect 10057 22933 10091 22967
rect 14381 22933 14415 22967
rect 18889 22933 18923 22967
rect 27169 22933 27203 22967
rect 27629 22933 27663 22967
rect 29653 22933 29687 22967
rect 33885 22933 33919 22967
rect 39313 22933 39347 22967
rect 41153 22933 41187 22967
rect 41429 22933 41463 22967
rect 44833 22933 44867 22967
rect 49433 22933 49467 22967
rect 4169 22729 4203 22763
rect 6469 22729 6503 22763
rect 9321 22729 9355 22763
rect 22477 22729 22511 22763
rect 24041 22729 24075 22763
rect 32321 22729 32355 22763
rect 36093 22729 36127 22763
rect 36461 22729 36495 22763
rect 39681 22729 39715 22763
rect 40049 22729 40083 22763
rect 40877 22729 40911 22763
rect 41245 22729 41279 22763
rect 45753 22729 45787 22763
rect 46857 22729 46891 22763
rect 6653 22661 6687 22695
rect 6837 22661 6871 22695
rect 7021 22661 7055 22695
rect 9505 22661 9539 22695
rect 15853 22661 15887 22695
rect 22937 22661 22971 22695
rect 25145 22661 25179 22695
rect 27445 22661 27479 22695
rect 30757 22661 30791 22695
rect 44465 22661 44499 22695
rect 49157 22661 49191 22695
rect 1777 22593 1811 22627
rect 3525 22593 3559 22627
rect 4629 22593 4663 22627
rect 7665 22593 7699 22627
rect 9781 22593 9815 22627
rect 11989 22593 12023 22627
rect 13093 22593 13127 22627
rect 15117 22593 15151 22627
rect 19257 22593 19291 22627
rect 22845 22593 22879 22627
rect 24133 22593 24167 22627
rect 30665 22593 30699 22627
rect 31585 22593 31619 22627
rect 31769 22593 31803 22627
rect 32689 22593 32723 22627
rect 33609 22593 33643 22627
rect 37473 22593 37507 22627
rect 42625 22593 42659 22627
rect 43729 22593 43763 22627
rect 45109 22593 45143 22627
rect 46213 22593 46247 22627
rect 47777 22593 47811 22627
rect 48881 22593 48915 22627
rect 2789 22525 2823 22559
rect 5089 22525 5123 22559
rect 7941 22525 7975 22559
rect 10241 22525 10275 22559
rect 11713 22525 11747 22559
rect 13829 22525 13863 22559
rect 16865 22525 16899 22559
rect 17141 22525 17175 22559
rect 19533 22525 19567 22559
rect 21281 22525 21315 22559
rect 23029 22525 23063 22559
rect 24225 22525 24259 22559
rect 24869 22525 24903 22559
rect 28089 22525 28123 22559
rect 28365 22525 28399 22559
rect 30941 22525 30975 22559
rect 32781 22525 32815 22559
rect 32873 22525 32907 22559
rect 35357 22525 35391 22559
rect 36553 22525 36587 22559
rect 36645 22525 36679 22559
rect 37749 22525 37783 22559
rect 40141 22525 40175 22559
rect 40325 22525 40359 22559
rect 41337 22525 41371 22559
rect 41521 22525 41555 22559
rect 22109 22457 22143 22491
rect 26985 22457 27019 22491
rect 27629 22457 27663 22491
rect 30297 22457 30331 22491
rect 35725 22457 35759 22491
rect 39221 22457 39255 22491
rect 41889 22457 41923 22491
rect 47317 22457 47351 22491
rect 18613 22389 18647 22423
rect 18889 22389 18923 22423
rect 21557 22389 21591 22423
rect 22017 22389 22051 22423
rect 23673 22389 23707 22423
rect 26617 22389 26651 22423
rect 29837 22389 29871 22423
rect 33872 22389 33906 22423
rect 42073 22389 42107 22423
rect 43269 22389 43303 22423
rect 47133 22389 47167 22423
rect 48421 22389 48455 22423
rect 15282 22185 15316 22219
rect 23305 22185 23339 22219
rect 31112 22185 31146 22219
rect 38577 22185 38611 22219
rect 14565 22117 14599 22151
rect 33149 22117 33183 22151
rect 34437 22117 34471 22151
rect 37381 22117 37415 22151
rect 2053 22049 2087 22083
rect 4445 22049 4479 22083
rect 6285 22049 6319 22083
rect 9781 22049 9815 22083
rect 12449 22049 12483 22083
rect 15025 22049 15059 22083
rect 17969 22049 18003 22083
rect 20177 22049 20211 22083
rect 21373 22049 21407 22083
rect 22569 22049 22603 22083
rect 23765 22049 23799 22083
rect 23857 22049 23891 22083
rect 25329 22049 25363 22083
rect 26433 22049 26467 22083
rect 26525 22049 26559 22083
rect 30389 22049 30423 22083
rect 30849 22049 30883 22083
rect 33793 22049 33827 22083
rect 35541 22049 35575 22083
rect 36093 22049 36127 22083
rect 36829 22049 36863 22083
rect 38025 22049 38059 22083
rect 39129 22049 39163 22083
rect 40693 22049 40727 22083
rect 41797 22049 41831 22083
rect 43085 22049 43119 22083
rect 44189 22049 44223 22083
rect 44557 22049 44591 22083
rect 49433 22049 49467 22083
rect 1777 21981 1811 22015
rect 3985 21981 4019 22015
rect 5825 21981 5859 22015
rect 7941 21981 7975 22015
rect 9137 21981 9171 22015
rect 10977 21981 11011 22015
rect 11989 21981 12023 22015
rect 14841 21981 14875 22015
rect 17509 21981 17543 22015
rect 19993 21981 20027 22015
rect 22385 21981 22419 22015
rect 25145 21981 25179 22015
rect 27169 21981 27203 22015
rect 28549 21981 28583 22015
rect 29193 21981 29227 22015
rect 29745 21981 29779 22015
rect 36645 21981 36679 22015
rect 37749 21981 37783 22015
rect 41705 21981 41739 22015
rect 42441 21981 42475 22015
rect 43545 21981 43579 22015
rect 45201 21981 45235 22015
rect 46305 21981 46339 22015
rect 47409 21981 47443 22015
rect 48513 21981 48547 22015
rect 3617 21913 3651 21947
rect 11345 21913 11379 21947
rect 14381 21913 14415 21947
rect 21189 21913 21223 21947
rect 22477 21913 22511 21947
rect 25237 21913 25271 21947
rect 27905 21913 27939 21947
rect 35357 21913 35391 21947
rect 39037 21913 39071 21947
rect 40417 21913 40451 21947
rect 41613 21913 41647 21947
rect 3433 21845 3467 21879
rect 7665 21845 7699 21879
rect 8585 21845 8619 21879
rect 11437 21845 11471 21879
rect 13737 21845 13771 21879
rect 13829 21845 13863 21879
rect 16773 21845 16807 21879
rect 17141 21845 17175 21879
rect 19349 21845 19383 21879
rect 19625 21845 19659 21879
rect 20085 21845 20119 21879
rect 20821 21845 20855 21879
rect 21281 21845 21315 21879
rect 22017 21845 22051 21879
rect 23673 21845 23707 21879
rect 24501 21845 24535 21879
rect 24777 21845 24811 21879
rect 25973 21845 26007 21879
rect 26341 21845 26375 21879
rect 32597 21845 32631 21879
rect 33517 21845 33551 21879
rect 33609 21845 33643 21879
rect 34161 21845 34195 21879
rect 34897 21845 34931 21879
rect 35265 21845 35299 21879
rect 36185 21845 36219 21879
rect 36553 21845 36587 21879
rect 37841 21845 37875 21879
rect 38945 21845 38979 21879
rect 39589 21845 39623 21879
rect 40049 21845 40083 21879
rect 40509 21845 40543 21879
rect 41245 21845 41279 21879
rect 44649 21845 44683 21879
rect 45845 21845 45879 21879
rect 46949 21845 46983 21879
rect 48053 21845 48087 21879
rect 49157 21845 49191 21879
rect 6009 21641 6043 21675
rect 10149 21641 10183 21675
rect 12817 21641 12851 21675
rect 13921 21641 13955 21675
rect 14381 21641 14415 21675
rect 15945 21641 15979 21675
rect 16037 21641 16071 21675
rect 27169 21641 27203 21675
rect 28549 21641 28583 21675
rect 32321 21641 32355 21675
rect 32689 21641 32723 21675
rect 33425 21641 33459 21675
rect 36093 21641 36127 21675
rect 40509 21641 40543 21675
rect 40877 21641 40911 21675
rect 44373 21641 44407 21675
rect 46581 21641 46615 21675
rect 47041 21641 47075 21675
rect 49065 21641 49099 21675
rect 4353 21573 4387 21607
rect 18153 21573 18187 21607
rect 22293 21573 22327 21607
rect 26709 21573 26743 21607
rect 27629 21573 27663 21607
rect 30113 21573 30147 21607
rect 32781 21573 32815 21607
rect 34069 21573 34103 21607
rect 38577 21573 38611 21607
rect 40969 21573 41003 21607
rect 42073 21573 42107 21607
rect 1777 21505 1811 21539
rect 3433 21505 3467 21539
rect 5365 21505 5399 21539
rect 6561 21505 6595 21539
rect 8401 21505 8435 21539
rect 10517 21505 10551 21539
rect 12265 21505 12299 21539
rect 13277 21505 13311 21539
rect 14749 21505 14783 21539
rect 14841 21505 14875 21539
rect 16957 21505 16991 21539
rect 20453 21505 20487 21539
rect 21465 21505 21499 21539
rect 24317 21505 24351 21539
rect 26525 21505 26559 21539
rect 27537 21505 27571 21539
rect 28917 21505 28951 21539
rect 30205 21505 30239 21539
rect 31309 21505 31343 21539
rect 33793 21505 33827 21539
rect 36461 21505 36495 21539
rect 37657 21505 37691 21539
rect 37841 21505 37875 21539
rect 41889 21505 41923 21539
rect 42625 21505 42659 21539
rect 43729 21505 43763 21539
rect 44833 21505 44867 21539
rect 45937 21505 45971 21539
rect 47225 21505 47259 21539
rect 47777 21505 47811 21539
rect 48973 21505 49007 21539
rect 2789 21437 2823 21471
rect 7021 21437 7055 21471
rect 8861 21437 8895 21471
rect 11161 21437 11195 21471
rect 14933 21437 14967 21471
rect 16129 21437 16163 21471
rect 17233 21437 17267 21471
rect 17877 21437 17911 21471
rect 19625 21437 19659 21471
rect 20545 21437 20579 21471
rect 20729 21437 20763 21471
rect 22017 21437 22051 21471
rect 24593 21437 24627 21471
rect 27721 21437 27755 21471
rect 29009 21437 29043 21471
rect 29101 21437 29135 21471
rect 30297 21437 30331 21471
rect 31401 21437 31435 21471
rect 31493 21437 31527 21471
rect 32873 21437 32907 21471
rect 36553 21437 36587 21471
rect 36645 21437 36679 21471
rect 38301 21437 38335 21471
rect 41061 21437 41095 21471
rect 11805 21369 11839 21403
rect 23765 21369 23799 21403
rect 40049 21369 40083 21403
rect 45477 21369 45511 21403
rect 11621 21301 11655 21335
rect 15577 21301 15611 21335
rect 20085 21301 20119 21335
rect 21281 21301 21315 21335
rect 26065 21301 26099 21335
rect 26341 21301 26375 21335
rect 28273 21301 28307 21335
rect 29745 21301 29779 21335
rect 30941 21301 30975 21335
rect 35541 21301 35575 21335
rect 43269 21301 43303 21335
rect 48421 21301 48455 21335
rect 10333 21097 10367 21131
rect 11437 21097 11471 21131
rect 12541 21097 12575 21131
rect 23305 21097 23339 21131
rect 24685 21097 24719 21131
rect 28825 21097 28859 21131
rect 30941 21097 30975 21131
rect 40049 21097 40083 21131
rect 41889 21097 41923 21131
rect 49433 21097 49467 21131
rect 3433 21029 3467 21063
rect 9045 21029 9079 21063
rect 48053 21029 48087 21063
rect 4445 20961 4479 20995
rect 6745 20961 6779 20995
rect 8585 20961 8619 20995
rect 13553 20961 13587 20995
rect 14473 20961 14507 20995
rect 17417 20961 17451 20995
rect 17509 20961 17543 20995
rect 18797 20961 18831 20995
rect 19993 20961 20027 20995
rect 20177 20961 20211 20995
rect 21373 20961 21407 20995
rect 23857 20961 23891 20995
rect 25237 20961 25271 20995
rect 26341 20961 26375 20995
rect 26433 20961 26467 20995
rect 27997 20961 28031 20995
rect 30297 20961 30331 20995
rect 31585 20961 31619 20995
rect 32597 20961 32631 20995
rect 32781 20961 32815 20995
rect 33885 20961 33919 20995
rect 34897 20961 34931 20995
rect 35173 20961 35207 20995
rect 37749 20961 37783 20995
rect 38025 20961 38059 20995
rect 40693 20961 40727 20995
rect 44373 20961 44407 20995
rect 45845 20961 45879 20995
rect 1777 20893 1811 20927
rect 4077 20893 4111 20927
rect 5825 20893 5859 20927
rect 7941 20893 7975 20927
rect 9321 20893 9355 20927
rect 9689 20893 9723 20927
rect 10793 20893 10827 20927
rect 11897 20893 11931 20927
rect 14105 20893 14139 20927
rect 17325 20893 17359 20927
rect 18613 20893 18647 20927
rect 21097 20893 21131 20927
rect 23673 20893 23707 20927
rect 28733 20893 28767 20927
rect 30113 20893 30147 20927
rect 41245 20893 41279 20927
rect 42349 20893 42383 20927
rect 43453 20893 43487 20927
rect 44649 20893 44683 20927
rect 45201 20893 45235 20927
rect 46305 20893 46339 20927
rect 47409 20893 47443 20927
rect 48513 20893 48547 20927
rect 2789 20825 2823 20859
rect 12817 20825 12851 20859
rect 13369 20825 13403 20859
rect 13461 20825 13495 20859
rect 14749 20825 14783 20859
rect 18521 20825 18555 20859
rect 19901 20825 19935 20859
rect 27813 20825 27847 20859
rect 29193 20825 29227 20859
rect 31309 20825 31343 20859
rect 33701 20825 33735 20859
rect 44097 20825 44131 20859
rect 3617 20757 3651 20791
rect 7665 20757 7699 20791
rect 9229 20757 9263 20791
rect 13001 20757 13035 20791
rect 16221 20757 16255 20791
rect 16681 20757 16715 20791
rect 16957 20757 16991 20791
rect 18153 20757 18187 20791
rect 19533 20757 19567 20791
rect 20545 20757 20579 20791
rect 20729 20757 20763 20791
rect 22845 20757 22879 20791
rect 23765 20757 23799 20791
rect 25053 20757 25087 20791
rect 25145 20757 25179 20791
rect 25881 20757 25915 20791
rect 26249 20757 26283 20791
rect 26985 20757 27019 20791
rect 27077 20757 27111 20791
rect 27445 20757 27479 20791
rect 27905 20757 27939 20791
rect 29745 20757 29779 20791
rect 30205 20757 30239 20791
rect 31401 20757 31435 20791
rect 32137 20757 32171 20791
rect 32505 20757 32539 20791
rect 33333 20757 33367 20791
rect 33793 20757 33827 20791
rect 34437 20757 34471 20791
rect 36645 20757 36679 20791
rect 37105 20757 37139 20791
rect 39497 20757 39531 20791
rect 40417 20757 40451 20791
rect 40509 20757 40543 20791
rect 42993 20757 43027 20791
rect 44741 20757 44775 20791
rect 46949 20757 46983 20791
rect 49157 20757 49191 20791
rect 6009 20553 6043 20587
rect 11161 20553 11195 20587
rect 22017 20553 22051 20587
rect 25789 20553 25823 20587
rect 27169 20553 27203 20587
rect 29469 20553 29503 20587
rect 30297 20553 30331 20587
rect 37565 20553 37599 20587
rect 42073 20553 42107 20587
rect 43269 20553 43303 20587
rect 45477 20553 45511 20587
rect 47041 20553 47075 20587
rect 8401 20485 8435 20519
rect 8953 20485 8987 20519
rect 12081 20485 12115 20519
rect 15761 20485 15795 20519
rect 16313 20485 16347 20519
rect 23489 20485 23523 20519
rect 32597 20485 32631 20519
rect 34345 20485 34379 20519
rect 36553 20485 36587 20519
rect 38301 20485 38335 20519
rect 46581 20485 46615 20519
rect 1777 20417 1811 20451
rect 3617 20417 3651 20451
rect 5365 20417 5399 20451
rect 6561 20417 6595 20451
rect 8769 20417 8803 20451
rect 9413 20417 9447 20451
rect 10517 20417 10551 20451
rect 11897 20417 11931 20451
rect 12541 20417 12575 20451
rect 13645 20417 13679 20451
rect 16129 20417 16163 20451
rect 17141 20417 17175 20451
rect 19625 20417 19659 20451
rect 22385 20417 22419 20451
rect 23213 20417 23247 20451
rect 26157 20417 26191 20451
rect 27537 20417 27571 20451
rect 28365 20417 28399 20451
rect 31125 20417 31159 20451
rect 35265 20417 35299 20451
rect 36461 20417 36495 20451
rect 38025 20417 38059 20451
rect 40601 20417 40635 20451
rect 40693 20417 40727 20451
rect 41429 20417 41463 20451
rect 42625 20417 42659 20451
rect 43729 20417 43763 20451
rect 44833 20417 44867 20451
rect 45937 20417 45971 20451
rect 48053 20417 48087 20451
rect 49065 20417 49099 20451
rect 2789 20349 2823 20383
rect 3893 20349 3927 20383
rect 7021 20349 7055 20383
rect 13185 20349 13219 20383
rect 13921 20349 13955 20383
rect 17417 20349 17451 20383
rect 19901 20349 19935 20383
rect 22477 20349 22511 20383
rect 22569 20349 22603 20383
rect 26249 20349 26283 20383
rect 26341 20349 26375 20383
rect 27629 20349 27663 20383
rect 27721 20349 27755 20383
rect 30389 20349 30423 20383
rect 30481 20349 30515 20383
rect 32321 20349 32355 20383
rect 34069 20349 34103 20383
rect 35357 20349 35391 20383
rect 35541 20349 35575 20383
rect 36645 20349 36679 20383
rect 40877 20349 40911 20383
rect 44373 20349 44407 20383
rect 47777 20349 47811 20383
rect 15393 20281 15427 20315
rect 19349 20281 19383 20315
rect 25237 20281 25271 20315
rect 25421 20281 25455 20315
rect 34529 20281 34563 20315
rect 39773 20281 39807 20315
rect 46857 20281 46891 20315
rect 10057 20213 10091 20247
rect 16865 20213 16899 20247
rect 18889 20213 18923 20247
rect 21373 20213 21407 20247
rect 24961 20213 24995 20247
rect 29009 20213 29043 20247
rect 29285 20213 29319 20247
rect 29929 20213 29963 20247
rect 31769 20213 31803 20247
rect 34897 20213 34931 20247
rect 36093 20213 36127 20247
rect 37289 20213 37323 20247
rect 37657 20213 37691 20247
rect 40233 20213 40267 20247
rect 47225 20213 47259 20247
rect 49249 20213 49283 20247
rect 3433 20009 3467 20043
rect 3617 20009 3651 20043
rect 23213 20009 23247 20043
rect 29745 20009 29779 20043
rect 42993 20009 43027 20043
rect 44097 20009 44131 20043
rect 44741 20009 44775 20043
rect 45845 20009 45879 20043
rect 49157 20009 49191 20043
rect 11529 19941 11563 19975
rect 19533 19941 19567 19975
rect 22477 19941 22511 19975
rect 22937 19941 22971 19975
rect 28917 19941 28951 19975
rect 30941 19941 30975 19975
rect 36093 19941 36127 19975
rect 4905 19873 4939 19907
rect 6285 19873 6319 19907
rect 10425 19873 10459 19907
rect 16497 19873 16531 19907
rect 17049 19873 17083 19907
rect 18797 19873 18831 19907
rect 20177 19873 20211 19907
rect 20729 19873 20763 19907
rect 23765 19873 23799 19907
rect 24961 19873 24995 19907
rect 25237 19873 25271 19907
rect 27445 19873 27479 19907
rect 30389 19873 30423 19907
rect 32413 19873 32447 19907
rect 33517 19873 33551 19907
rect 36553 19873 36587 19907
rect 36737 19873 36771 19907
rect 39221 19873 39255 19907
rect 39313 19873 39347 19907
rect 40693 19873 40727 19907
rect 46949 19873 46983 19907
rect 1777 19805 1811 19839
rect 3985 19805 4019 19839
rect 6009 19805 6043 19839
rect 7941 19805 7975 19839
rect 9781 19805 9815 19839
rect 10885 19805 10919 19839
rect 11989 19805 12023 19839
rect 14565 19805 14599 19839
rect 19901 19805 19935 19839
rect 23673 19805 23707 19839
rect 27169 19805 27203 19839
rect 31125 19805 31159 19839
rect 34161 19805 34195 19839
rect 34989 19805 35023 19839
rect 39129 19805 39163 19839
rect 40417 19805 40451 19839
rect 41245 19805 41279 19839
rect 41889 19805 41923 19839
rect 42349 19805 42383 19839
rect 43453 19805 43487 19839
rect 45201 19805 45235 19839
rect 46305 19805 46339 19839
rect 47409 19805 47443 19839
rect 48513 19805 48547 19839
rect 2789 19737 2823 19771
rect 10701 19737 10735 19771
rect 12265 19737 12299 19771
rect 14289 19737 14323 19771
rect 15669 19737 15703 19771
rect 17325 19737 17359 19771
rect 21005 19737 21039 19771
rect 24593 19737 24627 19771
rect 30113 19737 30147 19771
rect 31585 19737 31619 19771
rect 33333 19737 33367 19771
rect 35357 19737 35391 19771
rect 36461 19737 36495 19771
rect 37381 19737 37415 19771
rect 38209 19737 38243 19771
rect 44373 19737 44407 19771
rect 44649 19737 44683 19771
rect 7665 19669 7699 19703
rect 8585 19669 8619 19703
rect 9137 19669 9171 19703
rect 13737 19669 13771 19703
rect 15209 19669 15243 19703
rect 19993 19669 20027 19703
rect 23581 19669 23615 19703
rect 24501 19669 24535 19703
rect 26709 19669 26743 19703
rect 29285 19669 29319 19703
rect 30205 19669 30239 19703
rect 32965 19669 32999 19703
rect 33425 19669 33459 19703
rect 38761 19669 38795 19703
rect 40049 19669 40083 19703
rect 40509 19669 40543 19703
rect 48053 19669 48087 19703
rect 49525 19669 49559 19703
rect 9965 19465 9999 19499
rect 10425 19465 10459 19499
rect 10885 19465 10919 19499
rect 12909 19465 12943 19499
rect 15577 19465 15611 19499
rect 22017 19465 22051 19499
rect 22385 19465 22419 19499
rect 24593 19465 24627 19499
rect 27905 19465 27939 19499
rect 28917 19465 28951 19499
rect 29285 19465 29319 19499
rect 30573 19465 30607 19499
rect 30941 19465 30975 19499
rect 32597 19465 32631 19499
rect 32965 19465 32999 19499
rect 34253 19465 34287 19499
rect 40785 19465 40819 19499
rect 43269 19465 43303 19499
rect 46581 19465 46615 19499
rect 4537 19397 4571 19431
rect 8861 19397 8895 19431
rect 11805 19397 11839 19431
rect 13829 19397 13863 19431
rect 20545 19397 20579 19431
rect 22477 19397 22511 19431
rect 30113 19397 30147 19431
rect 36001 19397 36035 19431
rect 38853 19397 38887 19431
rect 41153 19397 41187 19431
rect 45477 19397 45511 19431
rect 1777 19329 1811 19363
rect 3617 19329 3651 19363
rect 5365 19329 5399 19363
rect 6009 19329 6043 19363
rect 7113 19329 7147 19363
rect 7757 19329 7791 19363
rect 8217 19329 8251 19363
rect 9321 19329 9355 19363
rect 10333 19329 10367 19363
rect 10793 19329 10827 19363
rect 12817 19329 12851 19363
rect 14473 19329 14507 19363
rect 15117 19329 15151 19363
rect 15945 19329 15979 19363
rect 16037 19329 16071 19363
rect 16865 19329 16899 19363
rect 17969 19329 18003 19363
rect 19993 19329 20027 19363
rect 21281 19329 21315 19363
rect 23765 19329 23799 19363
rect 24961 19329 24995 19363
rect 25053 19329 25087 19363
rect 25973 19329 26007 19363
rect 26617 19329 26651 19363
rect 27077 19329 27111 19363
rect 29377 19329 29411 19363
rect 31309 19329 31343 19363
rect 31401 19329 31435 19363
rect 34161 19329 34195 19363
rect 34805 19329 34839 19363
rect 35265 19329 35299 19363
rect 36737 19329 36771 19363
rect 37461 19329 37495 19363
rect 38577 19329 38611 19363
rect 41245 19329 41279 19363
rect 42625 19329 42659 19363
rect 43717 19329 43751 19363
rect 44833 19329 44867 19363
rect 45937 19329 45971 19363
rect 48053 19329 48087 19363
rect 49157 19329 49191 19363
rect 2053 19261 2087 19295
rect 10977 19261 11011 19295
rect 11989 19261 12023 19295
rect 13001 19261 13035 19295
rect 14013 19261 14047 19295
rect 16129 19261 16163 19295
rect 18245 19261 18279 19295
rect 22569 19261 22603 19295
rect 23857 19261 23891 19295
rect 24041 19261 24075 19295
rect 25145 19261 25179 19295
rect 27997 19261 28031 19295
rect 28181 19261 28215 19295
rect 29561 19261 29595 19295
rect 31585 19261 31619 19295
rect 33057 19261 33091 19295
rect 33241 19261 33275 19295
rect 34345 19261 34379 19295
rect 41429 19261 41463 19295
rect 41981 19261 42015 19295
rect 47225 19261 47259 19295
rect 47777 19261 47811 19295
rect 6469 19193 6503 19227
rect 23397 19193 23431 19227
rect 25605 19193 25639 19227
rect 27169 19193 27203 19227
rect 28641 19193 28675 19227
rect 33793 19193 33827 19227
rect 35449 19193 35483 19227
rect 44373 19193 44407 19227
rect 46857 19193 46891 19227
rect 49341 19193 49375 19227
rect 6561 19125 6595 19159
rect 6837 19125 6871 19159
rect 11253 19125 11287 19159
rect 12265 19125 12299 19159
rect 12449 19125 12483 19159
rect 17509 19125 17543 19159
rect 23121 19125 23155 19159
rect 27537 19125 27571 19159
rect 32229 19125 32263 19159
rect 38117 19125 38151 19159
rect 40325 19125 40359 19159
rect 41889 19125 41923 19159
rect 42257 19125 42291 19159
rect 47041 19125 47075 19159
rect 47685 19125 47719 19159
rect 48697 19125 48731 19159
rect 3433 18921 3467 18955
rect 6285 18921 6319 18955
rect 7481 18921 7515 18955
rect 9045 18921 9079 18955
rect 10866 18921 10900 18955
rect 19625 18921 19659 18955
rect 20177 18921 20211 18955
rect 25513 18921 25547 18955
rect 29009 18921 29043 18955
rect 29745 18921 29779 18955
rect 44465 18921 44499 18955
rect 45845 18921 45879 18955
rect 47409 18921 47443 18955
rect 48421 18921 48455 18955
rect 49065 18921 49099 18955
rect 23121 18853 23155 18887
rect 24869 18853 24903 18887
rect 27905 18853 27939 18887
rect 32781 18853 32815 18887
rect 38025 18853 38059 18887
rect 39589 18853 39623 18887
rect 49433 18853 49467 18887
rect 4445 18785 4479 18819
rect 10149 18785 10183 18819
rect 14289 18785 14323 18819
rect 18429 18785 18463 18819
rect 20637 18785 20671 18819
rect 20821 18785 20855 18819
rect 23765 18785 23799 18819
rect 26065 18785 26099 18819
rect 27353 18785 27387 18819
rect 28549 18785 28583 18819
rect 30205 18785 30239 18819
rect 30297 18785 30331 18819
rect 32229 18785 32263 18819
rect 33241 18785 33275 18819
rect 33425 18785 33459 18819
rect 34345 18785 34379 18819
rect 35449 18785 35483 18819
rect 36001 18785 36035 18819
rect 36277 18785 36311 18819
rect 39129 18785 39163 18819
rect 46949 18785 46983 18819
rect 1777 18717 1811 18751
rect 3985 18717 4019 18751
rect 6837 18717 6871 18751
rect 7941 18717 7975 18751
rect 9505 18717 9539 18751
rect 10609 18717 10643 18751
rect 13093 18717 13127 18751
rect 18337 18717 18371 18751
rect 21373 18717 21407 18751
rect 23581 18717 23615 18751
rect 25881 18717 25915 18751
rect 27169 18717 27203 18751
rect 28273 18717 28307 18751
rect 29285 18717 29319 18751
rect 30113 18717 30147 18751
rect 31401 18717 31435 18751
rect 40049 18717 40083 18751
rect 42257 18717 42291 18751
rect 43361 18717 43395 18751
rect 44649 18717 44683 18751
rect 45201 18717 45235 18751
rect 46305 18717 46339 18751
rect 47777 18717 47811 18751
rect 2789 18649 2823 18683
rect 6193 18649 6227 18683
rect 14565 18649 14599 18683
rect 16497 18649 16531 18683
rect 17325 18649 17359 18683
rect 18245 18649 18279 18683
rect 19533 18649 19567 18683
rect 20545 18649 20579 18683
rect 22201 18649 22235 18683
rect 24685 18649 24719 18683
rect 25973 18649 26007 18683
rect 28365 18649 28399 18683
rect 30941 18649 30975 18683
rect 33149 18649 33183 18683
rect 34161 18649 34195 18683
rect 35265 18649 35299 18683
rect 35357 18649 35391 18683
rect 36553 18649 36587 18683
rect 40312 18649 40346 18683
rect 48973 18649 49007 18683
rect 3617 18581 3651 18615
rect 5825 18581 5859 18615
rect 8585 18581 8619 18615
rect 9137 18581 9171 18615
rect 12357 18581 12391 18615
rect 12817 18581 12851 18615
rect 13737 18581 13771 18615
rect 16037 18581 16071 18615
rect 17877 18581 17911 18615
rect 18981 18581 19015 18615
rect 22569 18581 22603 18615
rect 22753 18581 22787 18615
rect 23489 18581 23523 18615
rect 24133 18581 24167 18615
rect 25237 18581 25271 18615
rect 26709 18581 26743 18615
rect 27077 18581 27111 18615
rect 29193 18581 29227 18615
rect 30757 18581 30791 18615
rect 34897 18581 34931 18615
rect 38485 18581 38519 18615
rect 38853 18581 38887 18615
rect 38945 18581 38979 18615
rect 41797 18581 41831 18615
rect 42901 18581 42935 18615
rect 44005 18581 44039 18615
rect 47225 18581 47259 18615
rect 3341 18377 3375 18411
rect 3617 18377 3651 18411
rect 10977 18377 11011 18411
rect 16865 18377 16899 18411
rect 17325 18377 17359 18411
rect 18245 18377 18279 18411
rect 19165 18377 19199 18411
rect 22201 18377 22235 18411
rect 25513 18377 25547 18411
rect 25881 18377 25915 18411
rect 26801 18377 26835 18411
rect 30021 18377 30055 18411
rect 31033 18377 31067 18411
rect 33793 18377 33827 18411
rect 36185 18377 36219 18411
rect 36829 18377 36863 18411
rect 47225 18377 47259 18411
rect 49249 18377 49283 18411
rect 8769 18309 8803 18343
rect 10885 18309 10919 18343
rect 12909 18309 12943 18343
rect 19901 18309 19935 18343
rect 23121 18309 23155 18343
rect 33885 18309 33919 18343
rect 34713 18309 34747 18343
rect 41245 18309 41279 18343
rect 1777 18241 1811 18275
rect 3801 18241 3835 18275
rect 4261 18241 4295 18275
rect 5365 18241 5399 18275
rect 6929 18241 6963 18275
rect 7389 18241 7423 18275
rect 8493 18241 8527 18275
rect 11805 18241 11839 18275
rect 15209 18241 15243 18275
rect 16129 18241 16163 18275
rect 17233 18241 17267 18275
rect 18521 18241 18555 18275
rect 19625 18241 19659 18275
rect 22109 18241 22143 18275
rect 25237 18241 25271 18275
rect 26617 18241 26651 18275
rect 27169 18241 27203 18275
rect 29377 18241 29411 18275
rect 30941 18241 30975 18275
rect 32229 18241 32263 18275
rect 33057 18241 33091 18275
rect 36737 18241 36771 18275
rect 37473 18241 37507 18275
rect 41337 18241 41371 18275
rect 42625 18241 42659 18275
rect 43729 18241 43763 18275
rect 44373 18241 44407 18275
rect 44833 18241 44867 18275
rect 45937 18241 45971 18275
rect 48053 18241 48087 18275
rect 49065 18241 49099 18275
rect 2053 18173 2087 18207
rect 10241 18173 10275 18207
rect 12633 18173 12667 18207
rect 14381 18173 14415 18207
rect 15301 18173 15335 18207
rect 15485 18173 15519 18207
rect 17417 18173 17451 18207
rect 22845 18173 22879 18207
rect 24593 18173 24627 18207
rect 25973 18173 26007 18207
rect 26157 18173 26191 18207
rect 27445 18173 27479 18207
rect 31217 18173 31251 18207
rect 32321 18173 32355 18207
rect 33149 18173 33183 18207
rect 33241 18173 33275 18207
rect 34161 18173 34195 18207
rect 34437 18173 34471 18207
rect 38577 18173 38611 18207
rect 38853 18173 38887 18207
rect 41429 18173 41463 18207
rect 42073 18173 42107 18207
rect 47685 18173 47719 18207
rect 47777 18173 47811 18207
rect 6745 18105 6779 18139
rect 12357 18105 12391 18139
rect 40325 18105 40359 18139
rect 46581 18105 46615 18139
rect 46949 18105 46983 18139
rect 4905 18037 4939 18071
rect 6009 18037 6043 18071
rect 6469 18037 6503 18071
rect 8033 18037 8067 18071
rect 11897 18037 11931 18071
rect 14841 18037 14875 18071
rect 16221 18037 16255 18071
rect 18061 18037 18095 18071
rect 21373 18037 21407 18071
rect 24961 18037 24995 18071
rect 28917 18037 28951 18071
rect 30573 18037 30607 18071
rect 31585 18037 31619 18071
rect 31769 18037 31803 18071
rect 32689 18037 32723 18071
rect 38117 18037 38151 18071
rect 40877 18037 40911 18071
rect 41981 18037 42015 18071
rect 43269 18037 43303 18071
rect 45477 18037 45511 18071
rect 47041 18037 47075 18071
rect 3525 17833 3559 17867
rect 6377 17833 6411 17867
rect 8585 17833 8619 17867
rect 20526 17833 20560 17867
rect 22477 17833 22511 17867
rect 27629 17833 27663 17867
rect 33609 17833 33643 17867
rect 34897 17833 34931 17867
rect 36001 17833 36035 17867
rect 36724 17833 36758 17867
rect 44281 17833 44315 17867
rect 48053 17833 48087 17867
rect 33057 17765 33091 17799
rect 36185 17765 36219 17799
rect 41797 17765 41831 17799
rect 2053 17697 2087 17731
rect 3985 17697 4019 17731
rect 5273 17697 5307 17731
rect 7481 17697 7515 17731
rect 11161 17697 11195 17731
rect 13737 17697 13771 17731
rect 17877 17697 17911 17731
rect 18797 17697 18831 17731
rect 23029 17697 23063 17731
rect 24593 17697 24627 17731
rect 25697 17697 25731 17731
rect 28089 17697 28123 17731
rect 29009 17697 29043 17731
rect 30297 17697 30331 17731
rect 31309 17697 31343 17731
rect 34069 17697 34103 17731
rect 34161 17697 34195 17731
rect 35357 17697 35391 17731
rect 35541 17697 35575 17731
rect 39313 17697 39347 17731
rect 40049 17697 40083 17731
rect 40325 17697 40359 17731
rect 44465 17697 44499 17731
rect 1777 17629 1811 17663
rect 3433 17629 3467 17663
rect 4629 17629 4663 17663
rect 5733 17629 5767 17663
rect 6837 17629 6871 17663
rect 7941 17629 7975 17663
rect 10057 17629 10091 17663
rect 14289 17629 14323 17663
rect 17785 17629 17819 17663
rect 19717 17629 19751 17663
rect 20269 17629 20303 17663
rect 25421 17629 25455 17663
rect 27813 17629 27847 17663
rect 28825 17629 28859 17663
rect 30941 17629 30975 17663
rect 36461 17629 36495 17663
rect 42257 17629 42291 17663
rect 43395 17629 43429 17663
rect 45201 17629 45235 17663
rect 46305 17629 46339 17663
rect 47409 17629 47443 17663
rect 48513 17629 48547 17663
rect 9413 17561 9447 17595
rect 11437 17561 11471 17595
rect 13553 17561 13587 17595
rect 14565 17561 14599 17595
rect 16589 17561 16623 17595
rect 18613 17561 18647 17595
rect 19533 17561 19567 17595
rect 22937 17561 22971 17595
rect 23765 17561 23799 17595
rect 28917 17561 28951 17595
rect 31585 17561 31619 17595
rect 39037 17561 39071 17595
rect 49433 17561 49467 17595
rect 8953 17493 8987 17527
rect 9505 17493 9539 17527
rect 10701 17493 10735 17527
rect 12909 17493 12943 17527
rect 16037 17493 16071 17527
rect 16681 17493 16715 17527
rect 17325 17493 17359 17527
rect 17693 17493 17727 17527
rect 22017 17493 22051 17527
rect 22845 17493 22879 17527
rect 23857 17493 23891 17527
rect 25053 17493 25087 17527
rect 27169 17493 27203 17527
rect 28457 17493 28491 17527
rect 29745 17493 29779 17527
rect 30113 17493 30147 17527
rect 30205 17493 30239 17527
rect 30849 17493 30883 17527
rect 33977 17493 34011 17527
rect 35265 17493 35299 17527
rect 38209 17493 38243 17527
rect 38669 17493 38703 17527
rect 39129 17493 39163 17527
rect 42901 17493 42935 17527
rect 44005 17493 44039 17527
rect 45845 17493 45879 17527
rect 46949 17493 46983 17527
rect 49157 17493 49191 17527
rect 3617 17289 3651 17323
rect 6009 17289 6043 17323
rect 6745 17289 6779 17323
rect 7757 17289 7791 17323
rect 12449 17289 12483 17323
rect 14013 17289 14047 17323
rect 15577 17289 15611 17323
rect 18889 17289 18923 17323
rect 25329 17289 25363 17323
rect 26617 17289 26651 17323
rect 31585 17289 31619 17323
rect 35265 17289 35299 17323
rect 38117 17289 38151 17323
rect 40877 17289 40911 17323
rect 46581 17289 46615 17323
rect 48421 17289 48455 17323
rect 4905 17221 4939 17255
rect 6469 17221 6503 17255
rect 9965 17221 9999 17255
rect 11529 17221 11563 17255
rect 19625 17221 19659 17255
rect 32873 17221 32907 17255
rect 35173 17221 35207 17255
rect 41337 17221 41371 17255
rect 48973 17221 49007 17255
rect 1777 17153 1811 17187
rect 3801 17153 3835 17187
rect 4261 17153 4295 17187
rect 5365 17153 5399 17187
rect 6561 17153 6595 17187
rect 7113 17153 7147 17187
rect 8217 17153 8251 17187
rect 9321 17153 9355 17187
rect 10793 17153 10827 17187
rect 12541 17153 12575 17187
rect 13369 17153 13403 17187
rect 14473 17153 14507 17187
rect 15945 17153 15979 17187
rect 17141 17153 17175 17187
rect 19349 17153 19383 17187
rect 22017 17153 22051 17187
rect 23121 17153 23155 17187
rect 25697 17153 25731 17187
rect 25789 17153 25823 17187
rect 27169 17153 27203 17187
rect 28273 17153 28307 17187
rect 30849 17153 30883 17187
rect 30941 17153 30975 17187
rect 32597 17153 32631 17187
rect 36369 17153 36403 17187
rect 37473 17153 37507 17187
rect 38577 17153 38611 17187
rect 41245 17153 41279 17187
rect 42165 17153 42199 17187
rect 42625 17153 42659 17187
rect 43729 17153 43763 17187
rect 44833 17153 44867 17187
rect 45937 17153 45971 17187
rect 47777 17153 47811 17187
rect 2053 17085 2087 17119
rect 10885 17085 10919 17119
rect 11069 17085 11103 17119
rect 12633 17085 12667 17119
rect 16037 17085 16071 17119
rect 16129 17085 16163 17119
rect 17417 17085 17451 17119
rect 21465 17085 21499 17119
rect 21649 17085 21683 17119
rect 23397 17085 23431 17119
rect 25881 17085 25915 17119
rect 26433 17085 26467 17119
rect 26709 17085 26743 17119
rect 28549 17085 28583 17119
rect 31033 17085 31067 17119
rect 31769 17085 31803 17119
rect 35449 17085 35483 17119
rect 36461 17085 36495 17119
rect 36645 17085 36679 17119
rect 37013 17085 37047 17119
rect 38853 17085 38887 17119
rect 41521 17085 41555 17119
rect 43269 17085 43303 17119
rect 46949 17085 46983 17119
rect 47041 17085 47075 17119
rect 3341 17017 3375 17051
rect 11805 17017 11839 17051
rect 44373 17017 44407 17051
rect 45477 17017 45511 17051
rect 49433 17017 49467 17051
rect 8861 16949 8895 16983
rect 10425 16949 10459 16983
rect 12081 16949 12115 16983
rect 15117 16949 15151 16983
rect 16865 16949 16899 16983
rect 21097 16949 21131 16983
rect 22661 16949 22695 16983
rect 24869 16949 24903 16983
rect 27813 16949 27847 16983
rect 30021 16949 30055 16983
rect 30481 16949 30515 16983
rect 31861 16949 31895 16983
rect 32229 16949 32263 16983
rect 34345 16949 34379 16983
rect 34805 16949 34839 16983
rect 36001 16949 36035 16983
rect 40325 16949 40359 16983
rect 41889 16949 41923 16983
rect 49065 16949 49099 16983
rect 13829 16745 13863 16779
rect 15393 16745 15427 16779
rect 17877 16745 17911 16779
rect 18981 16745 19015 16779
rect 20545 16745 20579 16779
rect 24593 16745 24627 16779
rect 25224 16745 25258 16779
rect 27169 16745 27203 16779
rect 29561 16745 29595 16779
rect 29745 16745 29779 16779
rect 37105 16745 37139 16779
rect 41889 16745 41923 16779
rect 42993 16745 43027 16779
rect 49433 16745 49467 16779
rect 3617 16677 3651 16711
rect 7573 16677 7607 16711
rect 8769 16677 8803 16711
rect 27077 16677 27111 16711
rect 32321 16677 32355 16711
rect 3433 16609 3467 16643
rect 8033 16609 8067 16643
rect 8125 16609 8159 16643
rect 11989 16609 12023 16643
rect 13093 16609 13127 16643
rect 13277 16609 13311 16643
rect 14841 16609 14875 16643
rect 18429 16609 18463 16643
rect 20085 16609 20119 16643
rect 20729 16609 20763 16643
rect 21005 16609 21039 16643
rect 23949 16609 23983 16643
rect 24961 16609 24995 16643
rect 27997 16609 28031 16643
rect 28181 16609 28215 16643
rect 30113 16609 30147 16643
rect 32781 16609 32815 16643
rect 32965 16609 32999 16643
rect 33977 16609 34011 16643
rect 34161 16609 34195 16643
rect 35173 16609 35207 16643
rect 37749 16609 37783 16643
rect 38945 16609 38979 16643
rect 39497 16609 39531 16643
rect 40509 16609 40543 16643
rect 40693 16609 40727 16643
rect 1777 16541 1811 16575
rect 4261 16541 4295 16575
rect 5365 16541 5399 16575
rect 6469 16541 6503 16575
rect 7113 16541 7147 16575
rect 9229 16541 9263 16575
rect 9873 16541 9907 16575
rect 10333 16541 10367 16575
rect 10977 16541 11011 16575
rect 14657 16541 14691 16575
rect 14749 16541 14783 16575
rect 15657 16541 15691 16575
rect 16313 16541 16347 16575
rect 16773 16541 16807 16575
rect 17417 16541 17451 16575
rect 19901 16541 19935 16575
rect 24409 16541 24443 16575
rect 27905 16541 27939 16575
rect 34897 16541 34931 16575
rect 41245 16541 41279 16575
rect 42349 16541 42383 16575
rect 43453 16541 43487 16575
rect 44741 16541 44775 16575
rect 45201 16541 45235 16575
rect 45845 16541 45879 16575
rect 46305 16541 46339 16575
rect 47409 16541 47443 16575
rect 48513 16541 48547 16575
rect 2513 16473 2547 16507
rect 13737 16473 13771 16507
rect 18337 16473 18371 16507
rect 21281 16473 21315 16507
rect 30389 16473 30423 16507
rect 37013 16473 37047 16507
rect 37473 16473 37507 16507
rect 40417 16473 40451 16507
rect 44557 16473 44591 16507
rect 3893 16405 3927 16439
rect 4905 16405 4939 16439
rect 6009 16405 6043 16439
rect 7941 16405 7975 16439
rect 11437 16405 11471 16439
rect 11805 16405 11839 16439
rect 11897 16405 11931 16439
rect 12633 16405 12667 16439
rect 13001 16405 13035 16439
rect 14289 16405 14323 16439
rect 18245 16405 18279 16439
rect 19441 16405 19475 16439
rect 19809 16405 19843 16439
rect 22753 16405 22787 16439
rect 23305 16405 23339 16439
rect 23673 16405 23707 16439
rect 23765 16405 23799 16439
rect 26709 16405 26743 16439
rect 27537 16405 27571 16439
rect 28549 16405 28583 16439
rect 28917 16405 28951 16439
rect 31861 16405 31895 16439
rect 32689 16405 32723 16439
rect 33517 16405 33551 16439
rect 33885 16405 33919 16439
rect 36645 16405 36679 16439
rect 37565 16405 37599 16439
rect 38301 16405 38335 16439
rect 38669 16405 38703 16439
rect 38761 16405 38795 16439
rect 39405 16405 39439 16439
rect 40049 16405 40083 16439
rect 44097 16405 44131 16439
rect 44465 16405 44499 16439
rect 46949 16405 46983 16439
rect 48053 16405 48087 16439
rect 49157 16405 49191 16439
rect 6009 16201 6043 16235
rect 11989 16201 12023 16235
rect 12449 16201 12483 16235
rect 13185 16201 13219 16235
rect 13553 16201 13587 16235
rect 14841 16201 14875 16235
rect 15945 16201 15979 16235
rect 16037 16201 16071 16235
rect 24777 16201 24811 16235
rect 27629 16201 27663 16235
rect 29929 16201 29963 16235
rect 31217 16201 31251 16235
rect 31953 16201 31987 16235
rect 32321 16201 32355 16235
rect 32781 16201 32815 16235
rect 33517 16201 33551 16235
rect 41245 16201 41279 16235
rect 42257 16201 42291 16235
rect 44373 16201 44407 16235
rect 47777 16201 47811 16235
rect 48789 16201 48823 16235
rect 49525 16201 49559 16235
rect 3801 16133 3835 16167
rect 7297 16133 7331 16167
rect 12357 16133 12391 16167
rect 16865 16133 16899 16167
rect 17693 16133 17727 16167
rect 19441 16133 19475 16167
rect 35265 16133 35299 16167
rect 38577 16133 38611 16167
rect 49341 16133 49375 16167
rect 1777 16065 1811 16099
rect 3617 16065 3651 16099
rect 4261 16065 4295 16099
rect 5365 16065 5399 16099
rect 6653 16065 6687 16099
rect 8125 16065 8159 16099
rect 9413 16065 9447 16099
rect 10517 16065 10551 16099
rect 13645 16065 13679 16099
rect 14749 16065 14783 16099
rect 16773 16065 16807 16099
rect 17601 16065 17635 16099
rect 18521 16065 18555 16099
rect 18705 16065 18739 16099
rect 19165 16065 19199 16099
rect 21373 16065 21407 16099
rect 22385 16065 22419 16099
rect 23581 16065 23615 16099
rect 24869 16065 24903 16099
rect 25973 16065 26007 16099
rect 26065 16065 26099 16099
rect 26709 16065 26743 16099
rect 27537 16065 27571 16099
rect 28365 16065 28399 16099
rect 32689 16065 32723 16099
rect 33885 16065 33919 16099
rect 34989 16065 35023 16099
rect 37657 16065 37691 16099
rect 38301 16065 38335 16099
rect 40417 16065 40451 16099
rect 41153 16065 41187 16099
rect 42625 16065 42659 16099
rect 43729 16065 43763 16099
rect 44833 16065 44867 16099
rect 45937 16065 45971 16099
rect 47593 16065 47627 16099
rect 48145 16065 48179 16099
rect 2053 15997 2087 16031
rect 8217 15997 8251 16031
rect 8401 15997 8435 16031
rect 12633 15997 12667 16031
rect 13737 15997 13771 16031
rect 14933 15997 14967 16031
rect 16129 15997 16163 16031
rect 17785 15997 17819 16031
rect 22477 15997 22511 16031
rect 22569 15997 22603 16031
rect 23673 15997 23707 16031
rect 23765 15997 23799 16031
rect 25053 15997 25087 16031
rect 26157 15997 26191 16031
rect 27721 15997 27755 16031
rect 29009 15997 29043 16031
rect 30021 15997 30055 16031
rect 30205 15997 30239 16031
rect 31309 15997 31343 16031
rect 31401 15997 31435 16031
rect 32965 15997 32999 16031
rect 33977 15997 34011 16031
rect 34069 15997 34103 16031
rect 41337 15997 41371 16031
rect 41889 15997 41923 16031
rect 47041 15997 47075 16031
rect 7757 15929 7791 15963
rect 11161 15929 11195 15963
rect 22017 15929 22051 15963
rect 23213 15929 23247 15963
rect 29561 15929 29595 15963
rect 36737 15929 36771 15963
rect 40785 15929 40819 15963
rect 4905 15861 4939 15895
rect 8861 15861 8895 15895
rect 9045 15861 9079 15895
rect 10057 15861 10091 15895
rect 11713 15861 11747 15895
rect 14381 15861 14415 15895
rect 15577 15861 15611 15895
rect 17233 15861 17267 15895
rect 20913 15861 20947 15895
rect 21557 15861 21591 15895
rect 24409 15861 24443 15895
rect 25605 15861 25639 15895
rect 27169 15861 27203 15895
rect 30849 15861 30883 15895
rect 34621 15861 34655 15895
rect 37749 15861 37783 15895
rect 40049 15861 40083 15895
rect 42073 15861 42107 15895
rect 43269 15861 43303 15895
rect 45477 15861 45511 15895
rect 46581 15861 46615 15895
rect 49065 15861 49099 15895
rect 3617 15657 3651 15691
rect 3985 15657 4019 15691
rect 5273 15657 5307 15691
rect 7481 15657 7515 15691
rect 12357 15657 12391 15691
rect 16773 15657 16807 15691
rect 19349 15657 19383 15691
rect 20913 15657 20947 15691
rect 24593 15657 24627 15691
rect 25513 15657 25547 15691
rect 26617 15657 26651 15691
rect 29285 15657 29319 15691
rect 31769 15657 31803 15691
rect 35173 15657 35207 15691
rect 37736 15657 37770 15691
rect 3433 15589 3467 15623
rect 8585 15589 8619 15623
rect 14289 15589 14323 15623
rect 27077 15589 27111 15623
rect 29745 15589 29779 15623
rect 39497 15589 39531 15623
rect 41797 15589 41831 15623
rect 42901 15589 42935 15623
rect 2053 15521 2087 15555
rect 9137 15521 9171 15555
rect 10149 15521 10183 15555
rect 12817 15521 12851 15555
rect 13001 15521 13035 15555
rect 14749 15521 14783 15555
rect 14933 15521 14967 15555
rect 15945 15521 15979 15555
rect 16037 15521 16071 15555
rect 17233 15521 17267 15555
rect 17325 15521 17359 15555
rect 18521 15521 18555 15555
rect 20453 15521 20487 15555
rect 21373 15521 21407 15555
rect 21465 15521 21499 15555
rect 23489 15521 23523 15555
rect 27629 15521 27663 15555
rect 30297 15521 30331 15555
rect 32413 15521 32447 15555
rect 33425 15521 33459 15555
rect 33609 15521 33643 15555
rect 34161 15521 34195 15555
rect 35817 15521 35851 15555
rect 40049 15521 40083 15555
rect 40325 15521 40359 15555
rect 45201 15521 45235 15555
rect 45477 15521 45511 15555
rect 1777 15453 1811 15487
rect 4169 15453 4203 15487
rect 4629 15453 4663 15487
rect 5733 15453 5767 15487
rect 6837 15453 6871 15487
rect 7941 15453 7975 15487
rect 18337 15453 18371 15487
rect 18981 15453 19015 15487
rect 19809 15453 19843 15487
rect 22293 15453 22327 15487
rect 23305 15453 23339 15487
rect 23397 15453 23431 15487
rect 24869 15453 24903 15487
rect 25973 15453 26007 15487
rect 28273 15453 28307 15487
rect 30113 15453 30147 15487
rect 30205 15453 30239 15487
rect 32137 15453 32171 15487
rect 32229 15453 32263 15487
rect 34713 15453 34747 15487
rect 36369 15453 36403 15487
rect 37473 15453 37507 15487
rect 42257 15453 42291 15487
rect 43361 15453 43395 15487
rect 44649 15453 44683 15487
rect 46673 15453 46707 15487
rect 47133 15453 47167 15487
rect 48237 15453 48271 15487
rect 6377 15385 6411 15419
rect 9505 15385 9539 15419
rect 10425 15385 10459 15419
rect 14657 15385 14691 15419
rect 21281 15385 21315 15419
rect 27445 15385 27479 15419
rect 27537 15385 27571 15419
rect 28917 15385 28951 15419
rect 49249 15385 49283 15419
rect 49433 15385 49467 15419
rect 9597 15317 9631 15351
rect 11897 15317 11931 15351
rect 12725 15317 12759 15351
rect 13553 15317 13587 15351
rect 15485 15317 15519 15351
rect 15853 15317 15887 15351
rect 17141 15317 17175 15351
rect 17969 15317 18003 15351
rect 18429 15317 18463 15351
rect 19533 15317 19567 15351
rect 21925 15317 21959 15351
rect 22937 15317 22971 15351
rect 23949 15317 23983 15351
rect 24225 15317 24259 15351
rect 30849 15317 30883 15351
rect 31125 15317 31159 15351
rect 32965 15317 32999 15351
rect 33333 15317 33367 15351
rect 35081 15317 35115 15351
rect 35541 15317 35575 15351
rect 35633 15317 35667 15351
rect 37013 15317 37047 15351
rect 39221 15317 39255 15351
rect 44005 15317 44039 15351
rect 44465 15317 44499 15351
rect 46489 15317 46523 15351
rect 47777 15317 47811 15351
rect 48881 15317 48915 15351
rect 3617 15113 3651 15147
rect 7573 15113 7607 15147
rect 9505 15113 9539 15147
rect 10425 15113 10459 15147
rect 10793 15113 10827 15147
rect 11897 15113 11931 15147
rect 16037 15113 16071 15147
rect 18245 15113 18279 15147
rect 19441 15113 19475 15147
rect 20269 15113 20303 15147
rect 21465 15113 21499 15147
rect 21649 15113 21683 15147
rect 23581 15113 23615 15147
rect 24133 15113 24167 15147
rect 25421 15113 25455 15147
rect 27169 15113 27203 15147
rect 27537 15113 27571 15147
rect 27629 15113 27663 15147
rect 28733 15113 28767 15147
rect 28825 15113 28859 15147
rect 29929 15113 29963 15147
rect 32321 15113 32355 15147
rect 33517 15113 33551 15147
rect 35265 15113 35299 15147
rect 35357 15113 35391 15147
rect 37657 15113 37691 15147
rect 40233 15113 40267 15147
rect 45845 15113 45879 15147
rect 47961 15113 47995 15147
rect 49249 15113 49283 15147
rect 3341 15045 3375 15079
rect 8677 15045 8711 15079
rect 9597 15045 9631 15079
rect 10885 15045 10919 15079
rect 12265 15045 12299 15079
rect 14565 15045 14599 15079
rect 17601 15045 17635 15079
rect 25789 15045 25823 15079
rect 32781 15045 32815 15079
rect 40601 15045 40635 15079
rect 44925 15045 44959 15079
rect 1777 14977 1811 15011
rect 3801 14977 3835 15011
rect 4261 14977 4295 15011
rect 5365 14977 5399 15011
rect 6929 14977 6963 15011
rect 8033 14977 8067 15011
rect 13461 14977 13495 15011
rect 13553 14977 13587 15011
rect 16405 14977 16439 15011
rect 16957 14977 16991 15011
rect 17141 14977 17175 15011
rect 18337 14977 18371 15011
rect 20637 14977 20671 15011
rect 22017 14977 22051 15011
rect 23305 14977 23339 15011
rect 23857 14977 23891 15011
rect 24501 14977 24535 15011
rect 31217 14977 31251 15011
rect 32689 14977 32723 15011
rect 33885 14977 33919 15011
rect 33977 14977 34011 15011
rect 36461 14977 36495 15011
rect 36553 14977 36587 15011
rect 38025 14977 38059 15011
rect 41429 14977 41463 15011
rect 42625 14977 42659 15011
rect 43269 14977 43303 15011
rect 43729 14977 43763 15011
rect 45201 14977 45235 15011
rect 46581 14977 46615 15011
rect 47777 14977 47811 15011
rect 48605 14977 48639 15011
rect 2053 14909 2087 14943
rect 6469 14909 6503 14943
rect 9781 14909 9815 14943
rect 10977 14909 11011 14943
rect 12357 14909 12391 14943
rect 12449 14909 12483 14943
rect 13737 14909 13771 14943
rect 14289 14909 14323 14943
rect 18429 14909 18463 14943
rect 19533 14909 19567 14943
rect 19625 14909 19659 14943
rect 20729 14909 20763 14943
rect 20821 14909 20855 14943
rect 22753 14909 22787 14943
rect 24593 14909 24627 14943
rect 24685 14909 24719 14943
rect 25881 14909 25915 14943
rect 26065 14909 26099 14943
rect 26433 14909 26467 14943
rect 26617 14909 26651 14943
rect 27813 14909 27847 14943
rect 28917 14909 28951 14943
rect 30021 14909 30055 14943
rect 30205 14909 30239 14943
rect 31309 14909 31343 14943
rect 31401 14909 31435 14943
rect 32965 14909 32999 14943
rect 34161 14909 34195 14943
rect 35541 14909 35575 14943
rect 36737 14909 36771 14943
rect 37381 14909 37415 14943
rect 38301 14909 38335 14943
rect 40693 14909 40727 14943
rect 40785 14909 40819 14943
rect 4905 14841 4939 14875
rect 17877 14841 17911 14875
rect 28365 14841 28399 14875
rect 30849 14841 30883 14875
rect 46397 14841 46431 14875
rect 47225 14841 47259 14875
rect 47317 14841 47351 14875
rect 6009 14773 6043 14807
rect 6653 14773 6687 14807
rect 9137 14773 9171 14807
rect 11529 14773 11563 14807
rect 13093 14773 13127 14807
rect 19073 14773 19107 14807
rect 23489 14773 23523 14807
rect 29561 14773 29595 14807
rect 31953 14773 31987 14807
rect 34529 14773 34563 14807
rect 34897 14773 34931 14807
rect 36093 14773 36127 14807
rect 37565 14773 37599 14807
rect 39773 14773 39807 14807
rect 42073 14773 42107 14807
rect 44373 14773 44407 14807
rect 44741 14773 44775 14807
rect 46121 14773 46155 14807
rect 3525 14569 3559 14603
rect 7481 14569 7515 14603
rect 8585 14569 8619 14603
rect 10057 14569 10091 14603
rect 13921 14569 13955 14603
rect 16773 14569 16807 14603
rect 18153 14569 18187 14603
rect 19625 14569 19659 14603
rect 23305 14569 23339 14603
rect 25513 14569 25547 14603
rect 27997 14569 28031 14603
rect 28273 14569 28307 14603
rect 28457 14569 28491 14603
rect 33149 14569 33183 14603
rect 35160 14569 35194 14603
rect 45845 14569 45879 14603
rect 46949 14569 46983 14603
rect 49341 14569 49375 14603
rect 3985 14501 4019 14535
rect 6377 14501 6411 14535
rect 24501 14501 24535 14535
rect 31493 14501 31527 14535
rect 38853 14501 38887 14535
rect 39313 14501 39347 14535
rect 44005 14501 44039 14535
rect 48053 14501 48087 14535
rect 2053 14433 2087 14467
rect 14841 14433 14875 14467
rect 16129 14433 16163 14467
rect 17693 14433 17727 14467
rect 18797 14433 18831 14467
rect 20177 14433 20211 14467
rect 22845 14433 22879 14467
rect 23949 14433 23983 14467
rect 26249 14433 26283 14467
rect 29101 14433 29135 14467
rect 29745 14433 29779 14467
rect 32413 14433 32447 14467
rect 32597 14433 32631 14467
rect 33701 14433 33735 14467
rect 34161 14433 34195 14467
rect 36645 14433 36679 14467
rect 37105 14433 37139 14467
rect 41797 14433 41831 14467
rect 44281 14433 44315 14467
rect 44465 14433 44499 14467
rect 48329 14433 48363 14467
rect 1777 14365 1811 14399
rect 3433 14365 3467 14399
rect 4169 14365 4203 14399
rect 4629 14365 4663 14399
rect 5733 14365 5767 14399
rect 6825 14365 6859 14399
rect 7941 14365 7975 14399
rect 9413 14365 9447 14399
rect 10517 14365 10551 14399
rect 11621 14365 11655 14399
rect 15853 14365 15887 14399
rect 17049 14365 17083 14399
rect 20821 14365 20855 14399
rect 23765 14365 23799 14399
rect 24869 14365 24903 14399
rect 25973 14365 26007 14399
rect 32321 14365 32355 14399
rect 33609 14365 33643 14399
rect 34897 14365 34931 14399
rect 39497 14365 39531 14399
rect 40049 14365 40083 14399
rect 41153 14365 41187 14399
rect 42257 14365 42291 14399
rect 43361 14365 43395 14399
rect 45201 14365 45235 14399
rect 46305 14365 46339 14399
rect 47409 14365 47443 14399
rect 48697 14365 48731 14399
rect 5273 14297 5307 14331
rect 11897 14297 11931 14331
rect 14749 14297 14783 14331
rect 18521 14297 18555 14331
rect 21097 14297 21131 14331
rect 23673 14297 23707 14331
rect 28825 14297 28859 14331
rect 30021 14297 30055 14331
rect 37381 14297 37415 14331
rect 40693 14297 40727 14331
rect 42901 14297 42935 14331
rect 9045 14229 9079 14263
rect 11161 14229 11195 14263
rect 13369 14229 13403 14263
rect 14289 14229 14323 14263
rect 14657 14229 14691 14263
rect 15485 14229 15519 14263
rect 15945 14229 15979 14263
rect 16589 14229 16623 14263
rect 18613 14229 18647 14263
rect 19349 14229 19383 14263
rect 19993 14229 20027 14263
rect 20085 14229 20119 14263
rect 27721 14229 27755 14263
rect 28917 14229 28951 14263
rect 31953 14229 31987 14263
rect 33517 14229 33551 14263
rect 34529 14229 34563 14263
rect 3617 14025 3651 14059
rect 4905 14025 4939 14059
rect 6009 14025 6043 14059
rect 6561 14025 6595 14059
rect 7849 14025 7883 14059
rect 10057 14025 10091 14059
rect 11161 14025 11195 14059
rect 12357 14025 12391 14059
rect 14473 14025 14507 14059
rect 15209 14025 15243 14059
rect 15669 14025 15703 14059
rect 16221 14025 16255 14059
rect 17233 14025 17267 14059
rect 17601 14025 17635 14059
rect 21465 14025 21499 14059
rect 22017 14025 22051 14059
rect 22477 14025 22511 14059
rect 23305 14025 23339 14059
rect 23765 14025 23799 14059
rect 26617 14025 26651 14059
rect 32781 14025 32815 14059
rect 34897 14025 34931 14059
rect 35357 14025 35391 14059
rect 37473 14025 37507 14059
rect 38669 14025 38703 14059
rect 41613 14025 41647 14059
rect 43269 14025 43303 14059
rect 44373 14025 44407 14059
rect 44649 14025 44683 14059
rect 46949 14025 46983 14059
rect 47225 14025 47259 14059
rect 47961 14025 47995 14059
rect 49341 14025 49375 14059
rect 13185 13957 13219 13991
rect 15577 13957 15611 13991
rect 17693 13957 17727 13991
rect 18337 13957 18371 13991
rect 28917 13957 28951 13991
rect 32321 13957 32355 13991
rect 36001 13957 36035 13991
rect 36829 13957 36863 13991
rect 44833 13957 44867 13991
rect 1777 13889 1811 13923
rect 3801 13889 3835 13923
rect 4261 13889 4295 13923
rect 5365 13889 5399 13923
rect 6745 13889 6779 13923
rect 7205 13889 7239 13923
rect 8309 13889 8343 13923
rect 8953 13889 8987 13923
rect 9413 13889 9447 13923
rect 10517 13889 10551 13923
rect 11713 13889 11747 13923
rect 13277 13889 13311 13923
rect 14381 13889 14415 13923
rect 16497 13889 16531 13923
rect 18613 13889 18647 13923
rect 19717 13889 19751 13923
rect 22385 13889 22419 13923
rect 23673 13889 23707 13923
rect 24409 13889 24443 13923
rect 24869 13889 24903 13923
rect 27169 13889 27203 13923
rect 29377 13889 29411 13923
rect 33149 13889 33183 13923
rect 35541 13889 35575 13923
rect 37841 13889 37875 13923
rect 39037 13889 39071 13923
rect 39865 13889 39899 13923
rect 40969 13889 41003 13923
rect 42625 13889 42659 13923
rect 43729 13889 43763 13923
rect 45201 13889 45235 13923
rect 46305 13889 46339 13923
rect 47777 13889 47811 13923
rect 48697 13889 48731 13923
rect 2053 13821 2087 13855
rect 3341 13821 3375 13855
rect 13461 13821 13495 13855
rect 14565 13821 14599 13855
rect 15761 13821 15795 13855
rect 16957 13821 16991 13855
rect 17785 13821 17819 13855
rect 22569 13821 22603 13855
rect 23857 13821 23891 13855
rect 31125 13821 31159 13855
rect 31585 13821 31619 13855
rect 37933 13821 37967 13855
rect 38117 13821 38151 13855
rect 39129 13821 39163 13855
rect 39313 13821 39347 13855
rect 40509 13821 40543 13855
rect 41981 13821 42015 13855
rect 42165 13821 42199 13855
rect 48329 13821 48363 13855
rect 12817 13685 12851 13719
rect 14013 13685 14047 13719
rect 16681 13685 16715 13719
rect 19257 13685 19291 13719
rect 19980 13685 20014 13719
rect 24593 13685 24627 13719
rect 25132 13685 25166 13719
rect 29640 13685 29674 13719
rect 33412 13685 33446 13719
rect 45845 13685 45879 13719
rect 3433 13481 3467 13515
rect 7481 13481 7515 13515
rect 8585 13481 8619 13515
rect 17877 13481 17911 13515
rect 18337 13481 18371 13515
rect 19441 13481 19475 13515
rect 19717 13481 19751 13515
rect 26341 13481 26375 13515
rect 30113 13481 30147 13515
rect 34897 13481 34931 13515
rect 38209 13481 38243 13515
rect 39681 13481 39715 13515
rect 40693 13481 40727 13515
rect 42901 13481 42935 13515
rect 45017 13481 45051 13515
rect 46397 13481 46431 13515
rect 9045 13413 9079 13447
rect 9965 13413 9999 13447
rect 13921 13413 13955 13447
rect 18521 13413 18555 13447
rect 29561 13413 29595 13447
rect 29929 13413 29963 13447
rect 30389 13413 30423 13447
rect 32505 13413 32539 13447
rect 35265 13413 35299 13447
rect 45201 13413 45235 13447
rect 47501 13413 47535 13447
rect 2789 13345 2823 13379
rect 3617 13345 3651 13379
rect 10425 13345 10459 13379
rect 13185 13345 13219 13379
rect 13369 13345 13403 13379
rect 16405 13345 16439 13379
rect 18705 13345 18739 13379
rect 18889 13345 18923 13379
rect 19073 13345 19107 13379
rect 20269 13345 20303 13379
rect 20913 13345 20947 13379
rect 22661 13345 22695 13379
rect 23029 13345 23063 13379
rect 23765 13345 23799 13379
rect 23949 13345 23983 13379
rect 24593 13345 24627 13379
rect 26893 13345 26927 13379
rect 30757 13345 30791 13379
rect 35817 13345 35851 13379
rect 36461 13345 36495 13379
rect 45385 13345 45419 13379
rect 1777 13277 1811 13311
rect 4629 13277 4663 13311
rect 5733 13277 5767 13311
rect 6837 13277 6871 13311
rect 7941 13277 7975 13311
rect 9321 13277 9355 13311
rect 13093 13277 13127 13311
rect 15485 13277 15519 13311
rect 16129 13277 16163 13311
rect 28917 13277 28951 13311
rect 33793 13277 33827 13311
rect 34713 13277 34747 13311
rect 35725 13277 35759 13311
rect 38669 13277 38703 13311
rect 40049 13277 40083 13311
rect 41153 13277 41187 13311
rect 42257 13277 42291 13311
rect 43361 13277 43395 13311
rect 45753 13277 45787 13311
rect 46857 13277 46891 13311
rect 47961 13277 47995 13311
rect 49157 13277 49191 13311
rect 3985 13209 4019 13243
rect 10701 13209 10735 13243
rect 14381 13209 14415 13243
rect 14749 13209 14783 13243
rect 20085 13209 20119 13243
rect 21189 13209 21223 13243
rect 24869 13209 24903 13243
rect 27169 13209 27203 13243
rect 31033 13209 31067 13243
rect 33057 13209 33091 13243
rect 34437 13209 34471 13243
rect 35633 13209 35667 13243
rect 36737 13209 36771 13243
rect 44465 13209 44499 13243
rect 5273 13141 5307 13175
rect 6377 13141 6411 13175
rect 12173 13141 12207 13175
rect 12725 13141 12759 13175
rect 14197 13141 14231 13175
rect 20177 13141 20211 13175
rect 23305 13141 23339 13175
rect 23673 13141 23707 13175
rect 29193 13141 29227 13175
rect 29837 13141 29871 13175
rect 39313 13141 39347 13175
rect 41797 13141 41831 13175
rect 44005 13141 44039 13175
rect 3801 12937 3835 12971
rect 4905 12937 4939 12971
rect 6009 12937 6043 12971
rect 6469 12937 6503 12971
rect 6837 12937 6871 12971
rect 8861 12937 8895 12971
rect 10885 12937 10919 12971
rect 12081 12937 12115 12971
rect 13461 12937 13495 12971
rect 14105 12937 14139 12971
rect 16313 12937 16347 12971
rect 17601 12937 17635 12971
rect 27813 12937 27847 12971
rect 31861 12937 31895 12971
rect 34069 12937 34103 12971
rect 40601 12937 40635 12971
rect 41705 12937 41739 12971
rect 43269 12937 43303 12971
rect 44925 12937 44959 12971
rect 45385 12937 45419 12971
rect 47593 12937 47627 12971
rect 2881 12869 2915 12903
rect 7757 12869 7791 12903
rect 14841 12869 14875 12903
rect 18705 12869 18739 12903
rect 22201 12869 22235 12903
rect 23305 12869 23339 12903
rect 24317 12869 24351 12903
rect 30573 12869 30607 12903
rect 35265 12869 35299 12903
rect 41981 12869 42015 12903
rect 42257 12869 42291 12903
rect 47225 12869 47259 12903
rect 1593 12801 1627 12835
rect 1869 12801 1903 12835
rect 3157 12801 3191 12835
rect 4261 12801 4295 12835
rect 5365 12801 5399 12835
rect 7113 12801 7147 12835
rect 8217 12801 8251 12835
rect 9321 12801 9355 12835
rect 10793 12801 10827 12835
rect 13369 12801 13403 12835
rect 14565 12801 14599 12835
rect 16681 12801 16715 12835
rect 17325 12801 17359 12835
rect 17969 12801 18003 12835
rect 19717 12801 19751 12835
rect 21097 12801 21131 12835
rect 23213 12801 23247 12835
rect 24041 12801 24075 12835
rect 26709 12801 26743 12835
rect 27169 12801 27203 12835
rect 32321 12801 32355 12835
rect 36645 12801 36679 12835
rect 37473 12801 37507 12835
rect 39957 12801 39991 12835
rect 41061 12801 41095 12835
rect 42625 12801 42659 12835
rect 43729 12801 43763 12835
rect 45293 12801 45327 12835
rect 46121 12801 46155 12835
rect 46581 12801 46615 12835
rect 47961 12801 47995 12835
rect 49157 12801 49191 12835
rect 10977 12733 11011 12767
rect 12173 12733 12207 12767
rect 12357 12733 12391 12767
rect 13553 12733 13587 12767
rect 19809 12733 19843 12767
rect 19993 12733 20027 12767
rect 21189 12733 21223 12767
rect 21373 12733 21407 12767
rect 21925 12733 21959 12767
rect 23397 12733 23431 12767
rect 26249 12733 26283 12767
rect 28365 12733 28399 12767
rect 28641 12733 28675 12767
rect 31309 12733 31343 12767
rect 32597 12733 32631 12767
rect 34529 12733 34563 12767
rect 36001 12733 36035 12767
rect 37749 12733 37783 12767
rect 39497 12733 39531 12767
rect 17141 12665 17175 12699
rect 19349 12665 19383 12699
rect 20453 12665 20487 12699
rect 22845 12665 22879 12699
rect 25789 12665 25823 12699
rect 44373 12665 44407 12699
rect 45937 12665 45971 12699
rect 9965 12597 9999 12631
rect 10425 12597 10459 12631
rect 11713 12597 11747 12631
rect 13001 12597 13035 12631
rect 14197 12597 14231 12631
rect 20729 12597 20763 12631
rect 30113 12597 30147 12631
rect 36829 12597 36863 12631
rect 44649 12597 44683 12631
rect 2329 12393 2363 12427
rect 2789 12393 2823 12427
rect 6377 12393 6411 12427
rect 7481 12393 7515 12427
rect 9873 12393 9907 12427
rect 13001 12393 13035 12427
rect 19625 12393 19659 12427
rect 30205 12393 30239 12427
rect 30928 12393 30962 12427
rect 40693 12393 40727 12427
rect 44465 12393 44499 12427
rect 3985 12325 4019 12359
rect 12725 12325 12759 12359
rect 16037 12325 16071 12359
rect 23673 12325 23707 12359
rect 3433 12257 3467 12291
rect 10333 12257 10367 12291
rect 13553 12257 13587 12291
rect 18521 12257 18555 12291
rect 20177 12257 20211 12291
rect 24133 12257 24167 12291
rect 24869 12257 24903 12291
rect 27445 12257 27479 12291
rect 27997 12257 28031 12291
rect 29101 12257 29135 12291
rect 33425 12257 33459 12291
rect 36645 12257 36679 12291
rect 37749 12257 37783 12291
rect 38761 12257 38795 12291
rect 38945 12257 38979 12291
rect 45477 12257 45511 12291
rect 46765 12257 46799 12291
rect 49157 12257 49191 12291
rect 1685 12189 1719 12223
rect 3249 12189 3283 12223
rect 4169 12189 4203 12223
rect 4629 12189 4663 12223
rect 5733 12189 5767 12223
rect 6837 12189 6871 12223
rect 7941 12189 7975 12223
rect 9229 12189 9263 12223
rect 12541 12189 12575 12223
rect 14289 12189 14323 12223
rect 16589 12189 16623 12223
rect 19349 12189 19383 12223
rect 20913 12189 20947 12223
rect 22293 12189 22327 12223
rect 23857 12189 23891 12223
rect 24593 12189 24627 12223
rect 30665 12189 30699 12223
rect 34897 12189 34931 12223
rect 37473 12189 37507 12223
rect 39405 12189 39439 12223
rect 40049 12189 40083 12223
rect 41153 12189 41187 12223
rect 42257 12189 42291 12223
rect 43361 12189 43395 12223
rect 44649 12189 44683 12223
rect 45201 12189 45235 12223
rect 46489 12189 46523 12223
rect 47961 12189 47995 12223
rect 10609 12121 10643 12155
rect 13369 12121 13403 12155
rect 14565 12121 14599 12155
rect 17325 12121 17359 12155
rect 18337 12121 18371 12155
rect 19993 12121 20027 12155
rect 21649 12121 21683 12155
rect 23121 12121 23155 12155
rect 28917 12121 28951 12155
rect 29745 12121 29779 12155
rect 33333 12121 33367 12155
rect 35173 12121 35207 12155
rect 42901 12121 42935 12155
rect 5273 12053 5307 12087
rect 8585 12053 8619 12087
rect 12081 12053 12115 12087
rect 13461 12053 13495 12087
rect 17969 12053 18003 12087
rect 18429 12053 18463 12087
rect 18981 12053 19015 12087
rect 20085 12053 20119 12087
rect 26341 12053 26375 12087
rect 26801 12053 26835 12087
rect 27169 12053 27203 12087
rect 27261 12053 27295 12087
rect 27905 12053 27939 12087
rect 28457 12053 28491 12087
rect 28825 12053 28859 12087
rect 32413 12053 32447 12087
rect 32873 12053 32907 12087
rect 33241 12053 33275 12087
rect 33977 12053 34011 12087
rect 34161 12053 34195 12087
rect 34437 12053 34471 12087
rect 37105 12053 37139 12087
rect 37565 12053 37599 12087
rect 38301 12053 38335 12087
rect 38669 12053 38703 12087
rect 39497 12053 39531 12087
rect 41797 12053 41831 12087
rect 44005 12053 44039 12087
rect 47593 12053 47627 12087
rect 1777 11849 1811 11883
rect 2605 11849 2639 11883
rect 4905 11849 4939 11883
rect 5457 11849 5491 11883
rect 14105 11849 14139 11883
rect 15945 11849 15979 11883
rect 19441 11849 19475 11883
rect 19809 11849 19843 11883
rect 24593 11849 24627 11883
rect 25421 11849 25455 11883
rect 25789 11849 25823 11883
rect 30113 11849 30147 11883
rect 31953 11849 31987 11883
rect 36277 11849 36311 11883
rect 37013 11849 37047 11883
rect 39221 11849 39255 11883
rect 40325 11849 40359 11883
rect 41429 11849 41463 11883
rect 41889 11849 41923 11883
rect 44373 11849 44407 11883
rect 45109 11849 45143 11883
rect 47133 11849 47167 11883
rect 2513 11781 2547 11815
rect 3249 11781 3283 11815
rect 3433 11781 3467 11815
rect 8953 11781 8987 11815
rect 11161 11781 11195 11815
rect 11989 11781 12023 11815
rect 13737 11781 13771 11815
rect 17049 11781 17083 11815
rect 20085 11781 20119 11815
rect 24685 11781 24719 11815
rect 26709 11781 26743 11815
rect 28641 11781 28675 11815
rect 30665 11781 30699 11815
rect 36829 11781 36863 11815
rect 37749 11781 37783 11815
rect 47593 11781 47627 11815
rect 49157 11781 49191 11815
rect 1593 11713 1627 11747
rect 4261 11713 4295 11747
rect 5825 11713 5859 11747
rect 6469 11713 6503 11747
rect 6745 11713 6779 11747
rect 7205 11713 7239 11747
rect 8309 11713 8343 11747
rect 9413 11713 9447 11747
rect 10517 11713 10551 11747
rect 14749 11713 14783 11747
rect 14841 11713 14875 11747
rect 21097 11713 21131 11747
rect 27537 11713 27571 11747
rect 31401 11713 31435 11747
rect 32689 11713 32723 11747
rect 36185 11713 36219 11747
rect 39681 11713 39715 11747
rect 40785 11713 40819 11747
rect 42073 11713 42107 11747
rect 42717 11713 42751 11747
rect 42901 11713 42935 11747
rect 43453 11713 43487 11747
rect 44189 11713 44223 11747
rect 44925 11713 44959 11747
rect 45937 11713 45971 11747
rect 46949 11713 46983 11747
rect 47961 11713 47995 11747
rect 6009 11645 6043 11679
rect 7849 11645 7883 11679
rect 11713 11645 11747 11679
rect 15025 11645 15059 11679
rect 16037 11645 16071 11679
rect 16221 11645 16255 11679
rect 17693 11645 17727 11679
rect 17969 11645 18003 11679
rect 21189 11645 21223 11679
rect 21373 11645 21407 11679
rect 22017 11645 22051 11679
rect 22293 11645 22327 11679
rect 24777 11645 24811 11679
rect 25881 11645 25915 11679
rect 25973 11645 26007 11679
rect 27629 11645 27663 11679
rect 27813 11645 27847 11679
rect 28365 11645 28399 11679
rect 32781 11645 32815 11679
rect 32873 11645 32907 11679
rect 33517 11645 33551 11679
rect 33793 11645 33827 11679
rect 35265 11645 35299 11679
rect 36461 11645 36495 11679
rect 37473 11645 37507 11679
rect 45661 11645 45695 11679
rect 3801 11577 3835 11611
rect 5273 11577 5307 11611
rect 14381 11577 14415 11611
rect 20729 11577 20763 11611
rect 24225 11577 24259 11611
rect 3893 11509 3927 11543
rect 6561 11509 6595 11543
rect 10057 11509 10091 11543
rect 15577 11509 15611 11543
rect 16773 11509 16807 11543
rect 23765 11509 23799 11543
rect 26525 11509 26559 11543
rect 27169 11509 27203 11543
rect 32321 11509 32355 11543
rect 35817 11509 35851 11543
rect 43637 11509 43671 11543
rect 1777 11305 1811 11339
rect 3341 11305 3375 11339
rect 3801 11305 3835 11339
rect 4445 11305 4479 11339
rect 5181 11305 5215 11339
rect 5733 11305 5767 11339
rect 6285 11305 6319 11339
rect 8953 11305 8987 11339
rect 9321 11305 9355 11339
rect 10333 11305 10367 11339
rect 14289 11305 14323 11339
rect 18153 11305 18187 11339
rect 19901 11305 19935 11339
rect 20085 11305 20119 11339
rect 20453 11305 20487 11339
rect 26341 11305 26375 11339
rect 27156 11305 27190 11339
rect 30389 11305 30423 11339
rect 35081 11305 35115 11339
rect 35265 11305 35299 11339
rect 35541 11305 35575 11339
rect 39129 11305 39163 11339
rect 39497 11305 39531 11339
rect 42993 11305 43027 11339
rect 44833 11305 44867 11339
rect 46765 11305 46799 11339
rect 47409 11305 47443 11339
rect 2697 11237 2731 11271
rect 5641 11237 5675 11271
rect 13001 11237 13035 11271
rect 16957 11237 16991 11271
rect 23397 11237 23431 11271
rect 28641 11237 28675 11271
rect 33057 11237 33091 11271
rect 45017 11237 45051 11271
rect 8585 11169 8619 11203
rect 9137 11169 9171 11203
rect 12541 11169 12575 11203
rect 13461 11169 13495 11203
rect 13645 11169 13679 11203
rect 15025 11169 15059 11203
rect 15117 11169 15151 11203
rect 16313 11169 16347 11203
rect 17601 11169 17635 11203
rect 18613 11169 18647 11203
rect 18705 11169 18739 11203
rect 21097 11169 21131 11203
rect 24593 11169 24627 11203
rect 26893 11169 26927 11203
rect 33517 11169 33551 11203
rect 33609 11169 33643 11203
rect 35633 11169 35667 11203
rect 36001 11169 36035 11203
rect 36277 11169 36311 11203
rect 41797 11169 41831 11203
rect 43913 11169 43947 11203
rect 45937 11169 45971 11203
rect 49157 11169 49191 11203
rect 1593 11101 1627 11135
rect 2513 11101 2547 11135
rect 4353 11101 4387 11135
rect 5089 11101 5123 11135
rect 6193 11101 6227 11135
rect 6837 11101 6871 11135
rect 7941 11101 7975 11135
rect 9689 11101 9723 11135
rect 10793 11101 10827 11135
rect 13369 11101 13403 11135
rect 14933 11101 14967 11135
rect 19625 11101 19659 11135
rect 21649 11101 21683 11135
rect 29745 11101 29779 11135
rect 30849 11101 30883 11135
rect 33425 11101 33459 11135
rect 34161 11101 34195 11135
rect 38485 11101 38519 11135
rect 39681 11101 39715 11135
rect 40049 11101 40083 11135
rect 40693 11101 40727 11135
rect 41153 11101 41187 11135
rect 42349 11101 42383 11135
rect 43177 11101 43211 11135
rect 43637 11101 43671 11135
rect 45569 11101 45603 11135
rect 45661 11101 45695 11135
rect 47225 11101 47259 11135
rect 47961 11101 47995 11135
rect 3249 11033 3283 11067
rect 7481 11033 7515 11067
rect 11069 11033 11103 11067
rect 16129 11033 16163 11067
rect 17325 11033 17359 11067
rect 20821 11033 20855 11067
rect 20913 11033 20947 11067
rect 21925 11033 21959 11067
rect 23857 11033 23891 11067
rect 24869 11033 24903 11067
rect 31125 11033 31159 11067
rect 38025 11033 38059 11067
rect 42533 11033 42567 11067
rect 45201 11033 45235 11067
rect 14565 10965 14599 10999
rect 15761 10965 15795 10999
rect 16221 10965 16255 10999
rect 17417 10965 17451 10999
rect 18521 10965 18555 10999
rect 19441 10965 19475 10999
rect 32597 10965 32631 10999
rect 2881 10761 2915 10795
rect 3157 10761 3191 10795
rect 5641 10761 5675 10795
rect 7757 10761 7791 10795
rect 8953 10761 8987 10795
rect 11621 10761 11655 10795
rect 12357 10761 12391 10795
rect 18153 10761 18187 10795
rect 19441 10761 19475 10795
rect 22109 10761 22143 10795
rect 26525 10761 26559 10795
rect 28273 10761 28307 10795
rect 29285 10761 29319 10795
rect 32965 10761 32999 10795
rect 35541 10761 35575 10795
rect 36461 10761 36495 10795
rect 37105 10761 37139 10795
rect 42073 10761 42107 10795
rect 46949 10761 46983 10795
rect 47685 10761 47719 10795
rect 6101 10693 6135 10727
rect 7113 10693 7147 10727
rect 16313 10693 16347 10727
rect 22477 10693 22511 10727
rect 33057 10693 33091 10727
rect 47409 10693 47443 10727
rect 49157 10693 49191 10727
rect 1593 10625 1627 10659
rect 2329 10625 2363 10659
rect 3709 10625 3743 10659
rect 4445 10625 4479 10659
rect 5549 10625 5583 10659
rect 6929 10625 6963 10659
rect 7665 10625 7699 10659
rect 8309 10625 8343 10659
rect 9413 10625 9447 10659
rect 10517 10625 10551 10659
rect 12449 10625 12483 10659
rect 13185 10625 13219 10659
rect 15669 10625 15703 10659
rect 17325 10625 17359 10659
rect 17417 10625 17451 10659
rect 18521 10625 18555 10659
rect 24225 10625 24259 10659
rect 27629 10625 27663 10659
rect 28641 10625 28675 10659
rect 36369 10625 36403 10659
rect 37841 10625 37875 10659
rect 37933 10625 37967 10659
rect 38669 10625 38703 10659
rect 39773 10625 39807 10659
rect 40877 10625 40911 10659
rect 42809 10625 42843 10659
rect 43545 10625 43579 10659
rect 44557 10625 44591 10659
rect 45845 10625 45879 10659
rect 46121 10625 46155 10659
rect 47961 10625 47995 10659
rect 4169 10557 4203 10591
rect 6561 10557 6595 10591
rect 12541 10557 12575 10591
rect 13461 10557 13495 10591
rect 15209 10557 15243 10591
rect 17601 10557 17635 10591
rect 18613 10557 18647 10591
rect 18705 10557 18739 10591
rect 19717 10557 19751 10591
rect 19993 10557 20027 10591
rect 21465 10557 21499 10591
rect 22569 10557 22603 10591
rect 22753 10557 22787 10591
rect 23305 10557 23339 10591
rect 24501 10557 24535 10591
rect 26249 10557 26283 10591
rect 26801 10557 26835 10591
rect 27721 10557 27755 10591
rect 27905 10557 27939 10591
rect 29929 10557 29963 10591
rect 30205 10557 30239 10591
rect 33149 10557 33183 10591
rect 33793 10557 33827 10591
rect 34069 10557 34103 10591
rect 36645 10557 36679 10591
rect 38025 10557 38059 10591
rect 41797 10557 41831 10591
rect 42165 10557 42199 10591
rect 43269 10557 43303 10591
rect 44833 10557 44867 10591
rect 47225 10557 47259 10591
rect 1777 10489 1811 10523
rect 2513 10489 2547 10523
rect 11161 10489 11195 10523
rect 27261 10489 27295 10523
rect 31677 10489 31711 10523
rect 37473 10489 37507 10523
rect 41521 10489 41555 10523
rect 3525 10421 3559 10455
rect 10057 10421 10091 10455
rect 11989 10421 12023 10455
rect 16957 10421 16991 10455
rect 19165 10421 19199 10455
rect 23949 10421 23983 10455
rect 25973 10421 26007 10455
rect 29561 10421 29595 10455
rect 32597 10421 32631 10455
rect 36001 10421 36035 10455
rect 39313 10421 39347 10455
rect 40417 10421 40451 10455
rect 42625 10421 42659 10455
rect 3341 10217 3375 10251
rect 3617 10217 3651 10251
rect 5181 10217 5215 10251
rect 5917 10217 5951 10251
rect 7389 10217 7423 10251
rect 9137 10217 9171 10251
rect 10241 10217 10275 10251
rect 11345 10217 11379 10251
rect 16497 10217 16531 10251
rect 16957 10217 16991 10251
rect 22937 10217 22971 10251
rect 24041 10217 24075 10251
rect 25605 10217 25639 10251
rect 26065 10217 26099 10251
rect 28549 10217 28583 10251
rect 36921 10217 36955 10251
rect 37473 10217 37507 10251
rect 40693 10217 40727 10251
rect 43729 10217 43763 10251
rect 45109 10217 45143 10251
rect 45569 10217 45603 10251
rect 6745 10149 6779 10183
rect 9229 10149 9263 10183
rect 13001 10149 13035 10183
rect 16037 10149 16071 10183
rect 21741 10149 21775 10183
rect 24593 10149 24627 10183
rect 32597 10149 32631 10183
rect 41429 10149 41463 10183
rect 1869 10081 1903 10115
rect 4261 10081 4295 10115
rect 12265 10081 12299 10115
rect 12357 10081 12391 10115
rect 13461 10081 13495 10115
rect 13645 10081 13679 10115
rect 14289 10081 14323 10115
rect 17417 10081 17451 10115
rect 17601 10081 17635 10115
rect 18613 10081 18647 10115
rect 18797 10081 18831 10115
rect 19441 10081 19475 10115
rect 21189 10081 21223 10115
rect 22385 10081 22419 10115
rect 23397 10081 23431 10115
rect 23489 10081 23523 10115
rect 25237 10081 25271 10115
rect 25881 10081 25915 10115
rect 26801 10081 26835 10115
rect 30205 10081 30239 10115
rect 30389 10081 30423 10115
rect 31769 10081 31803 10115
rect 33149 10081 33183 10115
rect 34897 10081 34931 10115
rect 35173 10081 35207 10115
rect 37933 10081 37967 10115
rect 38025 10081 38059 10115
rect 39313 10081 39347 10115
rect 42901 10081 42935 10115
rect 46857 10081 46891 10115
rect 49157 10081 49191 10115
rect 1593 10013 1627 10047
rect 3985 10013 4019 10047
rect 7297 10013 7331 10047
rect 7941 10013 7975 10047
rect 9597 10013 9631 10047
rect 10701 10013 10735 10047
rect 12173 10013 12207 10047
rect 17325 10013 17359 10047
rect 22109 10013 22143 10047
rect 24961 10013 24995 10047
rect 25053 10013 25087 10047
rect 30113 10013 30147 10047
rect 32965 10013 32999 10047
rect 38669 10013 38703 10047
rect 40049 10013 40083 10047
rect 41981 10013 42015 10047
rect 42625 10013 42659 10047
rect 44465 10013 44499 10047
rect 45385 10013 45419 10047
rect 46121 10013 46155 10047
rect 47961 10013 47995 10047
rect 2697 9945 2731 9979
rect 5825 9945 5859 9979
rect 6561 9945 6595 9979
rect 8585 9945 8619 9979
rect 14565 9945 14599 9979
rect 19717 9945 19751 9979
rect 27077 9945 27111 9979
rect 31585 9945 31619 9979
rect 33057 9945 33091 9979
rect 37841 9945 37875 9979
rect 41245 9945 41279 9979
rect 43913 9945 43947 9979
rect 44649 9945 44683 9979
rect 2881 9877 2915 9911
rect 11805 9877 11839 9911
rect 13369 9877 13403 9911
rect 16589 9877 16623 9911
rect 18153 9877 18187 9911
rect 18521 9877 18555 9911
rect 22201 9877 22235 9911
rect 23305 9877 23339 9911
rect 29009 9877 29043 9911
rect 29745 9877 29779 9911
rect 31217 9877 31251 9911
rect 31677 9877 31711 9911
rect 36645 9877 36679 9911
rect 37105 9877 37139 9911
rect 39589 9877 39623 9911
rect 42073 9877 42107 9911
rect 2421 9673 2455 9707
rect 3433 9673 3467 9707
rect 4077 9673 4111 9707
rect 22017 9673 22051 9707
rect 23213 9673 23247 9707
rect 39221 9673 39255 9707
rect 4721 9605 4755 9639
rect 7941 9605 7975 9639
rect 8677 9605 8711 9639
rect 8769 9605 8803 9639
rect 13553 9605 13587 9639
rect 21557 9605 21591 9639
rect 30113 9605 30147 9639
rect 32597 9605 32631 9639
rect 34989 9605 35023 9639
rect 36461 9605 36495 9639
rect 46305 9605 46339 9639
rect 47317 9605 47351 9639
rect 47685 9605 47719 9639
rect 49157 9605 49191 9639
rect 1593 9537 1627 9571
rect 2329 9537 2363 9571
rect 2973 9537 3007 9571
rect 3617 9537 3651 9571
rect 4261 9537 4295 9571
rect 4537 9537 4571 9571
rect 5365 9537 5399 9571
rect 6009 9537 6043 9571
rect 6561 9537 6595 9571
rect 9413 9537 9447 9571
rect 10517 9537 10551 9571
rect 12173 9537 12207 9571
rect 13277 9537 13311 9571
rect 15853 9537 15887 9571
rect 16865 9537 16899 9571
rect 22385 9537 22419 9571
rect 22477 9537 22511 9571
rect 23489 9537 23523 9571
rect 26249 9537 26283 9571
rect 27905 9537 27939 9571
rect 30665 9537 30699 9571
rect 31401 9537 31435 9571
rect 32321 9537 32355 9571
rect 34897 9537 34931 9571
rect 36369 9537 36403 9571
rect 37473 9537 37507 9571
rect 38577 9537 38611 9571
rect 39773 9537 39807 9571
rect 40601 9537 40635 9571
rect 41521 9537 41555 9571
rect 42901 9537 42935 9571
rect 44189 9537 44223 9571
rect 45477 9537 45511 9571
rect 46765 9537 46799 9571
rect 47961 9537 47995 9571
rect 6837 9469 6871 9503
rect 10057 9469 10091 9503
rect 15945 9469 15979 9503
rect 16037 9469 16071 9503
rect 17141 9469 17175 9503
rect 18889 9469 18923 9503
rect 19349 9469 19383 9503
rect 19625 9469 19659 9503
rect 22569 9469 22603 9503
rect 23765 9469 23799 9503
rect 25513 9469 25547 9503
rect 26341 9469 26375 9503
rect 26525 9469 26559 9503
rect 27261 9469 27295 9503
rect 28181 9469 28215 9503
rect 31493 9469 31527 9503
rect 31677 9469 31711 9503
rect 35081 9469 35115 9503
rect 35541 9469 35575 9503
rect 36553 9469 36587 9503
rect 41245 9469 41279 9503
rect 42625 9469 42659 9503
rect 43913 9469 43947 9503
rect 45201 9469 45235 9503
rect 1777 9401 1811 9435
rect 2789 9401 2823 9435
rect 11161 9401 11195 9435
rect 11897 9401 11931 9435
rect 21465 9401 21499 9435
rect 34529 9401 34563 9435
rect 46949 9401 46983 9435
rect 5181 9333 5215 9367
rect 5825 9333 5859 9367
rect 8033 9333 8067 9367
rect 11713 9333 11747 9367
rect 12817 9333 12851 9367
rect 15025 9333 15059 9367
rect 15485 9333 15519 9367
rect 21097 9333 21131 9367
rect 25237 9333 25271 9367
rect 25881 9333 25915 9367
rect 29653 9333 29687 9367
rect 31033 9333 31067 9367
rect 34069 9333 34103 9367
rect 36001 9333 36035 9367
rect 37013 9333 37047 9367
rect 38117 9333 38151 9367
rect 39865 9333 39899 9367
rect 40693 9333 40727 9367
rect 3617 9129 3651 9163
rect 10333 9129 10367 9163
rect 11437 9129 11471 9163
rect 13001 9129 13035 9163
rect 18245 9129 18279 9163
rect 19349 9129 19383 9163
rect 23949 9129 23983 9163
rect 27721 9129 27755 9163
rect 28273 9129 28307 9163
rect 37013 9129 37047 9163
rect 38761 9129 38795 9163
rect 43821 9129 43855 9163
rect 45201 9129 45235 9163
rect 46673 9129 46707 9163
rect 47409 9129 47443 9163
rect 2513 9061 2547 9095
rect 18705 9061 18739 9095
rect 31493 9061 31527 9095
rect 33701 9061 33735 9095
rect 39589 9061 39623 9095
rect 6193 8993 6227 9027
rect 7757 8993 7791 9027
rect 13461 8993 13495 9027
rect 13645 8993 13679 9027
rect 15485 8993 15519 9027
rect 15577 8993 15611 9027
rect 16221 8993 16255 9027
rect 19533 8993 19567 9027
rect 19993 8993 20027 9027
rect 22201 8993 22235 9027
rect 25605 8993 25639 9027
rect 28733 8993 28767 9027
rect 28917 8993 28951 9027
rect 30021 8993 30055 9027
rect 31953 8993 31987 9027
rect 34161 8993 34195 9027
rect 35357 8993 35391 9027
rect 35449 8993 35483 9027
rect 38117 8993 38151 9027
rect 40785 8993 40819 9027
rect 42349 8993 42383 9027
rect 45569 8993 45603 9027
rect 49157 8993 49191 9027
rect 1593 8925 1627 8959
rect 2329 8925 2363 8959
rect 3249 8925 3283 8959
rect 3801 8925 3835 8959
rect 5917 8925 5951 8959
rect 8033 8925 8067 8959
rect 9689 8925 9723 8959
rect 10793 8925 10827 8959
rect 11897 8925 11931 8959
rect 14381 8925 14415 8959
rect 15393 8925 15427 8959
rect 18889 8925 18923 8959
rect 19717 8925 19751 8959
rect 24593 8925 24627 8959
rect 25973 8925 26007 8959
rect 27077 8925 27111 8959
rect 29745 8925 29779 8959
rect 35265 8925 35299 8959
rect 36093 8925 36127 8959
rect 36737 8925 36771 8959
rect 37473 8925 37507 8959
rect 41061 8925 41095 8959
rect 42073 8925 42107 8959
rect 43545 8925 43579 8959
rect 44373 8925 44407 8959
rect 45845 8925 45879 8959
rect 47225 8925 47259 8959
rect 47961 8925 47995 8959
rect 12541 8857 12575 8891
rect 16497 8857 16531 8891
rect 20269 8857 20303 8891
rect 22477 8857 22511 8891
rect 28641 8857 28675 8891
rect 32229 8857 32263 8891
rect 39129 8857 39163 8891
rect 39313 8857 39347 8891
rect 40141 8857 40175 8891
rect 40325 8857 40359 8891
rect 44557 8857 44591 8891
rect 1777 8789 1811 8823
rect 3065 8789 3099 8823
rect 5549 8789 5583 8823
rect 13369 8789 13403 8823
rect 15025 8789 15059 8823
rect 17969 8789 18003 8823
rect 21741 8789 21775 8823
rect 25237 8789 25271 8823
rect 26617 8789 26651 8823
rect 34897 8789 34931 8823
rect 38485 8789 38519 8823
rect 43361 8789 43395 8823
rect 45017 8789 45051 8823
rect 46949 8789 46983 8823
rect 3249 8585 3283 8619
rect 7481 8585 7515 8619
rect 13001 8585 13035 8619
rect 14105 8585 14139 8619
rect 14289 8585 14323 8619
rect 16957 8585 16991 8619
rect 18061 8585 18095 8619
rect 21189 8585 21223 8619
rect 25145 8585 25179 8619
rect 26617 8585 26651 8619
rect 30665 8585 30699 8619
rect 31033 8585 31067 8619
rect 32413 8585 32447 8619
rect 32781 8585 32815 8619
rect 33977 8585 34011 8619
rect 34069 8585 34103 8619
rect 34897 8585 34931 8619
rect 38117 8585 38151 8619
rect 38577 8585 38611 8619
rect 39037 8585 39071 8619
rect 41521 8585 41555 8619
rect 41797 8585 41831 8619
rect 42625 8585 42659 8619
rect 44649 8585 44683 8619
rect 3433 8517 3467 8551
rect 6101 8517 6135 8551
rect 15209 8517 15243 8551
rect 31493 8517 31527 8551
rect 35265 8517 35299 8551
rect 35357 8517 35391 8551
rect 42073 8517 42107 8551
rect 45201 8517 45235 8551
rect 45385 8517 45419 8551
rect 49157 8517 49191 8551
rect 1869 8449 1903 8483
rect 3157 8449 3191 8483
rect 7665 8449 7699 8483
rect 8309 8449 8343 8483
rect 9413 8449 9447 8483
rect 10517 8449 10551 8483
rect 11897 8449 11931 8483
rect 13369 8449 13403 8483
rect 14565 8449 14599 8483
rect 15669 8449 15703 8483
rect 17325 8449 17359 8483
rect 17417 8449 17451 8483
rect 18245 8449 18279 8483
rect 24041 8449 24075 8483
rect 24501 8449 24535 8483
rect 25973 8449 26007 8483
rect 27353 8449 27387 8483
rect 31401 8449 31435 8483
rect 36093 8449 36127 8483
rect 36737 8449 36771 8483
rect 37473 8449 37507 8483
rect 38761 8449 38795 8483
rect 39681 8449 39715 8483
rect 39957 8449 39991 8483
rect 41061 8449 41095 8483
rect 42809 8449 42843 8483
rect 44189 8449 44223 8483
rect 44373 8449 44407 8483
rect 45845 8449 45879 8483
rect 47961 8449 47995 8483
rect 1593 8381 1627 8415
rect 9137 8381 9171 8415
rect 11621 8381 11655 8415
rect 13461 8381 13495 8415
rect 13645 8381 13679 8415
rect 17601 8381 17635 8415
rect 18981 8381 19015 8415
rect 20729 8381 20763 8415
rect 22017 8381 22051 8415
rect 23765 8381 23799 8415
rect 28457 8381 28491 8415
rect 28733 8381 28767 8415
rect 31677 8381 31711 8415
rect 32873 8381 32907 8415
rect 33057 8381 33091 8415
rect 34253 8381 34287 8415
rect 35541 8381 35575 8415
rect 39313 8381 39347 8415
rect 41245 8381 41279 8415
rect 43085 8381 43119 8415
rect 43453 8381 43487 8415
rect 46857 8381 46891 8415
rect 2789 8313 2823 8347
rect 8125 8313 8159 8347
rect 11161 8313 11195 8347
rect 16313 8313 16347 8347
rect 30205 8313 30239 8347
rect 33609 8313 33643 8347
rect 41889 8313 41923 8347
rect 47593 8313 47627 8347
rect 2881 8245 2915 8279
rect 12541 8245 12575 8279
rect 18337 8245 18371 8279
rect 18613 8245 18647 8279
rect 19238 8245 19272 8279
rect 22280 8245 22314 8279
rect 27997 8245 28031 8279
rect 2145 8041 2179 8075
rect 8401 8041 8435 8075
rect 11345 8041 11379 8075
rect 13737 8041 13771 8075
rect 14565 8041 14599 8075
rect 15853 8041 15887 8075
rect 18981 8041 19015 8075
rect 21281 8041 21315 8075
rect 24041 8041 24075 8075
rect 24409 8041 24443 8075
rect 26801 8041 26835 8075
rect 28089 8041 28123 8075
rect 32965 8041 32999 8075
rect 34253 8041 34287 8075
rect 44741 8041 44775 8075
rect 45201 8041 45235 8075
rect 45569 8041 45603 8075
rect 1777 7973 1811 8007
rect 18061 7973 18095 8007
rect 22385 7973 22419 8007
rect 22753 7973 22787 8007
rect 29193 7973 29227 8007
rect 40601 7973 40635 8007
rect 40877 7973 40911 8007
rect 41061 7973 41095 8007
rect 41245 7973 41279 8007
rect 41705 7973 41739 8007
rect 41981 7973 42015 8007
rect 42165 7973 42199 8007
rect 44005 7973 44039 8007
rect 47501 7973 47535 8007
rect 10057 7905 10091 7939
rect 10701 7905 10735 7939
rect 12633 7905 12667 7939
rect 31861 7905 31895 7939
rect 39313 7905 39347 7939
rect 42349 7905 42383 7939
rect 44557 7905 44591 7939
rect 49157 7905 49191 7939
rect 1593 7837 1627 7871
rect 2329 7837 2363 7871
rect 8585 7837 8619 7871
rect 9321 7837 9355 7871
rect 9597 7837 9631 7871
rect 11529 7837 11563 7871
rect 11989 7837 12023 7871
rect 13093 7837 13127 7871
rect 14749 7837 14783 7871
rect 15209 7837 15243 7871
rect 16313 7837 16347 7871
rect 19533 7837 19567 7871
rect 20637 7837 20671 7871
rect 21741 7837 21775 7871
rect 23397 7837 23431 7871
rect 25053 7837 25087 7871
rect 25697 7837 25731 7871
rect 26157 7837 26191 7871
rect 27445 7837 27479 7871
rect 28549 7837 28583 7871
rect 29745 7837 29779 7871
rect 30849 7837 30883 7871
rect 32321 7837 32355 7871
rect 33333 7837 33367 7871
rect 33609 7837 33643 7871
rect 34897 7837 34931 7871
rect 37381 7837 37415 7871
rect 37933 7837 37967 7871
rect 38853 7837 38887 7871
rect 42901 7837 42935 7871
rect 43545 7837 43579 7871
rect 44189 7837 44223 7871
rect 45753 7837 45787 7871
rect 46213 7837 46247 7871
rect 46949 7837 46983 7871
rect 47961 7837 47995 7871
rect 16589 7769 16623 7803
rect 30389 7769 30423 7803
rect 35541 7769 35575 7803
rect 38669 7769 38703 7803
rect 40141 7769 40175 7803
rect 40325 7769 40359 7803
rect 9413 7701 9447 7735
rect 14197 7701 14231 7735
rect 18521 7701 18555 7735
rect 20177 7701 20211 7735
rect 22937 7701 22971 7735
rect 31493 7701 31527 7735
rect 37197 7701 37231 7735
rect 38025 7701 38059 7735
rect 41521 7701 41555 7735
rect 42717 7701 42751 7735
rect 43361 7701 43395 7735
rect 45017 7701 45051 7735
rect 46397 7701 46431 7735
rect 47133 7701 47167 7735
rect 9781 7497 9815 7531
rect 10333 7497 10367 7531
rect 10425 7497 10459 7531
rect 11345 7497 11379 7531
rect 11805 7497 11839 7531
rect 12449 7497 12483 7531
rect 14105 7497 14139 7531
rect 16313 7497 16347 7531
rect 16681 7497 16715 7531
rect 17325 7497 17359 7531
rect 18981 7497 19015 7531
rect 20361 7497 20395 7531
rect 28181 7497 28215 7531
rect 29377 7497 29411 7531
rect 31585 7497 31619 7531
rect 34253 7497 34287 7531
rect 34529 7497 34563 7531
rect 39773 7497 39807 7531
rect 45569 7497 45603 7531
rect 46397 7497 46431 7531
rect 16957 7429 16991 7463
rect 18889 7429 18923 7463
rect 33149 7429 33183 7463
rect 40233 7429 40267 7463
rect 44925 7429 44959 7463
rect 47225 7429 47259 7463
rect 49157 7429 49191 7463
rect 1593 7361 1627 7395
rect 2145 7361 2179 7395
rect 9137 7361 9171 7395
rect 9965 7361 9999 7395
rect 11161 7361 11195 7395
rect 11989 7361 12023 7395
rect 12633 7361 12667 7395
rect 13093 7361 13127 7395
rect 14565 7361 14599 7395
rect 15669 7361 15703 7395
rect 17693 7361 17727 7395
rect 19717 7361 19751 7395
rect 20821 7361 20855 7395
rect 22753 7361 22787 7395
rect 23857 7361 23891 7395
rect 24961 7361 24995 7395
rect 27537 7361 27571 7395
rect 28733 7361 28767 7395
rect 29837 7361 29871 7395
rect 30941 7361 30975 7395
rect 32505 7361 32539 7395
rect 33609 7361 33643 7395
rect 34897 7361 34931 7395
rect 38025 7361 38059 7395
rect 38485 7361 38519 7395
rect 39313 7361 39347 7395
rect 39957 7361 39991 7395
rect 43177 7361 43211 7395
rect 43729 7361 43763 7395
rect 44373 7361 44407 7395
rect 45753 7361 45787 7395
rect 46213 7361 46247 7395
rect 47041 7361 47075 7395
rect 47961 7361 47995 7395
rect 13737 7293 13771 7327
rect 15209 7293 15243 7327
rect 17785 7293 17819 7327
rect 17877 7293 17911 7327
rect 19073 7293 19107 7327
rect 30481 7293 30515 7327
rect 37749 7293 37783 7327
rect 38669 7293 38703 7327
rect 47593 7293 47627 7327
rect 9321 7225 9355 7259
rect 39129 7225 39163 7259
rect 43545 7225 43579 7259
rect 45109 7225 45143 7259
rect 1777 7157 1811 7191
rect 18521 7157 18555 7191
rect 21465 7157 21499 7191
rect 21833 7157 21867 7191
rect 23397 7157 23431 7191
rect 24501 7157 24535 7191
rect 25605 7157 25639 7191
rect 35541 7157 35575 7191
rect 42901 7157 42935 7191
rect 43085 7157 43119 7191
rect 44189 7157 44223 7191
rect 9505 6953 9539 6987
rect 12817 6953 12851 6987
rect 18613 6953 18647 6987
rect 17601 6885 17635 6919
rect 11069 6817 11103 6851
rect 13737 6817 13771 6851
rect 15945 6817 15979 6851
rect 17141 6817 17175 6851
rect 18153 6817 18187 6851
rect 19441 6817 19475 6851
rect 22017 6817 22051 6851
rect 24041 6817 24075 6851
rect 25881 6817 25915 6851
rect 28457 6817 28491 6851
rect 35541 6817 35575 6851
rect 43453 6817 43487 6851
rect 43821 6817 43855 6851
rect 44741 6817 44775 6851
rect 49157 6817 49191 6851
rect 1593 6749 1627 6783
rect 2513 6749 2547 6783
rect 2789 6749 2823 6783
rect 11345 6749 11379 6783
rect 14473 6745 14507 6779
rect 15301 6749 15335 6783
rect 16497 6749 16531 6783
rect 17969 6749 18003 6783
rect 18889 6749 18923 6783
rect 20269 6749 20303 6783
rect 21373 6749 21407 6783
rect 23397 6749 23431 6783
rect 25237 6749 25271 6783
rect 26341 6749 26375 6783
rect 27813 6749 27847 6783
rect 29745 6749 29779 6783
rect 30849 6749 30883 6783
rect 32321 6749 32355 6783
rect 33425 6749 33459 6783
rect 34897 6749 34931 6783
rect 43545 6749 43579 6783
rect 45661 6749 45695 6783
rect 46121 6749 46155 6783
rect 47961 6749 47995 6783
rect 13553 6681 13587 6715
rect 20913 6681 20947 6715
rect 32965 6681 32999 6715
rect 34069 6681 34103 6715
rect 44189 6681 44223 6715
rect 44373 6681 44407 6715
rect 47317 6681 47351 6715
rect 1777 6613 1811 6647
rect 2329 6613 2363 6647
rect 12357 6613 12391 6647
rect 14289 6613 14323 6647
rect 18061 6613 18095 6647
rect 18981 6613 19015 6647
rect 26985 6613 27019 6647
rect 30389 6613 30423 6647
rect 31493 6613 31527 6647
rect 45017 6613 45051 6647
rect 45477 6613 45511 6647
rect 2145 6409 2179 6443
rect 16313 6409 16347 6443
rect 18153 6409 18187 6443
rect 19257 6409 19291 6443
rect 20361 6409 20395 6443
rect 22661 6409 22695 6443
rect 24225 6409 24259 6443
rect 25329 6409 25363 6443
rect 29285 6409 29319 6443
rect 30481 6409 30515 6443
rect 31585 6409 31619 6443
rect 32965 6409 32999 6443
rect 33425 6409 33459 6443
rect 44005 6409 44039 6443
rect 44189 6409 44223 6443
rect 44373 6409 44407 6443
rect 44649 6409 44683 6443
rect 45109 6409 45143 6443
rect 46029 6409 46063 6443
rect 47225 6409 47259 6443
rect 47409 6409 47443 6443
rect 13553 6341 13587 6375
rect 38209 6341 38243 6375
rect 38669 6341 38703 6375
rect 49157 6341 49191 6375
rect 1593 6273 1627 6307
rect 2329 6273 2363 6307
rect 11805 6273 11839 6307
rect 14473 6273 14507 6307
rect 15209 6273 15243 6307
rect 15669 6273 15703 6307
rect 16865 6273 16899 6307
rect 17509 6273 17543 6307
rect 18613 6273 18647 6307
rect 19717 6273 19751 6307
rect 20821 6273 20855 6307
rect 21465 6273 21499 6307
rect 22017 6273 22051 6307
rect 23581 6273 23615 6307
rect 24685 6273 24719 6307
rect 28641 6273 28675 6307
rect 29837 6273 29871 6307
rect 30941 6273 30975 6307
rect 32321 6273 32355 6307
rect 44465 6273 44499 6307
rect 45569 6273 45603 6307
rect 46213 6273 46247 6307
rect 46857 6273 46891 6307
rect 47685 6273 47719 6307
rect 47961 6273 47995 6307
rect 12357 6205 12391 6239
rect 38393 6205 38427 6239
rect 1777 6137 1811 6171
rect 11989 6137 12023 6171
rect 14289 6137 14323 6171
rect 46673 6137 46707 6171
rect 15025 6069 15059 6103
rect 44925 6069 44959 6103
rect 45385 6069 45419 6103
rect 18889 5865 18923 5899
rect 21005 5865 21039 5899
rect 24041 5865 24075 5899
rect 30389 5865 30423 5899
rect 32965 5865 32999 5899
rect 44649 5865 44683 5899
rect 45201 5865 45235 5899
rect 45385 5865 45419 5899
rect 46029 5865 46063 5899
rect 46397 5865 46431 5899
rect 47041 5865 47075 5899
rect 47317 5865 47351 5899
rect 2513 5797 2547 5831
rect 44833 5797 44867 5831
rect 45753 5797 45787 5831
rect 3065 5729 3099 5763
rect 15853 5729 15887 5763
rect 16497 5729 16531 5763
rect 19441 5729 19475 5763
rect 25237 5729 25271 5763
rect 31677 5729 31711 5763
rect 49157 5729 49191 5763
rect 1593 5661 1627 5695
rect 2329 5661 2363 5695
rect 2881 5661 2915 5695
rect 17141 5661 17175 5695
rect 18245 5661 18279 5695
rect 20361 5661 20395 5695
rect 21684 5661 21718 5695
rect 22293 5661 22327 5695
rect 23397 5661 23431 5695
rect 24593 5661 24627 5695
rect 29745 5661 29779 5695
rect 32321 5661 32355 5695
rect 43729 5661 43763 5695
rect 46581 5661 46615 5695
rect 47501 5661 47535 5695
rect 47961 5661 47995 5695
rect 21787 5593 21821 5627
rect 43913 5593 43947 5627
rect 45937 5593 45971 5627
rect 1777 5525 1811 5559
rect 17785 5525 17819 5559
rect 22937 5525 22971 5559
rect 45569 5525 45603 5559
rect 20177 5321 20211 5355
rect 23581 5321 23615 5355
rect 32321 5321 32355 5355
rect 45569 5321 45603 5355
rect 47685 5321 47719 5355
rect 19073 5253 19107 5287
rect 39313 5253 39347 5287
rect 39773 5253 39807 5287
rect 49157 5253 49191 5287
rect 1869 5185 1903 5219
rect 16957 5185 16991 5219
rect 17969 5185 18003 5219
rect 18429 5185 18463 5219
rect 19533 5185 19567 5219
rect 20821 5185 20855 5219
rect 22328 5185 22362 5219
rect 22937 5185 22971 5219
rect 24076 5185 24110 5219
rect 24685 5185 24719 5219
rect 38117 5185 38151 5219
rect 38577 5185 38611 5219
rect 45845 5185 45879 5219
rect 47961 5185 47995 5219
rect 1593 5117 1627 5151
rect 17141 5117 17175 5151
rect 17509 5117 17543 5151
rect 22431 5117 22465 5151
rect 39497 5117 39531 5151
rect 46857 5117 46891 5151
rect 17785 5049 17819 5083
rect 38761 5049 38795 5083
rect 21465 4981 21499 5015
rect 24179 4981 24213 5015
rect 25329 4981 25363 5015
rect 2145 4777 2179 4811
rect 20177 4777 20211 4811
rect 24041 4777 24075 4811
rect 45845 4777 45879 4811
rect 46489 4777 46523 4811
rect 46765 4777 46799 4811
rect 47041 4777 47075 4811
rect 47593 4777 47627 4811
rect 18705 4709 18739 4743
rect 46121 4709 46155 4743
rect 21005 4641 21039 4675
rect 23029 4641 23063 4675
rect 25421 4641 25455 4675
rect 25697 4641 25731 4675
rect 49157 4641 49191 4675
rect 2329 4573 2363 4607
rect 18889 4573 18923 4607
rect 19533 4573 19567 4607
rect 23397 4573 23431 4607
rect 24628 4573 24662 4607
rect 25237 4573 25271 4607
rect 38117 4573 38151 4607
rect 38577 4573 38611 4607
rect 46305 4573 46339 4607
rect 47225 4573 47259 4607
rect 47961 4573 47995 4607
rect 1685 4505 1719 4539
rect 1869 4505 1903 4539
rect 21281 4505 21315 4539
rect 37381 4505 37415 4539
rect 38301 4505 38335 4539
rect 20729 4437 20763 4471
rect 22753 4437 22787 4471
rect 24731 4437 24765 4471
rect 36921 4437 36955 4471
rect 37473 4437 37507 4471
rect 21097 4233 21131 4267
rect 27353 4165 27387 4199
rect 37565 4165 37599 4199
rect 38025 4165 38059 4199
rect 1593 4097 1627 4131
rect 2329 4097 2363 4131
rect 3065 4097 3099 4131
rect 9689 4097 9723 4131
rect 18153 4097 18187 4131
rect 20453 4097 20487 4131
rect 22017 4097 22051 4131
rect 23121 4097 23155 4131
rect 37749 4097 37783 4131
rect 45845 4097 45879 4131
rect 47961 4097 47995 4131
rect 49157 4097 49191 4131
rect 18337 4029 18371 4063
rect 19993 4029 20027 4063
rect 22661 4029 22695 4063
rect 24133 4029 24167 4063
rect 24317 4029 24351 4063
rect 24961 4029 24995 4063
rect 27169 4029 27203 4063
rect 27629 4029 27663 4063
rect 46673 4029 46707 4063
rect 47685 4029 47719 4063
rect 1777 3961 1811 3995
rect 2513 3961 2547 3995
rect 2881 3893 2915 3927
rect 10333 3893 10367 3927
rect 23213 3893 23247 3927
rect 23581 3893 23615 3927
rect 20085 3689 20119 3723
rect 1869 3553 1903 3587
rect 24593 3553 24627 3587
rect 24869 3553 24903 3587
rect 49157 3553 49191 3587
rect 1593 3485 1627 3519
rect 9597 3485 9631 3519
rect 10057 3485 10091 3519
rect 11161 3485 11195 3519
rect 16221 3485 16255 3519
rect 17141 3485 17175 3519
rect 17601 3485 17635 3519
rect 18245 3485 18279 3519
rect 19441 3485 19475 3519
rect 21005 3485 21039 3519
rect 23397 3485 23431 3519
rect 24041 3485 24075 3519
rect 27169 3485 27203 3519
rect 27813 3485 27847 3519
rect 28273 3485 28307 3519
rect 28917 3485 28951 3519
rect 29745 3485 29779 3519
rect 46121 3485 46155 3519
rect 47961 3485 47995 3519
rect 21189 3417 21223 3451
rect 22845 3417 22879 3451
rect 47317 3417 47351 3451
rect 8769 3349 8803 3383
rect 9413 3349 9447 3383
rect 10701 3349 10735 3383
rect 11805 3349 11839 3383
rect 16313 3349 16347 3383
rect 16957 3349 16991 3383
rect 26341 3349 26375 3383
rect 30389 3349 30423 3383
rect 2145 3145 2179 3179
rect 10057 3145 10091 3179
rect 11161 3145 11195 3179
rect 18705 3145 18739 3179
rect 22753 3145 22787 3179
rect 23305 3145 23339 3179
rect 27997 3145 28031 3179
rect 19533 3077 19567 3111
rect 23857 3077 23891 3111
rect 29101 3077 29135 3111
rect 49157 3077 49191 3111
rect 1593 3009 1627 3043
rect 2513 3009 2547 3043
rect 8309 3009 8343 3043
rect 9413 3009 9447 3043
rect 10517 3009 10551 3043
rect 12357 3009 12391 3043
rect 13001 3009 13035 3043
rect 13461 3009 13495 3043
rect 14565 3009 14599 3043
rect 17049 3009 17083 3043
rect 18889 3009 18923 3043
rect 22293 3009 22327 3043
rect 27537 3009 27571 3043
rect 28825 3009 28859 3043
rect 44005 3009 44039 3043
rect 45845 3009 45879 3043
rect 47961 3009 47995 3043
rect 14105 2941 14139 2975
rect 14841 2941 14875 2975
rect 17325 2941 17359 2975
rect 19349 2941 19383 2975
rect 21189 2941 21223 2975
rect 23673 2941 23707 2975
rect 24133 2941 24167 2975
rect 30573 2941 30607 2975
rect 45201 2941 45235 2975
rect 46857 2941 46891 2975
rect 1777 2873 1811 2907
rect 2329 2805 2363 2839
rect 2789 2805 2823 2839
rect 8953 2805 8987 2839
rect 16313 2805 16347 2839
rect 22385 2805 22419 2839
rect 27813 2805 27847 2839
rect 3065 2601 3099 2635
rect 9781 2601 9815 2635
rect 10885 2601 10919 2635
rect 24501 2601 24535 2635
rect 25145 2601 25179 2635
rect 30849 2601 30883 2635
rect 32965 2601 32999 2635
rect 35081 2601 35115 2635
rect 2513 2533 2547 2567
rect 28733 2533 28767 2567
rect 8585 2465 8619 2499
rect 12265 2465 12299 2499
rect 14749 2465 14783 2499
rect 22201 2465 22235 2499
rect 22385 2465 22419 2499
rect 25329 2465 25363 2499
rect 37749 2465 37783 2499
rect 41429 2465 41463 2499
rect 49157 2465 49191 2499
rect 1593 2397 1627 2431
rect 2329 2397 2363 2431
rect 3249 2397 3283 2431
rect 3525 2397 3559 2431
rect 7941 2397 7975 2431
rect 9137 2397 9171 2431
rect 10241 2397 10275 2431
rect 11989 2397 12023 2431
rect 14473 2397 14507 2431
rect 17693 2397 17727 2431
rect 20453 2397 20487 2431
rect 24869 2397 24903 2431
rect 28917 2397 28951 2431
rect 29193 2397 29227 2431
rect 31033 2397 31067 2431
rect 31309 2397 31343 2431
rect 33149 2397 33183 2431
rect 33425 2397 33459 2431
rect 35265 2397 35299 2431
rect 35541 2397 35575 2431
rect 37473 2397 37507 2431
rect 40693 2397 40727 2431
rect 45845 2397 45879 2431
rect 47961 2397 47995 2431
rect 18429 2329 18463 2363
rect 24041 2329 24075 2363
rect 47041 2329 47075 2363
rect 1777 2261 1811 2295
rect 20269 2261 20303 2295
rect 37105 2261 37139 2295
<< metal1 >>
rect 24210 26324 24216 26376
rect 24268 26364 24274 26376
rect 43806 26364 43812 26376
rect 24268 26336 43812 26364
rect 24268 26324 24274 26336
rect 43806 26324 43812 26336
rect 43864 26324 43870 26376
rect 12250 26256 12256 26308
rect 12308 26296 12314 26308
rect 26326 26296 26332 26308
rect 12308 26268 26332 26296
rect 12308 26256 12314 26268
rect 26326 26256 26332 26268
rect 26384 26256 26390 26308
rect 33502 26188 33508 26240
rect 33560 26228 33566 26240
rect 47210 26228 47216 26240
rect 33560 26200 47216 26228
rect 33560 26188 33566 26200
rect 47210 26188 47216 26200
rect 47268 26188 47274 26240
rect 35802 26120 35808 26172
rect 35860 26160 35866 26172
rect 47486 26160 47492 26172
rect 35860 26132 47492 26160
rect 35860 26120 35866 26132
rect 47486 26120 47492 26132
rect 47544 26120 47550 26172
rect 28350 26052 28356 26104
rect 28408 26092 28414 26104
rect 43346 26092 43352 26104
rect 28408 26064 43352 26092
rect 28408 26052 28414 26064
rect 43346 26052 43352 26064
rect 43404 26052 43410 26104
rect 21174 25984 21180 26036
rect 21232 26024 21238 26036
rect 47118 26024 47124 26036
rect 21232 25996 47124 26024
rect 21232 25984 21238 25996
rect 47118 25984 47124 25996
rect 47176 25984 47182 26036
rect 19702 25916 19708 25968
rect 19760 25956 19766 25968
rect 45554 25956 45560 25968
rect 19760 25928 45560 25956
rect 19760 25916 19766 25928
rect 45554 25916 45560 25928
rect 45612 25916 45618 25968
rect 26878 25848 26884 25900
rect 26936 25888 26942 25900
rect 45186 25888 45192 25900
rect 26936 25860 45192 25888
rect 26936 25848 26942 25860
rect 45186 25848 45192 25860
rect 45244 25848 45250 25900
rect 24302 25780 24308 25832
rect 24360 25820 24366 25832
rect 40862 25820 40868 25832
rect 24360 25792 40868 25820
rect 24360 25780 24366 25792
rect 40862 25780 40868 25792
rect 40920 25780 40926 25832
rect 21726 25712 21732 25764
rect 21784 25752 21790 25764
rect 49234 25752 49240 25764
rect 21784 25724 49240 25752
rect 21784 25712 21790 25724
rect 49234 25712 49240 25724
rect 49292 25712 49298 25764
rect 4338 25644 4344 25696
rect 4396 25684 4402 25696
rect 44174 25684 44180 25696
rect 4396 25656 44180 25684
rect 4396 25644 4402 25656
rect 44174 25644 44180 25656
rect 44232 25644 44238 25696
rect 20346 25576 20352 25628
rect 20404 25616 20410 25628
rect 48774 25616 48780 25628
rect 20404 25588 48780 25616
rect 20404 25576 20410 25588
rect 48774 25576 48780 25588
rect 48832 25576 48838 25628
rect 12066 25508 12072 25560
rect 12124 25548 12130 25560
rect 44450 25548 44456 25560
rect 12124 25520 44456 25548
rect 12124 25508 12130 25520
rect 44450 25508 44456 25520
rect 44508 25508 44514 25560
rect 25130 25440 25136 25492
rect 25188 25480 25194 25492
rect 41874 25480 41880 25492
rect 25188 25452 41880 25480
rect 25188 25440 25194 25452
rect 41874 25440 41880 25452
rect 41932 25440 41938 25492
rect 27246 25372 27252 25424
rect 27304 25412 27310 25424
rect 44358 25412 44364 25424
rect 27304 25384 44364 25412
rect 27304 25372 27310 25384
rect 44358 25372 44364 25384
rect 44416 25372 44422 25424
rect 30558 25304 30564 25356
rect 30616 25344 30622 25356
rect 49050 25344 49056 25356
rect 30616 25316 49056 25344
rect 30616 25304 30622 25316
rect 49050 25304 49056 25316
rect 49108 25304 49114 25356
rect 17310 25236 17316 25288
rect 17368 25276 17374 25288
rect 40310 25276 40316 25288
rect 17368 25248 40316 25276
rect 17368 25236 17374 25248
rect 40310 25236 40316 25248
rect 40368 25236 40374 25288
rect 4062 25168 4068 25220
rect 4120 25208 4126 25220
rect 8846 25208 8852 25220
rect 4120 25180 8852 25208
rect 4120 25168 4126 25180
rect 8846 25168 8852 25180
rect 8904 25168 8910 25220
rect 35894 25168 35900 25220
rect 35952 25208 35958 25220
rect 42518 25208 42524 25220
rect 35952 25180 42524 25208
rect 35952 25168 35958 25180
rect 42518 25168 42524 25180
rect 42576 25168 42582 25220
rect 28258 25100 28264 25152
rect 28316 25140 28322 25152
rect 41414 25140 41420 25152
rect 28316 25112 41420 25140
rect 28316 25100 28322 25112
rect 41414 25100 41420 25112
rect 41472 25100 41478 25152
rect 15010 25032 15016 25084
rect 15068 25072 15074 25084
rect 31754 25072 31760 25084
rect 15068 25044 31760 25072
rect 15068 25032 15074 25044
rect 31754 25032 31760 25044
rect 31812 25032 31818 25084
rect 32214 25032 32220 25084
rect 32272 25072 32278 25084
rect 41966 25072 41972 25084
rect 32272 25044 41972 25072
rect 32272 25032 32278 25044
rect 41966 25032 41972 25044
rect 42024 25032 42030 25084
rect 15194 24964 15200 25016
rect 15252 25004 15258 25016
rect 27062 25004 27068 25016
rect 15252 24976 27068 25004
rect 15252 24964 15258 24976
rect 27062 24964 27068 24976
rect 27120 24964 27126 25016
rect 41322 24964 41328 25016
rect 41380 25004 41386 25016
rect 45830 25004 45836 25016
rect 41380 24976 45836 25004
rect 41380 24964 41386 24976
rect 45830 24964 45836 24976
rect 45888 24964 45894 25016
rect 4706 24896 4712 24948
rect 4764 24936 4770 24948
rect 4764 24908 12434 24936
rect 4764 24896 4770 24908
rect 3418 24828 3424 24880
rect 3476 24868 3482 24880
rect 9858 24868 9864 24880
rect 3476 24840 9864 24868
rect 3476 24828 3482 24840
rect 9858 24828 9864 24840
rect 9916 24828 9922 24880
rect 12406 24868 12434 24908
rect 12710 24896 12716 24948
rect 12768 24936 12774 24948
rect 33502 24936 33508 24948
rect 12768 24908 33508 24936
rect 12768 24896 12774 24908
rect 33502 24896 33508 24908
rect 33560 24896 33566 24948
rect 19886 24868 19892 24880
rect 12406 24840 19892 24868
rect 19886 24828 19892 24840
rect 19944 24828 19950 24880
rect 24578 24828 24584 24880
rect 24636 24868 24642 24880
rect 24636 24840 35848 24868
rect 24636 24828 24642 24840
rect 3694 24760 3700 24812
rect 3752 24800 3758 24812
rect 6270 24800 6276 24812
rect 3752 24772 6276 24800
rect 3752 24760 3758 24772
rect 6270 24760 6276 24772
rect 6328 24760 6334 24812
rect 30926 24760 30932 24812
rect 30984 24800 30990 24812
rect 33962 24800 33968 24812
rect 30984 24772 33968 24800
rect 30984 24760 30990 24772
rect 33962 24760 33968 24772
rect 34020 24760 34026 24812
rect 35820 24800 35848 24840
rect 36814 24828 36820 24880
rect 36872 24868 36878 24880
rect 43438 24868 43444 24880
rect 36872 24840 43444 24868
rect 36872 24828 36878 24840
rect 43438 24828 43444 24840
rect 43496 24828 43502 24880
rect 47762 24800 47768 24812
rect 35820 24772 47768 24800
rect 47762 24760 47768 24772
rect 47820 24760 47826 24812
rect 11790 24692 11796 24744
rect 11848 24732 11854 24744
rect 23382 24732 23388 24744
rect 11848 24704 23388 24732
rect 11848 24692 11854 24704
rect 23382 24692 23388 24704
rect 23440 24692 23446 24744
rect 30006 24692 30012 24744
rect 30064 24732 30070 24744
rect 42794 24732 42800 24744
rect 30064 24704 42800 24732
rect 30064 24692 30070 24704
rect 42794 24692 42800 24704
rect 42852 24692 42858 24744
rect 14182 24624 14188 24676
rect 14240 24664 14246 24676
rect 24854 24664 24860 24676
rect 14240 24636 24860 24664
rect 14240 24624 14246 24636
rect 24854 24624 24860 24636
rect 24912 24624 24918 24676
rect 34146 24664 34152 24676
rect 24964 24636 34152 24664
rect 1762 24556 1768 24608
rect 1820 24596 1826 24608
rect 11330 24596 11336 24608
rect 1820 24568 11336 24596
rect 1820 24556 1826 24568
rect 11330 24556 11336 24568
rect 11388 24556 11394 24608
rect 14826 24556 14832 24608
rect 14884 24596 14890 24608
rect 21358 24596 21364 24608
rect 14884 24568 21364 24596
rect 14884 24556 14890 24568
rect 21358 24556 21364 24568
rect 21416 24556 21422 24608
rect 23658 24556 23664 24608
rect 23716 24596 23722 24608
rect 24964 24596 24992 24636
rect 34146 24624 34152 24636
rect 34204 24624 34210 24676
rect 35526 24624 35532 24676
rect 35584 24664 35590 24676
rect 37550 24664 37556 24676
rect 35584 24636 37556 24664
rect 35584 24624 35590 24636
rect 37550 24624 37556 24636
rect 37608 24664 37614 24676
rect 40678 24664 40684 24676
rect 37608 24636 40684 24664
rect 37608 24624 37614 24636
rect 40678 24624 40684 24636
rect 40736 24624 40742 24676
rect 23716 24568 24992 24596
rect 23716 24556 23722 24568
rect 25958 24556 25964 24608
rect 26016 24596 26022 24608
rect 30834 24596 30840 24608
rect 26016 24568 30840 24596
rect 26016 24556 26022 24568
rect 30834 24556 30840 24568
rect 30892 24556 30898 24608
rect 31294 24556 31300 24608
rect 31352 24596 31358 24608
rect 37458 24596 37464 24608
rect 31352 24568 37464 24596
rect 31352 24556 31358 24568
rect 37458 24556 37464 24568
rect 37516 24556 37522 24608
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 1762 24352 1768 24404
rect 1820 24352 1826 24404
rect 2314 24352 2320 24404
rect 2372 24392 2378 24404
rect 6549 24395 6607 24401
rect 2372 24364 5764 24392
rect 2372 24352 2378 24364
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 3510 24256 3516 24268
rect 3283 24228 3516 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 2130 24148 2136 24200
rect 2188 24148 2194 24200
rect 2406 24148 2412 24200
rect 2464 24188 2470 24200
rect 4157 24191 4215 24197
rect 2464 24160 3740 24188
rect 2464 24148 2470 24160
rect 1581 24123 1639 24129
rect 1581 24089 1593 24123
rect 1627 24120 1639 24123
rect 3602 24120 3608 24132
rect 1627 24092 3608 24120
rect 1627 24089 1639 24092
rect 1581 24083 1639 24089
rect 3602 24080 3608 24092
rect 3660 24080 3666 24132
rect 3712 24120 3740 24160
rect 4157 24157 4169 24191
rect 4203 24188 4215 24191
rect 4246 24188 4252 24200
rect 4203 24160 4252 24188
rect 4203 24157 4215 24160
rect 4157 24151 4215 24157
rect 4246 24148 4252 24160
rect 4304 24148 4310 24200
rect 4617 24191 4675 24197
rect 4617 24157 4629 24191
rect 4663 24157 4675 24191
rect 5736 24188 5764 24364
rect 6549 24361 6561 24395
rect 6595 24392 6607 24395
rect 10502 24392 10508 24404
rect 6595 24364 10508 24392
rect 6595 24361 6607 24364
rect 6549 24355 6607 24361
rect 10502 24352 10508 24364
rect 10560 24352 10566 24404
rect 19426 24392 19432 24404
rect 16224 24364 19432 24392
rect 6730 24324 6736 24336
rect 5828 24296 6736 24324
rect 5828 24265 5856 24296
rect 6730 24284 6736 24296
rect 6788 24284 6794 24336
rect 10134 24324 10140 24336
rect 6840 24296 10140 24324
rect 5813 24259 5871 24265
rect 5813 24225 5825 24259
rect 5859 24225 5871 24259
rect 6840 24256 6868 24296
rect 10134 24284 10140 24296
rect 10192 24284 10198 24336
rect 11606 24284 11612 24336
rect 11664 24324 11670 24336
rect 16224 24324 16252 24364
rect 19426 24352 19432 24364
rect 19484 24352 19490 24404
rect 27341 24395 27399 24401
rect 27341 24392 27353 24395
rect 19536 24364 27353 24392
rect 11664 24296 16252 24324
rect 11664 24284 11670 24296
rect 5813 24219 5871 24225
rect 5920 24228 6868 24256
rect 8205 24259 8263 24265
rect 5920 24188 5948 24228
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 8662 24256 8668 24268
rect 8251 24228 8668 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 8662 24216 8668 24228
rect 8720 24216 8726 24268
rect 8938 24216 8944 24268
rect 8996 24256 9002 24268
rect 10965 24259 11023 24265
rect 8996 24228 9812 24256
rect 8996 24216 9002 24228
rect 5736 24160 5948 24188
rect 6733 24191 6791 24197
rect 4617 24151 4675 24157
rect 6733 24157 6745 24191
rect 6779 24157 6791 24191
rect 6733 24151 6791 24157
rect 7377 24191 7435 24197
rect 7377 24157 7389 24191
rect 7423 24157 7435 24191
rect 7377 24151 7435 24157
rect 4632 24120 4660 24151
rect 3712 24092 4660 24120
rect 3694 24012 3700 24064
rect 3752 24052 3758 24064
rect 3973 24055 4031 24061
rect 3973 24052 3985 24055
rect 3752 24024 3985 24052
rect 3752 24012 3758 24024
rect 3973 24021 3985 24024
rect 4019 24021 4031 24055
rect 3973 24015 4031 24021
rect 4062 24012 4068 24064
rect 4120 24052 4126 24064
rect 6748 24052 6776 24151
rect 7392 24120 7420 24151
rect 9030 24148 9036 24200
rect 9088 24188 9094 24200
rect 9784 24197 9812 24228
rect 10965 24225 10977 24259
rect 11011 24256 11023 24259
rect 12434 24256 12440 24268
rect 11011 24228 12440 24256
rect 11011 24225 11023 24228
rect 10965 24219 11023 24225
rect 12434 24216 12440 24228
rect 12492 24216 12498 24268
rect 13541 24259 13599 24265
rect 13541 24225 13553 24259
rect 13587 24256 13599 24259
rect 14458 24256 14464 24268
rect 13587 24228 14464 24256
rect 13587 24225 13599 24228
rect 13541 24219 13599 24225
rect 14458 24216 14464 24228
rect 14516 24216 14522 24268
rect 18693 24259 18751 24265
rect 18693 24225 18705 24259
rect 18739 24256 18751 24259
rect 19242 24256 19248 24268
rect 18739 24228 19248 24256
rect 18739 24225 18751 24228
rect 18693 24219 18751 24225
rect 19242 24216 19248 24228
rect 19300 24216 19306 24268
rect 19536 24256 19564 24364
rect 27341 24361 27353 24364
rect 27387 24361 27399 24395
rect 27341 24355 27399 24361
rect 27522 24352 27528 24404
rect 27580 24392 27586 24404
rect 31846 24392 31852 24404
rect 27580 24364 31852 24392
rect 27580 24352 27586 24364
rect 31846 24352 31852 24364
rect 31904 24352 31910 24404
rect 32122 24352 32128 24404
rect 32180 24392 32186 24404
rect 32180 24364 33732 24392
rect 32180 24352 32186 24364
rect 21174 24284 21180 24336
rect 21232 24284 21238 24336
rect 24394 24284 24400 24336
rect 24452 24324 24458 24336
rect 27893 24327 27951 24333
rect 27893 24324 27905 24327
rect 24452 24296 27905 24324
rect 24452 24284 24458 24296
rect 27893 24293 27905 24296
rect 27939 24293 27951 24327
rect 33704 24324 33732 24364
rect 34146 24352 34152 24404
rect 34204 24352 34210 24404
rect 36081 24395 36139 24401
rect 36081 24392 36093 24395
rect 34256 24364 36093 24392
rect 34256 24324 34284 24364
rect 36081 24361 36093 24364
rect 36127 24361 36139 24395
rect 36081 24355 36139 24361
rect 37458 24352 37464 24404
rect 37516 24352 37522 24404
rect 40678 24352 40684 24404
rect 40736 24392 40742 24404
rect 40736 24364 42288 24392
rect 40736 24352 40742 24364
rect 27893 24287 27951 24293
rect 32968 24296 33640 24324
rect 33704 24296 34284 24324
rect 34885 24327 34943 24333
rect 19352 24228 19564 24256
rect 9217 24191 9275 24197
rect 9217 24188 9229 24191
rect 9088 24160 9229 24188
rect 9088 24148 9094 24160
rect 9217 24157 9229 24160
rect 9263 24157 9275 24191
rect 9217 24151 9275 24157
rect 9769 24191 9827 24197
rect 9769 24157 9781 24191
rect 9815 24157 9827 24191
rect 9769 24151 9827 24157
rect 12529 24191 12587 24197
rect 12529 24157 12541 24191
rect 12575 24188 12587 24191
rect 13998 24188 14004 24200
rect 12575 24160 14004 24188
rect 12575 24157 12587 24160
rect 12529 24151 12587 24157
rect 13998 24148 14004 24160
rect 14056 24148 14062 24200
rect 15105 24191 15163 24197
rect 15105 24157 15117 24191
rect 15151 24188 15163 24191
rect 15194 24188 15200 24200
rect 15151 24160 15200 24188
rect 15151 24157 15163 24160
rect 15105 24151 15163 24157
rect 15194 24148 15200 24160
rect 15252 24148 15258 24200
rect 16942 24188 16948 24200
rect 16040 24160 16948 24188
rect 10778 24120 10784 24132
rect 7392 24092 10784 24120
rect 10778 24080 10784 24092
rect 10836 24080 10842 24132
rect 11698 24080 11704 24132
rect 11756 24080 11762 24132
rect 11885 24123 11943 24129
rect 11885 24089 11897 24123
rect 11931 24120 11943 24123
rect 12158 24120 12164 24132
rect 11931 24092 12164 24120
rect 11931 24089 11943 24092
rect 11885 24083 11943 24089
rect 12158 24080 12164 24092
rect 12216 24080 12222 24132
rect 16040 24120 16068 24160
rect 16942 24148 16948 24160
rect 17000 24148 17006 24200
rect 17037 24191 17095 24197
rect 17037 24157 17049 24191
rect 17083 24188 17095 24191
rect 17126 24188 17132 24200
rect 17083 24160 17132 24188
rect 17083 24157 17095 24160
rect 17037 24151 17095 24157
rect 17126 24148 17132 24160
rect 17184 24148 17190 24200
rect 17681 24191 17739 24197
rect 17681 24157 17693 24191
rect 17727 24188 17739 24191
rect 19352 24188 19380 24228
rect 21266 24216 21272 24268
rect 21324 24256 21330 24268
rect 22465 24259 22523 24265
rect 22465 24256 22477 24259
rect 21324 24228 22477 24256
rect 21324 24216 21330 24228
rect 22465 24225 22477 24228
rect 22511 24225 22523 24259
rect 25406 24256 25412 24268
rect 22465 24219 22523 24225
rect 24044 24228 25412 24256
rect 17727 24160 19380 24188
rect 19429 24191 19487 24197
rect 17727 24157 17739 24160
rect 17681 24151 17739 24157
rect 19429 24157 19441 24191
rect 19475 24157 19487 24191
rect 19429 24151 19487 24157
rect 14200 24092 16068 24120
rect 16117 24123 16175 24129
rect 4120 24024 6776 24052
rect 9125 24055 9183 24061
rect 4120 24012 4126 24024
rect 9125 24021 9137 24055
rect 9171 24052 9183 24055
rect 9306 24052 9312 24064
rect 9171 24024 9312 24052
rect 9171 24021 9183 24024
rect 9125 24015 9183 24021
rect 9306 24012 9312 24024
rect 9364 24012 9370 24064
rect 9398 24012 9404 24064
rect 9456 24052 9462 24064
rect 11422 24052 11428 24064
rect 9456 24024 11428 24052
rect 9456 24012 9462 24024
rect 11422 24012 11428 24024
rect 11480 24012 11486 24064
rect 12069 24055 12127 24061
rect 12069 24021 12081 24055
rect 12115 24052 12127 24055
rect 14200 24052 14228 24092
rect 16117 24089 16129 24123
rect 16163 24120 16175 24123
rect 18322 24120 18328 24132
rect 16163 24092 18328 24120
rect 16163 24089 16175 24092
rect 16117 24083 16175 24089
rect 18322 24080 18328 24092
rect 18380 24080 18386 24132
rect 19242 24080 19248 24132
rect 19300 24120 19306 24132
rect 19444 24120 19472 24151
rect 22094 24148 22100 24200
rect 22152 24148 22158 24200
rect 24044 24197 24072 24228
rect 25406 24216 25412 24228
rect 25464 24216 25470 24268
rect 28442 24216 28448 24268
rect 28500 24216 28506 24268
rect 28718 24216 28724 24268
rect 28776 24256 28782 24268
rect 32968 24265 32996 24296
rect 32953 24259 33011 24265
rect 28776 24228 30972 24256
rect 28776 24216 28782 24228
rect 24029 24191 24087 24197
rect 24029 24157 24041 24191
rect 24075 24157 24087 24191
rect 24029 24151 24087 24157
rect 24854 24148 24860 24200
rect 24912 24148 24918 24200
rect 25958 24148 25964 24200
rect 26016 24148 26022 24200
rect 26605 24191 26663 24197
rect 26605 24157 26617 24191
rect 26651 24188 26663 24191
rect 27430 24188 27436 24200
rect 26651 24160 27436 24188
rect 26651 24157 26663 24160
rect 26605 24151 26663 24157
rect 27430 24148 27436 24160
rect 27488 24148 27494 24200
rect 28258 24148 28264 24200
rect 28316 24148 28322 24200
rect 29178 24148 29184 24200
rect 29236 24148 29242 24200
rect 29454 24148 29460 24200
rect 29512 24188 29518 24200
rect 29733 24191 29791 24197
rect 29733 24188 29745 24191
rect 29512 24160 29745 24188
rect 29512 24148 29518 24160
rect 29733 24157 29745 24160
rect 29779 24157 29791 24191
rect 29733 24151 29791 24157
rect 30006 24148 30012 24200
rect 30064 24188 30070 24200
rect 30837 24191 30895 24197
rect 30837 24188 30849 24191
rect 30064 24160 30849 24188
rect 30064 24148 30070 24160
rect 30837 24157 30849 24160
rect 30883 24157 30895 24191
rect 30837 24151 30895 24157
rect 19300 24092 19472 24120
rect 19300 24080 19306 24092
rect 19702 24080 19708 24132
rect 19760 24080 19766 24132
rect 19978 24080 19984 24132
rect 20036 24120 20042 24132
rect 27249 24123 27307 24129
rect 27249 24120 27261 24123
rect 20036 24092 20194 24120
rect 21192 24092 24624 24120
rect 20036 24080 20042 24092
rect 12115 24024 14228 24052
rect 14277 24055 14335 24061
rect 12115 24021 12127 24024
rect 12069 24015 12127 24021
rect 14277 24021 14289 24055
rect 14323 24052 14335 24055
rect 16758 24052 16764 24064
rect 14323 24024 16764 24052
rect 14323 24021 14335 24024
rect 14277 24015 14335 24021
rect 16758 24012 16764 24024
rect 16816 24012 16822 24064
rect 16853 24055 16911 24061
rect 16853 24021 16865 24055
rect 16899 24052 16911 24055
rect 21192 24052 21220 24092
rect 16899 24024 21220 24052
rect 16899 24021 16911 24024
rect 16853 24015 16911 24021
rect 21266 24012 21272 24064
rect 21324 24052 21330 24064
rect 21545 24055 21603 24061
rect 21545 24052 21557 24055
rect 21324 24024 21557 24052
rect 21324 24012 21330 24024
rect 21545 24021 21557 24024
rect 21591 24021 21603 24055
rect 21545 24015 21603 24021
rect 23842 24012 23848 24064
rect 23900 24012 23906 24064
rect 24486 24012 24492 24064
rect 24544 24012 24550 24064
rect 24596 24052 24624 24092
rect 24872 24092 27261 24120
rect 24872 24052 24900 24092
rect 27249 24089 27261 24092
rect 27295 24089 27307 24123
rect 27249 24083 27307 24089
rect 28353 24123 28411 24129
rect 28353 24089 28365 24123
rect 28399 24120 28411 24123
rect 30466 24120 30472 24132
rect 28399 24092 30472 24120
rect 28399 24089 28411 24092
rect 28353 24083 28411 24089
rect 30466 24080 30472 24092
rect 30524 24080 30530 24132
rect 30944 24120 30972 24228
rect 32953 24225 32965 24259
rect 32999 24225 33011 24259
rect 33612 24256 33640 24296
rect 34885 24293 34897 24327
rect 34931 24324 34943 24327
rect 34931 24296 39160 24324
rect 34931 24293 34943 24296
rect 34885 24287 34943 24293
rect 34974 24256 34980 24268
rect 33612 24228 34980 24256
rect 32953 24219 33011 24225
rect 34974 24216 34980 24228
rect 35032 24216 35038 24268
rect 35526 24216 35532 24268
rect 35584 24216 35590 24268
rect 35802 24216 35808 24268
rect 35860 24256 35866 24268
rect 36725 24259 36783 24265
rect 36725 24256 36737 24259
rect 35860 24228 36737 24256
rect 35860 24216 35866 24228
rect 36725 24225 36737 24228
rect 36771 24256 36783 24259
rect 36814 24256 36820 24268
rect 36771 24228 36820 24256
rect 36771 24225 36783 24228
rect 36725 24219 36783 24225
rect 36814 24216 36820 24228
rect 36872 24216 36878 24268
rect 38105 24259 38163 24265
rect 38105 24225 38117 24259
rect 38151 24256 38163 24259
rect 38654 24256 38660 24268
rect 38151 24228 38660 24256
rect 38151 24225 38163 24228
rect 38105 24219 38163 24225
rect 38654 24216 38660 24228
rect 38712 24216 38718 24268
rect 39132 24265 39160 24296
rect 39942 24284 39948 24336
rect 40000 24324 40006 24336
rect 40000 24296 41287 24324
rect 40000 24284 40006 24296
rect 39117 24259 39175 24265
rect 39117 24225 39129 24259
rect 39163 24225 39175 24259
rect 39117 24219 39175 24225
rect 39301 24259 39359 24265
rect 39301 24225 39313 24259
rect 39347 24256 39359 24259
rect 39390 24256 39396 24268
rect 39347 24228 39396 24256
rect 39347 24225 39359 24228
rect 39301 24219 39359 24225
rect 39390 24216 39396 24228
rect 39448 24216 39454 24268
rect 40678 24216 40684 24268
rect 40736 24216 40742 24268
rect 33502 24148 33508 24200
rect 33560 24148 33566 24200
rect 35250 24148 35256 24200
rect 35308 24188 35314 24200
rect 35345 24191 35403 24197
rect 35345 24188 35357 24191
rect 35308 24160 35357 24188
rect 35308 24148 35314 24160
rect 35345 24157 35357 24160
rect 35391 24157 35403 24191
rect 35345 24151 35403 24157
rect 35618 24148 35624 24200
rect 35676 24188 35682 24200
rect 36541 24191 36599 24197
rect 36541 24188 36553 24191
rect 35676 24160 36553 24188
rect 35676 24148 35682 24160
rect 36541 24157 36553 24160
rect 36587 24157 36599 24191
rect 36541 24151 36599 24157
rect 37921 24191 37979 24197
rect 37921 24157 37933 24191
rect 37967 24188 37979 24191
rect 39666 24188 39672 24200
rect 37967 24160 39672 24188
rect 37967 24157 37979 24160
rect 37921 24151 37979 24157
rect 39666 24148 39672 24160
rect 39724 24148 39730 24200
rect 41259 24197 41287 24296
rect 41414 24216 41420 24268
rect 41472 24256 41478 24268
rect 42153 24259 42211 24265
rect 42153 24256 42165 24259
rect 41472 24228 42165 24256
rect 41472 24216 41478 24228
rect 42153 24225 42165 24228
rect 42199 24225 42211 24259
rect 42260 24256 42288 24364
rect 42794 24352 42800 24404
rect 42852 24392 42858 24404
rect 44637 24395 44695 24401
rect 44637 24392 44649 24395
rect 42852 24364 44649 24392
rect 42852 24352 42858 24364
rect 44637 24361 44649 24364
rect 44683 24361 44695 24395
rect 44637 24355 44695 24361
rect 45738 24352 45744 24404
rect 45796 24392 45802 24404
rect 45833 24395 45891 24401
rect 45833 24392 45845 24395
rect 45796 24364 45845 24392
rect 45796 24352 45802 24364
rect 45833 24361 45845 24364
rect 45879 24361 45891 24395
rect 45833 24355 45891 24361
rect 47210 24352 47216 24404
rect 47268 24352 47274 24404
rect 44082 24284 44088 24336
rect 44140 24324 44146 24336
rect 48041 24327 48099 24333
rect 48041 24324 48053 24327
rect 44140 24296 48053 24324
rect 44140 24284 44146 24296
rect 48041 24293 48053 24296
rect 48087 24293 48099 24327
rect 48041 24287 48099 24293
rect 46198 24256 46204 24268
rect 42260 24228 46204 24256
rect 42153 24219 42211 24225
rect 46198 24216 46204 24228
rect 46256 24216 46262 24268
rect 46937 24259 46995 24265
rect 46937 24256 46949 24259
rect 46400 24228 46949 24256
rect 41249 24191 41307 24197
rect 41249 24157 41261 24191
rect 41295 24157 41307 24191
rect 41249 24151 41307 24157
rect 42613 24191 42671 24197
rect 42613 24157 42625 24191
rect 42659 24157 42671 24191
rect 42613 24151 42671 24157
rect 31757 24123 31815 24129
rect 31757 24120 31769 24123
rect 30944 24092 31769 24120
rect 31757 24089 31769 24092
rect 31803 24089 31815 24123
rect 31757 24083 31815 24089
rect 32769 24123 32827 24129
rect 32769 24089 32781 24123
rect 32815 24120 32827 24123
rect 39025 24123 39083 24129
rect 32815 24092 33640 24120
rect 32815 24089 32827 24092
rect 32769 24083 32827 24089
rect 24596 24024 24900 24052
rect 25222 24012 25228 24064
rect 25280 24052 25286 24064
rect 25501 24055 25559 24061
rect 25501 24052 25513 24055
rect 25280 24024 25513 24052
rect 25280 24012 25286 24024
rect 25501 24021 25513 24024
rect 25547 24021 25559 24055
rect 25501 24015 25559 24021
rect 28994 24012 29000 24064
rect 29052 24012 29058 24064
rect 29365 24055 29423 24061
rect 29365 24021 29377 24055
rect 29411 24052 29423 24055
rect 30282 24052 30288 24064
rect 29411 24024 30288 24052
rect 29411 24021 29423 24024
rect 29365 24015 29423 24021
rect 30282 24012 30288 24024
rect 30340 24012 30346 24064
rect 30374 24012 30380 24064
rect 30432 24012 30438 24064
rect 31110 24012 31116 24064
rect 31168 24052 31174 24064
rect 31481 24055 31539 24061
rect 31481 24052 31493 24055
rect 31168 24024 31493 24052
rect 31168 24012 31174 24024
rect 31481 24021 31493 24024
rect 31527 24021 31539 24055
rect 31481 24015 31539 24021
rect 32306 24012 32312 24064
rect 32364 24012 32370 24064
rect 32677 24055 32735 24061
rect 32677 24021 32689 24055
rect 32723 24052 32735 24055
rect 33134 24052 33140 24064
rect 32723 24024 33140 24052
rect 32723 24021 32735 24024
rect 32677 24015 32735 24021
rect 33134 24012 33140 24024
rect 33192 24012 33198 24064
rect 33612 24052 33640 24092
rect 33888 24092 38700 24120
rect 33888 24052 33916 24092
rect 33612 24024 33916 24052
rect 33962 24012 33968 24064
rect 34020 24052 34026 24064
rect 34425 24055 34483 24061
rect 34425 24052 34437 24055
rect 34020 24024 34437 24052
rect 34020 24012 34026 24024
rect 34425 24021 34437 24024
rect 34471 24021 34483 24055
rect 34425 24015 34483 24021
rect 35253 24055 35311 24061
rect 35253 24021 35265 24055
rect 35299 24052 35311 24055
rect 35710 24052 35716 24064
rect 35299 24024 35716 24052
rect 35299 24021 35311 24024
rect 35253 24015 35311 24021
rect 35710 24012 35716 24024
rect 35768 24012 35774 24064
rect 36446 24012 36452 24064
rect 36504 24012 36510 24064
rect 36538 24012 36544 24064
rect 36596 24052 36602 24064
rect 38672 24061 38700 24092
rect 39025 24089 39037 24123
rect 39071 24120 39083 24123
rect 40497 24123 40555 24129
rect 39071 24092 40080 24120
rect 39071 24089 39083 24092
rect 39025 24083 39083 24089
rect 40052 24061 40080 24092
rect 40497 24089 40509 24123
rect 40543 24120 40555 24123
rect 41690 24120 41696 24132
rect 40543 24092 41696 24120
rect 40543 24089 40555 24092
rect 40497 24083 40555 24089
rect 41690 24080 41696 24092
rect 41748 24080 41754 24132
rect 42628 24120 42656 24151
rect 42702 24148 42708 24200
rect 42760 24188 42766 24200
rect 43717 24191 43775 24197
rect 43717 24188 43729 24191
rect 42760 24160 43729 24188
rect 42760 24148 42766 24160
rect 43717 24157 43729 24160
rect 43763 24157 43775 24191
rect 43717 24151 43775 24157
rect 45189 24191 45247 24197
rect 45189 24157 45201 24191
rect 45235 24188 45247 24191
rect 45646 24188 45652 24200
rect 45235 24160 45652 24188
rect 45235 24157 45247 24160
rect 45189 24151 45247 24157
rect 45646 24148 45652 24160
rect 45704 24148 45710 24200
rect 46290 24148 46296 24200
rect 46348 24148 46354 24200
rect 44361 24123 44419 24129
rect 44361 24120 44373 24123
rect 42628 24092 44373 24120
rect 44361 24089 44373 24092
rect 44407 24089 44419 24123
rect 44361 24083 44419 24089
rect 37829 24055 37887 24061
rect 37829 24052 37841 24055
rect 36596 24024 37841 24052
rect 36596 24012 36602 24024
rect 37829 24021 37841 24024
rect 37875 24021 37887 24055
rect 37829 24015 37887 24021
rect 38657 24055 38715 24061
rect 38657 24021 38669 24055
rect 38703 24021 38715 24055
rect 38657 24015 38715 24021
rect 40037 24055 40095 24061
rect 40037 24021 40049 24055
rect 40083 24021 40095 24055
rect 40037 24015 40095 24021
rect 40402 24012 40408 24064
rect 40460 24012 40466 24064
rect 41138 24012 41144 24064
rect 41196 24052 41202 24064
rect 41877 24055 41935 24061
rect 41877 24052 41889 24055
rect 41196 24024 41889 24052
rect 41196 24012 41202 24024
rect 41877 24021 41889 24024
rect 41923 24021 41935 24055
rect 41877 24015 41935 24021
rect 43257 24055 43315 24061
rect 43257 24021 43269 24055
rect 43303 24052 43315 24055
rect 43714 24052 43720 24064
rect 43303 24024 43720 24052
rect 43303 24021 43315 24024
rect 43257 24015 43315 24021
rect 43714 24012 43720 24024
rect 43772 24012 43778 24064
rect 43806 24012 43812 24064
rect 43864 24052 43870 24064
rect 46400 24052 46428 24228
rect 46937 24225 46949 24228
rect 46983 24225 46995 24259
rect 46937 24219 46995 24225
rect 48774 24216 48780 24268
rect 48832 24216 48838 24268
rect 48501 24191 48559 24197
rect 48501 24188 48513 24191
rect 48332 24160 48513 24188
rect 46842 24080 46848 24132
rect 46900 24120 46906 24132
rect 47857 24123 47915 24129
rect 47857 24120 47869 24123
rect 46900 24092 47869 24120
rect 46900 24080 46906 24092
rect 47857 24089 47869 24092
rect 47903 24089 47915 24123
rect 47857 24083 47915 24089
rect 43864 24024 46428 24052
rect 43864 24012 43870 24024
rect 46658 24012 46664 24064
rect 46716 24052 46722 24064
rect 48332 24061 48360 24160
rect 48501 24157 48513 24160
rect 48547 24157 48559 24191
rect 48501 24151 48559 24157
rect 48317 24055 48375 24061
rect 48317 24052 48329 24055
rect 46716 24024 48329 24052
rect 46716 24012 46722 24024
rect 48317 24021 48329 24024
rect 48363 24021 48375 24055
rect 48317 24015 48375 24021
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 2314 23808 2320 23860
rect 2372 23808 2378 23860
rect 3602 23808 3608 23860
rect 3660 23848 3666 23860
rect 3660 23820 4292 23848
rect 3660 23808 3666 23820
rect 3973 23783 4031 23789
rect 3973 23749 3985 23783
rect 4019 23780 4031 23783
rect 4154 23780 4160 23792
rect 4019 23752 4160 23780
rect 4019 23749 4031 23752
rect 3973 23743 4031 23749
rect 4154 23740 4160 23752
rect 4212 23740 4218 23792
rect 4264 23780 4292 23820
rect 6454 23808 6460 23860
rect 6512 23848 6518 23860
rect 18782 23848 18788 23860
rect 6512 23820 18788 23848
rect 6512 23808 6518 23820
rect 18782 23808 18788 23820
rect 18840 23808 18846 23860
rect 18892 23820 21220 23848
rect 8754 23780 8760 23792
rect 4264 23752 8760 23780
rect 8754 23740 8760 23752
rect 8812 23740 8818 23792
rect 9122 23740 9128 23792
rect 9180 23740 9186 23792
rect 10686 23740 10692 23792
rect 10744 23740 10750 23792
rect 14277 23783 14335 23789
rect 14277 23749 14289 23783
rect 14323 23780 14335 23783
rect 15102 23780 15108 23792
rect 14323 23752 15108 23780
rect 14323 23749 14335 23752
rect 14277 23743 14335 23749
rect 15102 23740 15108 23752
rect 15160 23740 15166 23792
rect 16117 23783 16175 23789
rect 16117 23749 16129 23783
rect 16163 23780 16175 23783
rect 17034 23780 17040 23792
rect 16163 23752 17040 23780
rect 16163 23749 16175 23752
rect 16117 23743 16175 23749
rect 17034 23740 17040 23752
rect 17092 23740 17098 23792
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23681 1731 23715
rect 1673 23675 1731 23681
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23712 3019 23715
rect 3878 23712 3884 23724
rect 3007 23684 3884 23712
rect 3007 23681 3019 23684
rect 2961 23675 3019 23681
rect 1688 23644 1716 23675
rect 3878 23672 3884 23684
rect 3936 23672 3942 23724
rect 4798 23672 4804 23724
rect 4856 23672 4862 23724
rect 6457 23715 6515 23721
rect 6457 23681 6469 23715
rect 6503 23712 6515 23715
rect 6546 23712 6552 23724
rect 6503 23684 6552 23712
rect 6503 23681 6515 23684
rect 6457 23675 6515 23681
rect 6546 23672 6552 23684
rect 6604 23672 6610 23724
rect 8113 23715 8171 23721
rect 8113 23681 8125 23715
rect 8159 23712 8171 23715
rect 9214 23712 9220 23724
rect 8159 23684 9220 23712
rect 8159 23681 8171 23684
rect 8113 23675 8171 23681
rect 9214 23672 9220 23684
rect 9272 23672 9278 23724
rect 9953 23715 10011 23721
rect 9953 23681 9965 23715
rect 9999 23681 10011 23715
rect 9953 23675 10011 23681
rect 4154 23644 4160 23656
rect 1688 23616 4160 23644
rect 4154 23604 4160 23616
rect 4212 23604 4218 23656
rect 5442 23604 5448 23656
rect 5500 23604 5506 23656
rect 6825 23647 6883 23653
rect 6825 23613 6837 23647
rect 6871 23644 6883 23647
rect 6914 23644 6920 23656
rect 6871 23616 6920 23644
rect 6871 23613 6883 23616
rect 6825 23607 6883 23613
rect 6914 23604 6920 23616
rect 6972 23604 6978 23656
rect 3694 23536 3700 23588
rect 3752 23576 3758 23588
rect 5626 23576 5632 23588
rect 3752 23548 5632 23576
rect 3752 23536 3758 23548
rect 5626 23536 5632 23548
rect 5684 23536 5690 23588
rect 9968 23576 9996 23675
rect 11790 23672 11796 23724
rect 11848 23672 11854 23724
rect 12066 23672 12072 23724
rect 12124 23672 12130 23724
rect 13265 23715 13323 23721
rect 13265 23681 13277 23715
rect 13311 23712 13323 23715
rect 14642 23712 14648 23724
rect 13311 23684 14648 23712
rect 13311 23681 13323 23684
rect 13265 23675 13323 23681
rect 14642 23672 14648 23684
rect 14700 23672 14706 23724
rect 15010 23672 15016 23724
rect 15068 23672 15074 23724
rect 16850 23672 16856 23724
rect 16908 23672 16914 23724
rect 17310 23672 17316 23724
rect 17368 23672 17374 23724
rect 17865 23715 17923 23721
rect 17865 23681 17877 23715
rect 17911 23712 17923 23715
rect 18892 23712 18920 23820
rect 18966 23740 18972 23792
rect 19024 23740 19030 23792
rect 19889 23783 19947 23789
rect 19889 23780 19901 23783
rect 19306 23752 19901 23780
rect 19306 23712 19334 23752
rect 19889 23749 19901 23752
rect 19935 23749 19947 23783
rect 19889 23743 19947 23749
rect 19978 23740 19984 23792
rect 20036 23780 20042 23792
rect 20036 23752 20378 23780
rect 20036 23740 20042 23752
rect 17911 23684 18920 23712
rect 18984 23684 19334 23712
rect 21192 23712 21220 23820
rect 21358 23808 21364 23860
rect 21416 23848 21422 23860
rect 23842 23848 23848 23860
rect 21416 23820 23848 23848
rect 21416 23808 21422 23820
rect 23842 23808 23848 23820
rect 23900 23808 23906 23860
rect 24946 23848 24952 23860
rect 24044 23820 24952 23848
rect 22189 23715 22247 23721
rect 21192 23684 22094 23712
rect 17911 23681 17923 23684
rect 17865 23675 17923 23681
rect 11422 23604 11428 23656
rect 11480 23644 11486 23656
rect 18984 23644 19012 23684
rect 11480 23616 19012 23644
rect 11480 23604 11486 23616
rect 19242 23604 19248 23656
rect 19300 23644 19306 23656
rect 19613 23647 19671 23653
rect 19613 23644 19625 23647
rect 19300 23616 19625 23644
rect 19300 23604 19306 23616
rect 19613 23613 19625 23616
rect 19659 23644 19671 23647
rect 21174 23644 21180 23656
rect 19659 23616 21180 23644
rect 19659 23613 19671 23616
rect 19613 23607 19671 23613
rect 21174 23604 21180 23616
rect 21232 23604 21238 23656
rect 16666 23576 16672 23588
rect 9968 23548 16672 23576
rect 16666 23536 16672 23548
rect 16724 23536 16730 23588
rect 16758 23536 16764 23588
rect 16816 23576 16822 23588
rect 19518 23576 19524 23588
rect 16816 23548 19524 23576
rect 16816 23536 16822 23548
rect 19518 23536 19524 23548
rect 19576 23536 19582 23588
rect 22066 23576 22094 23684
rect 22189 23681 22201 23715
rect 22235 23712 22247 23715
rect 23198 23712 23204 23724
rect 22235 23684 23204 23712
rect 22235 23681 22247 23684
rect 22189 23675 22247 23681
rect 23198 23672 23204 23684
rect 23256 23672 23262 23724
rect 22462 23604 22468 23656
rect 22520 23604 22526 23656
rect 23753 23647 23811 23653
rect 23753 23613 23765 23647
rect 23799 23644 23811 23647
rect 24044 23644 24072 23820
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 25038 23808 25044 23860
rect 25096 23848 25102 23860
rect 27617 23851 27675 23857
rect 27617 23848 27629 23851
rect 25096 23820 27629 23848
rect 25096 23808 25102 23820
rect 27617 23817 27629 23820
rect 27663 23817 27675 23851
rect 27617 23811 27675 23817
rect 27890 23808 27896 23860
rect 27948 23848 27954 23860
rect 30285 23851 30343 23857
rect 30285 23848 30297 23851
rect 27948 23820 30297 23848
rect 27948 23808 27954 23820
rect 30285 23817 30297 23820
rect 30331 23817 30343 23851
rect 30285 23811 30343 23817
rect 30650 23808 30656 23860
rect 30708 23808 30714 23860
rect 31386 23808 31392 23860
rect 31444 23848 31450 23860
rect 35345 23851 35403 23857
rect 35345 23848 35357 23851
rect 31444 23820 35357 23848
rect 31444 23808 31450 23820
rect 35345 23817 35357 23820
rect 35391 23817 35403 23851
rect 35345 23811 35403 23817
rect 35989 23851 36047 23857
rect 35989 23817 36001 23851
rect 36035 23848 36047 23851
rect 36538 23848 36544 23860
rect 36035 23820 36544 23848
rect 36035 23817 36047 23820
rect 35989 23811 36047 23817
rect 36538 23808 36544 23820
rect 36596 23808 36602 23860
rect 37826 23808 37832 23860
rect 37884 23808 37890 23860
rect 37918 23808 37924 23860
rect 37976 23848 37982 23860
rect 40037 23851 40095 23857
rect 40037 23848 40049 23851
rect 37976 23820 40049 23848
rect 37976 23808 37982 23820
rect 40037 23817 40049 23820
rect 40083 23817 40095 23851
rect 40037 23811 40095 23817
rect 41874 23808 41880 23860
rect 41932 23808 41938 23860
rect 42242 23808 42248 23860
rect 42300 23848 42306 23860
rect 42300 23820 42840 23848
rect 42300 23808 42306 23820
rect 25133 23783 25191 23789
rect 25133 23780 25145 23783
rect 23799 23616 24072 23644
rect 24136 23752 25145 23780
rect 23799 23613 23811 23616
rect 23753 23607 23811 23613
rect 22646 23576 22652 23588
rect 22066 23548 22652 23576
rect 22646 23536 22652 23548
rect 22704 23536 22710 23588
rect 2774 23468 2780 23520
rect 2832 23508 2838 23520
rect 6178 23508 6184 23520
rect 2832 23480 6184 23508
rect 2832 23468 2838 23480
rect 6178 23468 6184 23480
rect 6236 23468 6242 23520
rect 10778 23468 10784 23520
rect 10836 23508 10842 23520
rect 12526 23508 12532 23520
rect 10836 23480 12532 23508
rect 10836 23468 10842 23480
rect 12526 23468 12532 23480
rect 12584 23468 12590 23520
rect 17129 23511 17187 23517
rect 17129 23477 17141 23511
rect 17175 23508 17187 23511
rect 17494 23508 17500 23520
rect 17175 23480 17500 23508
rect 17175 23477 17187 23480
rect 17129 23471 17187 23477
rect 17494 23468 17500 23480
rect 17552 23468 17558 23520
rect 21358 23468 21364 23520
rect 21416 23468 21422 23520
rect 23566 23468 23572 23520
rect 23624 23508 23630 23520
rect 24136 23508 24164 23752
rect 25133 23749 25145 23752
rect 25179 23749 25191 23783
rect 26418 23780 26424 23792
rect 26358 23752 26424 23780
rect 25133 23743 25191 23749
rect 26418 23740 26424 23752
rect 26476 23740 26482 23792
rect 27522 23740 27528 23792
rect 27580 23780 27586 23792
rect 29457 23783 29515 23789
rect 29457 23780 29469 23783
rect 27580 23752 29469 23780
rect 27580 23740 27586 23752
rect 29457 23749 29469 23752
rect 29503 23749 29515 23783
rect 29457 23743 29515 23749
rect 31754 23740 31760 23792
rect 31812 23740 31818 23792
rect 32674 23740 32680 23792
rect 32732 23780 32738 23792
rect 33597 23783 33655 23789
rect 33597 23780 33609 23783
rect 32732 23752 33609 23780
rect 32732 23740 32738 23752
rect 33597 23749 33609 23752
rect 33643 23749 33655 23783
rect 33597 23743 33655 23749
rect 34054 23740 34060 23792
rect 34112 23740 34118 23792
rect 37737 23783 37795 23789
rect 37737 23749 37749 23783
rect 37783 23780 37795 23783
rect 37844 23780 37872 23808
rect 42812 23780 42840 23820
rect 45186 23808 45192 23860
rect 45244 23808 45250 23860
rect 47762 23808 47768 23860
rect 47820 23848 47826 23860
rect 48041 23851 48099 23857
rect 48041 23848 48053 23851
rect 47820 23820 48053 23848
rect 47820 23808 47826 23820
rect 48041 23817 48053 23820
rect 48087 23817 48099 23851
rect 48041 23811 48099 23817
rect 45462 23780 45468 23792
rect 37783 23752 37872 23780
rect 41248 23752 42748 23780
rect 42812 23752 45468 23780
rect 37783 23749 37795 23752
rect 37737 23743 37795 23749
rect 24210 23672 24216 23724
rect 24268 23672 24274 23724
rect 27798 23712 27804 23724
rect 27540 23684 27804 23712
rect 24854 23604 24860 23656
rect 24912 23604 24918 23656
rect 27540 23644 27568 23684
rect 27798 23672 27804 23684
rect 27856 23672 27862 23724
rect 27985 23715 28043 23721
rect 27985 23681 27997 23715
rect 28031 23712 28043 23715
rect 28813 23715 28871 23721
rect 28031 23684 28764 23712
rect 28031 23681 28043 23684
rect 27985 23675 28043 23681
rect 26252 23616 27568 23644
rect 23624 23480 24164 23508
rect 24305 23511 24363 23517
rect 23624 23468 23630 23480
rect 24305 23477 24317 23511
rect 24351 23508 24363 23511
rect 26252 23508 26280 23616
rect 27706 23604 27712 23656
rect 27764 23644 27770 23656
rect 28077 23647 28135 23653
rect 28077 23644 28089 23647
rect 27764 23616 28089 23644
rect 27764 23604 27770 23616
rect 28077 23613 28089 23616
rect 28123 23613 28135 23647
rect 28077 23607 28135 23613
rect 28261 23647 28319 23653
rect 28261 23613 28273 23647
rect 28307 23644 28319 23647
rect 28350 23644 28356 23656
rect 28307 23616 28356 23644
rect 28307 23613 28319 23616
rect 28261 23607 28319 23613
rect 28350 23604 28356 23616
rect 28408 23604 28414 23656
rect 28736 23644 28764 23684
rect 28813 23681 28825 23715
rect 28859 23712 28871 23715
rect 30374 23712 30380 23724
rect 28859 23684 30380 23712
rect 28859 23681 28871 23684
rect 28813 23675 28871 23681
rect 30374 23672 30380 23684
rect 30432 23672 30438 23724
rect 30484 23684 30972 23712
rect 30098 23644 30104 23656
rect 28736 23616 30104 23644
rect 30098 23604 30104 23616
rect 30156 23604 30162 23656
rect 26605 23579 26663 23585
rect 26605 23545 26617 23579
rect 26651 23576 26663 23579
rect 30484 23576 30512 23684
rect 30944 23656 30972 23684
rect 31570 23672 31576 23724
rect 31628 23672 31634 23724
rect 32398 23672 32404 23724
rect 32456 23712 32462 23724
rect 32493 23715 32551 23721
rect 32493 23712 32505 23715
rect 32456 23684 32505 23712
rect 32456 23672 32462 23684
rect 32493 23681 32505 23684
rect 32539 23681 32551 23715
rect 32493 23675 32551 23681
rect 33226 23672 33232 23724
rect 33284 23712 33290 23724
rect 33321 23715 33379 23721
rect 33321 23712 33333 23715
rect 33284 23684 33333 23712
rect 33284 23672 33290 23684
rect 33321 23681 33333 23684
rect 33367 23681 33379 23715
rect 33321 23675 33379 23681
rect 35897 23715 35955 23721
rect 35897 23681 35909 23715
rect 35943 23712 35955 23715
rect 36354 23712 36360 23724
rect 35943 23684 36360 23712
rect 35943 23681 35955 23684
rect 35897 23675 35955 23681
rect 36354 23672 36360 23684
rect 36412 23672 36418 23724
rect 38838 23672 38844 23724
rect 38896 23672 38902 23724
rect 39942 23712 39948 23724
rect 39132 23684 39948 23712
rect 30745 23647 30803 23653
rect 30745 23613 30757 23647
rect 30791 23613 30803 23647
rect 30745 23607 30803 23613
rect 26651 23548 28120 23576
rect 26651 23545 26663 23548
rect 26605 23539 26663 23545
rect 24351 23480 26280 23508
rect 24351 23477 24363 23480
rect 24305 23471 24363 23477
rect 26786 23468 26792 23520
rect 26844 23508 26850 23520
rect 26973 23511 27031 23517
rect 26973 23508 26985 23511
rect 26844 23480 26985 23508
rect 26844 23468 26850 23480
rect 26973 23477 26985 23480
rect 27019 23477 27031 23511
rect 26973 23471 27031 23477
rect 27154 23468 27160 23520
rect 27212 23468 27218 23520
rect 28092 23508 28120 23548
rect 28966 23548 30512 23576
rect 30760 23576 30788 23607
rect 30926 23604 30932 23656
rect 30984 23604 30990 23656
rect 33134 23604 33140 23656
rect 33192 23644 33198 23656
rect 34330 23644 34336 23656
rect 33192 23616 34336 23644
rect 33192 23604 33198 23616
rect 34330 23604 34336 23616
rect 34388 23604 34394 23656
rect 35066 23604 35072 23656
rect 35124 23644 35130 23656
rect 35529 23647 35587 23653
rect 35529 23644 35541 23647
rect 35124 23616 35541 23644
rect 35124 23604 35130 23616
rect 35529 23613 35541 23616
rect 35575 23613 35587 23647
rect 35529 23607 35587 23613
rect 36446 23604 36452 23656
rect 36504 23604 36510 23656
rect 36633 23647 36691 23653
rect 36633 23613 36645 23647
rect 36679 23644 36691 23647
rect 37182 23644 37188 23656
rect 36679 23616 37188 23644
rect 36679 23613 36691 23616
rect 36633 23607 36691 23613
rect 37182 23604 37188 23616
rect 37240 23604 37246 23656
rect 37458 23604 37464 23656
rect 37516 23604 37522 23656
rect 39132 23644 39160 23684
rect 39942 23672 39948 23684
rect 40000 23672 40006 23724
rect 40405 23715 40463 23721
rect 40405 23681 40417 23715
rect 40451 23712 40463 23715
rect 41046 23712 41052 23724
rect 40451 23684 41052 23712
rect 40451 23681 40463 23684
rect 40405 23675 40463 23681
rect 41046 23672 41052 23684
rect 41104 23672 41110 23724
rect 41248 23721 41276 23752
rect 41233 23715 41291 23721
rect 41233 23681 41245 23715
rect 41279 23681 41291 23715
rect 41233 23675 41291 23681
rect 42613 23715 42671 23721
rect 42613 23681 42625 23715
rect 42659 23681 42671 23715
rect 42613 23675 42671 23681
rect 37568 23616 39160 23644
rect 39485 23647 39543 23653
rect 33042 23576 33048 23588
rect 30760 23548 33048 23576
rect 28966 23508 28994 23548
rect 33042 23536 33048 23548
rect 33100 23536 33106 23588
rect 34698 23536 34704 23588
rect 34756 23576 34762 23588
rect 35618 23576 35624 23588
rect 34756 23548 35624 23576
rect 34756 23536 34762 23548
rect 35618 23536 35624 23548
rect 35676 23536 35682 23588
rect 37568 23576 37596 23616
rect 39485 23613 39497 23647
rect 39531 23644 39543 23647
rect 39850 23644 39856 23656
rect 39531 23616 39856 23644
rect 39531 23613 39543 23616
rect 39485 23607 39543 23613
rect 39850 23604 39856 23616
rect 39908 23604 39914 23656
rect 40497 23647 40555 23653
rect 40497 23613 40509 23647
rect 40543 23613 40555 23647
rect 40497 23607 40555 23613
rect 35728 23548 37596 23576
rect 40512 23576 40540 23607
rect 40678 23604 40684 23656
rect 40736 23604 40742 23656
rect 40770 23604 40776 23656
rect 40828 23644 40834 23656
rect 42628 23644 42656 23675
rect 40828 23616 42656 23644
rect 42720 23644 42748 23752
rect 45462 23740 45468 23752
rect 45520 23740 45526 23792
rect 46937 23783 46995 23789
rect 46937 23749 46949 23783
rect 46983 23780 46995 23783
rect 46983 23752 48728 23780
rect 46983 23749 46995 23752
rect 46937 23743 46995 23749
rect 43714 23672 43720 23724
rect 43772 23672 43778 23724
rect 44358 23672 44364 23724
rect 44416 23672 44422 23724
rect 44542 23672 44548 23724
rect 44600 23712 44606 23724
rect 44637 23715 44695 23721
rect 44637 23712 44649 23715
rect 44600 23684 44649 23712
rect 44600 23672 44606 23684
rect 44637 23681 44649 23684
rect 44683 23712 44695 23715
rect 44726 23712 44732 23724
rect 44683 23684 44732 23712
rect 44683 23681 44695 23684
rect 44637 23675 44695 23681
rect 44726 23672 44732 23684
rect 44784 23672 44790 23724
rect 45097 23715 45155 23721
rect 45097 23712 45109 23715
rect 44836 23684 45109 23712
rect 43257 23647 43315 23653
rect 43257 23644 43269 23647
rect 42720 23616 43269 23644
rect 40828 23604 40834 23616
rect 43257 23613 43269 23616
rect 43303 23613 43315 23647
rect 43257 23607 43315 23613
rect 41230 23576 41236 23588
rect 40512 23548 41236 23576
rect 28092 23480 28994 23508
rect 29730 23468 29736 23520
rect 29788 23468 29794 23520
rect 30006 23468 30012 23520
rect 30064 23468 30070 23520
rect 30374 23468 30380 23520
rect 30432 23508 30438 23520
rect 30834 23508 30840 23520
rect 30432 23480 30840 23508
rect 30432 23468 30438 23480
rect 30834 23468 30840 23480
rect 30892 23468 30898 23520
rect 32766 23468 32772 23520
rect 32824 23468 32830 23520
rect 33226 23468 33232 23520
rect 33284 23508 33290 23520
rect 34882 23508 34888 23520
rect 33284 23480 34888 23508
rect 33284 23468 33290 23480
rect 34882 23468 34888 23480
rect 34940 23468 34946 23520
rect 34974 23468 34980 23520
rect 35032 23508 35038 23520
rect 35069 23511 35127 23517
rect 35069 23508 35081 23511
rect 35032 23480 35081 23508
rect 35032 23468 35038 23480
rect 35069 23477 35081 23480
rect 35115 23508 35127 23511
rect 35728 23508 35756 23548
rect 41230 23536 41236 23548
rect 41288 23536 41294 23588
rect 44836 23585 44864 23684
rect 45097 23681 45109 23684
rect 45143 23681 45155 23715
rect 45097 23675 45155 23681
rect 45554 23672 45560 23724
rect 45612 23712 45618 23724
rect 46017 23715 46075 23721
rect 46017 23712 46029 23715
rect 45612 23684 46029 23712
rect 45612 23672 45618 23684
rect 46017 23681 46029 23684
rect 46063 23681 46075 23715
rect 46017 23675 46075 23681
rect 47210 23672 47216 23724
rect 47268 23672 47274 23724
rect 48700 23721 48728 23752
rect 47857 23715 47915 23721
rect 47857 23712 47869 23715
rect 47688 23684 47869 23712
rect 45738 23604 45744 23656
rect 45796 23604 45802 23656
rect 44821 23579 44879 23585
rect 44821 23576 44833 23579
rect 43824 23548 44833 23576
rect 35115 23480 35756 23508
rect 35115 23477 35127 23480
rect 35069 23471 35127 23477
rect 36906 23468 36912 23520
rect 36964 23508 36970 23520
rect 37001 23511 37059 23517
rect 37001 23508 37013 23511
rect 36964 23480 37013 23508
rect 36964 23468 36970 23480
rect 37001 23477 37013 23480
rect 37047 23477 37059 23511
rect 37001 23471 37059 23477
rect 37274 23468 37280 23520
rect 37332 23508 37338 23520
rect 40770 23508 40776 23520
rect 37332 23480 40776 23508
rect 37332 23468 37338 23480
rect 40770 23468 40776 23480
rect 40828 23468 40834 23520
rect 42702 23468 42708 23520
rect 42760 23508 42766 23520
rect 43824 23508 43852 23548
rect 44821 23545 44833 23548
rect 44867 23545 44879 23579
rect 44821 23539 44879 23545
rect 47121 23579 47179 23585
rect 47121 23545 47133 23579
rect 47167 23576 47179 23579
rect 47578 23576 47584 23588
rect 47167 23548 47584 23576
rect 47167 23545 47179 23548
rect 47121 23539 47179 23545
rect 47578 23536 47584 23548
rect 47636 23536 47642 23588
rect 42760 23480 43852 23508
rect 42760 23468 42766 23480
rect 47394 23468 47400 23520
rect 47452 23508 47458 23520
rect 47688 23517 47716 23684
rect 47857 23681 47869 23684
rect 47903 23681 47915 23715
rect 47857 23675 47915 23681
rect 48685 23715 48743 23721
rect 48685 23681 48697 23715
rect 48731 23712 48743 23715
rect 49142 23712 49148 23724
rect 48731 23684 49148 23712
rect 48731 23681 48743 23684
rect 48685 23675 48743 23681
rect 49142 23672 49148 23684
rect 49200 23672 49206 23724
rect 47762 23604 47768 23656
rect 47820 23644 47826 23656
rect 48961 23647 49019 23653
rect 48961 23644 48973 23647
rect 47820 23616 48973 23644
rect 47820 23604 47826 23616
rect 48961 23613 48973 23616
rect 49007 23613 49019 23647
rect 48961 23607 49019 23613
rect 47673 23511 47731 23517
rect 47673 23508 47685 23511
rect 47452 23480 47685 23508
rect 47452 23468 47458 23480
rect 47673 23477 47685 23480
rect 47719 23477 47731 23511
rect 47673 23471 47731 23477
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 3605 23307 3663 23313
rect 3605 23273 3617 23307
rect 3651 23304 3663 23307
rect 14550 23304 14556 23316
rect 3651 23276 14556 23304
rect 3651 23273 3663 23276
rect 3605 23267 3663 23273
rect 14550 23264 14556 23276
rect 14608 23264 14614 23316
rect 14642 23264 14648 23316
rect 14700 23264 14706 23316
rect 14734 23264 14740 23316
rect 14792 23304 14798 23316
rect 17218 23304 17224 23316
rect 14792 23276 17224 23304
rect 14792 23264 14798 23276
rect 17218 23264 17224 23276
rect 17276 23264 17282 23316
rect 17862 23264 17868 23316
rect 17920 23304 17926 23316
rect 17920 23276 19334 23304
rect 17920 23264 17926 23276
rect 3418 23196 3424 23248
rect 3476 23196 3482 23248
rect 3973 23239 4031 23245
rect 3973 23205 3985 23239
rect 4019 23236 4031 23239
rect 4798 23236 4804 23248
rect 4019 23208 4804 23236
rect 4019 23205 4031 23208
rect 3973 23199 4031 23205
rect 4798 23196 4804 23208
rect 4856 23236 4862 23248
rect 17034 23236 17040 23248
rect 4856 23208 12434 23236
rect 4856 23196 4862 23208
rect 2866 23128 2872 23180
rect 2924 23168 2930 23180
rect 4430 23168 4436 23180
rect 2924 23140 4436 23168
rect 2924 23128 2930 23140
rect 4430 23128 4436 23140
rect 4488 23128 4494 23180
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 11238 23128 11244 23180
rect 11296 23128 11302 23180
rect 1762 23060 1768 23112
rect 1820 23060 1826 23112
rect 4246 23060 4252 23112
rect 4304 23060 4310 23112
rect 4338 23060 4344 23112
rect 4396 23100 4402 23112
rect 5353 23103 5411 23109
rect 5353 23100 5365 23103
rect 4396 23072 5365 23100
rect 4396 23060 4402 23072
rect 5353 23069 5365 23072
rect 5399 23069 5411 23103
rect 5353 23063 5411 23069
rect 7377 23103 7435 23109
rect 7377 23069 7389 23103
rect 7423 23100 7435 23103
rect 7466 23100 7472 23112
rect 7423 23072 7472 23100
rect 7423 23069 7435 23072
rect 7377 23063 7435 23069
rect 7466 23060 7472 23072
rect 7524 23060 7530 23112
rect 8294 23060 8300 23112
rect 8352 23100 8358 23112
rect 9401 23103 9459 23109
rect 9401 23100 9413 23103
rect 8352 23072 9413 23100
rect 8352 23060 8358 23072
rect 9401 23069 9413 23072
rect 9447 23069 9459 23103
rect 9401 23063 9459 23069
rect 10502 23060 10508 23112
rect 10560 23060 10566 23112
rect 2774 22992 2780 23044
rect 2832 22992 2838 23044
rect 3234 22992 3240 23044
rect 3292 23032 3298 23044
rect 6730 23032 6736 23044
rect 3292 23004 6736 23032
rect 3292 22992 3298 23004
rect 6730 22992 6736 23004
rect 6788 22992 6794 23044
rect 9125 23035 9183 23041
rect 9125 23001 9137 23035
rect 9171 23032 9183 23035
rect 12406 23032 12434 23208
rect 14108 23208 17040 23236
rect 13354 23128 13360 23180
rect 13412 23128 13418 23180
rect 12529 23103 12587 23109
rect 12529 23069 12541 23103
rect 12575 23100 12587 23103
rect 14108 23100 14136 23208
rect 17034 23196 17040 23208
rect 17092 23196 17098 23248
rect 14185 23171 14243 23177
rect 14185 23137 14197 23171
rect 14231 23168 14243 23171
rect 15746 23168 15752 23180
rect 14231 23140 15752 23168
rect 14231 23137 14243 23140
rect 14185 23131 14243 23137
rect 15746 23128 15752 23140
rect 15804 23128 15810 23180
rect 16390 23128 16396 23180
rect 16448 23128 16454 23180
rect 16758 23128 16764 23180
rect 16816 23168 16822 23180
rect 16816 23140 18736 23168
rect 16816 23128 16822 23140
rect 12575 23072 14136 23100
rect 12575 23069 12587 23072
rect 12529 23063 12587 23069
rect 14550 23060 14556 23112
rect 14608 23100 14614 23112
rect 14829 23103 14887 23109
rect 14829 23100 14841 23103
rect 14608 23072 14841 23100
rect 14608 23060 14614 23072
rect 14829 23069 14841 23072
rect 14875 23069 14887 23103
rect 14829 23063 14887 23069
rect 15473 23103 15531 23109
rect 15473 23069 15485 23103
rect 15519 23100 15531 23103
rect 16574 23100 16580 23112
rect 15519 23072 16580 23100
rect 15519 23069 15531 23072
rect 15473 23063 15531 23069
rect 16574 23060 16580 23072
rect 16632 23060 16638 23112
rect 17126 23060 17132 23112
rect 17184 23060 17190 23112
rect 18506 23060 18512 23112
rect 18564 23060 18570 23112
rect 17405 23035 17463 23041
rect 17405 23032 17417 23035
rect 9171 23004 11560 23032
rect 12406 23004 17417 23032
rect 9171 23001 9183 23004
rect 9125 22995 9183 23001
rect 4893 22967 4951 22973
rect 4893 22933 4905 22967
rect 4939 22964 4951 22967
rect 7742 22964 7748 22976
rect 4939 22936 7748 22964
rect 4939 22933 4951 22936
rect 4893 22927 4951 22933
rect 7742 22924 7748 22936
rect 7800 22924 7806 22976
rect 9674 22924 9680 22976
rect 9732 22964 9738 22976
rect 10045 22967 10103 22973
rect 10045 22964 10057 22967
rect 9732 22936 10057 22964
rect 9732 22924 9738 22936
rect 10045 22933 10057 22936
rect 10091 22933 10103 22967
rect 11532 22964 11560 23004
rect 17405 23001 17417 23004
rect 17451 23001 17463 23035
rect 18708 23032 18736 23140
rect 19306 23100 19334 23276
rect 20254 23264 20260 23316
rect 20312 23304 20318 23316
rect 22462 23304 22468 23316
rect 20312 23276 22468 23304
rect 20312 23264 20318 23276
rect 22462 23264 22468 23276
rect 22520 23264 22526 23316
rect 22646 23264 22652 23316
rect 22704 23304 22710 23316
rect 24765 23307 24823 23313
rect 24765 23304 24777 23307
rect 22704 23276 24777 23304
rect 22704 23264 22710 23276
rect 24765 23273 24777 23276
rect 24811 23273 24823 23307
rect 24765 23267 24823 23273
rect 26050 23264 26056 23316
rect 26108 23304 26114 23316
rect 29270 23304 29276 23316
rect 26108 23276 29276 23304
rect 26108 23264 26114 23276
rect 29270 23264 29276 23276
rect 29328 23264 29334 23316
rect 30926 23264 30932 23316
rect 30984 23304 30990 23316
rect 36814 23304 36820 23316
rect 30984 23276 36820 23304
rect 30984 23264 30990 23276
rect 24118 23196 24124 23248
rect 24176 23236 24182 23248
rect 24486 23236 24492 23248
rect 24176 23208 24492 23236
rect 24176 23196 24182 23208
rect 24486 23196 24492 23208
rect 24544 23196 24550 23248
rect 26694 23196 26700 23248
rect 26752 23236 26758 23248
rect 26752 23208 27384 23236
rect 26752 23196 26758 23208
rect 20809 23171 20867 23177
rect 20809 23137 20821 23171
rect 20855 23168 20867 23171
rect 21174 23168 21180 23180
rect 20855 23140 21180 23168
rect 20855 23137 20867 23140
rect 20809 23131 20867 23137
rect 21174 23128 21180 23140
rect 21232 23128 21238 23180
rect 22370 23128 22376 23180
rect 22428 23168 22434 23180
rect 23661 23171 23719 23177
rect 23661 23168 23673 23171
rect 22428 23140 23673 23168
rect 22428 23128 22434 23140
rect 23661 23137 23673 23140
rect 23707 23168 23719 23171
rect 23934 23168 23940 23180
rect 23707 23140 23940 23168
rect 23707 23137 23719 23140
rect 23661 23131 23719 23137
rect 23934 23128 23940 23140
rect 23992 23128 23998 23180
rect 25685 23171 25743 23177
rect 25685 23137 25697 23171
rect 25731 23168 25743 23171
rect 27246 23168 27252 23180
rect 25731 23140 27252 23168
rect 25731 23137 25743 23140
rect 25685 23131 25743 23137
rect 27246 23128 27252 23140
rect 27304 23128 27310 23180
rect 27356 23168 27384 23208
rect 27614 23196 27620 23248
rect 27672 23236 27678 23248
rect 28810 23236 28816 23248
rect 27672 23208 28816 23236
rect 27672 23196 27678 23208
rect 28810 23196 28816 23208
rect 28868 23196 28874 23248
rect 31680 23245 31708 23276
rect 36814 23264 36820 23276
rect 36872 23264 36878 23316
rect 37001 23307 37059 23313
rect 37001 23273 37013 23307
rect 37047 23304 37059 23307
rect 37356 23307 37414 23313
rect 37356 23304 37368 23307
rect 37047 23276 37368 23304
rect 37047 23273 37059 23276
rect 37001 23267 37059 23273
rect 37356 23273 37368 23276
rect 37402 23304 37414 23307
rect 39025 23307 39083 23313
rect 39025 23304 39037 23307
rect 37402 23276 39037 23304
rect 37402 23273 37414 23276
rect 37356 23267 37414 23273
rect 39025 23273 39037 23276
rect 39071 23304 39083 23307
rect 42334 23304 42340 23316
rect 39071 23276 42340 23304
rect 39071 23273 39083 23276
rect 39025 23267 39083 23273
rect 42334 23264 42340 23276
rect 42392 23264 42398 23316
rect 44174 23264 44180 23316
rect 44232 23304 44238 23316
rect 44361 23307 44419 23313
rect 44361 23304 44373 23307
rect 44232 23276 44373 23304
rect 44232 23264 44238 23276
rect 44361 23273 44373 23276
rect 44407 23273 44419 23307
rect 44361 23267 44419 23273
rect 45833 23307 45891 23313
rect 45833 23273 45845 23307
rect 45879 23304 45891 23307
rect 46290 23304 46296 23316
rect 45879 23276 46296 23304
rect 45879 23273 45891 23276
rect 45833 23267 45891 23273
rect 46290 23264 46296 23276
rect 46348 23264 46354 23316
rect 46382 23264 46388 23316
rect 46440 23304 46446 23316
rect 47302 23304 47308 23316
rect 46440 23276 47308 23304
rect 46440 23264 46446 23276
rect 47302 23264 47308 23276
rect 47360 23264 47366 23316
rect 47854 23264 47860 23316
rect 47912 23304 47918 23316
rect 48774 23304 48780 23316
rect 47912 23276 48780 23304
rect 47912 23264 47918 23276
rect 48774 23264 48780 23276
rect 48832 23264 48838 23316
rect 31665 23239 31723 23245
rect 31665 23205 31677 23239
rect 31711 23236 31723 23239
rect 34054 23236 34060 23248
rect 31711 23208 31745 23236
rect 33520 23208 34060 23236
rect 31711 23205 31723 23208
rect 31665 23199 31723 23205
rect 27890 23168 27896 23180
rect 27356 23140 27896 23168
rect 27890 23128 27896 23140
rect 27948 23128 27954 23180
rect 28261 23171 28319 23177
rect 28261 23137 28273 23171
rect 28307 23168 28319 23171
rect 28442 23168 28448 23180
rect 28307 23140 28448 23168
rect 28307 23137 28319 23140
rect 28261 23131 28319 23137
rect 28442 23128 28448 23140
rect 28500 23128 28506 23180
rect 29086 23128 29092 23180
rect 29144 23128 29150 23180
rect 32125 23171 32183 23177
rect 32125 23168 32137 23171
rect 29932 23140 32137 23168
rect 20165 23103 20223 23109
rect 20165 23100 20177 23103
rect 19306 23072 20177 23100
rect 20165 23069 20177 23072
rect 20211 23069 20223 23103
rect 20165 23063 20223 23069
rect 22922 23060 22928 23112
rect 22980 23100 22986 23112
rect 23385 23103 23443 23109
rect 23385 23100 23397 23103
rect 22980 23072 23397 23100
rect 22980 23060 22986 23072
rect 23385 23069 23397 23072
rect 23431 23069 23443 23103
rect 23385 23063 23443 23069
rect 24762 23060 24768 23112
rect 24820 23100 24826 23112
rect 25409 23103 25467 23109
rect 25409 23100 25421 23103
rect 24820 23072 25421 23100
rect 24820 23060 24826 23072
rect 25409 23069 25421 23072
rect 25455 23069 25467 23103
rect 25409 23063 25467 23069
rect 28074 23060 28080 23112
rect 28132 23100 28138 23112
rect 28534 23100 28540 23112
rect 28132 23072 28540 23100
rect 28132 23060 28138 23072
rect 28534 23060 28540 23072
rect 28592 23060 28598 23112
rect 28626 23060 28632 23112
rect 28684 23100 28690 23112
rect 29932 23109 29960 23140
rect 32125 23137 32137 23140
rect 32171 23168 32183 23171
rect 33410 23168 33416 23180
rect 32171 23140 33416 23168
rect 32171 23137 32183 23140
rect 32125 23131 32183 23137
rect 33410 23128 33416 23140
rect 33468 23128 33474 23180
rect 29917 23103 29975 23109
rect 29917 23100 29929 23103
rect 28684 23072 29929 23100
rect 28684 23060 28690 23072
rect 29917 23069 29929 23072
rect 29963 23069 29975 23103
rect 29917 23063 29975 23069
rect 19429 23035 19487 23041
rect 19429 23032 19441 23035
rect 18708 23004 19441 23032
rect 17405 22995 17463 23001
rect 19429 23001 19441 23004
rect 19475 23032 19487 23035
rect 20806 23032 20812 23044
rect 19475 23004 20812 23032
rect 19475 23001 19487 23004
rect 19429 22995 19487 23001
rect 20806 22992 20812 23004
rect 20864 22992 20870 23044
rect 21082 22992 21088 23044
rect 21140 22992 21146 23044
rect 21468 23004 21574 23032
rect 14369 22967 14427 22973
rect 14369 22964 14381 22967
rect 11532 22936 14381 22964
rect 10045 22927 10103 22933
rect 14369 22933 14381 22936
rect 14415 22964 14427 22967
rect 16758 22964 16764 22976
rect 14415 22936 16764 22964
rect 14415 22933 14427 22936
rect 14369 22927 14427 22933
rect 16758 22924 16764 22936
rect 16816 22924 16822 22976
rect 18322 22924 18328 22976
rect 18380 22964 18386 22976
rect 18877 22967 18935 22973
rect 18877 22964 18889 22967
rect 18380 22936 18889 22964
rect 18380 22924 18386 22936
rect 18877 22933 18889 22936
rect 18923 22933 18935 22967
rect 18877 22927 18935 22933
rect 19978 22924 19984 22976
rect 20036 22964 20042 22976
rect 21468 22964 21496 23004
rect 22738 22992 22744 23044
rect 22796 23032 22802 23044
rect 22833 23035 22891 23041
rect 22833 23032 22845 23035
rect 22796 23004 22845 23032
rect 22796 22992 22802 23004
rect 22833 23001 22845 23004
rect 22879 23001 22891 23035
rect 22833 22995 22891 23001
rect 24673 23035 24731 23041
rect 24673 23001 24685 23035
rect 24719 23032 24731 23035
rect 25314 23032 25320 23044
rect 24719 23004 25320 23032
rect 24719 23001 24731 23004
rect 24673 22995 24731 23001
rect 25314 22992 25320 23004
rect 25372 22992 25378 23044
rect 27338 23032 27344 23044
rect 26910 23004 27344 23032
rect 27338 22992 27344 23004
rect 27396 22992 27402 23044
rect 27985 23035 28043 23041
rect 27985 23001 27997 23035
rect 28031 23032 28043 23035
rect 28031 23004 28856 23032
rect 28031 23001 28043 23004
rect 27985 22995 28043 23001
rect 20036 22936 21496 22964
rect 20036 22924 20042 22936
rect 26510 22924 26516 22976
rect 26568 22964 26574 22976
rect 27154 22964 27160 22976
rect 26568 22936 27160 22964
rect 26568 22924 26574 22936
rect 27154 22924 27160 22936
rect 27212 22924 27218 22976
rect 27614 22924 27620 22976
rect 27672 22924 27678 22976
rect 28828 22964 28856 23004
rect 28902 22992 28908 23044
rect 28960 22992 28966 23044
rect 29564 23004 30144 23032
rect 29564 22964 29592 23004
rect 28828 22936 29592 22964
rect 29638 22924 29644 22976
rect 29696 22924 29702 22976
rect 30116 22964 30144 23004
rect 30190 22992 30196 23044
rect 30248 22992 30254 23044
rect 32401 23035 32459 23041
rect 31418 23004 31524 23032
rect 30834 22964 30840 22976
rect 30116 22936 30840 22964
rect 30834 22924 30840 22936
rect 30892 22924 30898 22976
rect 31496 22964 31524 23004
rect 32401 23001 32413 23035
rect 32447 23032 32459 23035
rect 32674 23032 32680 23044
rect 32447 23004 32680 23032
rect 32447 23001 32459 23004
rect 32401 22995 32459 23001
rect 32674 22992 32680 23004
rect 32732 22992 32738 23044
rect 31754 22964 31760 22976
rect 31496 22936 31760 22964
rect 31754 22924 31760 22936
rect 31812 22964 31818 22976
rect 32766 22964 32772 22976
rect 31812 22936 32772 22964
rect 31812 22924 31818 22936
rect 32766 22924 32772 22936
rect 32824 22964 32830 22976
rect 33318 22964 33324 22976
rect 32824 22936 33324 22964
rect 32824 22924 32830 22936
rect 33318 22924 33324 22936
rect 33376 22964 33382 22976
rect 33520 22964 33548 23208
rect 34054 23196 34060 23208
rect 34112 23196 34118 23248
rect 34146 23196 34152 23248
rect 34204 23236 34210 23248
rect 34241 23239 34299 23245
rect 34241 23236 34253 23239
rect 34204 23208 34253 23236
rect 34204 23196 34210 23208
rect 34241 23205 34253 23208
rect 34287 23205 34299 23239
rect 34241 23199 34299 23205
rect 36262 23196 36268 23248
rect 36320 23236 36326 23248
rect 36633 23239 36691 23245
rect 36633 23236 36645 23239
rect 36320 23208 36645 23236
rect 36320 23196 36326 23208
rect 36633 23205 36645 23208
rect 36679 23205 36691 23239
rect 36633 23199 36691 23205
rect 38654 23196 38660 23248
rect 38712 23236 38718 23248
rect 38841 23239 38899 23245
rect 38841 23236 38853 23239
rect 38712 23208 38853 23236
rect 38712 23196 38718 23208
rect 38841 23205 38853 23208
rect 38887 23236 38899 23239
rect 39758 23236 39764 23248
rect 38887 23208 39764 23236
rect 38887 23205 38899 23208
rect 38841 23199 38899 23205
rect 39758 23196 39764 23208
rect 39816 23196 39822 23248
rect 40402 23196 40408 23248
rect 40460 23236 40466 23248
rect 40954 23236 40960 23248
rect 40460 23208 40960 23236
rect 40460 23196 40466 23208
rect 40954 23196 40960 23208
rect 41012 23196 41018 23248
rect 46934 23196 46940 23248
rect 46992 23196 46998 23248
rect 47118 23196 47124 23248
rect 47176 23236 47182 23248
rect 47213 23239 47271 23245
rect 47213 23236 47225 23239
rect 47176 23208 47225 23236
rect 47176 23196 47182 23208
rect 47213 23205 47225 23208
rect 47259 23205 47271 23239
rect 47213 23199 47271 23205
rect 34517 23171 34575 23177
rect 34517 23137 34529 23171
rect 34563 23168 34575 23171
rect 34606 23168 34612 23180
rect 34563 23140 34612 23168
rect 34563 23137 34575 23140
rect 34517 23131 34575 23137
rect 34606 23128 34612 23140
rect 34664 23128 34670 23180
rect 34882 23128 34888 23180
rect 34940 23168 34946 23180
rect 37093 23171 37151 23177
rect 37093 23168 37105 23171
rect 34940 23140 37105 23168
rect 34940 23128 34946 23140
rect 37093 23137 37105 23140
rect 37139 23168 37151 23171
rect 37458 23168 37464 23180
rect 37139 23140 37464 23168
rect 37139 23137 37151 23140
rect 37093 23131 37151 23137
rect 37458 23128 37464 23140
rect 37516 23168 37522 23180
rect 41693 23171 41751 23177
rect 41693 23168 41705 23171
rect 37516 23140 41705 23168
rect 37516 23128 37522 23140
rect 41693 23137 41705 23140
rect 41739 23137 41751 23171
rect 41693 23131 41751 23137
rect 41969 23171 42027 23177
rect 41969 23137 41981 23171
rect 42015 23168 42027 23171
rect 42610 23168 42616 23180
rect 42015 23140 42616 23168
rect 42015 23137 42027 23140
rect 41969 23131 42027 23137
rect 42610 23128 42616 23140
rect 42668 23128 42674 23180
rect 43438 23128 43444 23180
rect 43496 23168 43502 23180
rect 45094 23168 45100 23180
rect 43496 23140 45100 23168
rect 43496 23128 43502 23140
rect 45094 23128 45100 23140
rect 45152 23128 45158 23180
rect 46658 23128 46664 23180
rect 46716 23168 46722 23180
rect 48041 23171 48099 23177
rect 48041 23168 48053 23171
rect 46716 23140 48053 23168
rect 46716 23128 46722 23140
rect 48041 23137 48053 23140
rect 48087 23137 48099 23171
rect 48041 23131 48099 23137
rect 38838 23100 38844 23112
rect 38502 23072 38844 23100
rect 38838 23060 38844 23072
rect 38896 23060 38902 23112
rect 39482 23060 39488 23112
rect 39540 23060 39546 23112
rect 40034 23060 40040 23112
rect 40092 23060 40098 23112
rect 40310 23060 40316 23112
rect 40368 23060 40374 23112
rect 44269 23103 44327 23109
rect 44269 23069 44281 23103
rect 44315 23100 44327 23103
rect 44450 23100 44456 23112
rect 44315 23072 44456 23100
rect 44315 23069 44327 23072
rect 44269 23063 44327 23069
rect 44450 23060 44456 23072
rect 44508 23060 44514 23112
rect 45186 23060 45192 23112
rect 45244 23060 45250 23112
rect 46293 23103 46351 23109
rect 46293 23069 46305 23103
rect 46339 23100 46351 23103
rect 46842 23100 46848 23112
rect 46339 23072 46848 23100
rect 46339 23069 46351 23072
rect 46293 23063 46351 23069
rect 46842 23060 46848 23072
rect 46900 23060 46906 23112
rect 47118 23060 47124 23112
rect 47176 23100 47182 23112
rect 47397 23103 47455 23109
rect 47397 23100 47409 23103
rect 47176 23072 47409 23100
rect 47176 23060 47182 23072
rect 47397 23069 47409 23072
rect 47443 23069 47455 23103
rect 47397 23063 47455 23069
rect 48501 23103 48559 23109
rect 48501 23069 48513 23103
rect 48547 23100 48559 23103
rect 48866 23100 48872 23112
rect 48547 23072 48872 23100
rect 48547 23069 48559 23072
rect 48501 23063 48559 23069
rect 48866 23060 48872 23072
rect 48924 23060 48930 23112
rect 34514 22992 34520 23044
rect 34572 23032 34578 23044
rect 35161 23035 35219 23041
rect 35161 23032 35173 23035
rect 34572 23004 35173 23032
rect 34572 22992 34578 23004
rect 35161 23001 35173 23004
rect 35207 23001 35219 23035
rect 36538 23032 36544 23044
rect 36386 23004 36544 23032
rect 35161 22995 35219 23001
rect 36538 22992 36544 23004
rect 36596 23032 36602 23044
rect 36596 23004 37858 23032
rect 36596 22992 36602 23004
rect 38654 22992 38660 23044
rect 38712 23032 38718 23044
rect 43254 23032 43260 23044
rect 38712 23004 42380 23032
rect 43194 23004 43260 23032
rect 38712 22992 38718 23004
rect 33376 22936 33548 22964
rect 33376 22924 33382 22936
rect 33686 22924 33692 22976
rect 33744 22964 33750 22976
rect 33873 22967 33931 22973
rect 33873 22964 33885 22967
rect 33744 22936 33885 22964
rect 33744 22924 33750 22936
rect 33873 22933 33885 22936
rect 33919 22964 33931 22967
rect 35526 22964 35532 22976
rect 33919 22936 35532 22964
rect 33919 22933 33931 22936
rect 33873 22927 33931 22933
rect 35526 22924 35532 22936
rect 35584 22924 35590 22976
rect 37090 22924 37096 22976
rect 37148 22964 37154 22976
rect 38378 22964 38384 22976
rect 37148 22936 38384 22964
rect 37148 22924 37154 22936
rect 38378 22924 38384 22936
rect 38436 22924 38442 22976
rect 38930 22924 38936 22976
rect 38988 22964 38994 22976
rect 39301 22967 39359 22973
rect 39301 22964 39313 22967
rect 38988 22936 39313 22964
rect 38988 22924 38994 22936
rect 39301 22933 39313 22936
rect 39347 22933 39359 22967
rect 39301 22927 39359 22933
rect 40954 22924 40960 22976
rect 41012 22964 41018 22976
rect 41141 22967 41199 22973
rect 41141 22964 41153 22967
rect 41012 22936 41153 22964
rect 41012 22924 41018 22936
rect 41141 22933 41153 22936
rect 41187 22933 41199 22967
rect 41141 22927 41199 22933
rect 41417 22967 41475 22973
rect 41417 22933 41429 22967
rect 41463 22964 41475 22967
rect 42058 22964 42064 22976
rect 41463 22936 42064 22964
rect 41463 22933 41475 22936
rect 41417 22927 41475 22933
rect 42058 22924 42064 22936
rect 42116 22924 42122 22976
rect 42352 22964 42380 23004
rect 43254 22992 43260 23004
rect 43312 22992 43318 23044
rect 43714 22992 43720 23044
rect 43772 22992 43778 23044
rect 47026 22992 47032 23044
rect 47084 23032 47090 23044
rect 49145 23035 49203 23041
rect 49145 23032 49157 23035
rect 47084 23004 49157 23032
rect 47084 22992 47090 23004
rect 49145 23001 49157 23004
rect 49191 23001 49203 23035
rect 49145 22995 49203 23001
rect 43990 22964 43996 22976
rect 42352 22936 43996 22964
rect 43990 22924 43996 22936
rect 44048 22924 44054 22976
rect 44818 22924 44824 22976
rect 44876 22924 44882 22976
rect 49418 22924 49424 22976
rect 49476 22924 49482 22976
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 4154 22720 4160 22772
rect 4212 22720 4218 22772
rect 6457 22763 6515 22769
rect 6457 22729 6469 22763
rect 6503 22760 6515 22763
rect 7282 22760 7288 22772
rect 6503 22732 7288 22760
rect 6503 22729 6515 22732
rect 6457 22723 6515 22729
rect 7282 22720 7288 22732
rect 7340 22720 7346 22772
rect 7558 22720 7564 22772
rect 7616 22760 7622 22772
rect 9306 22760 9312 22772
rect 7616 22732 9312 22760
rect 7616 22720 7622 22732
rect 9306 22720 9312 22732
rect 9364 22720 9370 22772
rect 11164 22732 16528 22760
rect 6362 22692 6368 22704
rect 1780 22664 6368 22692
rect 1780 22633 1808 22664
rect 6362 22652 6368 22664
rect 6420 22652 6426 22704
rect 6641 22695 6699 22701
rect 6641 22661 6653 22695
rect 6687 22692 6699 22695
rect 6822 22692 6828 22704
rect 6687 22664 6828 22692
rect 6687 22661 6699 22664
rect 6641 22655 6699 22661
rect 6822 22652 6828 22664
rect 6880 22652 6886 22704
rect 7006 22652 7012 22704
rect 7064 22652 7070 22704
rect 9493 22695 9551 22701
rect 9493 22692 9505 22695
rect 7116 22664 9505 22692
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22593 1823 22627
rect 1765 22587 1823 22593
rect 3510 22584 3516 22636
rect 3568 22584 3574 22636
rect 4617 22627 4675 22633
rect 4617 22593 4629 22627
rect 4663 22593 4675 22627
rect 4617 22587 4675 22593
rect 2777 22559 2835 22565
rect 2777 22525 2789 22559
rect 2823 22556 2835 22559
rect 2866 22556 2872 22568
rect 2823 22528 2872 22556
rect 2823 22525 2835 22528
rect 2777 22519 2835 22525
rect 2866 22516 2872 22528
rect 2924 22516 2930 22568
rect 1946 22448 1952 22500
rect 2004 22488 2010 22500
rect 4632 22488 4660 22587
rect 5074 22516 5080 22568
rect 5132 22516 5138 22568
rect 6638 22516 6644 22568
rect 6696 22556 6702 22568
rect 7116 22556 7144 22664
rect 9493 22661 9505 22664
rect 9539 22692 9551 22695
rect 11054 22692 11060 22704
rect 9539 22664 11060 22692
rect 9539 22661 9551 22664
rect 9493 22655 9551 22661
rect 11054 22652 11060 22664
rect 11112 22652 11118 22704
rect 7653 22627 7711 22633
rect 7653 22593 7665 22627
rect 7699 22624 7711 22627
rect 7834 22624 7840 22636
rect 7699 22596 7840 22624
rect 7699 22593 7711 22596
rect 7653 22587 7711 22593
rect 7834 22584 7840 22596
rect 7892 22584 7898 22636
rect 9766 22584 9772 22636
rect 9824 22584 9830 22636
rect 11164 22624 11192 22732
rect 12406 22664 14964 22692
rect 9876 22596 11192 22624
rect 11977 22627 12035 22633
rect 6696 22528 7144 22556
rect 6696 22516 6702 22528
rect 7374 22516 7380 22568
rect 7432 22556 7438 22568
rect 7929 22559 7987 22565
rect 7929 22556 7941 22559
rect 7432 22528 7941 22556
rect 7432 22516 7438 22528
rect 7929 22525 7941 22528
rect 7975 22525 7987 22559
rect 7929 22519 7987 22525
rect 8018 22516 8024 22568
rect 8076 22556 8082 22568
rect 9876 22556 9904 22596
rect 11977 22593 11989 22627
rect 12023 22624 12035 22627
rect 12406 22624 12434 22664
rect 12023 22596 12434 22624
rect 12023 22593 12035 22596
rect 11977 22587 12035 22593
rect 12710 22584 12716 22636
rect 12768 22624 12774 22636
rect 13081 22627 13139 22633
rect 13081 22624 13093 22627
rect 12768 22596 13093 22624
rect 12768 22584 12774 22596
rect 13081 22593 13093 22596
rect 13127 22593 13139 22627
rect 13081 22587 13139 22593
rect 8076 22528 9904 22556
rect 8076 22516 8082 22528
rect 10226 22516 10232 22568
rect 10284 22516 10290 22568
rect 11698 22516 11704 22568
rect 11756 22556 11762 22568
rect 12250 22556 12256 22568
rect 11756 22528 12256 22556
rect 11756 22516 11762 22528
rect 12250 22516 12256 22528
rect 12308 22516 12314 22568
rect 13814 22516 13820 22568
rect 13872 22516 13878 22568
rect 14936 22556 14964 22664
rect 15838 22652 15844 22704
rect 15896 22652 15902 22704
rect 15102 22584 15108 22636
rect 15160 22584 15166 22636
rect 14936 22528 16436 22556
rect 2004 22460 4660 22488
rect 2004 22448 2010 22460
rect 4982 22448 4988 22500
rect 5040 22488 5046 22500
rect 5040 22460 12434 22488
rect 5040 22448 5046 22460
rect 1578 22380 1584 22432
rect 1636 22420 1642 22432
rect 4522 22420 4528 22432
rect 1636 22392 4528 22420
rect 1636 22380 1642 22392
rect 4522 22380 4528 22392
rect 4580 22380 4586 22432
rect 7374 22380 7380 22432
rect 7432 22420 7438 22432
rect 8018 22420 8024 22432
rect 7432 22392 8024 22420
rect 7432 22380 7438 22392
rect 8018 22380 8024 22392
rect 8076 22380 8082 22432
rect 12406 22420 12434 22460
rect 13906 22448 13912 22500
rect 13964 22488 13970 22500
rect 16022 22488 16028 22500
rect 13964 22460 16028 22488
rect 13964 22448 13970 22460
rect 16022 22448 16028 22460
rect 16080 22448 16086 22500
rect 16298 22420 16304 22432
rect 12406 22392 16304 22420
rect 16298 22380 16304 22392
rect 16356 22380 16362 22432
rect 16408 22420 16436 22528
rect 16500 22488 16528 22732
rect 17126 22720 17132 22772
rect 17184 22760 17190 22772
rect 19242 22760 19248 22772
rect 17184 22732 19248 22760
rect 17184 22720 17190 22732
rect 19242 22720 19248 22732
rect 19300 22720 19306 22772
rect 19610 22720 19616 22772
rect 19668 22760 19674 22772
rect 22465 22763 22523 22769
rect 22465 22760 22477 22763
rect 19668 22732 22477 22760
rect 19668 22720 19674 22732
rect 22465 22729 22477 22732
rect 22511 22729 22523 22763
rect 23014 22760 23020 22772
rect 22465 22723 22523 22729
rect 22572 22732 23020 22760
rect 17862 22652 17868 22704
rect 17920 22652 17926 22704
rect 19978 22692 19984 22704
rect 19076 22664 19984 22692
rect 18506 22584 18512 22636
rect 18564 22624 18570 22636
rect 19076 22624 19104 22664
rect 19978 22652 19984 22664
rect 20036 22652 20042 22704
rect 20806 22652 20812 22704
rect 20864 22692 20870 22704
rect 22572 22692 22600 22732
rect 23014 22720 23020 22732
rect 23072 22720 23078 22772
rect 24029 22763 24087 22769
rect 24029 22729 24041 22763
rect 24075 22760 24087 22763
rect 27614 22760 27620 22772
rect 24075 22732 27620 22760
rect 24075 22729 24087 22732
rect 24029 22723 24087 22729
rect 27614 22720 27620 22732
rect 27672 22720 27678 22772
rect 29178 22760 29184 22772
rect 28000 22732 29184 22760
rect 20864 22664 22600 22692
rect 22925 22695 22983 22701
rect 20864 22652 20870 22664
rect 22925 22661 22937 22695
rect 22971 22692 22983 22695
rect 25038 22692 25044 22704
rect 22971 22664 25044 22692
rect 22971 22661 22983 22664
rect 22925 22655 22983 22661
rect 25038 22652 25044 22664
rect 25096 22652 25102 22704
rect 25130 22652 25136 22704
rect 25188 22652 25194 22704
rect 26418 22692 26424 22704
rect 26358 22664 26424 22692
rect 26418 22652 26424 22664
rect 26476 22692 26482 22704
rect 27338 22692 27344 22704
rect 26476 22664 27344 22692
rect 26476 22652 26482 22664
rect 27338 22652 27344 22664
rect 27396 22652 27402 22704
rect 27433 22695 27491 22701
rect 27433 22661 27445 22695
rect 27479 22692 27491 22695
rect 28000 22692 28028 22732
rect 29178 22720 29184 22732
rect 29236 22720 29242 22772
rect 30006 22720 30012 22772
rect 30064 22760 30070 22772
rect 30190 22760 30196 22772
rect 30064 22732 30196 22760
rect 30064 22720 30070 22732
rect 30190 22720 30196 22732
rect 30248 22720 30254 22772
rect 30466 22720 30472 22772
rect 30524 22760 30530 22772
rect 32309 22763 32367 22769
rect 32309 22760 32321 22763
rect 30524 22732 32321 22760
rect 30524 22720 30530 22732
rect 32309 22729 32321 22732
rect 32355 22729 32367 22763
rect 32309 22723 32367 22729
rect 32582 22720 32588 22772
rect 32640 22760 32646 22772
rect 36081 22763 36139 22769
rect 36081 22760 36093 22763
rect 32640 22732 36093 22760
rect 32640 22720 32646 22732
rect 36081 22729 36093 22732
rect 36127 22729 36139 22763
rect 36081 22723 36139 22729
rect 36449 22763 36507 22769
rect 36449 22729 36461 22763
rect 36495 22760 36507 22763
rect 36495 22732 39620 22760
rect 36495 22729 36507 22732
rect 36449 22723 36507 22729
rect 28626 22692 28632 22704
rect 27479 22664 28028 22692
rect 28092 22664 28632 22692
rect 27479 22661 27491 22664
rect 27433 22655 27491 22661
rect 18564 22596 19104 22624
rect 18564 22584 18570 22596
rect 19242 22584 19248 22636
rect 19300 22584 19306 22636
rect 22833 22627 22891 22633
rect 22833 22593 22845 22627
rect 22879 22624 22891 22627
rect 23290 22624 23296 22636
rect 22879 22596 23296 22624
rect 22879 22593 22891 22596
rect 22833 22587 22891 22593
rect 23290 22584 23296 22596
rect 23348 22584 23354 22636
rect 24121 22627 24179 22633
rect 24121 22593 24133 22627
rect 24167 22624 24179 22627
rect 24394 22624 24400 22636
rect 24167 22596 24400 22624
rect 24167 22593 24179 22596
rect 24121 22587 24179 22593
rect 24394 22584 24400 22596
rect 24452 22584 24458 22636
rect 27614 22584 27620 22636
rect 27672 22624 27678 22636
rect 27798 22624 27804 22636
rect 27672 22596 27804 22624
rect 27672 22584 27678 22596
rect 27798 22584 27804 22596
rect 27856 22584 27862 22636
rect 16850 22516 16856 22568
rect 16908 22516 16914 22568
rect 17129 22559 17187 22565
rect 17129 22556 17141 22559
rect 16960 22528 17141 22556
rect 16960 22488 16988 22528
rect 17129 22525 17141 22528
rect 17175 22525 17187 22559
rect 17129 22519 17187 22525
rect 18138 22516 18144 22568
rect 18196 22556 18202 22568
rect 19521 22559 19579 22565
rect 19521 22556 19533 22559
rect 18196 22528 19533 22556
rect 18196 22516 18202 22528
rect 19521 22525 19533 22528
rect 19567 22525 19579 22559
rect 19521 22519 19579 22525
rect 20898 22516 20904 22568
rect 20956 22556 20962 22568
rect 21266 22556 21272 22568
rect 20956 22528 21272 22556
rect 20956 22516 20962 22528
rect 21266 22516 21272 22528
rect 21324 22516 21330 22568
rect 21358 22516 21364 22568
rect 21416 22556 21422 22568
rect 22186 22556 22192 22568
rect 21416 22528 22192 22556
rect 21416 22516 21422 22528
rect 22186 22516 22192 22528
rect 22244 22556 22250 22568
rect 23017 22559 23075 22565
rect 23017 22556 23029 22559
rect 22244 22528 23029 22556
rect 22244 22516 22250 22528
rect 23017 22525 23029 22528
rect 23063 22525 23075 22559
rect 23017 22519 23075 22525
rect 23382 22516 23388 22568
rect 23440 22556 23446 22568
rect 24213 22559 24271 22565
rect 24213 22556 24225 22559
rect 23440 22528 24225 22556
rect 23440 22516 23446 22528
rect 24213 22525 24225 22528
rect 24259 22525 24271 22559
rect 24213 22519 24271 22525
rect 22097 22491 22155 22497
rect 22097 22488 22109 22491
rect 16500 22460 16988 22488
rect 18156 22460 19012 22488
rect 18156 22420 18184 22460
rect 16408 22392 18184 22420
rect 18598 22380 18604 22432
rect 18656 22380 18662 22432
rect 18874 22380 18880 22432
rect 18932 22380 18938 22432
rect 18984 22420 19012 22460
rect 21284 22460 22109 22488
rect 21284 22420 21312 22460
rect 22097 22457 22109 22460
rect 22143 22488 22155 22491
rect 23474 22488 23480 22500
rect 22143 22460 23480 22488
rect 22143 22457 22155 22460
rect 22097 22451 22155 22457
rect 23474 22448 23480 22460
rect 23532 22448 23538 22500
rect 18984 22392 21312 22420
rect 21358 22380 21364 22432
rect 21416 22420 21422 22432
rect 21545 22423 21603 22429
rect 21545 22420 21557 22423
rect 21416 22392 21557 22420
rect 21416 22380 21422 22392
rect 21545 22389 21557 22392
rect 21591 22389 21603 22423
rect 21545 22383 21603 22389
rect 22005 22423 22063 22429
rect 22005 22389 22017 22423
rect 22051 22420 22063 22423
rect 22370 22420 22376 22432
rect 22051 22392 22376 22420
rect 22051 22389 22063 22392
rect 22005 22383 22063 22389
rect 22370 22380 22376 22392
rect 22428 22380 22434 22432
rect 23658 22380 23664 22432
rect 23716 22380 23722 22432
rect 24228 22420 24256 22519
rect 24302 22516 24308 22568
rect 24360 22556 24366 22568
rect 24762 22556 24768 22568
rect 24360 22528 24768 22556
rect 24360 22516 24366 22528
rect 24762 22516 24768 22528
rect 24820 22556 24826 22568
rect 28092 22565 28120 22664
rect 28626 22652 28632 22664
rect 28684 22652 28690 22704
rect 30745 22695 30803 22701
rect 30745 22661 30757 22695
rect 30791 22692 30803 22695
rect 32122 22692 32128 22704
rect 30791 22664 32128 22692
rect 30791 22661 30803 22664
rect 30745 22655 30803 22661
rect 32122 22652 32128 22664
rect 32180 22652 32186 22704
rect 35158 22692 35164 22704
rect 35098 22664 35164 22692
rect 35158 22652 35164 22664
rect 35216 22692 35222 22704
rect 36538 22692 36544 22704
rect 35216 22664 36544 22692
rect 35216 22652 35222 22664
rect 36538 22652 36544 22664
rect 36596 22652 36602 22704
rect 39022 22652 39028 22704
rect 39080 22692 39086 22704
rect 39390 22692 39396 22704
rect 39080 22664 39396 22692
rect 39080 22652 39086 22664
rect 39390 22652 39396 22664
rect 39448 22652 39454 22704
rect 39592 22692 39620 22732
rect 39666 22720 39672 22772
rect 39724 22720 39730 22772
rect 40037 22763 40095 22769
rect 40037 22729 40049 22763
rect 40083 22760 40095 22763
rect 40865 22763 40923 22769
rect 40865 22760 40877 22763
rect 40083 22732 40877 22760
rect 40083 22729 40095 22732
rect 40037 22723 40095 22729
rect 40865 22729 40877 22732
rect 40911 22729 40923 22763
rect 41233 22763 41291 22769
rect 41233 22760 41245 22763
rect 40865 22723 40923 22729
rect 40972 22732 41245 22760
rect 40126 22692 40132 22704
rect 39592 22664 40132 22692
rect 40126 22652 40132 22664
rect 40184 22652 40190 22704
rect 24857 22559 24915 22565
rect 24857 22556 24869 22559
rect 24820 22528 24869 22556
rect 24820 22516 24826 22528
rect 24857 22525 24869 22528
rect 24903 22556 24915 22559
rect 28077 22559 28135 22565
rect 28077 22556 28089 22559
rect 24903 22528 28089 22556
rect 24903 22525 24915 22528
rect 24857 22519 24915 22525
rect 28077 22525 28089 22528
rect 28123 22525 28135 22559
rect 28077 22519 28135 22525
rect 28350 22516 28356 22568
rect 28408 22516 28414 22568
rect 29086 22516 29092 22568
rect 29144 22556 29150 22568
rect 29472 22556 29500 22610
rect 30650 22584 30656 22636
rect 30708 22584 30714 22636
rect 30760 22596 31524 22624
rect 30760 22556 30788 22596
rect 29144 22528 30788 22556
rect 29144 22516 29150 22528
rect 30926 22516 30932 22568
rect 30984 22516 30990 22568
rect 31496 22556 31524 22596
rect 31570 22584 31576 22636
rect 31628 22584 31634 22636
rect 31757 22627 31815 22633
rect 31757 22593 31769 22627
rect 31803 22624 31815 22627
rect 31846 22624 31852 22636
rect 31803 22596 31852 22624
rect 31803 22593 31815 22596
rect 31757 22587 31815 22593
rect 31846 22584 31852 22596
rect 31904 22584 31910 22636
rect 32674 22584 32680 22636
rect 32732 22584 32738 22636
rect 33410 22584 33416 22636
rect 33468 22624 33474 22636
rect 33594 22624 33600 22636
rect 33468 22596 33600 22624
rect 33468 22584 33474 22596
rect 33594 22584 33600 22596
rect 33652 22584 33658 22636
rect 37274 22624 37280 22636
rect 35084 22596 37280 22624
rect 31662 22556 31668 22568
rect 31496 22528 31668 22556
rect 31662 22516 31668 22528
rect 31720 22516 31726 22568
rect 32766 22516 32772 22568
rect 32824 22516 32830 22568
rect 32858 22516 32864 22568
rect 32916 22516 32922 22568
rect 35084 22556 35112 22596
rect 37274 22584 37280 22596
rect 37332 22584 37338 22636
rect 37458 22584 37464 22636
rect 37516 22584 37522 22636
rect 38838 22584 38844 22636
rect 38896 22624 38902 22636
rect 40494 22624 40500 22636
rect 38896 22596 40500 22624
rect 38896 22584 38902 22596
rect 40494 22584 40500 22596
rect 40552 22584 40558 22636
rect 33704 22528 35112 22556
rect 26326 22448 26332 22500
rect 26384 22488 26390 22500
rect 26973 22491 27031 22497
rect 26973 22488 26985 22491
rect 26384 22460 26985 22488
rect 26384 22448 26390 22460
rect 26973 22457 26985 22460
rect 27019 22457 27031 22491
rect 26973 22451 27031 22457
rect 27062 22448 27068 22500
rect 27120 22488 27126 22500
rect 27617 22491 27675 22497
rect 27617 22488 27629 22491
rect 27120 22460 27629 22488
rect 27120 22448 27126 22460
rect 27617 22457 27629 22460
rect 27663 22457 27675 22491
rect 27617 22451 27675 22457
rect 30285 22491 30343 22497
rect 30285 22457 30297 22491
rect 30331 22488 30343 22491
rect 31570 22488 31576 22500
rect 30331 22460 31576 22488
rect 30331 22457 30343 22460
rect 30285 22451 30343 22457
rect 31570 22448 31576 22460
rect 31628 22448 31634 22500
rect 32306 22448 32312 22500
rect 32364 22488 32370 22500
rect 32876 22488 32904 22516
rect 33704 22488 33732 22528
rect 35342 22516 35348 22568
rect 35400 22516 35406 22568
rect 36538 22516 36544 22568
rect 36596 22516 36602 22568
rect 36630 22516 36636 22568
rect 36688 22516 36694 22568
rect 37734 22516 37740 22568
rect 37792 22516 37798 22568
rect 38470 22516 38476 22568
rect 38528 22556 38534 22568
rect 40129 22559 40187 22565
rect 40129 22556 40141 22559
rect 38528 22528 40141 22556
rect 38528 22516 38534 22528
rect 40129 22525 40141 22528
rect 40175 22525 40187 22559
rect 40310 22556 40316 22568
rect 40129 22519 40187 22525
rect 40236 22528 40316 22556
rect 32364 22460 32904 22488
rect 33244 22460 33732 22488
rect 35713 22491 35771 22497
rect 32364 22448 32370 22460
rect 26605 22423 26663 22429
rect 26605 22420 26617 22423
rect 24228 22392 26617 22420
rect 26605 22389 26617 22392
rect 26651 22389 26663 22423
rect 26605 22383 26663 22389
rect 28442 22380 28448 22432
rect 28500 22420 28506 22432
rect 29825 22423 29883 22429
rect 29825 22420 29837 22423
rect 28500 22392 29837 22420
rect 28500 22380 28506 22392
rect 29825 22389 29837 22392
rect 29871 22420 29883 22423
rect 33244 22420 33272 22460
rect 35713 22457 35725 22491
rect 35759 22488 35771 22491
rect 35986 22488 35992 22500
rect 35759 22460 35992 22488
rect 35759 22457 35771 22460
rect 35713 22451 35771 22457
rect 35986 22448 35992 22460
rect 36044 22448 36050 22500
rect 39209 22491 39267 22497
rect 39209 22457 39221 22491
rect 39255 22488 39267 22491
rect 40236 22488 40264 22528
rect 40310 22516 40316 22528
rect 40368 22516 40374 22568
rect 40678 22516 40684 22568
rect 40736 22556 40742 22568
rect 40972 22556 41000 22732
rect 41233 22729 41245 22732
rect 41279 22729 41291 22763
rect 41233 22723 41291 22729
rect 45646 22720 45652 22772
rect 45704 22760 45710 22772
rect 45741 22763 45799 22769
rect 45741 22760 45753 22763
rect 45704 22732 45753 22760
rect 45704 22720 45710 22732
rect 45741 22729 45753 22732
rect 45787 22729 45799 22763
rect 45741 22723 45799 22729
rect 46842 22720 46848 22772
rect 46900 22720 46906 22772
rect 47762 22720 47768 22772
rect 47820 22720 47826 22772
rect 43254 22652 43260 22704
rect 43312 22692 43318 22704
rect 44453 22695 44511 22701
rect 44453 22692 44465 22695
rect 43312 22664 44465 22692
rect 43312 22652 43318 22664
rect 44453 22661 44465 22664
rect 44499 22661 44511 22695
rect 46934 22692 46940 22704
rect 44453 22655 44511 22661
rect 44560 22664 46940 22692
rect 42426 22584 42432 22636
rect 42484 22624 42490 22636
rect 42613 22627 42671 22633
rect 42613 22624 42625 22627
rect 42484 22596 42625 22624
rect 42484 22584 42490 22596
rect 42613 22593 42625 22596
rect 42659 22593 42671 22627
rect 42613 22587 42671 22593
rect 43714 22584 43720 22636
rect 43772 22624 43778 22636
rect 44560 22624 44588 22664
rect 46934 22652 46940 22664
rect 46992 22692 46998 22704
rect 47780 22692 47808 22720
rect 46992 22664 47808 22692
rect 46992 22652 46998 22664
rect 48682 22652 48688 22704
rect 48740 22692 48746 22704
rect 49142 22692 49148 22704
rect 48740 22664 49148 22692
rect 48740 22652 48746 22664
rect 49142 22652 49148 22664
rect 49200 22652 49206 22704
rect 43772 22596 44588 22624
rect 43772 22584 43778 22596
rect 45094 22584 45100 22636
rect 45152 22584 45158 22636
rect 46198 22584 46204 22636
rect 46256 22584 46262 22636
rect 47762 22584 47768 22636
rect 47820 22584 47826 22636
rect 48869 22627 48927 22633
rect 48869 22593 48881 22627
rect 48915 22624 48927 22627
rect 50522 22624 50528 22636
rect 48915 22596 50528 22624
rect 48915 22593 48927 22596
rect 48869 22587 48927 22593
rect 50522 22584 50528 22596
rect 50580 22584 50586 22636
rect 40736 22528 41000 22556
rect 40736 22516 40742 22528
rect 41230 22516 41236 22568
rect 41288 22556 41294 22568
rect 41325 22559 41383 22565
rect 41325 22556 41337 22559
rect 41288 22528 41337 22556
rect 41288 22516 41294 22528
rect 41325 22525 41337 22528
rect 41371 22525 41383 22559
rect 41509 22559 41567 22565
rect 41509 22556 41521 22559
rect 41467 22528 41521 22556
rect 41325 22519 41383 22525
rect 41509 22525 41521 22528
rect 41555 22556 41567 22559
rect 41555 22528 42196 22556
rect 41555 22525 41567 22528
rect 41509 22519 41567 22525
rect 39255 22460 40264 22488
rect 40328 22460 41184 22488
rect 39255 22457 39267 22460
rect 39209 22451 39267 22457
rect 29871 22392 33272 22420
rect 33860 22423 33918 22429
rect 29871 22389 29883 22392
rect 29825 22383 29883 22389
rect 33860 22389 33872 22423
rect 33906 22420 33918 22423
rect 34422 22420 34428 22432
rect 33906 22392 34428 22420
rect 33906 22389 33918 22392
rect 33860 22383 33918 22389
rect 34422 22380 34428 22392
rect 34480 22380 34486 22432
rect 34974 22380 34980 22432
rect 35032 22420 35038 22432
rect 36170 22420 36176 22432
rect 35032 22392 36176 22420
rect 35032 22380 35038 22392
rect 36170 22380 36176 22392
rect 36228 22380 36234 22432
rect 37182 22380 37188 22432
rect 37240 22420 37246 22432
rect 39224 22420 39252 22451
rect 37240 22392 39252 22420
rect 37240 22380 37246 22392
rect 39390 22380 39396 22432
rect 39448 22420 39454 22432
rect 40328 22420 40356 22460
rect 39448 22392 40356 22420
rect 41156 22420 41184 22460
rect 41524 22420 41552 22519
rect 41874 22448 41880 22500
rect 41932 22448 41938 22500
rect 41156 22392 41552 22420
rect 39448 22380 39454 22392
rect 41598 22380 41604 22432
rect 41656 22420 41662 22432
rect 42061 22423 42119 22429
rect 42061 22420 42073 22423
rect 41656 22392 42073 22420
rect 41656 22380 41662 22392
rect 42061 22389 42073 22392
rect 42107 22389 42119 22423
rect 42168 22420 42196 22528
rect 43806 22516 43812 22568
rect 43864 22556 43870 22568
rect 46106 22556 46112 22568
rect 43864 22528 46112 22556
rect 43864 22516 43870 22528
rect 46106 22516 46112 22528
rect 46164 22516 46170 22568
rect 44174 22488 44180 22500
rect 42352 22460 44180 22488
rect 42352 22420 42380 22460
rect 44174 22448 44180 22460
rect 44232 22448 44238 22500
rect 44450 22448 44456 22500
rect 44508 22488 44514 22500
rect 45002 22488 45008 22500
rect 44508 22460 45008 22488
rect 44508 22448 44514 22460
rect 45002 22448 45008 22460
rect 45060 22448 45066 22500
rect 45278 22448 45284 22500
rect 45336 22488 45342 22500
rect 47305 22491 47363 22497
rect 47305 22488 47317 22491
rect 45336 22460 47317 22488
rect 45336 22448 45342 22460
rect 47305 22457 47317 22460
rect 47351 22457 47363 22491
rect 47305 22451 47363 22457
rect 42168 22392 42380 22420
rect 43257 22423 43315 22429
rect 42061 22383 42119 22389
rect 43257 22389 43269 22423
rect 43303 22420 43315 22423
rect 45186 22420 45192 22432
rect 43303 22392 45192 22420
rect 43303 22389 43315 22392
rect 43257 22383 43315 22389
rect 45186 22380 45192 22392
rect 45244 22380 45250 22432
rect 45370 22380 45376 22432
rect 45428 22420 45434 22432
rect 47121 22423 47179 22429
rect 47121 22420 47133 22423
rect 45428 22392 47133 22420
rect 45428 22380 45434 22392
rect 47121 22389 47133 22392
rect 47167 22389 47179 22423
rect 47121 22383 47179 22389
rect 48406 22380 48412 22432
rect 48464 22380 48470 22432
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 2222 22176 2228 22228
rect 2280 22216 2286 22228
rect 4890 22216 4896 22228
rect 2280 22188 4896 22216
rect 2280 22176 2286 22188
rect 4890 22176 4896 22188
rect 4948 22176 4954 22228
rect 6362 22176 6368 22228
rect 6420 22216 6426 22228
rect 9950 22216 9956 22228
rect 6420 22188 9956 22216
rect 6420 22176 6426 22188
rect 9950 22176 9956 22188
rect 10008 22176 10014 22228
rect 10318 22176 10324 22228
rect 10376 22216 10382 22228
rect 14458 22216 14464 22228
rect 10376 22188 14464 22216
rect 10376 22176 10382 22188
rect 14458 22176 14464 22188
rect 14516 22176 14522 22228
rect 15286 22225 15292 22228
rect 15270 22219 15292 22225
rect 15270 22185 15282 22219
rect 15270 22179 15292 22185
rect 15286 22176 15292 22179
rect 15344 22176 15350 22228
rect 16022 22176 16028 22228
rect 16080 22216 16086 22228
rect 18598 22216 18604 22228
rect 16080 22188 18604 22216
rect 16080 22176 16086 22188
rect 18598 22176 18604 22188
rect 18656 22216 18662 22228
rect 18656 22188 20208 22216
rect 18656 22176 18662 22188
rect 3694 22108 3700 22160
rect 3752 22148 3758 22160
rect 3752 22120 6316 22148
rect 3752 22108 3758 22120
rect 1302 22040 1308 22092
rect 1360 22080 1366 22092
rect 2041 22083 2099 22089
rect 2041 22080 2053 22083
rect 1360 22052 2053 22080
rect 1360 22040 1366 22052
rect 2041 22049 2053 22052
rect 2087 22049 2099 22083
rect 2041 22043 2099 22049
rect 3234 22040 3240 22092
rect 3292 22080 3298 22092
rect 6288 22089 6316 22120
rect 6822 22108 6828 22160
rect 6880 22148 6886 22160
rect 11698 22148 11704 22160
rect 6880 22120 11704 22148
rect 6880 22108 6886 22120
rect 11698 22108 11704 22120
rect 11756 22108 11762 22160
rect 11882 22108 11888 22160
rect 11940 22148 11946 22160
rect 11940 22120 12480 22148
rect 11940 22108 11946 22120
rect 4433 22083 4491 22089
rect 4433 22080 4445 22083
rect 3292 22052 4445 22080
rect 3292 22040 3298 22052
rect 4433 22049 4445 22052
rect 4479 22049 4491 22083
rect 4433 22043 4491 22049
rect 6273 22083 6331 22089
rect 6273 22049 6285 22083
rect 6319 22080 6331 22083
rect 6319 22052 6353 22080
rect 6472 22052 9168 22080
rect 6319 22049 6331 22052
rect 6273 22043 6331 22049
rect 1765 22015 1823 22021
rect 1765 21981 1777 22015
rect 1811 21981 1823 22015
rect 1765 21975 1823 21981
rect 1780 21944 1808 21975
rect 3142 21972 3148 22024
rect 3200 22012 3206 22024
rect 3973 22015 4031 22021
rect 3973 22012 3985 22015
rect 3200 21984 3985 22012
rect 3200 21972 3206 21984
rect 3973 21981 3985 21984
rect 4019 21981 4031 22015
rect 3973 21975 4031 21981
rect 5810 21972 5816 22024
rect 5868 21972 5874 22024
rect 6086 21972 6092 22024
rect 6144 22012 6150 22024
rect 6472 22012 6500 22052
rect 6144 21984 6500 22012
rect 6144 21972 6150 21984
rect 7650 21972 7656 22024
rect 7708 22012 7714 22024
rect 9140 22021 9168 22052
rect 9766 22040 9772 22092
rect 9824 22040 9830 22092
rect 12452 22089 12480 22120
rect 12526 22108 12532 22160
rect 12584 22148 12590 22160
rect 14553 22151 14611 22157
rect 14553 22148 14565 22151
rect 12584 22120 14565 22148
rect 12584 22108 12590 22120
rect 14553 22117 14565 22120
rect 14599 22117 14611 22151
rect 16850 22148 16856 22160
rect 14553 22111 14611 22117
rect 16546 22120 16856 22148
rect 12437 22083 12495 22089
rect 10888 22052 12112 22080
rect 7929 22015 7987 22021
rect 7929 22012 7941 22015
rect 7708 21984 7941 22012
rect 7708 21972 7714 21984
rect 7929 21981 7941 21984
rect 7975 21981 7987 22015
rect 7929 21975 7987 21981
rect 9125 22015 9183 22021
rect 9125 21981 9137 22015
rect 9171 21981 9183 22015
rect 10888 22012 10916 22052
rect 9125 21975 9183 21981
rect 9232 21984 10916 22012
rect 10965 22015 11023 22021
rect 3605 21947 3663 21953
rect 1780 21916 3556 21944
rect 3418 21836 3424 21888
rect 3476 21836 3482 21888
rect 3528 21876 3556 21916
rect 3605 21913 3617 21947
rect 3651 21944 3663 21947
rect 9232 21944 9260 21984
rect 10965 21981 10977 22015
rect 11011 22012 11023 22015
rect 11977 22015 12035 22021
rect 11011 21984 11652 22012
rect 11011 21981 11023 21984
rect 10965 21975 11023 21981
rect 3651 21916 9260 21944
rect 3651 21913 3663 21916
rect 3605 21907 3663 21913
rect 11330 21904 11336 21956
rect 11388 21904 11394 21956
rect 5534 21876 5540 21888
rect 3528 21848 5540 21876
rect 5534 21836 5540 21848
rect 5592 21836 5598 21888
rect 7650 21836 7656 21888
rect 7708 21836 7714 21888
rect 8573 21879 8631 21885
rect 8573 21845 8585 21879
rect 8619 21876 8631 21879
rect 9398 21876 9404 21888
rect 8619 21848 9404 21876
rect 8619 21845 8631 21848
rect 8573 21839 8631 21845
rect 9398 21836 9404 21848
rect 9456 21836 9462 21888
rect 9490 21836 9496 21888
rect 9548 21876 9554 21888
rect 11425 21879 11483 21885
rect 11425 21876 11437 21879
rect 9548 21848 11437 21876
rect 9548 21836 9554 21848
rect 11425 21845 11437 21848
rect 11471 21845 11483 21879
rect 11624 21876 11652 21984
rect 11977 21981 11989 22015
rect 12023 21981 12035 22015
rect 12084 22012 12112 22052
rect 12437 22049 12449 22083
rect 12483 22049 12495 22083
rect 12437 22043 12495 22049
rect 15010 22040 15016 22092
rect 15068 22080 15074 22092
rect 16546 22080 16574 22120
rect 16850 22108 16856 22120
rect 16908 22108 16914 22160
rect 17402 22108 17408 22160
rect 17460 22148 17466 22160
rect 19610 22148 19616 22160
rect 17460 22120 19616 22148
rect 17460 22108 17466 22120
rect 19610 22108 19616 22120
rect 19668 22108 19674 22160
rect 15068 22052 16574 22080
rect 16684 22052 17632 22080
rect 15068 22040 15074 22052
rect 16684 22024 16712 22052
rect 12084 21984 14044 22012
rect 11977 21975 12035 21981
rect 11992 21944 12020 21975
rect 12342 21944 12348 21956
rect 11992 21916 12348 21944
rect 12342 21904 12348 21916
rect 12400 21904 12406 21956
rect 12618 21904 12624 21956
rect 12676 21944 12682 21956
rect 14016 21944 14044 21984
rect 14642 21972 14648 22024
rect 14700 22012 14706 22024
rect 14829 22015 14887 22021
rect 14829 22012 14841 22015
rect 14700 21984 14841 22012
rect 14700 21972 14706 21984
rect 14829 21981 14841 21984
rect 14875 21981 14887 22015
rect 16666 22012 16672 22024
rect 16422 21984 16672 22012
rect 14829 21975 14887 21981
rect 16666 21972 16672 21984
rect 16724 21972 16730 22024
rect 16758 21972 16764 22024
rect 16816 22012 16822 22024
rect 17310 22012 17316 22024
rect 16816 21984 17316 22012
rect 16816 21972 16822 21984
rect 17310 21972 17316 21984
rect 17368 21972 17374 22024
rect 17494 21972 17500 22024
rect 17552 21972 17558 22024
rect 17604 22012 17632 22052
rect 17678 22040 17684 22092
rect 17736 22080 17742 22092
rect 20180 22089 20208 22188
rect 21266 22176 21272 22228
rect 21324 22216 21330 22228
rect 21324 22188 22784 22216
rect 21324 22176 21330 22188
rect 21082 22108 21088 22160
rect 21140 22148 21146 22160
rect 22756 22148 22784 22188
rect 23290 22176 23296 22228
rect 23348 22176 23354 22228
rect 23842 22216 23848 22228
rect 23768 22188 23848 22216
rect 23768 22148 23796 22188
rect 23842 22176 23848 22188
rect 23900 22176 23906 22228
rect 24210 22176 24216 22228
rect 24268 22216 24274 22228
rect 24578 22216 24584 22228
rect 24268 22188 24584 22216
rect 24268 22176 24274 22188
rect 24578 22176 24584 22188
rect 24636 22176 24642 22228
rect 27338 22176 27344 22228
rect 27396 22216 27402 22228
rect 28534 22216 28540 22228
rect 27396 22188 28540 22216
rect 27396 22176 27402 22188
rect 28534 22176 28540 22188
rect 28592 22176 28598 22228
rect 28810 22176 28816 22228
rect 28868 22216 28874 22228
rect 31100 22219 31158 22225
rect 28868 22188 30972 22216
rect 28868 22176 28874 22188
rect 21140 22120 21404 22148
rect 21140 22108 21146 22120
rect 21376 22089 21404 22120
rect 22480 22120 22692 22148
rect 22756 22120 23796 22148
rect 17957 22083 18015 22089
rect 17957 22080 17969 22083
rect 17736 22052 17969 22080
rect 17736 22040 17742 22052
rect 17957 22049 17969 22052
rect 18003 22049 18015 22083
rect 17957 22043 18015 22049
rect 20165 22083 20223 22089
rect 20165 22049 20177 22083
rect 20211 22049 20223 22083
rect 20165 22043 20223 22049
rect 21361 22083 21419 22089
rect 21361 22049 21373 22083
rect 21407 22049 21419 22083
rect 22480 22080 22508 22120
rect 21361 22043 21419 22049
rect 21560 22052 22508 22080
rect 17862 22012 17868 22024
rect 17604 21984 17868 22012
rect 17862 21972 17868 21984
rect 17920 21972 17926 22024
rect 19426 21972 19432 22024
rect 19484 22012 19490 22024
rect 19981 22015 20039 22021
rect 19981 22012 19993 22015
rect 19484 21984 19993 22012
rect 19484 21972 19490 21984
rect 19981 21981 19993 21984
rect 20027 21981 20039 22015
rect 21560 22012 21588 22052
rect 22554 22040 22560 22092
rect 22612 22040 22618 22092
rect 22664 22080 22692 22120
rect 23934 22108 23940 22160
rect 23992 22148 23998 22160
rect 26694 22148 26700 22160
rect 23992 22120 25360 22148
rect 23992 22108 23998 22120
rect 23382 22080 23388 22092
rect 22664 22052 23388 22080
rect 23382 22040 23388 22052
rect 23440 22040 23446 22092
rect 23750 22040 23756 22092
rect 23808 22040 23814 22092
rect 23842 22040 23848 22092
rect 23900 22040 23906 22092
rect 25332 22089 25360 22120
rect 26436 22120 26700 22148
rect 26436 22089 26464 22120
rect 26694 22108 26700 22120
rect 26752 22108 26758 22160
rect 28626 22108 28632 22160
rect 28684 22148 28690 22160
rect 28684 22120 30880 22148
rect 28684 22108 28690 22120
rect 25317 22083 25375 22089
rect 25317 22049 25329 22083
rect 25363 22080 25375 22083
rect 26421 22083 26479 22089
rect 25363 22052 25397 22080
rect 25363 22049 25375 22052
rect 25317 22043 25375 22049
rect 26421 22049 26433 22083
rect 26467 22049 26479 22083
rect 26421 22043 26479 22049
rect 26510 22040 26516 22092
rect 26568 22040 26574 22092
rect 29822 22080 29828 22092
rect 26620 22052 29828 22080
rect 19981 21975 20039 21981
rect 20088 21984 21588 22012
rect 14366 21944 14372 21956
rect 12676 21916 13952 21944
rect 14016 21916 14372 21944
rect 12676 21904 12682 21916
rect 13630 21876 13636 21888
rect 11624 21848 13636 21876
rect 11425 21839 11483 21845
rect 13630 21836 13636 21848
rect 13688 21836 13694 21888
rect 13722 21836 13728 21888
rect 13780 21836 13786 21888
rect 13814 21836 13820 21888
rect 13872 21836 13878 21888
rect 13924 21876 13952 21916
rect 14366 21904 14372 21916
rect 14424 21904 14430 21956
rect 15378 21944 15384 21956
rect 14844 21916 15384 21944
rect 14844 21876 14872 21916
rect 15378 21904 15384 21916
rect 15436 21904 15442 21956
rect 17218 21904 17224 21956
rect 17276 21944 17282 21956
rect 20088 21944 20116 21984
rect 22094 21972 22100 22024
rect 22152 22012 22158 22024
rect 22373 22015 22431 22021
rect 22373 22012 22385 22015
rect 22152 21984 22385 22012
rect 22152 21972 22158 21984
rect 22373 21981 22385 21984
rect 22419 21981 22431 22015
rect 22373 21975 22431 21981
rect 25130 21972 25136 22024
rect 25188 22012 25194 22024
rect 26620 22012 26648 22052
rect 29822 22040 29828 22052
rect 29880 22040 29886 22092
rect 30377 22083 30435 22089
rect 30377 22049 30389 22083
rect 30423 22080 30435 22083
rect 30466 22080 30472 22092
rect 30423 22052 30472 22080
rect 30423 22049 30435 22052
rect 30377 22043 30435 22049
rect 30466 22040 30472 22052
rect 30524 22040 30530 22092
rect 30852 22089 30880 22120
rect 30837 22083 30895 22089
rect 30837 22049 30849 22083
rect 30883 22049 30895 22083
rect 30944 22080 30972 22188
rect 31100 22185 31112 22219
rect 31146 22216 31158 22219
rect 31478 22216 31484 22228
rect 31146 22188 31484 22216
rect 31146 22185 31158 22188
rect 31100 22179 31158 22185
rect 31478 22176 31484 22188
rect 31536 22176 31542 22228
rect 34974 22216 34980 22228
rect 32232 22188 34980 22216
rect 32232 22148 32260 22188
rect 34974 22176 34980 22188
rect 35032 22176 35038 22228
rect 35342 22176 35348 22228
rect 35400 22216 35406 22228
rect 35400 22188 38424 22216
rect 35400 22176 35406 22188
rect 32140 22120 32260 22148
rect 33137 22151 33195 22157
rect 32140 22080 32168 22120
rect 33137 22117 33149 22151
rect 33183 22148 33195 22151
rect 34238 22148 34244 22160
rect 33183 22120 33640 22148
rect 33183 22117 33195 22120
rect 33137 22111 33195 22117
rect 30944 22052 32168 22080
rect 30837 22043 30895 22049
rect 32398 22040 32404 22092
rect 32456 22080 32462 22092
rect 32858 22080 32864 22092
rect 32456 22052 32864 22080
rect 32456 22040 32462 22052
rect 32858 22040 32864 22052
rect 32916 22040 32922 22092
rect 25188 21984 26648 22012
rect 25188 21972 25194 21984
rect 27154 21972 27160 22024
rect 27212 21972 27218 22024
rect 27614 21972 27620 22024
rect 27672 22012 27678 22024
rect 27672 21984 28028 22012
rect 27672 21972 27678 21984
rect 17276 21916 20116 21944
rect 21177 21947 21235 21953
rect 17276 21904 17282 21916
rect 21177 21913 21189 21947
rect 21223 21944 21235 21947
rect 21818 21944 21824 21956
rect 21223 21916 21824 21944
rect 21223 21913 21235 21916
rect 21177 21907 21235 21913
rect 21818 21904 21824 21916
rect 21876 21904 21882 21956
rect 22462 21904 22468 21956
rect 22520 21904 22526 21956
rect 24946 21904 24952 21956
rect 25004 21944 25010 21956
rect 25225 21947 25283 21953
rect 25225 21944 25237 21947
rect 25004 21916 25237 21944
rect 25004 21904 25010 21916
rect 25225 21913 25237 21916
rect 25271 21944 25283 21947
rect 25498 21944 25504 21956
rect 25271 21916 25504 21944
rect 25271 21913 25283 21916
rect 25225 21907 25283 21913
rect 25498 21904 25504 21916
rect 25556 21904 25562 21956
rect 25866 21904 25872 21956
rect 25924 21944 25930 21956
rect 27893 21947 27951 21953
rect 27893 21944 27905 21947
rect 25924 21916 27905 21944
rect 25924 21904 25930 21916
rect 27893 21913 27905 21916
rect 27939 21913 27951 21947
rect 28000 21944 28028 21984
rect 28442 21972 28448 22024
rect 28500 22012 28506 22024
rect 28537 22015 28595 22021
rect 28537 22012 28549 22015
rect 28500 21984 28549 22012
rect 28500 21972 28506 21984
rect 28537 21981 28549 21984
rect 28583 21981 28595 22015
rect 28537 21975 28595 21981
rect 29181 22015 29239 22021
rect 29181 21981 29193 22015
rect 29227 22012 29239 22015
rect 29733 22015 29791 22021
rect 29733 22012 29745 22015
rect 29227 21984 29745 22012
rect 29227 21981 29239 21984
rect 29181 21975 29239 21981
rect 29733 21981 29745 21984
rect 29779 21981 29791 22015
rect 29733 21975 29791 21981
rect 30006 21972 30012 22024
rect 30064 22012 30070 22024
rect 30282 22012 30288 22024
rect 30064 21984 30288 22012
rect 30064 21972 30070 21984
rect 30282 21972 30288 21984
rect 30340 21972 30346 22024
rect 33612 22012 33640 22120
rect 33888 22120 34244 22148
rect 33781 22083 33839 22089
rect 33781 22049 33793 22083
rect 33827 22080 33839 22083
rect 33888 22080 33916 22120
rect 34238 22108 34244 22120
rect 34296 22108 34302 22160
rect 34422 22108 34428 22160
rect 34480 22108 34486 22160
rect 35544 22094 35572 22188
rect 37369 22151 37427 22157
rect 37369 22117 37381 22151
rect 37415 22148 37427 22151
rect 38396 22148 38424 22188
rect 38470 22176 38476 22228
rect 38528 22216 38534 22228
rect 38565 22219 38623 22225
rect 38565 22216 38577 22219
rect 38528 22188 38577 22216
rect 38528 22176 38534 22188
rect 38565 22185 38577 22188
rect 38611 22185 38623 22219
rect 39022 22216 39028 22228
rect 38565 22179 38623 22185
rect 38672 22188 39028 22216
rect 38672 22148 38700 22188
rect 39022 22176 39028 22188
rect 39080 22176 39086 22228
rect 39390 22216 39396 22228
rect 39132 22188 39396 22216
rect 37415 22120 37872 22148
rect 38396 22120 38700 22148
rect 37415 22117 37427 22120
rect 37369 22111 37427 22117
rect 33827 22052 33916 22080
rect 35452 22089 35572 22094
rect 35452 22083 35587 22089
rect 35452 22052 35541 22083
rect 33827 22049 33839 22052
rect 33781 22043 33839 22049
rect 35529 22049 35541 22052
rect 35575 22049 35587 22083
rect 35529 22043 35587 22049
rect 36081 22083 36139 22089
rect 36081 22049 36093 22083
rect 36127 22080 36139 22083
rect 36354 22080 36360 22092
rect 36127 22052 36360 22080
rect 36127 22049 36139 22052
rect 36081 22043 36139 22049
rect 36354 22040 36360 22052
rect 36412 22040 36418 22092
rect 36814 22040 36820 22092
rect 36872 22040 36878 22092
rect 34606 22012 34612 22024
rect 33612 21984 34612 22012
rect 34606 21972 34612 21984
rect 34664 21972 34670 22024
rect 34974 21972 34980 22024
rect 35032 22012 35038 22024
rect 36633 22015 36691 22021
rect 36633 22012 36645 22015
rect 35032 21984 36645 22012
rect 35032 21972 35038 21984
rect 36633 21981 36645 21984
rect 36679 21981 36691 22015
rect 37737 22015 37795 22021
rect 37737 22012 37749 22015
rect 36633 21975 36691 21981
rect 36740 21984 37749 22012
rect 29086 21944 29092 21956
rect 28000 21916 29092 21944
rect 27893 21907 27951 21913
rect 29086 21904 29092 21916
rect 29144 21944 29150 21956
rect 31386 21944 31392 21956
rect 29144 21916 31392 21944
rect 29144 21904 29150 21916
rect 31386 21904 31392 21916
rect 31444 21904 31450 21956
rect 31754 21904 31760 21956
rect 31812 21904 31818 21956
rect 32490 21904 32496 21956
rect 32548 21944 32554 21956
rect 35345 21947 35403 21953
rect 35345 21944 35357 21947
rect 32548 21916 35357 21944
rect 32548 21904 32554 21916
rect 35345 21913 35357 21916
rect 35391 21913 35403 21947
rect 36740 21944 36768 21984
rect 37737 21981 37749 21984
rect 37783 21981 37795 22015
rect 37844 22012 37872 22120
rect 38838 22108 38844 22160
rect 38896 22148 38902 22160
rect 39132 22148 39160 22188
rect 39390 22176 39396 22188
rect 39448 22176 39454 22228
rect 39574 22176 39580 22228
rect 39632 22216 39638 22228
rect 44818 22216 44824 22228
rect 39632 22188 44824 22216
rect 39632 22176 39638 22188
rect 44818 22176 44824 22188
rect 44876 22176 44882 22228
rect 38896 22120 39160 22148
rect 38896 22108 38902 22120
rect 38013 22083 38071 22089
rect 38013 22049 38025 22083
rect 38059 22080 38071 22083
rect 38654 22080 38660 22092
rect 38059 22052 38660 22080
rect 38059 22049 38071 22052
rect 38013 22043 38071 22049
rect 38654 22040 38660 22052
rect 38712 22040 38718 22092
rect 39132 22089 39160 22120
rect 39206 22108 39212 22160
rect 39264 22148 39270 22160
rect 48498 22148 48504 22160
rect 39264 22120 39896 22148
rect 39264 22108 39270 22120
rect 39868 22092 39896 22120
rect 41800 22120 48504 22148
rect 39117 22083 39175 22089
rect 39117 22049 39129 22083
rect 39163 22080 39175 22083
rect 39163 22052 39197 22080
rect 39163 22049 39175 22052
rect 39117 22043 39175 22049
rect 39850 22040 39856 22092
rect 39908 22080 39914 22092
rect 41800 22089 41828 22120
rect 48498 22108 48504 22120
rect 48556 22108 48562 22160
rect 40681 22083 40739 22089
rect 40681 22080 40693 22083
rect 39908 22052 40693 22080
rect 39908 22040 39914 22052
rect 40681 22049 40693 22052
rect 40727 22080 40739 22083
rect 41785 22083 41843 22089
rect 41785 22080 41797 22083
rect 40727 22052 41797 22080
rect 40727 22049 40739 22052
rect 40681 22043 40739 22049
rect 41785 22049 41797 22052
rect 41831 22049 41843 22083
rect 41785 22043 41843 22049
rect 42242 22040 42248 22092
rect 42300 22080 42306 22092
rect 43073 22083 43131 22089
rect 42300 22052 42564 22080
rect 42300 22040 42306 22052
rect 41506 22012 41512 22024
rect 37844 21984 41512 22012
rect 37737 21975 37795 21981
rect 41506 21972 41512 21984
rect 41564 21972 41570 22024
rect 41690 21972 41696 22024
rect 41748 21972 41754 22024
rect 41874 21972 41880 22024
rect 41932 22012 41938 22024
rect 42429 22015 42487 22021
rect 42429 22012 42441 22015
rect 41932 21984 42441 22012
rect 41932 21972 41938 21984
rect 42429 21981 42441 21984
rect 42475 21981 42487 22015
rect 42536 22012 42564 22052
rect 43073 22049 43085 22083
rect 43119 22080 43131 22083
rect 43346 22080 43352 22092
rect 43119 22052 43352 22080
rect 43119 22049 43131 22052
rect 43073 22043 43131 22049
rect 43346 22040 43352 22052
rect 43404 22040 43410 22092
rect 44177 22083 44235 22089
rect 43456 22052 43760 22080
rect 42886 22012 42892 22024
rect 42536 21984 42892 22012
rect 42429 21975 42487 21981
rect 42886 21972 42892 21984
rect 42944 22012 42950 22024
rect 43456 22012 43484 22052
rect 42944 21984 43484 22012
rect 43533 22015 43591 22021
rect 42944 21972 42950 21984
rect 43533 21981 43545 22015
rect 43579 22012 43591 22015
rect 43622 22012 43628 22024
rect 43579 21984 43628 22012
rect 43579 21981 43591 21984
rect 43533 21975 43591 21981
rect 43622 21972 43628 21984
rect 43680 21972 43686 22024
rect 43732 22012 43760 22052
rect 44177 22049 44189 22083
rect 44223 22080 44235 22083
rect 44450 22080 44456 22092
rect 44223 22052 44456 22080
rect 44223 22049 44235 22052
rect 44177 22043 44235 22049
rect 44450 22040 44456 22052
rect 44508 22040 44514 22092
rect 44542 22040 44548 22092
rect 44600 22080 44606 22092
rect 44600 22052 46060 22080
rect 44600 22040 44606 22052
rect 46032 22024 46060 22052
rect 46198 22040 46204 22092
rect 46256 22080 46262 22092
rect 49421 22083 49479 22089
rect 49421 22080 49433 22083
rect 46256 22052 49433 22080
rect 46256 22040 46262 22052
rect 49421 22049 49433 22052
rect 49467 22049 49479 22083
rect 49421 22043 49479 22049
rect 44726 22012 44732 22024
rect 43732 21984 44732 22012
rect 44726 21972 44732 21984
rect 44784 21972 44790 22024
rect 45186 21972 45192 22024
rect 45244 21972 45250 22024
rect 46014 21972 46020 22024
rect 46072 21972 46078 22024
rect 46293 22015 46351 22021
rect 46293 21981 46305 22015
rect 46339 21981 46351 22015
rect 46293 21975 46351 21981
rect 35345 21907 35403 21913
rect 36188 21916 36768 21944
rect 13924 21848 14872 21876
rect 14918 21836 14924 21888
rect 14976 21876 14982 21888
rect 16761 21879 16819 21885
rect 16761 21876 16773 21879
rect 14976 21848 16773 21876
rect 14976 21836 14982 21848
rect 16761 21845 16773 21848
rect 16807 21845 16819 21879
rect 16761 21839 16819 21845
rect 17129 21879 17187 21885
rect 17129 21845 17141 21879
rect 17175 21876 17187 21879
rect 17494 21876 17500 21888
rect 17175 21848 17500 21876
rect 17175 21845 17187 21848
rect 17129 21839 17187 21845
rect 17494 21836 17500 21848
rect 17552 21836 17558 21888
rect 19334 21836 19340 21888
rect 19392 21836 19398 21888
rect 19610 21836 19616 21888
rect 19668 21836 19674 21888
rect 19978 21836 19984 21888
rect 20036 21876 20042 21888
rect 20073 21879 20131 21885
rect 20073 21876 20085 21879
rect 20036 21848 20085 21876
rect 20036 21836 20042 21848
rect 20073 21845 20085 21848
rect 20119 21876 20131 21879
rect 20346 21876 20352 21888
rect 20119 21848 20352 21876
rect 20119 21845 20131 21848
rect 20073 21839 20131 21845
rect 20346 21836 20352 21848
rect 20404 21836 20410 21888
rect 20806 21836 20812 21888
rect 20864 21836 20870 21888
rect 21269 21879 21327 21885
rect 21269 21845 21281 21879
rect 21315 21876 21327 21879
rect 21634 21876 21640 21888
rect 21315 21848 21640 21876
rect 21315 21845 21327 21848
rect 21269 21839 21327 21845
rect 21634 21836 21640 21848
rect 21692 21836 21698 21888
rect 22002 21836 22008 21888
rect 22060 21836 22066 21888
rect 23661 21879 23719 21885
rect 23661 21845 23673 21879
rect 23707 21876 23719 21879
rect 24118 21876 24124 21888
rect 23707 21848 24124 21876
rect 23707 21845 23719 21848
rect 23661 21839 23719 21845
rect 24118 21836 24124 21848
rect 24176 21836 24182 21888
rect 24486 21836 24492 21888
rect 24544 21836 24550 21888
rect 24762 21836 24768 21888
rect 24820 21836 24826 21888
rect 25958 21836 25964 21888
rect 26016 21836 26022 21888
rect 26326 21836 26332 21888
rect 26384 21836 26390 21888
rect 28902 21836 28908 21888
rect 28960 21876 28966 21888
rect 32585 21879 32643 21885
rect 32585 21876 32597 21879
rect 28960 21848 32597 21876
rect 28960 21836 28966 21848
rect 32585 21845 32597 21848
rect 32631 21876 32643 21879
rect 33410 21876 33416 21888
rect 32631 21848 33416 21876
rect 32631 21845 32643 21848
rect 32585 21839 32643 21845
rect 33410 21836 33416 21848
rect 33468 21836 33474 21888
rect 33502 21836 33508 21888
rect 33560 21836 33566 21888
rect 33597 21879 33655 21885
rect 33597 21845 33609 21879
rect 33643 21876 33655 21879
rect 33778 21876 33784 21888
rect 33643 21848 33784 21876
rect 33643 21845 33655 21848
rect 33597 21839 33655 21845
rect 33778 21836 33784 21848
rect 33836 21836 33842 21888
rect 33962 21836 33968 21888
rect 34020 21876 34026 21888
rect 34149 21879 34207 21885
rect 34149 21876 34161 21879
rect 34020 21848 34161 21876
rect 34020 21836 34026 21848
rect 34149 21845 34161 21848
rect 34195 21845 34207 21879
rect 34149 21839 34207 21845
rect 34330 21836 34336 21888
rect 34388 21876 34394 21888
rect 34885 21879 34943 21885
rect 34885 21876 34897 21879
rect 34388 21848 34897 21876
rect 34388 21836 34394 21848
rect 34885 21845 34897 21848
rect 34931 21845 34943 21879
rect 34885 21839 34943 21845
rect 35250 21836 35256 21888
rect 35308 21836 35314 21888
rect 36188 21885 36216 21916
rect 37274 21904 37280 21956
rect 37332 21944 37338 21956
rect 39025 21947 39083 21953
rect 39025 21944 39037 21947
rect 37332 21916 39037 21944
rect 37332 21904 37338 21916
rect 39025 21913 39037 21916
rect 39071 21944 39083 21947
rect 40310 21944 40316 21956
rect 39071 21916 40316 21944
rect 39071 21913 39083 21916
rect 39025 21907 39083 21913
rect 40310 21904 40316 21916
rect 40368 21904 40374 21956
rect 40402 21904 40408 21956
rect 40460 21944 40466 21956
rect 40862 21944 40868 21956
rect 40460 21916 40868 21944
rect 40460 21904 40466 21916
rect 40862 21904 40868 21916
rect 40920 21904 40926 21956
rect 41601 21947 41659 21953
rect 41601 21913 41613 21947
rect 41647 21944 41659 21947
rect 41782 21944 41788 21956
rect 41647 21916 41788 21944
rect 41647 21913 41659 21916
rect 41601 21907 41659 21913
rect 41782 21904 41788 21916
rect 41840 21904 41846 21956
rect 44174 21904 44180 21956
rect 44232 21944 44238 21956
rect 46308 21944 46336 21975
rect 46474 21972 46480 22024
rect 46532 22012 46538 22024
rect 47397 22015 47455 22021
rect 47397 22012 47409 22015
rect 46532 21984 47409 22012
rect 46532 21972 46538 21984
rect 47397 21981 47409 21984
rect 47443 21981 47455 22015
rect 47397 21975 47455 21981
rect 48314 21972 48320 22024
rect 48372 22012 48378 22024
rect 48501 22015 48559 22021
rect 48501 22012 48513 22015
rect 48372 21984 48513 22012
rect 48372 21972 48378 21984
rect 48501 21981 48513 21984
rect 48547 21981 48559 22015
rect 48501 21975 48559 21981
rect 48682 21972 48688 22024
rect 48740 22012 48746 22024
rect 49694 22012 49700 22024
rect 48740 21984 49700 22012
rect 48740 21972 48746 21984
rect 49694 21972 49700 21984
rect 49752 21972 49758 22024
rect 44232 21916 46336 21944
rect 44232 21904 44238 21916
rect 47118 21904 47124 21956
rect 47176 21944 47182 21956
rect 47670 21944 47676 21956
rect 47176 21916 47676 21944
rect 47176 21904 47182 21916
rect 47670 21904 47676 21916
rect 47728 21904 47734 21956
rect 36173 21879 36231 21885
rect 36173 21845 36185 21879
rect 36219 21845 36231 21879
rect 36173 21839 36231 21845
rect 36354 21836 36360 21888
rect 36412 21876 36418 21888
rect 36541 21879 36599 21885
rect 36541 21876 36553 21879
rect 36412 21848 36553 21876
rect 36412 21836 36418 21848
rect 36541 21845 36553 21848
rect 36587 21876 36599 21879
rect 36906 21876 36912 21888
rect 36587 21848 36912 21876
rect 36587 21845 36599 21848
rect 36541 21839 36599 21845
rect 36906 21836 36912 21848
rect 36964 21836 36970 21888
rect 37826 21836 37832 21888
rect 37884 21836 37890 21888
rect 37918 21836 37924 21888
rect 37976 21876 37982 21888
rect 38838 21876 38844 21888
rect 37976 21848 38844 21876
rect 37976 21836 37982 21848
rect 38838 21836 38844 21848
rect 38896 21876 38902 21888
rect 38933 21879 38991 21885
rect 38933 21876 38945 21879
rect 38896 21848 38945 21876
rect 38896 21836 38902 21848
rect 38933 21845 38945 21848
rect 38979 21845 38991 21879
rect 38933 21839 38991 21845
rect 39390 21836 39396 21888
rect 39448 21876 39454 21888
rect 39577 21879 39635 21885
rect 39577 21876 39589 21879
rect 39448 21848 39589 21876
rect 39448 21836 39454 21848
rect 39577 21845 39589 21848
rect 39623 21845 39635 21879
rect 39577 21839 39635 21845
rect 40034 21836 40040 21888
rect 40092 21836 40098 21888
rect 40494 21836 40500 21888
rect 40552 21836 40558 21888
rect 41230 21836 41236 21888
rect 41288 21836 41294 21888
rect 42150 21836 42156 21888
rect 42208 21876 42214 21888
rect 43714 21876 43720 21888
rect 42208 21848 43720 21876
rect 42208 21836 42214 21848
rect 43714 21836 43720 21848
rect 43772 21836 43778 21888
rect 44542 21836 44548 21888
rect 44600 21876 44606 21888
rect 44637 21879 44695 21885
rect 44637 21876 44649 21879
rect 44600 21848 44649 21876
rect 44600 21836 44606 21848
rect 44637 21845 44649 21848
rect 44683 21845 44695 21879
rect 44637 21839 44695 21845
rect 45554 21836 45560 21888
rect 45612 21876 45618 21888
rect 45833 21879 45891 21885
rect 45833 21876 45845 21879
rect 45612 21848 45845 21876
rect 45612 21836 45618 21848
rect 45833 21845 45845 21848
rect 45879 21845 45891 21879
rect 45833 21839 45891 21845
rect 46937 21879 46995 21885
rect 46937 21845 46949 21879
rect 46983 21876 46995 21879
rect 47302 21876 47308 21888
rect 46983 21848 47308 21876
rect 46983 21845 46995 21848
rect 46937 21839 46995 21845
rect 47302 21836 47308 21848
rect 47360 21836 47366 21888
rect 48041 21879 48099 21885
rect 48041 21845 48053 21879
rect 48087 21876 48099 21879
rect 48682 21876 48688 21888
rect 48087 21848 48688 21876
rect 48087 21845 48099 21848
rect 48041 21839 48099 21845
rect 48682 21836 48688 21848
rect 48740 21836 48746 21888
rect 49142 21836 49148 21888
rect 49200 21836 49206 21888
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 5994 21632 6000 21684
rect 6052 21632 6058 21684
rect 10134 21632 10140 21684
rect 10192 21632 10198 21684
rect 12710 21672 12716 21684
rect 10244 21644 12716 21672
rect 4338 21564 4344 21616
rect 4396 21564 4402 21616
rect 4430 21564 4436 21616
rect 4488 21604 4494 21616
rect 4488 21576 6592 21604
rect 4488 21564 4494 21576
rect 1765 21539 1823 21545
rect 1765 21505 1777 21539
rect 1811 21505 1823 21539
rect 1765 21499 1823 21505
rect 1780 21400 1808 21499
rect 2590 21496 2596 21548
rect 2648 21536 2654 21548
rect 3421 21539 3479 21545
rect 3421 21536 3433 21539
rect 2648 21508 3433 21536
rect 2648 21496 2654 21508
rect 3421 21505 3433 21508
rect 3467 21505 3479 21539
rect 3421 21499 3479 21505
rect 5353 21539 5411 21545
rect 5353 21505 5365 21539
rect 5399 21536 5411 21539
rect 5902 21536 5908 21548
rect 5399 21508 5908 21536
rect 5399 21505 5411 21508
rect 5353 21499 5411 21505
rect 5902 21496 5908 21508
rect 5960 21496 5966 21548
rect 6564 21545 6592 21576
rect 7926 21564 7932 21616
rect 7984 21604 7990 21616
rect 10244 21604 10272 21644
rect 12710 21632 12716 21644
rect 12768 21632 12774 21684
rect 12802 21632 12808 21684
rect 12860 21632 12866 21684
rect 13909 21675 13967 21681
rect 13909 21641 13921 21675
rect 13955 21672 13967 21675
rect 14182 21672 14188 21684
rect 13955 21644 14188 21672
rect 13955 21641 13967 21644
rect 13909 21635 13967 21641
rect 14182 21632 14188 21644
rect 14240 21632 14246 21684
rect 14274 21632 14280 21684
rect 14332 21672 14338 21684
rect 14369 21675 14427 21681
rect 14369 21672 14381 21675
rect 14332 21644 14381 21672
rect 14332 21632 14338 21644
rect 14369 21641 14381 21644
rect 14415 21641 14427 21675
rect 14369 21635 14427 21641
rect 14458 21632 14464 21684
rect 14516 21672 14522 21684
rect 15010 21672 15016 21684
rect 14516 21644 15016 21672
rect 14516 21632 14522 21644
rect 15010 21632 15016 21644
rect 15068 21632 15074 21684
rect 15102 21632 15108 21684
rect 15160 21672 15166 21684
rect 15933 21675 15991 21681
rect 15933 21672 15945 21675
rect 15160 21644 15945 21672
rect 15160 21632 15166 21644
rect 15933 21641 15945 21644
rect 15979 21641 15991 21675
rect 15933 21635 15991 21641
rect 16025 21675 16083 21681
rect 16025 21641 16037 21675
rect 16071 21672 16083 21675
rect 19610 21672 19616 21684
rect 16071 21644 19616 21672
rect 16071 21641 16083 21644
rect 16025 21635 16083 21641
rect 19610 21632 19616 21644
rect 19668 21632 19674 21684
rect 21634 21632 21640 21684
rect 21692 21672 21698 21684
rect 27157 21675 27215 21681
rect 27157 21672 27169 21675
rect 21692 21644 27169 21672
rect 21692 21632 21698 21644
rect 27157 21641 27169 21644
rect 27203 21641 27215 21675
rect 27157 21635 27215 21641
rect 28537 21675 28595 21681
rect 28537 21641 28549 21675
rect 28583 21672 28595 21675
rect 30650 21672 30656 21684
rect 28583 21644 30656 21672
rect 28583 21641 28595 21644
rect 28537 21635 28595 21641
rect 30650 21632 30656 21644
rect 30708 21632 30714 21684
rect 31570 21632 31576 21684
rect 31628 21672 31634 21684
rect 31754 21672 31760 21684
rect 31628 21644 31760 21672
rect 31628 21632 31634 21644
rect 31754 21632 31760 21644
rect 31812 21632 31818 21684
rect 31846 21632 31852 21684
rect 31904 21672 31910 21684
rect 32309 21675 32367 21681
rect 32309 21672 32321 21675
rect 31904 21644 32321 21672
rect 31904 21632 31910 21644
rect 32309 21641 32321 21644
rect 32355 21641 32367 21675
rect 32309 21635 32367 21641
rect 32490 21632 32496 21684
rect 32548 21632 32554 21684
rect 32677 21675 32735 21681
rect 32677 21641 32689 21675
rect 32723 21672 32735 21675
rect 32723 21644 33364 21672
rect 32723 21641 32735 21644
rect 32677 21635 32735 21641
rect 11698 21604 11704 21616
rect 7984 21576 10272 21604
rect 10428 21576 11704 21604
rect 7984 21564 7990 21576
rect 6549 21539 6607 21545
rect 6549 21505 6561 21539
rect 6595 21505 6607 21539
rect 6549 21499 6607 21505
rect 8389 21539 8447 21545
rect 8389 21505 8401 21539
rect 8435 21505 8447 21539
rect 8389 21499 8447 21505
rect 2777 21471 2835 21477
rect 2777 21437 2789 21471
rect 2823 21468 2835 21471
rect 3326 21468 3332 21480
rect 2823 21440 3332 21468
rect 2823 21437 2835 21440
rect 2777 21431 2835 21437
rect 3326 21428 3332 21440
rect 3384 21428 3390 21480
rect 5626 21428 5632 21480
rect 5684 21468 5690 21480
rect 7009 21471 7067 21477
rect 7009 21468 7021 21471
rect 5684 21440 7021 21468
rect 5684 21428 5690 21440
rect 7009 21437 7021 21440
rect 7055 21437 7067 21471
rect 7009 21431 7067 21437
rect 7558 21400 7564 21412
rect 1780 21372 7564 21400
rect 7558 21360 7564 21372
rect 7616 21360 7622 21412
rect 3142 21292 3148 21344
rect 3200 21332 3206 21344
rect 3970 21332 3976 21344
rect 3200 21304 3976 21332
rect 3200 21292 3206 21304
rect 3970 21292 3976 21304
rect 4028 21292 4034 21344
rect 5626 21292 5632 21344
rect 5684 21332 5690 21344
rect 8404 21332 8432 21499
rect 9030 21496 9036 21548
rect 9088 21536 9094 21548
rect 10428 21536 10456 21576
rect 11698 21564 11704 21576
rect 11756 21564 11762 21616
rect 17218 21604 17224 21616
rect 12176 21576 17224 21604
rect 9088 21508 10456 21536
rect 10505 21539 10563 21545
rect 9088 21496 9094 21508
rect 10505 21505 10517 21539
rect 10551 21536 10563 21539
rect 12176 21536 12204 21576
rect 17218 21564 17224 21576
rect 17276 21564 17282 21616
rect 18138 21564 18144 21616
rect 18196 21564 18202 21616
rect 18598 21564 18604 21616
rect 18656 21564 18662 21616
rect 20346 21564 20352 21616
rect 20404 21604 20410 21616
rect 22002 21604 22008 21616
rect 20404 21576 22008 21604
rect 20404 21564 20410 21576
rect 22002 21564 22008 21576
rect 22060 21564 22066 21616
rect 22278 21564 22284 21616
rect 22336 21564 22342 21616
rect 22370 21564 22376 21616
rect 22428 21604 22434 21616
rect 25866 21604 25872 21616
rect 22428 21576 22770 21604
rect 25806 21576 25872 21604
rect 22428 21564 22434 21576
rect 25866 21564 25872 21576
rect 25924 21564 25930 21616
rect 26142 21564 26148 21616
rect 26200 21604 26206 21616
rect 26697 21607 26755 21613
rect 26697 21604 26709 21607
rect 26200 21576 26709 21604
rect 26200 21564 26206 21576
rect 26697 21573 26709 21576
rect 26743 21604 26755 21607
rect 27338 21604 27344 21616
rect 26743 21576 27344 21604
rect 26743 21573 26755 21576
rect 26697 21567 26755 21573
rect 27338 21564 27344 21576
rect 27396 21564 27402 21616
rect 27617 21607 27675 21613
rect 27617 21573 27629 21607
rect 27663 21604 27675 21607
rect 28994 21604 29000 21616
rect 27663 21576 29000 21604
rect 27663 21573 27675 21576
rect 27617 21567 27675 21573
rect 28994 21564 29000 21576
rect 29052 21564 29058 21616
rect 30101 21607 30159 21613
rect 30101 21573 30113 21607
rect 30147 21604 30159 21607
rect 30374 21604 30380 21616
rect 30147 21576 30380 21604
rect 30147 21573 30159 21576
rect 30101 21567 30159 21573
rect 30374 21564 30380 21576
rect 30432 21564 30438 21616
rect 32030 21564 32036 21616
rect 32088 21604 32094 21616
rect 32508 21604 32536 21632
rect 32088 21576 32536 21604
rect 32769 21607 32827 21613
rect 32088 21564 32094 21576
rect 32769 21573 32781 21607
rect 32815 21604 32827 21607
rect 32950 21604 32956 21616
rect 32815 21576 32956 21604
rect 32815 21573 32827 21576
rect 32769 21567 32827 21573
rect 32950 21564 32956 21576
rect 33008 21564 33014 21616
rect 33336 21604 33364 21644
rect 33410 21632 33416 21684
rect 33468 21672 33474 21684
rect 35802 21672 35808 21684
rect 33468 21644 35808 21672
rect 33468 21632 33474 21644
rect 35802 21632 35808 21644
rect 35860 21632 35866 21684
rect 36081 21675 36139 21681
rect 36081 21641 36093 21675
rect 36127 21672 36139 21675
rect 36538 21672 36544 21684
rect 36127 21644 36544 21672
rect 36127 21641 36139 21644
rect 36081 21635 36139 21641
rect 36538 21632 36544 21644
rect 36596 21632 36602 21684
rect 37826 21632 37832 21684
rect 37884 21672 37890 21684
rect 40497 21675 40555 21681
rect 40497 21672 40509 21675
rect 37884 21644 40509 21672
rect 37884 21632 37890 21644
rect 40497 21641 40509 21644
rect 40543 21641 40555 21675
rect 40497 21635 40555 21641
rect 40865 21675 40923 21681
rect 40865 21641 40877 21675
rect 40911 21672 40923 21675
rect 41230 21672 41236 21684
rect 40911 21644 41236 21672
rect 40911 21641 40923 21644
rect 40865 21635 40923 21641
rect 41230 21632 41236 21644
rect 41288 21632 41294 21684
rect 41340 21644 42196 21672
rect 33336 21576 33548 21604
rect 10551 21508 12204 21536
rect 10551 21505 10563 21508
rect 10505 21499 10563 21505
rect 12250 21496 12256 21548
rect 12308 21496 12314 21548
rect 12526 21496 12532 21548
rect 12584 21536 12590 21548
rect 13265 21539 13323 21545
rect 13265 21536 13277 21539
rect 12584 21508 13277 21536
rect 12584 21496 12590 21508
rect 13265 21505 13277 21508
rect 13311 21505 13323 21539
rect 13265 21499 13323 21505
rect 14734 21496 14740 21548
rect 14792 21496 14798 21548
rect 14829 21539 14887 21545
rect 14829 21505 14841 21539
rect 14875 21536 14887 21539
rect 15562 21536 15568 21548
rect 14875 21508 15568 21536
rect 14875 21505 14887 21508
rect 14829 21499 14887 21505
rect 15562 21496 15568 21508
rect 15620 21496 15626 21548
rect 15838 21496 15844 21548
rect 15896 21536 15902 21548
rect 16666 21536 16672 21548
rect 15896 21508 16672 21536
rect 15896 21496 15902 21508
rect 16666 21496 16672 21508
rect 16724 21496 16730 21548
rect 16942 21496 16948 21548
rect 17000 21496 17006 21548
rect 20441 21539 20499 21545
rect 17052 21508 17816 21536
rect 8846 21428 8852 21480
rect 8904 21428 8910 21480
rect 11149 21471 11207 21477
rect 11149 21437 11161 21471
rect 11195 21468 11207 21471
rect 12066 21468 12072 21480
rect 11195 21440 12072 21468
rect 11195 21437 11207 21440
rect 11149 21431 11207 21437
rect 12066 21428 12072 21440
rect 12124 21428 12130 21480
rect 13906 21468 13912 21480
rect 12176 21440 13912 21468
rect 11793 21403 11851 21409
rect 11793 21400 11805 21403
rect 8864 21372 11805 21400
rect 8864 21344 8892 21372
rect 11793 21369 11805 21372
rect 11839 21400 11851 21403
rect 12176 21400 12204 21440
rect 13906 21428 13912 21440
rect 13964 21428 13970 21480
rect 14918 21428 14924 21480
rect 14976 21428 14982 21480
rect 15378 21428 15384 21480
rect 15436 21468 15442 21480
rect 16117 21471 16175 21477
rect 16117 21468 16129 21471
rect 15436 21440 16129 21468
rect 15436 21428 15442 21440
rect 16117 21437 16129 21440
rect 16163 21468 16175 21471
rect 17052 21468 17080 21508
rect 16163 21440 17080 21468
rect 17221 21471 17279 21477
rect 16163 21437 16175 21440
rect 16117 21431 16175 21437
rect 17221 21437 17233 21471
rect 17267 21468 17279 21471
rect 17310 21468 17316 21480
rect 17267 21440 17316 21468
rect 17267 21437 17279 21440
rect 17221 21431 17279 21437
rect 17310 21428 17316 21440
rect 17368 21468 17374 21480
rect 17678 21468 17684 21480
rect 17368 21440 17684 21468
rect 17368 21428 17374 21440
rect 17678 21428 17684 21440
rect 17736 21428 17742 21480
rect 11839 21372 12204 21400
rect 11839 21369 11851 21372
rect 11793 21363 11851 21369
rect 12250 21360 12256 21412
rect 12308 21400 12314 21412
rect 14936 21400 14964 21428
rect 17586 21400 17592 21412
rect 12308 21372 14964 21400
rect 15028 21372 17592 21400
rect 12308 21360 12314 21372
rect 5684 21304 8432 21332
rect 5684 21292 5690 21304
rect 8846 21292 8852 21344
rect 8904 21292 8910 21344
rect 11054 21292 11060 21344
rect 11112 21332 11118 21344
rect 11606 21332 11612 21344
rect 11112 21304 11612 21332
rect 11112 21292 11118 21304
rect 11606 21292 11612 21304
rect 11664 21292 11670 21344
rect 11698 21292 11704 21344
rect 11756 21332 11762 21344
rect 12618 21332 12624 21344
rect 11756 21304 12624 21332
rect 11756 21292 11762 21304
rect 12618 21292 12624 21304
rect 12676 21292 12682 21344
rect 12710 21292 12716 21344
rect 12768 21332 12774 21344
rect 15028 21332 15056 21372
rect 17586 21360 17592 21372
rect 17644 21360 17650 21412
rect 17788 21400 17816 21508
rect 20441 21505 20453 21539
rect 20487 21505 20499 21539
rect 20441 21499 20499 21505
rect 17862 21428 17868 21480
rect 17920 21428 17926 21480
rect 18230 21468 18236 21480
rect 17972 21440 18236 21468
rect 17972 21400 18000 21440
rect 18230 21428 18236 21440
rect 18288 21428 18294 21480
rect 18782 21428 18788 21480
rect 18840 21468 18846 21480
rect 19613 21471 19671 21477
rect 19613 21468 19625 21471
rect 18840 21440 19625 21468
rect 18840 21428 18846 21440
rect 19613 21437 19625 21440
rect 19659 21437 19671 21471
rect 20456 21468 20484 21499
rect 21082 21496 21088 21548
rect 21140 21536 21146 21548
rect 21453 21539 21511 21545
rect 21453 21536 21465 21539
rect 21140 21508 21465 21536
rect 21140 21496 21146 21508
rect 21453 21505 21465 21508
rect 21499 21536 21511 21539
rect 21910 21536 21916 21548
rect 21499 21508 21916 21536
rect 21499 21505 21511 21508
rect 21453 21499 21511 21505
rect 21910 21496 21916 21508
rect 21968 21496 21974 21548
rect 23750 21496 23756 21548
rect 23808 21536 23814 21548
rect 24118 21536 24124 21548
rect 23808 21508 24124 21536
rect 23808 21496 23814 21508
rect 24118 21496 24124 21508
rect 24176 21496 24182 21548
rect 24302 21496 24308 21548
rect 24360 21496 24366 21548
rect 26513 21539 26571 21545
rect 26513 21536 26525 21539
rect 25792 21508 26525 21536
rect 19613 21431 19671 21437
rect 19720 21440 20484 21468
rect 17788 21372 18000 21400
rect 19150 21360 19156 21412
rect 19208 21400 19214 21412
rect 19720 21400 19748 21440
rect 20530 21428 20536 21480
rect 20588 21428 20594 21480
rect 20717 21471 20775 21477
rect 20717 21437 20729 21471
rect 20763 21437 20775 21471
rect 20717 21431 20775 21437
rect 19208 21372 19748 21400
rect 19208 21360 19214 21372
rect 19794 21360 19800 21412
rect 19852 21400 19858 21412
rect 20732 21400 20760 21431
rect 21266 21428 21272 21480
rect 21324 21468 21330 21480
rect 22005 21471 22063 21477
rect 22005 21468 22017 21471
rect 21324 21440 22017 21468
rect 21324 21428 21330 21440
rect 22005 21437 22017 21440
rect 22051 21437 22063 21471
rect 22278 21468 22284 21480
rect 22005 21431 22063 21437
rect 22112 21440 22284 21468
rect 21634 21400 21640 21412
rect 19852 21372 21640 21400
rect 19852 21360 19858 21372
rect 21634 21360 21640 21372
rect 21692 21400 21698 21412
rect 22112 21400 22140 21440
rect 22278 21428 22284 21440
rect 22336 21428 22342 21480
rect 22646 21428 22652 21480
rect 22704 21468 22710 21480
rect 24581 21471 24639 21477
rect 24581 21468 24593 21471
rect 22704 21440 24593 21468
rect 22704 21428 22710 21440
rect 24581 21437 24593 21440
rect 24627 21437 24639 21471
rect 24581 21431 24639 21437
rect 25130 21428 25136 21480
rect 25188 21468 25194 21480
rect 25792 21468 25820 21508
rect 26513 21505 26525 21508
rect 26559 21536 26571 21539
rect 27525 21539 27583 21545
rect 26559 21508 27016 21536
rect 26559 21505 26571 21508
rect 26513 21499 26571 21505
rect 25188 21440 25820 21468
rect 25188 21428 25194 21440
rect 26326 21428 26332 21480
rect 26384 21468 26390 21480
rect 26878 21468 26884 21480
rect 26384 21440 26884 21468
rect 26384 21428 26390 21440
rect 26878 21428 26884 21440
rect 26936 21428 26942 21480
rect 26988 21468 27016 21508
rect 27525 21505 27537 21539
rect 27571 21536 27583 21539
rect 28810 21536 28816 21548
rect 27571 21508 28816 21536
rect 27571 21505 27583 21508
rect 27525 21499 27583 21505
rect 28810 21496 28816 21508
rect 28868 21496 28874 21548
rect 28905 21539 28963 21545
rect 28905 21505 28917 21539
rect 28951 21536 28963 21539
rect 29730 21536 29736 21548
rect 28951 21508 29736 21536
rect 28951 21505 28963 21508
rect 28905 21499 28963 21505
rect 29730 21496 29736 21508
rect 29788 21496 29794 21548
rect 30193 21539 30251 21545
rect 30193 21505 30205 21539
rect 30239 21536 30251 21539
rect 30926 21536 30932 21548
rect 30239 21508 30932 21536
rect 30239 21505 30251 21508
rect 30193 21499 30251 21505
rect 30926 21496 30932 21508
rect 30984 21496 30990 21548
rect 31297 21539 31355 21545
rect 31297 21505 31309 21539
rect 31343 21536 31355 21539
rect 31570 21536 31576 21548
rect 31343 21508 31576 21536
rect 31343 21505 31355 21508
rect 31297 21499 31355 21505
rect 31570 21496 31576 21508
rect 31628 21496 31634 21548
rect 27709 21471 27767 21477
rect 27709 21468 27721 21471
rect 26988 21440 27721 21468
rect 27709 21437 27721 21440
rect 27755 21437 27767 21471
rect 27709 21431 27767 21437
rect 27798 21428 27804 21480
rect 27856 21468 27862 21480
rect 28997 21471 29055 21477
rect 28997 21468 29009 21471
rect 27856 21440 29009 21468
rect 27856 21428 27862 21440
rect 28997 21437 29009 21440
rect 29043 21437 29055 21471
rect 28997 21431 29055 21437
rect 29089 21471 29147 21477
rect 29089 21437 29101 21471
rect 29135 21437 29147 21471
rect 29089 21431 29147 21437
rect 21692 21372 22140 21400
rect 21692 21360 21698 21372
rect 23382 21360 23388 21412
rect 23440 21400 23446 21412
rect 23658 21400 23664 21412
rect 23440 21372 23664 21400
rect 23440 21360 23446 21372
rect 23658 21360 23664 21372
rect 23716 21360 23722 21412
rect 23753 21403 23811 21409
rect 23753 21369 23765 21403
rect 23799 21400 23811 21403
rect 24302 21400 24308 21412
rect 23799 21372 24308 21400
rect 23799 21369 23811 21372
rect 23753 21363 23811 21369
rect 24302 21360 24308 21372
rect 24360 21360 24366 21412
rect 26418 21400 26424 21412
rect 26068 21372 26424 21400
rect 12768 21304 15056 21332
rect 15565 21335 15623 21341
rect 12768 21292 12774 21304
rect 15565 21301 15577 21335
rect 15611 21332 15623 21335
rect 15654 21332 15660 21344
rect 15611 21304 15660 21332
rect 15611 21301 15623 21304
rect 15565 21295 15623 21301
rect 15654 21292 15660 21304
rect 15712 21292 15718 21344
rect 15746 21292 15752 21344
rect 15804 21332 15810 21344
rect 17218 21332 17224 21344
rect 15804 21304 17224 21332
rect 15804 21292 15810 21304
rect 17218 21292 17224 21304
rect 17276 21292 17282 21344
rect 17310 21292 17316 21344
rect 17368 21332 17374 21344
rect 20073 21335 20131 21341
rect 20073 21332 20085 21335
rect 17368 21304 20085 21332
rect 17368 21292 17374 21304
rect 20073 21301 20085 21304
rect 20119 21301 20131 21335
rect 20073 21295 20131 21301
rect 21269 21335 21327 21341
rect 21269 21301 21281 21335
rect 21315 21332 21327 21335
rect 22094 21332 22100 21344
rect 21315 21304 22100 21332
rect 21315 21301 21327 21304
rect 21269 21295 21327 21301
rect 22094 21292 22100 21304
rect 22152 21292 22158 21344
rect 22738 21292 22744 21344
rect 22796 21332 22802 21344
rect 22922 21332 22928 21344
rect 22796 21304 22928 21332
rect 22796 21292 22802 21304
rect 22922 21292 22928 21304
rect 22980 21292 22986 21344
rect 23676 21332 23704 21360
rect 26068 21341 26096 21372
rect 26418 21360 26424 21372
rect 26476 21360 26482 21412
rect 27614 21360 27620 21412
rect 27672 21400 27678 21412
rect 28902 21400 28908 21412
rect 27672 21372 28908 21400
rect 27672 21360 27678 21372
rect 28902 21360 28908 21372
rect 28960 21400 28966 21412
rect 29104 21400 29132 21431
rect 29270 21428 29276 21480
rect 29328 21468 29334 21480
rect 30006 21468 30012 21480
rect 29328 21440 30012 21468
rect 29328 21428 29334 21440
rect 30006 21428 30012 21440
rect 30064 21468 30070 21480
rect 30285 21471 30343 21477
rect 30285 21468 30297 21471
rect 30064 21440 30297 21468
rect 30064 21428 30070 21440
rect 30285 21437 30297 21440
rect 30331 21437 30343 21471
rect 30285 21431 30343 21437
rect 30374 21428 30380 21480
rect 30432 21468 30438 21480
rect 30650 21468 30656 21480
rect 30432 21440 30656 21468
rect 30432 21428 30438 21440
rect 30650 21428 30656 21440
rect 30708 21428 30714 21480
rect 31386 21428 31392 21480
rect 31444 21428 31450 21480
rect 31478 21428 31484 21480
rect 31536 21428 31542 21480
rect 32861 21471 32919 21477
rect 32861 21468 32873 21471
rect 31588 21440 32873 21468
rect 28960 21372 29132 21400
rect 28960 21360 28966 21372
rect 29454 21360 29460 21412
rect 29512 21400 29518 21412
rect 31588 21400 31616 21440
rect 32861 21437 32873 21440
rect 32907 21437 32919 21471
rect 33520 21468 33548 21576
rect 34054 21564 34060 21616
rect 34112 21564 34118 21616
rect 36262 21564 36268 21616
rect 36320 21604 36326 21616
rect 38470 21604 38476 21616
rect 36320 21576 38476 21604
rect 36320 21564 36326 21576
rect 33594 21496 33600 21548
rect 33652 21536 33658 21548
rect 33781 21539 33839 21545
rect 33781 21536 33793 21539
rect 33652 21508 33793 21536
rect 33652 21496 33658 21508
rect 33781 21505 33793 21508
rect 33827 21505 33839 21539
rect 33781 21499 33839 21505
rect 35158 21496 35164 21548
rect 35216 21536 35222 21548
rect 35618 21536 35624 21548
rect 35216 21508 35624 21536
rect 35216 21496 35222 21508
rect 35618 21496 35624 21508
rect 35676 21496 35682 21548
rect 36354 21496 36360 21548
rect 36412 21536 36418 21548
rect 36449 21539 36507 21545
rect 36449 21536 36461 21539
rect 36412 21508 36461 21536
rect 36412 21496 36418 21508
rect 36449 21505 36461 21508
rect 36495 21505 36507 21539
rect 36449 21499 36507 21505
rect 35250 21468 35256 21480
rect 33520 21440 35256 21468
rect 32861 21431 32919 21437
rect 35250 21428 35256 21440
rect 35308 21428 35314 21480
rect 36262 21428 36268 21480
rect 36320 21468 36326 21480
rect 36648 21477 36676 21576
rect 38470 21564 38476 21576
rect 38528 21564 38534 21616
rect 38562 21564 38568 21616
rect 38620 21564 38626 21616
rect 40034 21564 40040 21616
rect 40092 21604 40098 21616
rect 40957 21607 41015 21613
rect 40957 21604 40969 21607
rect 40092 21576 40969 21604
rect 40092 21564 40098 21576
rect 40957 21573 40969 21576
rect 41003 21573 41015 21607
rect 40957 21567 41015 21573
rect 37642 21496 37648 21548
rect 37700 21496 37706 21548
rect 37826 21496 37832 21548
rect 37884 21496 37890 21548
rect 36541 21471 36599 21477
rect 36541 21468 36553 21471
rect 36320 21440 36553 21468
rect 36320 21428 36326 21440
rect 36541 21437 36553 21440
rect 36587 21437 36599 21471
rect 36541 21431 36599 21437
rect 36633 21471 36691 21477
rect 36633 21437 36645 21471
rect 36679 21437 36691 21471
rect 37274 21468 37280 21480
rect 36633 21431 36691 21437
rect 36740 21440 37280 21468
rect 29512 21372 31616 21400
rect 29512 21360 29518 21372
rect 32398 21360 32404 21412
rect 32456 21400 32462 21412
rect 33594 21400 33600 21412
rect 32456 21372 33600 21400
rect 32456 21360 32462 21372
rect 33594 21360 33600 21372
rect 33652 21360 33658 21412
rect 36740 21400 36768 21440
rect 37274 21428 37280 21440
rect 37332 21428 37338 21480
rect 37458 21428 37464 21480
rect 37516 21468 37522 21480
rect 38289 21471 38347 21477
rect 38289 21468 38301 21471
rect 37516 21440 38301 21468
rect 37516 21428 37522 21440
rect 38289 21437 38301 21440
rect 38335 21437 38347 21471
rect 38289 21431 38347 21437
rect 38562 21428 38568 21480
rect 38620 21468 38626 21480
rect 39022 21468 39028 21480
rect 38620 21440 39028 21468
rect 38620 21428 38626 21440
rect 39022 21428 39028 21440
rect 39080 21428 39086 21480
rect 39114 21428 39120 21480
rect 39172 21468 39178 21480
rect 39684 21468 39712 21522
rect 39942 21496 39948 21548
rect 40000 21536 40006 21548
rect 40000 21508 40264 21536
rect 40000 21496 40006 21508
rect 40236 21468 40264 21508
rect 40402 21496 40408 21548
rect 40460 21536 40466 21548
rect 41340 21536 41368 21644
rect 41598 21564 41604 21616
rect 41656 21604 41662 21616
rect 42061 21607 42119 21613
rect 42061 21604 42073 21607
rect 41656 21576 42073 21604
rect 41656 21564 41662 21576
rect 42061 21573 42073 21576
rect 42107 21573 42119 21607
rect 42168 21604 42196 21644
rect 42518 21632 42524 21684
rect 42576 21672 42582 21684
rect 44361 21675 44419 21681
rect 44361 21672 44373 21675
rect 42576 21644 44373 21672
rect 42576 21632 42582 21644
rect 44361 21641 44373 21644
rect 44407 21641 44419 21675
rect 44361 21635 44419 21641
rect 45462 21632 45468 21684
rect 45520 21672 45526 21684
rect 46474 21672 46480 21684
rect 45520 21644 46480 21672
rect 45520 21632 45526 21644
rect 46474 21632 46480 21644
rect 46532 21632 46538 21684
rect 46566 21632 46572 21684
rect 46624 21632 46630 21684
rect 47026 21632 47032 21684
rect 47084 21632 47090 21684
rect 47394 21632 47400 21684
rect 47452 21672 47458 21684
rect 47670 21672 47676 21684
rect 47452 21644 47676 21672
rect 47452 21632 47458 21644
rect 47670 21632 47676 21644
rect 47728 21632 47734 21684
rect 49050 21632 49056 21684
rect 49108 21632 49114 21684
rect 44450 21604 44456 21616
rect 42168 21576 44456 21604
rect 42061 21567 42119 21573
rect 44450 21564 44456 21576
rect 44508 21564 44514 21616
rect 49142 21604 49148 21616
rect 45940 21576 49148 21604
rect 40460 21508 41368 21536
rect 41877 21539 41935 21545
rect 42518 21540 42524 21548
rect 40460 21496 40466 21508
rect 41877 21505 41889 21539
rect 41923 21536 41935 21539
rect 42444 21536 42524 21540
rect 41923 21512 42524 21536
rect 41923 21508 42472 21512
rect 41923 21505 41935 21508
rect 41877 21499 41935 21505
rect 42518 21496 42524 21512
rect 42576 21496 42582 21548
rect 42613 21540 42671 21545
rect 42613 21539 42748 21540
rect 42613 21505 42625 21539
rect 42659 21536 42748 21539
rect 42794 21536 42800 21548
rect 42659 21512 42800 21536
rect 42659 21505 42671 21512
rect 42720 21508 42800 21512
rect 42613 21499 42671 21505
rect 42794 21496 42800 21508
rect 42852 21496 42858 21548
rect 43714 21496 43720 21548
rect 43772 21496 43778 21548
rect 44818 21496 44824 21548
rect 44876 21496 44882 21548
rect 45940 21545 45968 21576
rect 49142 21564 49148 21576
rect 49200 21564 49206 21616
rect 45925 21539 45983 21545
rect 45925 21505 45937 21539
rect 45971 21505 45983 21539
rect 47213 21539 47271 21545
rect 47213 21536 47225 21539
rect 45925 21499 45983 21505
rect 46032 21508 47225 21536
rect 41049 21471 41107 21477
rect 39172 21440 40172 21468
rect 40236 21440 40908 21468
rect 39172 21428 39178 21440
rect 35452 21372 36768 21400
rect 26053 21335 26111 21341
rect 26053 21332 26065 21335
rect 23676 21304 26065 21332
rect 26053 21301 26065 21304
rect 26099 21301 26111 21335
rect 26053 21295 26111 21301
rect 26326 21292 26332 21344
rect 26384 21292 26390 21344
rect 26602 21292 26608 21344
rect 26660 21332 26666 21344
rect 28166 21332 28172 21344
rect 26660 21304 28172 21332
rect 26660 21292 26666 21304
rect 28166 21292 28172 21304
rect 28224 21292 28230 21344
rect 28261 21335 28319 21341
rect 28261 21301 28273 21335
rect 28307 21332 28319 21335
rect 28350 21332 28356 21344
rect 28307 21304 28356 21332
rect 28307 21301 28319 21304
rect 28261 21295 28319 21301
rect 28350 21292 28356 21304
rect 28408 21292 28414 21344
rect 28626 21292 28632 21344
rect 28684 21332 28690 21344
rect 29733 21335 29791 21341
rect 29733 21332 29745 21335
rect 28684 21304 29745 21332
rect 28684 21292 28690 21304
rect 29733 21301 29745 21304
rect 29779 21301 29791 21335
rect 29733 21295 29791 21301
rect 30374 21292 30380 21344
rect 30432 21332 30438 21344
rect 30929 21335 30987 21341
rect 30929 21332 30941 21335
rect 30432 21304 30941 21332
rect 30432 21292 30438 21304
rect 30929 21301 30941 21304
rect 30975 21301 30987 21335
rect 30929 21295 30987 21301
rect 33778 21292 33784 21344
rect 33836 21332 33842 21344
rect 35452 21332 35480 21372
rect 36814 21360 36820 21412
rect 36872 21400 36878 21412
rect 36872 21372 38424 21400
rect 36872 21360 36878 21372
rect 33836 21304 35480 21332
rect 33836 21292 33842 21304
rect 35526 21292 35532 21344
rect 35584 21292 35590 21344
rect 36354 21292 36360 21344
rect 36412 21332 36418 21344
rect 37182 21332 37188 21344
rect 36412 21304 37188 21332
rect 36412 21292 36418 21304
rect 37182 21292 37188 21304
rect 37240 21292 37246 21344
rect 38396 21332 38424 21372
rect 39942 21360 39948 21412
rect 40000 21400 40006 21412
rect 40037 21403 40095 21409
rect 40037 21400 40049 21403
rect 40000 21372 40049 21400
rect 40000 21360 40006 21372
rect 40037 21369 40049 21372
rect 40083 21369 40095 21403
rect 40144 21400 40172 21440
rect 40880 21400 40908 21440
rect 41049 21437 41061 21471
rect 41095 21437 41107 21471
rect 41049 21431 41107 21437
rect 41064 21400 41092 21431
rect 41506 21428 41512 21480
rect 41564 21468 41570 21480
rect 46032 21468 46060 21508
rect 47213 21505 47225 21508
rect 47259 21505 47271 21539
rect 47213 21499 47271 21505
rect 47486 21496 47492 21548
rect 47544 21536 47550 21548
rect 47765 21539 47823 21545
rect 47765 21536 47777 21539
rect 47544 21508 47777 21536
rect 47544 21496 47550 21508
rect 47765 21505 47777 21508
rect 47811 21505 47823 21539
rect 47765 21499 47823 21505
rect 48961 21539 49019 21545
rect 48961 21505 48973 21539
rect 49007 21505 49019 21539
rect 48961 21499 49019 21505
rect 41564 21440 46060 21468
rect 41564 21428 41570 21440
rect 47946 21428 47952 21480
rect 48004 21468 48010 21480
rect 48976 21468 49004 21499
rect 48004 21440 49004 21468
rect 48004 21428 48010 21440
rect 41230 21400 41236 21412
rect 40144 21372 40356 21400
rect 40880 21372 41236 21400
rect 40037 21363 40095 21369
rect 39960 21332 39988 21360
rect 38396 21304 39988 21332
rect 40328 21332 40356 21372
rect 41230 21360 41236 21372
rect 41288 21360 41294 21412
rect 42150 21400 42156 21412
rect 41340 21372 42156 21400
rect 41340 21332 41368 21372
rect 42150 21360 42156 21372
rect 42208 21360 42214 21412
rect 42518 21360 42524 21412
rect 42576 21400 42582 21412
rect 45186 21400 45192 21412
rect 42576 21372 45192 21400
rect 42576 21360 42582 21372
rect 45186 21360 45192 21372
rect 45244 21360 45250 21412
rect 45465 21403 45523 21409
rect 45465 21369 45477 21403
rect 45511 21400 45523 21403
rect 47762 21400 47768 21412
rect 45511 21372 47768 21400
rect 45511 21369 45523 21372
rect 45465 21363 45523 21369
rect 47762 21360 47768 21372
rect 47820 21360 47826 21412
rect 40328 21304 41368 21332
rect 42058 21292 42064 21344
rect 42116 21332 42122 21344
rect 43257 21335 43315 21341
rect 43257 21332 43269 21335
rect 42116 21304 43269 21332
rect 42116 21292 42122 21304
rect 43257 21301 43269 21304
rect 43303 21301 43315 21335
rect 43257 21295 43315 21301
rect 47394 21292 47400 21344
rect 47452 21332 47458 21344
rect 48409 21335 48467 21341
rect 48409 21332 48421 21335
rect 47452 21304 48421 21332
rect 47452 21292 47458 21304
rect 48409 21301 48421 21304
rect 48455 21301 48467 21335
rect 48409 21295 48467 21301
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 9490 21128 9496 21140
rect 2746 21100 9496 21128
rect 2746 20992 2774 21100
rect 9490 21088 9496 21100
rect 9548 21088 9554 21140
rect 10318 21088 10324 21140
rect 10376 21088 10382 21140
rect 11425 21131 11483 21137
rect 11425 21097 11437 21131
rect 11471 21128 11483 21131
rect 11514 21128 11520 21140
rect 11471 21100 11520 21128
rect 11471 21097 11483 21100
rect 11425 21091 11483 21097
rect 11514 21088 11520 21100
rect 11572 21088 11578 21140
rect 12526 21088 12532 21140
rect 12584 21088 12590 21140
rect 16942 21128 16948 21140
rect 12636 21100 16948 21128
rect 3421 21063 3479 21069
rect 3421 21029 3433 21063
rect 3467 21060 3479 21063
rect 6362 21060 6368 21072
rect 3467 21032 6368 21060
rect 3467 21029 3479 21032
rect 3421 21023 3479 21029
rect 6362 21020 6368 21032
rect 6420 21020 6426 21072
rect 9033 21063 9091 21069
rect 9033 21029 9045 21063
rect 9079 21060 9091 21063
rect 12636 21060 12664 21100
rect 16942 21088 16948 21100
rect 17000 21088 17006 21140
rect 17218 21088 17224 21140
rect 17276 21128 17282 21140
rect 19794 21128 19800 21140
rect 17276 21100 19800 21128
rect 17276 21088 17282 21100
rect 19794 21088 19800 21100
rect 19852 21088 19858 21140
rect 19978 21088 19984 21140
rect 20036 21128 20042 21140
rect 21726 21128 21732 21140
rect 20036 21100 21732 21128
rect 20036 21088 20042 21100
rect 21726 21088 21732 21100
rect 21784 21088 21790 21140
rect 22002 21088 22008 21140
rect 22060 21128 22066 21140
rect 23293 21131 23351 21137
rect 23293 21128 23305 21131
rect 22060 21100 23305 21128
rect 22060 21088 22066 21100
rect 23293 21097 23305 21100
rect 23339 21097 23351 21131
rect 23293 21091 23351 21097
rect 24673 21131 24731 21137
rect 24673 21097 24685 21131
rect 24719 21128 24731 21131
rect 27798 21128 27804 21140
rect 24719 21100 27804 21128
rect 24719 21097 24731 21100
rect 24673 21091 24731 21097
rect 27798 21088 27804 21100
rect 27856 21088 27862 21140
rect 28166 21088 28172 21140
rect 28224 21128 28230 21140
rect 28224 21100 28764 21128
rect 28224 21088 28230 21100
rect 21082 21060 21088 21072
rect 9079 21032 12664 21060
rect 13740 21032 14596 21060
rect 9079 21029 9091 21032
rect 9033 21023 9091 21029
rect 1780 20964 2774 20992
rect 1780 20933 1808 20964
rect 4154 20952 4160 21004
rect 4212 20992 4218 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 4212 20964 4445 20992
rect 4212 20952 4218 20964
rect 4433 20961 4445 20964
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 6730 20952 6736 21004
rect 6788 20952 6794 21004
rect 8573 20995 8631 21001
rect 8573 20961 8585 20995
rect 8619 20992 8631 20995
rect 8619 20964 10824 20992
rect 8619 20961 8631 20964
rect 8573 20955 8631 20961
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20893 1823 20927
rect 1765 20887 1823 20893
rect 4065 20927 4123 20933
rect 4065 20893 4077 20927
rect 4111 20924 4123 20927
rect 4706 20924 4712 20936
rect 4111 20896 4712 20924
rect 4111 20893 4123 20896
rect 4065 20887 4123 20893
rect 4706 20884 4712 20896
rect 4764 20884 4770 20936
rect 5166 20884 5172 20936
rect 5224 20924 5230 20936
rect 5813 20927 5871 20933
rect 5813 20924 5825 20927
rect 5224 20896 5825 20924
rect 5224 20884 5230 20896
rect 5813 20893 5825 20896
rect 5859 20893 5871 20927
rect 7926 20924 7932 20936
rect 5813 20887 5871 20893
rect 6748 20896 7932 20924
rect 6748 20868 6776 20896
rect 7926 20884 7932 20896
rect 7984 20884 7990 20936
rect 9309 20927 9367 20933
rect 9309 20893 9321 20927
rect 9355 20924 9367 20927
rect 9355 20896 9628 20924
rect 9355 20893 9367 20896
rect 9309 20887 9367 20893
rect 2777 20859 2835 20865
rect 2777 20825 2789 20859
rect 2823 20856 2835 20859
rect 2866 20856 2872 20868
rect 2823 20828 2872 20856
rect 2823 20825 2835 20828
rect 2777 20819 2835 20825
rect 2866 20816 2872 20828
rect 2924 20816 2930 20868
rect 6730 20816 6736 20868
rect 6788 20816 6794 20868
rect 9600 20856 9628 20896
rect 9674 20884 9680 20936
rect 9732 20884 9738 20936
rect 10796 20933 10824 20964
rect 11330 20952 11336 21004
rect 11388 20992 11394 21004
rect 13538 20992 13544 21004
rect 11388 20964 13544 20992
rect 11388 20952 11394 20964
rect 13538 20952 13544 20964
rect 13596 20952 13602 21004
rect 10781 20927 10839 20933
rect 10781 20893 10793 20927
rect 10827 20893 10839 20927
rect 10781 20887 10839 20893
rect 11885 20927 11943 20933
rect 11885 20893 11897 20927
rect 11931 20924 11943 20927
rect 13740 20924 13768 21032
rect 13814 20952 13820 21004
rect 13872 20992 13878 21004
rect 14458 20992 14464 21004
rect 13872 20964 14464 20992
rect 13872 20952 13878 20964
rect 14458 20952 14464 20964
rect 14516 20952 14522 21004
rect 14568 20992 14596 21032
rect 16132 21032 21088 21060
rect 16022 20992 16028 21004
rect 14568 20964 16028 20992
rect 16022 20952 16028 20964
rect 16080 20952 16086 21004
rect 11931 20896 13768 20924
rect 11931 20893 11943 20896
rect 11885 20887 11943 20893
rect 14090 20884 14096 20936
rect 14148 20884 14154 20936
rect 15838 20884 15844 20936
rect 15896 20884 15902 20936
rect 11146 20856 11152 20868
rect 7576 20828 9444 20856
rect 9600 20828 11152 20856
rect 3605 20791 3663 20797
rect 3605 20757 3617 20791
rect 3651 20788 3663 20791
rect 7576 20788 7604 20828
rect 3651 20760 7604 20788
rect 3651 20757 3663 20760
rect 3605 20751 3663 20757
rect 7650 20748 7656 20800
rect 7708 20748 7714 20800
rect 9217 20791 9275 20797
rect 9217 20757 9229 20791
rect 9263 20788 9275 20791
rect 9306 20788 9312 20800
rect 9263 20760 9312 20788
rect 9263 20757 9275 20760
rect 9217 20751 9275 20757
rect 9306 20748 9312 20760
rect 9364 20748 9370 20800
rect 9416 20788 9444 20828
rect 11146 20816 11152 20828
rect 11204 20816 11210 20868
rect 11606 20816 11612 20868
rect 11664 20856 11670 20868
rect 12805 20859 12863 20865
rect 12805 20856 12817 20859
rect 11664 20828 12817 20856
rect 11664 20816 11670 20828
rect 12805 20825 12817 20828
rect 12851 20856 12863 20859
rect 13357 20859 13415 20865
rect 13357 20856 13369 20859
rect 12851 20828 13369 20856
rect 12851 20825 12863 20828
rect 12805 20819 12863 20825
rect 13357 20825 13369 20828
rect 13403 20825 13415 20859
rect 13357 20819 13415 20825
rect 13449 20859 13507 20865
rect 13449 20825 13461 20859
rect 13495 20856 13507 20859
rect 14642 20856 14648 20868
rect 13495 20828 14648 20856
rect 13495 20825 13507 20828
rect 13449 20819 13507 20825
rect 14642 20816 14648 20828
rect 14700 20816 14706 20868
rect 14737 20859 14795 20865
rect 14737 20825 14749 20859
rect 14783 20856 14795 20859
rect 15010 20856 15016 20868
rect 14783 20828 15016 20856
rect 14783 20825 14795 20828
rect 14737 20819 14795 20825
rect 15010 20816 15016 20828
rect 15068 20816 15074 20868
rect 9766 20788 9772 20800
rect 9416 20760 9772 20788
rect 9766 20748 9772 20760
rect 9824 20748 9830 20800
rect 10318 20748 10324 20800
rect 10376 20788 10382 20800
rect 12250 20788 12256 20800
rect 10376 20760 12256 20788
rect 10376 20748 10382 20760
rect 12250 20748 12256 20760
rect 12308 20748 12314 20800
rect 12986 20748 12992 20800
rect 13044 20748 13050 20800
rect 13906 20748 13912 20800
rect 13964 20788 13970 20800
rect 16132 20788 16160 21032
rect 21082 21020 21088 21032
rect 21140 21020 21146 21072
rect 25958 21060 25964 21072
rect 23768 21032 25964 21060
rect 17402 20952 17408 21004
rect 17460 20952 17466 21004
rect 17497 20995 17555 21001
rect 17497 20961 17509 20995
rect 17543 20992 17555 20995
rect 18690 20992 18696 21004
rect 17543 20964 18696 20992
rect 17543 20961 17555 20964
rect 17497 20955 17555 20961
rect 17310 20884 17316 20936
rect 17368 20884 17374 20936
rect 16758 20816 16764 20868
rect 16816 20856 16822 20868
rect 17512 20856 17540 20955
rect 18690 20952 18696 20964
rect 18748 20952 18754 21004
rect 18782 20952 18788 21004
rect 18840 20952 18846 21004
rect 19978 20952 19984 21004
rect 20036 20952 20042 21004
rect 20070 20952 20076 21004
rect 20128 20992 20134 21004
rect 20165 20995 20223 21001
rect 20165 20992 20177 20995
rect 20128 20964 20177 20992
rect 20128 20952 20134 20964
rect 20165 20961 20177 20964
rect 20211 20992 20223 20995
rect 21361 20995 21419 21001
rect 20211 20964 20944 20992
rect 20211 20961 20223 20964
rect 20165 20955 20223 20961
rect 18601 20927 18659 20933
rect 18601 20893 18613 20927
rect 18647 20924 18659 20927
rect 20806 20924 20812 20936
rect 18647 20896 20812 20924
rect 18647 20893 18659 20896
rect 18601 20887 18659 20893
rect 20806 20884 20812 20896
rect 20864 20884 20870 20936
rect 16816 20828 17540 20856
rect 18509 20859 18567 20865
rect 16816 20816 16822 20828
rect 18509 20825 18521 20859
rect 18555 20856 18567 20859
rect 19242 20856 19248 20868
rect 18555 20828 19248 20856
rect 18555 20825 18567 20828
rect 18509 20819 18567 20825
rect 19242 20816 19248 20828
rect 19300 20816 19306 20868
rect 19889 20859 19947 20865
rect 19889 20825 19901 20859
rect 19935 20856 19947 20859
rect 19935 20828 20852 20856
rect 19935 20825 19947 20828
rect 19889 20819 19947 20825
rect 20824 20800 20852 20828
rect 13964 20760 16160 20788
rect 13964 20748 13970 20760
rect 16206 20748 16212 20800
rect 16264 20748 16270 20800
rect 16666 20748 16672 20800
rect 16724 20748 16730 20800
rect 16942 20748 16948 20800
rect 17000 20748 17006 20800
rect 18141 20791 18199 20797
rect 18141 20757 18153 20791
rect 18187 20788 18199 20791
rect 19058 20788 19064 20800
rect 18187 20760 19064 20788
rect 18187 20757 18199 20760
rect 18141 20751 18199 20757
rect 19058 20748 19064 20760
rect 19116 20748 19122 20800
rect 19426 20748 19432 20800
rect 19484 20788 19490 20800
rect 19521 20791 19579 20797
rect 19521 20788 19533 20791
rect 19484 20760 19533 20788
rect 19484 20748 19490 20760
rect 19521 20757 19533 20760
rect 19567 20757 19579 20791
rect 19521 20751 19579 20757
rect 20254 20748 20260 20800
rect 20312 20788 20318 20800
rect 20533 20791 20591 20797
rect 20533 20788 20545 20791
rect 20312 20760 20545 20788
rect 20312 20748 20318 20760
rect 20533 20757 20545 20760
rect 20579 20757 20591 20791
rect 20533 20751 20591 20757
rect 20622 20748 20628 20800
rect 20680 20788 20686 20800
rect 20717 20791 20775 20797
rect 20717 20788 20729 20791
rect 20680 20760 20729 20788
rect 20680 20748 20686 20760
rect 20717 20757 20729 20760
rect 20763 20757 20775 20791
rect 20717 20751 20775 20757
rect 20806 20748 20812 20800
rect 20864 20748 20870 20800
rect 20916 20788 20944 20964
rect 21361 20961 21373 20995
rect 21407 20992 21419 20995
rect 21450 20992 21456 21004
rect 21407 20964 21456 20992
rect 21407 20961 21419 20964
rect 21361 20955 21419 20961
rect 21450 20952 21456 20964
rect 21508 20952 21514 21004
rect 21726 20952 21732 21004
rect 21784 20992 21790 21004
rect 23768 20992 23796 21032
rect 25958 21020 25964 21032
rect 26016 21020 26022 21072
rect 28626 21060 28632 21072
rect 26344 21032 28632 21060
rect 21784 20964 23796 20992
rect 21784 20952 21790 20964
rect 23842 20952 23848 21004
rect 23900 20952 23906 21004
rect 24486 20952 24492 21004
rect 24544 20992 24550 21004
rect 25225 20995 25283 21001
rect 25225 20992 25237 20995
rect 24544 20964 25237 20992
rect 24544 20952 24550 20964
rect 25225 20961 25237 20964
rect 25271 20961 25283 20995
rect 25225 20955 25283 20961
rect 21082 20884 21088 20936
rect 21140 20884 21146 20936
rect 22646 20884 22652 20936
rect 22704 20924 22710 20936
rect 23661 20927 23719 20933
rect 23661 20924 23673 20927
rect 22704 20896 23673 20924
rect 22704 20884 22710 20896
rect 23661 20893 23673 20896
rect 23707 20924 23719 20927
rect 24578 20924 24584 20936
rect 23707 20896 24584 20924
rect 23707 20893 23719 20896
rect 23661 20887 23719 20893
rect 24578 20884 24584 20896
rect 24636 20884 24642 20936
rect 25130 20924 25136 20936
rect 24688 20896 25136 20924
rect 22738 20856 22744 20868
rect 22586 20828 22744 20856
rect 22738 20816 22744 20828
rect 22796 20816 22802 20868
rect 23290 20816 23296 20868
rect 23348 20856 23354 20868
rect 23842 20856 23848 20868
rect 23348 20828 23848 20856
rect 23348 20816 23354 20828
rect 23842 20816 23848 20828
rect 23900 20856 23906 20868
rect 24210 20856 24216 20868
rect 23900 20828 24216 20856
rect 23900 20816 23906 20828
rect 24210 20816 24216 20828
rect 24268 20856 24274 20868
rect 24688 20856 24716 20896
rect 25130 20884 25136 20896
rect 25188 20884 25194 20936
rect 25240 20924 25268 20955
rect 25314 20952 25320 21004
rect 25372 20992 25378 21004
rect 25590 20992 25596 21004
rect 25372 20964 25596 20992
rect 25372 20952 25378 20964
rect 25590 20952 25596 20964
rect 25648 20952 25654 21004
rect 26344 21001 26372 21032
rect 28626 21020 28632 21032
rect 28684 21020 28690 21072
rect 28736 21060 28764 21100
rect 28810 21088 28816 21140
rect 28868 21088 28874 21140
rect 30190 21128 30196 21140
rect 28920 21100 30196 21128
rect 28920 21060 28948 21100
rect 30190 21088 30196 21100
rect 30248 21088 30254 21140
rect 30929 21131 30987 21137
rect 30929 21097 30941 21131
rect 30975 21128 30987 21131
rect 32030 21128 32036 21140
rect 30975 21100 32036 21128
rect 30975 21097 30987 21100
rect 30929 21091 30987 21097
rect 32030 21088 32036 21100
rect 32088 21088 32094 21140
rect 33778 21128 33784 21140
rect 32140 21100 33784 21128
rect 28736 21032 28948 21060
rect 30208 21060 30236 21088
rect 30208 21032 30328 21060
rect 26329 20995 26387 21001
rect 26329 20961 26341 20995
rect 26375 20961 26387 20995
rect 26329 20955 26387 20961
rect 26418 20952 26424 21004
rect 26476 20952 26482 21004
rect 27338 20952 27344 21004
rect 27396 20992 27402 21004
rect 27985 20995 28043 21001
rect 27985 20992 27997 20995
rect 27396 20964 27997 20992
rect 27396 20952 27402 20964
rect 27985 20961 27997 20964
rect 28031 20961 28043 20995
rect 30190 20992 30196 21004
rect 27985 20955 28043 20961
rect 28644 20964 30196 20992
rect 28644 20924 28672 20964
rect 30190 20952 30196 20964
rect 30248 20952 30254 21004
rect 30300 21001 30328 21032
rect 31386 21020 31392 21072
rect 31444 21060 31450 21072
rect 32140 21060 32168 21100
rect 33778 21088 33784 21100
rect 33836 21088 33842 21140
rect 34054 21088 34060 21140
rect 34112 21128 34118 21140
rect 40037 21131 40095 21137
rect 34112 21100 39988 21128
rect 34112 21088 34118 21100
rect 33686 21060 33692 21072
rect 31444 21032 32168 21060
rect 32508 21032 33692 21060
rect 31444 21020 31450 21032
rect 30285 20995 30343 21001
rect 30285 20961 30297 20995
rect 30331 20961 30343 20995
rect 30285 20955 30343 20961
rect 31573 20995 31631 21001
rect 31573 20961 31585 20995
rect 31619 20961 31631 20995
rect 31573 20955 31631 20961
rect 25240 20896 26464 20924
rect 24268 20828 24716 20856
rect 24268 20816 24274 20828
rect 24762 20816 24768 20868
rect 24820 20856 24826 20868
rect 25774 20856 25780 20868
rect 24820 20828 25780 20856
rect 24820 20816 24826 20828
rect 25774 20816 25780 20828
rect 25832 20816 25838 20868
rect 22833 20791 22891 20797
rect 22833 20788 22845 20791
rect 20916 20760 22845 20788
rect 22833 20757 22845 20760
rect 22879 20757 22891 20791
rect 22833 20751 22891 20757
rect 22922 20748 22928 20800
rect 22980 20788 22986 20800
rect 23382 20788 23388 20800
rect 22980 20760 23388 20788
rect 22980 20748 22986 20760
rect 23382 20748 23388 20760
rect 23440 20788 23446 20800
rect 23753 20791 23811 20797
rect 23753 20788 23765 20791
rect 23440 20760 23765 20788
rect 23440 20748 23446 20760
rect 23753 20757 23765 20760
rect 23799 20757 23811 20791
rect 23753 20751 23811 20757
rect 24302 20748 24308 20800
rect 24360 20788 24366 20800
rect 25041 20791 25099 20797
rect 25041 20788 25053 20791
rect 24360 20760 25053 20788
rect 24360 20748 24366 20760
rect 25041 20757 25053 20760
rect 25087 20757 25099 20791
rect 25041 20751 25099 20757
rect 25130 20748 25136 20800
rect 25188 20748 25194 20800
rect 25314 20748 25320 20800
rect 25372 20788 25378 20800
rect 25869 20791 25927 20797
rect 25869 20788 25881 20791
rect 25372 20760 25881 20788
rect 25372 20748 25378 20760
rect 25869 20757 25881 20760
rect 25915 20757 25927 20791
rect 25869 20751 25927 20757
rect 26234 20748 26240 20800
rect 26292 20748 26298 20800
rect 26436 20788 26464 20896
rect 26896 20896 28672 20924
rect 26896 20788 26924 20896
rect 28718 20884 28724 20936
rect 28776 20884 28782 20936
rect 29822 20884 29828 20936
rect 29880 20924 29886 20936
rect 30101 20927 30159 20933
rect 30101 20924 30113 20927
rect 29880 20896 30113 20924
rect 29880 20884 29886 20896
rect 30101 20893 30113 20896
rect 30147 20893 30159 20927
rect 31588 20924 31616 20955
rect 32508 20924 32536 21032
rect 33686 21020 33692 21032
rect 33744 21020 33750 21072
rect 39960 21060 39988 21100
rect 40037 21097 40049 21131
rect 40083 21128 40095 21131
rect 40126 21128 40132 21140
rect 40083 21100 40132 21128
rect 40083 21097 40095 21100
rect 40037 21091 40095 21097
rect 40126 21088 40132 21100
rect 40184 21088 40190 21140
rect 41230 21088 41236 21140
rect 41288 21128 41294 21140
rect 41288 21100 41552 21128
rect 41288 21088 41294 21100
rect 41414 21060 41420 21072
rect 39960 21032 41420 21060
rect 41414 21020 41420 21032
rect 41472 21020 41478 21072
rect 41524 21060 41552 21100
rect 41874 21088 41880 21140
rect 41932 21088 41938 21140
rect 47854 21128 47860 21140
rect 41984 21100 47860 21128
rect 41984 21060 42012 21100
rect 47854 21088 47860 21100
rect 47912 21128 47918 21140
rect 49421 21131 49479 21137
rect 49421 21128 49433 21131
rect 47912 21100 49433 21128
rect 47912 21088 47918 21100
rect 49421 21097 49433 21100
rect 49467 21097 49479 21131
rect 49421 21091 49479 21097
rect 41524 21032 42012 21060
rect 44266 21020 44272 21072
rect 44324 21060 44330 21072
rect 48041 21063 48099 21069
rect 48041 21060 48053 21063
rect 44324 21032 48053 21060
rect 44324 21020 44330 21032
rect 48041 21029 48053 21032
rect 48087 21029 48099 21063
rect 48041 21023 48099 21029
rect 32582 20952 32588 21004
rect 32640 20952 32646 21004
rect 32769 20995 32827 21001
rect 32769 20961 32781 20995
rect 32815 20961 32827 20995
rect 32769 20955 32827 20961
rect 31588 20896 32536 20924
rect 32784 20924 32812 20955
rect 33502 20952 33508 21004
rect 33560 20992 33566 21004
rect 33873 20995 33931 21001
rect 33873 20992 33885 20995
rect 33560 20964 33885 20992
rect 33560 20952 33566 20964
rect 33873 20961 33885 20964
rect 33919 20961 33931 20995
rect 33873 20955 33931 20961
rect 34882 20952 34888 21004
rect 34940 20952 34946 21004
rect 35161 20995 35219 21001
rect 35161 20961 35173 20995
rect 35207 20992 35219 20995
rect 36170 20992 36176 21004
rect 35207 20964 36176 20992
rect 35207 20961 35219 20964
rect 35161 20955 35219 20961
rect 36170 20952 36176 20964
rect 36228 20952 36234 21004
rect 37458 20952 37464 21004
rect 37516 20992 37522 21004
rect 37737 20995 37795 21001
rect 37737 20992 37749 20995
rect 37516 20964 37749 20992
rect 37516 20952 37522 20964
rect 37737 20961 37749 20964
rect 37783 20961 37795 20995
rect 37737 20955 37795 20961
rect 38013 20995 38071 21001
rect 38013 20961 38025 20995
rect 38059 20992 38071 20995
rect 38746 20992 38752 21004
rect 38059 20964 38752 20992
rect 38059 20961 38071 20964
rect 38013 20955 38071 20961
rect 38746 20952 38752 20964
rect 38804 20952 38810 21004
rect 39022 20952 39028 21004
rect 39080 20992 39086 21004
rect 40681 20995 40739 21001
rect 40681 20992 40693 20995
rect 39080 20964 40693 20992
rect 39080 20952 39086 20964
rect 40681 20961 40693 20964
rect 40727 20992 40739 20995
rect 40727 20964 42472 20992
rect 40727 20961 40739 20964
rect 40681 20955 40739 20961
rect 34054 20924 34060 20936
rect 32784 20896 34060 20924
rect 30101 20887 30159 20893
rect 34054 20884 34060 20896
rect 34112 20884 34118 20936
rect 39114 20884 39120 20936
rect 39172 20884 39178 20936
rect 41138 20884 41144 20936
rect 41196 20924 41202 20936
rect 41233 20927 41291 20933
rect 41233 20924 41245 20927
rect 41196 20896 41245 20924
rect 41196 20884 41202 20896
rect 41233 20893 41245 20896
rect 41279 20893 41291 20927
rect 41233 20887 41291 20893
rect 41414 20884 41420 20936
rect 41472 20924 41478 20936
rect 42337 20927 42395 20933
rect 42337 20924 42349 20927
rect 41472 20896 42349 20924
rect 41472 20884 41478 20896
rect 42337 20893 42349 20896
rect 42383 20893 42395 20927
rect 42444 20924 42472 20964
rect 42518 20952 42524 21004
rect 42576 20992 42582 21004
rect 44361 20995 44419 21001
rect 44361 20992 44373 20995
rect 42576 20964 44373 20992
rect 42576 20952 42582 20964
rect 44361 20961 44373 20964
rect 44407 20961 44419 20995
rect 45278 20992 45284 21004
rect 44361 20955 44419 20961
rect 44468 20964 45284 20992
rect 42444 20896 43392 20924
rect 42337 20887 42395 20893
rect 27801 20859 27859 20865
rect 27801 20825 27813 20859
rect 27847 20856 27859 20859
rect 29181 20859 29239 20865
rect 29181 20856 29193 20859
rect 27847 20828 29193 20856
rect 27847 20825 27859 20828
rect 27801 20819 27859 20825
rect 29181 20825 29193 20828
rect 29227 20856 29239 20859
rect 30926 20856 30932 20868
rect 29227 20828 30932 20856
rect 29227 20825 29239 20828
rect 29181 20819 29239 20825
rect 30926 20816 30932 20828
rect 30984 20816 30990 20868
rect 31202 20816 31208 20868
rect 31260 20856 31266 20868
rect 31297 20859 31355 20865
rect 31297 20856 31309 20859
rect 31260 20828 31309 20856
rect 31260 20816 31266 20828
rect 31297 20825 31309 20828
rect 31343 20856 31355 20859
rect 31343 20828 31524 20856
rect 31343 20825 31355 20828
rect 31297 20819 31355 20825
rect 26436 20760 26924 20788
rect 26970 20748 26976 20800
rect 27028 20748 27034 20800
rect 27062 20748 27068 20800
rect 27120 20748 27126 20800
rect 27154 20748 27160 20800
rect 27212 20788 27218 20800
rect 27433 20791 27491 20797
rect 27433 20788 27445 20791
rect 27212 20760 27445 20788
rect 27212 20748 27218 20760
rect 27433 20757 27445 20760
rect 27479 20757 27491 20791
rect 27433 20751 27491 20757
rect 27893 20791 27951 20797
rect 27893 20757 27905 20791
rect 27939 20788 27951 20791
rect 28902 20788 28908 20800
rect 27939 20760 28908 20788
rect 27939 20757 27951 20760
rect 27893 20751 27951 20757
rect 28902 20748 28908 20760
rect 28960 20748 28966 20800
rect 28994 20748 29000 20800
rect 29052 20788 29058 20800
rect 29362 20788 29368 20800
rect 29052 20760 29368 20788
rect 29052 20748 29058 20760
rect 29362 20748 29368 20760
rect 29420 20748 29426 20800
rect 29546 20748 29552 20800
rect 29604 20788 29610 20800
rect 29733 20791 29791 20797
rect 29733 20788 29745 20791
rect 29604 20760 29745 20788
rect 29604 20748 29610 20760
rect 29733 20757 29745 20760
rect 29779 20757 29791 20791
rect 29733 20751 29791 20757
rect 30193 20791 30251 20797
rect 30193 20757 30205 20791
rect 30239 20788 30251 20791
rect 30282 20788 30288 20800
rect 30239 20760 30288 20788
rect 30239 20757 30251 20760
rect 30193 20751 30251 20757
rect 30282 20748 30288 20760
rect 30340 20748 30346 20800
rect 31386 20748 31392 20800
rect 31444 20748 31450 20800
rect 31496 20788 31524 20828
rect 31570 20816 31576 20868
rect 31628 20856 31634 20868
rect 33689 20859 33747 20865
rect 33689 20856 33701 20859
rect 31628 20828 33701 20856
rect 31628 20816 31634 20828
rect 33689 20825 33701 20828
rect 33735 20856 33747 20859
rect 33735 20828 35572 20856
rect 33735 20825 33747 20828
rect 33689 20819 33747 20825
rect 31662 20788 31668 20800
rect 31496 20760 31668 20788
rect 31662 20748 31668 20760
rect 31720 20748 31726 20800
rect 32122 20748 32128 20800
rect 32180 20748 32186 20800
rect 32490 20748 32496 20800
rect 32548 20748 32554 20800
rect 33318 20748 33324 20800
rect 33376 20748 33382 20800
rect 33778 20748 33784 20800
rect 33836 20748 33842 20800
rect 34422 20748 34428 20800
rect 34480 20748 34486 20800
rect 35544 20788 35572 20828
rect 35618 20816 35624 20868
rect 35676 20816 35682 20868
rect 38286 20856 38292 20868
rect 36556 20828 38292 20856
rect 36556 20788 36584 20828
rect 38286 20816 38292 20828
rect 38344 20816 38350 20868
rect 43364 20856 43392 20896
rect 43438 20884 43444 20936
rect 43496 20884 43502 20936
rect 44468 20924 44496 20964
rect 45278 20952 45284 20964
rect 45336 20952 45342 21004
rect 45830 20952 45836 21004
rect 45888 20952 45894 21004
rect 43548 20896 44496 20924
rect 44637 20927 44695 20933
rect 43548 20856 43576 20896
rect 44637 20893 44649 20927
rect 44683 20924 44695 20927
rect 45002 20924 45008 20936
rect 44683 20896 45008 20924
rect 44683 20893 44695 20896
rect 44637 20887 44695 20893
rect 45002 20884 45008 20896
rect 45060 20884 45066 20936
rect 45094 20884 45100 20936
rect 45152 20924 45158 20936
rect 45189 20927 45247 20933
rect 45189 20924 45201 20927
rect 45152 20896 45201 20924
rect 45152 20884 45158 20896
rect 45189 20893 45201 20896
rect 45235 20893 45247 20927
rect 45189 20887 45247 20893
rect 45462 20884 45468 20936
rect 45520 20924 45526 20936
rect 46293 20927 46351 20933
rect 46293 20924 46305 20927
rect 45520 20896 46305 20924
rect 45520 20884 45526 20896
rect 46293 20893 46305 20896
rect 46339 20893 46351 20927
rect 46293 20887 46351 20893
rect 46658 20884 46664 20936
rect 46716 20924 46722 20936
rect 46934 20924 46940 20936
rect 46716 20896 46940 20924
rect 46716 20884 46722 20896
rect 46934 20884 46940 20896
rect 46992 20884 46998 20936
rect 47394 20884 47400 20936
rect 47452 20884 47458 20936
rect 48498 20884 48504 20936
rect 48556 20924 48562 20936
rect 50430 20924 50436 20936
rect 48556 20896 50436 20924
rect 48556 20884 48562 20896
rect 50430 20884 50436 20896
rect 50488 20884 50494 20936
rect 39500 20828 43300 20856
rect 43364 20828 43576 20856
rect 44085 20859 44143 20865
rect 35544 20760 36584 20788
rect 36630 20748 36636 20800
rect 36688 20748 36694 20800
rect 37090 20748 37096 20800
rect 37148 20748 37154 20800
rect 38654 20748 38660 20800
rect 38712 20788 38718 20800
rect 39500 20797 39528 20828
rect 39485 20791 39543 20797
rect 39485 20788 39497 20791
rect 38712 20760 39497 20788
rect 38712 20748 38718 20760
rect 39485 20757 39497 20760
rect 39531 20757 39543 20791
rect 39485 20751 39543 20757
rect 39758 20748 39764 20800
rect 39816 20788 39822 20800
rect 40405 20791 40463 20797
rect 40405 20788 40417 20791
rect 39816 20760 40417 20788
rect 39816 20748 39822 20760
rect 40405 20757 40417 20760
rect 40451 20757 40463 20791
rect 40405 20751 40463 20757
rect 40497 20791 40555 20797
rect 40497 20757 40509 20791
rect 40543 20788 40555 20791
rect 41506 20788 41512 20800
rect 40543 20760 41512 20788
rect 40543 20757 40555 20760
rect 40497 20751 40555 20757
rect 41506 20748 41512 20760
rect 41564 20748 41570 20800
rect 42978 20748 42984 20800
rect 43036 20748 43042 20800
rect 43272 20788 43300 20828
rect 44085 20825 44097 20859
rect 44131 20856 44143 20859
rect 45922 20856 45928 20868
rect 44131 20828 44496 20856
rect 44131 20825 44143 20828
rect 44085 20819 44143 20825
rect 44174 20788 44180 20800
rect 43272 20760 44180 20788
rect 44174 20748 44180 20760
rect 44232 20748 44238 20800
rect 44468 20788 44496 20828
rect 44652 20828 45928 20856
rect 44652 20788 44680 20828
rect 45922 20816 45928 20828
rect 45980 20816 45986 20868
rect 46566 20816 46572 20868
rect 46624 20856 46630 20868
rect 47946 20856 47952 20868
rect 46624 20828 47952 20856
rect 46624 20816 46630 20828
rect 47946 20816 47952 20828
rect 48004 20816 48010 20868
rect 44468 20760 44680 20788
rect 44726 20748 44732 20800
rect 44784 20748 44790 20800
rect 46934 20748 46940 20800
rect 46992 20748 46998 20800
rect 48498 20748 48504 20800
rect 48556 20788 48562 20800
rect 49145 20791 49203 20797
rect 49145 20788 49157 20791
rect 48556 20760 49157 20788
rect 48556 20748 48562 20760
rect 49145 20757 49157 20760
rect 49191 20757 49203 20791
rect 49145 20751 49203 20757
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 50062 20680 50068 20732
rect 50120 20720 50126 20732
rect 50246 20720 50252 20732
rect 50120 20692 50252 20720
rect 50120 20680 50126 20692
rect 50246 20680 50252 20692
rect 50304 20680 50310 20732
rect 1104 20624 49864 20646
rect 3510 20544 3516 20596
rect 3568 20584 3574 20596
rect 5997 20587 6055 20593
rect 5997 20584 6009 20587
rect 3568 20556 6009 20584
rect 3568 20544 3574 20556
rect 5997 20553 6009 20556
rect 6043 20553 6055 20587
rect 9674 20584 9680 20596
rect 5997 20547 6055 20553
rect 6196 20556 9680 20584
rect 4982 20516 4988 20528
rect 1780 20488 4988 20516
rect 1780 20457 1808 20488
rect 4982 20476 4988 20488
rect 5040 20476 5046 20528
rect 6196 20516 6224 20556
rect 9674 20544 9680 20556
rect 9732 20544 9738 20596
rect 11149 20587 11207 20593
rect 11149 20553 11161 20587
rect 11195 20584 11207 20587
rect 20714 20584 20720 20596
rect 11195 20556 18736 20584
rect 11195 20553 11207 20556
rect 11149 20547 11207 20553
rect 5368 20488 6224 20516
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20417 1823 20451
rect 1765 20411 1823 20417
rect 3602 20408 3608 20460
rect 3660 20408 3666 20460
rect 5368 20457 5396 20488
rect 6270 20476 6276 20528
rect 6328 20516 6334 20528
rect 6328 20488 7052 20516
rect 6328 20476 6334 20488
rect 5353 20451 5411 20457
rect 5353 20417 5365 20451
rect 5399 20417 5411 20451
rect 5353 20411 5411 20417
rect 6549 20451 6607 20457
rect 6549 20417 6561 20451
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 2774 20340 2780 20392
rect 2832 20340 2838 20392
rect 3878 20340 3884 20392
rect 3936 20340 3942 20392
rect 2682 20272 2688 20324
rect 2740 20312 2746 20324
rect 6564 20312 6592 20411
rect 7024 20389 7052 20488
rect 8386 20476 8392 20528
rect 8444 20476 8450 20528
rect 8938 20476 8944 20528
rect 8996 20476 9002 20528
rect 9950 20476 9956 20528
rect 10008 20516 10014 20528
rect 12069 20519 12127 20525
rect 12069 20516 12081 20519
rect 10008 20488 12081 20516
rect 10008 20476 10014 20488
rect 12069 20485 12081 20488
rect 12115 20485 12127 20519
rect 13814 20516 13820 20528
rect 12069 20479 12127 20485
rect 13648 20488 13820 20516
rect 8754 20408 8760 20460
rect 8812 20408 8818 20460
rect 9398 20408 9404 20460
rect 9456 20408 9462 20460
rect 10505 20451 10563 20457
rect 10505 20417 10517 20451
rect 10551 20448 10563 20451
rect 11514 20448 11520 20460
rect 10551 20420 11520 20448
rect 10551 20417 10563 20420
rect 10505 20411 10563 20417
rect 11514 20408 11520 20420
rect 11572 20408 11578 20460
rect 11882 20408 11888 20460
rect 11940 20408 11946 20460
rect 13648 20457 13676 20488
rect 13814 20476 13820 20488
rect 13872 20476 13878 20528
rect 15746 20476 15752 20528
rect 15804 20476 15810 20528
rect 16298 20476 16304 20528
rect 16356 20476 16362 20528
rect 12529 20451 12587 20457
rect 12529 20448 12541 20451
rect 12406 20420 12541 20448
rect 7009 20383 7067 20389
rect 7009 20349 7021 20383
rect 7055 20349 7067 20383
rect 7009 20343 7067 20349
rect 9950 20340 9956 20392
rect 10008 20380 10014 20392
rect 12406 20380 12434 20420
rect 12529 20417 12541 20420
rect 12575 20417 12587 20451
rect 12529 20411 12587 20417
rect 13633 20451 13691 20457
rect 13633 20417 13645 20451
rect 13679 20417 13691 20451
rect 13633 20411 13691 20417
rect 15010 20408 15016 20460
rect 15068 20448 15074 20460
rect 15838 20448 15844 20460
rect 15068 20420 15844 20448
rect 15068 20408 15074 20420
rect 15838 20408 15844 20420
rect 15896 20408 15902 20460
rect 16114 20408 16120 20460
rect 16172 20408 16178 20460
rect 16850 20408 16856 20460
rect 16908 20448 16914 20460
rect 17129 20451 17187 20457
rect 17129 20448 17141 20451
rect 16908 20420 17141 20448
rect 16908 20408 16914 20420
rect 17129 20417 17141 20420
rect 17175 20417 17187 20451
rect 17129 20411 17187 20417
rect 18506 20408 18512 20460
rect 18564 20408 18570 20460
rect 10008 20352 12434 20380
rect 13173 20383 13231 20389
rect 10008 20340 10014 20352
rect 13173 20349 13185 20383
rect 13219 20380 13231 20383
rect 13446 20380 13452 20392
rect 13219 20352 13452 20380
rect 13219 20349 13231 20352
rect 13173 20343 13231 20349
rect 13446 20340 13452 20352
rect 13504 20340 13510 20392
rect 13906 20340 13912 20392
rect 13964 20340 13970 20392
rect 17405 20383 17463 20389
rect 17405 20380 17417 20383
rect 14936 20352 17417 20380
rect 2740 20284 6592 20312
rect 2740 20272 2746 20284
rect 7742 20272 7748 20324
rect 7800 20312 7806 20324
rect 7800 20284 13768 20312
rect 7800 20272 7806 20284
rect 9766 20204 9772 20256
rect 9824 20244 9830 20256
rect 10045 20247 10103 20253
rect 10045 20244 10057 20247
rect 9824 20216 10057 20244
rect 9824 20204 9830 20216
rect 10045 20213 10057 20216
rect 10091 20213 10103 20247
rect 10045 20207 10103 20213
rect 10134 20204 10140 20256
rect 10192 20244 10198 20256
rect 13630 20244 13636 20256
rect 10192 20216 13636 20244
rect 10192 20204 10198 20216
rect 13630 20204 13636 20216
rect 13688 20204 13694 20256
rect 13740 20244 13768 20284
rect 14936 20244 14964 20352
rect 17405 20349 17417 20352
rect 17451 20349 17463 20383
rect 18708 20380 18736 20556
rect 19628 20556 20720 20584
rect 19628 20457 19656 20556
rect 20714 20544 20720 20556
rect 20772 20544 20778 20596
rect 20806 20544 20812 20596
rect 20864 20584 20870 20596
rect 22005 20587 22063 20593
rect 22005 20584 22017 20587
rect 20864 20556 22017 20584
rect 20864 20544 20870 20556
rect 22005 20553 22017 20556
rect 22051 20553 22063 20587
rect 22005 20547 22063 20553
rect 22094 20544 22100 20596
rect 22152 20584 22158 20596
rect 22922 20584 22928 20596
rect 22152 20556 22928 20584
rect 22152 20544 22158 20556
rect 22922 20544 22928 20556
rect 22980 20544 22986 20596
rect 24854 20584 24860 20596
rect 23216 20556 24860 20584
rect 22830 20516 22836 20528
rect 22066 20488 22836 20516
rect 19613 20451 19671 20457
rect 19613 20417 19625 20451
rect 19659 20417 19671 20451
rect 22066 20448 22094 20488
rect 22830 20476 22836 20488
rect 22888 20476 22894 20528
rect 21022 20434 22094 20448
rect 19613 20411 19671 20417
rect 21008 20420 22094 20434
rect 22373 20451 22431 20457
rect 19889 20383 19947 20389
rect 19889 20380 19901 20383
rect 18708 20352 19901 20380
rect 17405 20343 17463 20349
rect 19889 20349 19901 20352
rect 19935 20349 19947 20383
rect 19889 20343 19947 20349
rect 15378 20272 15384 20324
rect 15436 20272 15442 20324
rect 18506 20272 18512 20324
rect 18564 20312 18570 20324
rect 18564 20284 19288 20312
rect 18564 20272 18570 20284
rect 13740 20216 14964 20244
rect 16853 20247 16911 20253
rect 16853 20213 16865 20247
rect 16899 20244 16911 20247
rect 17586 20244 17592 20256
rect 16899 20216 17592 20244
rect 16899 20213 16911 20216
rect 16853 20207 16911 20213
rect 17586 20204 17592 20216
rect 17644 20204 17650 20256
rect 18874 20204 18880 20256
rect 18932 20204 18938 20256
rect 19260 20244 19288 20284
rect 19334 20272 19340 20324
rect 19392 20272 19398 20324
rect 21008 20244 21036 20420
rect 22373 20417 22385 20451
rect 22419 20448 22431 20451
rect 22646 20448 22652 20460
rect 22419 20420 22652 20448
rect 22419 20417 22431 20420
rect 22373 20411 22431 20417
rect 22646 20408 22652 20420
rect 22704 20408 22710 20460
rect 23216 20457 23244 20556
rect 24854 20544 24860 20556
rect 24912 20544 24918 20596
rect 25777 20587 25835 20593
rect 25777 20584 25789 20587
rect 24964 20556 25789 20584
rect 23477 20519 23535 20525
rect 23477 20485 23489 20519
rect 23523 20516 23535 20519
rect 23566 20516 23572 20528
rect 23523 20488 23572 20516
rect 23523 20485 23535 20488
rect 23477 20479 23535 20485
rect 23566 20476 23572 20488
rect 23624 20476 23630 20528
rect 24762 20516 24768 20528
rect 24702 20488 24768 20516
rect 24762 20476 24768 20488
rect 24820 20476 24826 20528
rect 23201 20451 23259 20457
rect 23201 20417 23213 20451
rect 23247 20417 23259 20451
rect 23201 20411 23259 20417
rect 22462 20340 22468 20392
rect 22520 20340 22526 20392
rect 22557 20383 22615 20389
rect 22557 20349 22569 20383
rect 22603 20380 22615 20383
rect 22922 20380 22928 20392
rect 22603 20352 22928 20380
rect 22603 20349 22615 20352
rect 22557 20343 22615 20349
rect 22922 20340 22928 20352
rect 22980 20340 22986 20392
rect 21082 20272 21088 20324
rect 21140 20312 21146 20324
rect 23216 20312 23244 20411
rect 24118 20340 24124 20392
rect 24176 20380 24182 20392
rect 24964 20380 24992 20556
rect 25777 20553 25789 20556
rect 25823 20553 25835 20587
rect 25777 20547 25835 20553
rect 26234 20544 26240 20596
rect 26292 20584 26298 20596
rect 27157 20587 27215 20593
rect 27157 20584 27169 20587
rect 26292 20556 27169 20584
rect 26292 20544 26298 20556
rect 27157 20553 27169 20556
rect 27203 20553 27215 20587
rect 27157 20547 27215 20553
rect 28350 20544 28356 20596
rect 28408 20584 28414 20596
rect 28718 20584 28724 20596
rect 28408 20556 28724 20584
rect 28408 20544 28414 20556
rect 28718 20544 28724 20556
rect 28776 20544 28782 20596
rect 28902 20544 28908 20596
rect 28960 20584 28966 20596
rect 29457 20587 29515 20593
rect 29457 20584 29469 20587
rect 28960 20556 29469 20584
rect 28960 20544 28966 20556
rect 29457 20553 29469 20556
rect 29503 20584 29515 20587
rect 30006 20584 30012 20596
rect 29503 20556 30012 20584
rect 29503 20553 29515 20556
rect 29457 20547 29515 20553
rect 30006 20544 30012 20556
rect 30064 20544 30070 20596
rect 30098 20544 30104 20596
rect 30156 20584 30162 20596
rect 30285 20587 30343 20593
rect 30285 20584 30297 20587
rect 30156 20556 30297 20584
rect 30156 20544 30162 20556
rect 30285 20553 30297 20556
rect 30331 20553 30343 20587
rect 30285 20547 30343 20553
rect 30834 20544 30840 20596
rect 30892 20584 30898 20596
rect 37090 20584 37096 20596
rect 30892 20556 37096 20584
rect 30892 20544 30898 20556
rect 37090 20544 37096 20556
rect 37148 20544 37154 20596
rect 37550 20544 37556 20596
rect 37608 20544 37614 20596
rect 41874 20584 41880 20596
rect 38304 20556 41880 20584
rect 29270 20516 29276 20528
rect 24176 20352 24992 20380
rect 25240 20488 29276 20516
rect 24176 20340 24182 20352
rect 21140 20284 23244 20312
rect 21140 20272 21146 20284
rect 24486 20272 24492 20324
rect 24544 20312 24550 20324
rect 25240 20321 25268 20488
rect 26145 20451 26203 20457
rect 26145 20417 26157 20451
rect 26191 20417 26203 20451
rect 26145 20411 26203 20417
rect 25225 20315 25283 20321
rect 25225 20312 25237 20315
rect 24544 20284 25237 20312
rect 24544 20272 24550 20284
rect 25225 20281 25237 20284
rect 25271 20281 25283 20315
rect 25225 20275 25283 20281
rect 25409 20315 25467 20321
rect 25409 20281 25421 20315
rect 25455 20312 25467 20315
rect 25682 20312 25688 20324
rect 25455 20284 25688 20312
rect 25455 20281 25467 20284
rect 25409 20275 25467 20281
rect 25682 20272 25688 20284
rect 25740 20272 25746 20324
rect 26160 20312 26188 20411
rect 26786 20408 26792 20460
rect 26844 20448 26850 20460
rect 26844 20420 27292 20448
rect 26844 20408 26850 20420
rect 26234 20340 26240 20392
rect 26292 20340 26298 20392
rect 26326 20340 26332 20392
rect 26384 20340 26390 20392
rect 27264 20380 27292 20420
rect 27338 20408 27344 20460
rect 27396 20448 27402 20460
rect 27525 20451 27583 20457
rect 27525 20448 27537 20451
rect 27396 20420 27537 20448
rect 27396 20408 27402 20420
rect 27525 20417 27537 20420
rect 27571 20417 27583 20451
rect 27632 20448 27660 20488
rect 29270 20476 29276 20488
rect 29328 20476 29334 20528
rect 32306 20476 32312 20528
rect 32364 20516 32370 20528
rect 32585 20519 32643 20525
rect 32585 20516 32597 20519
rect 32364 20488 32597 20516
rect 32364 20476 32370 20488
rect 32585 20485 32597 20488
rect 32631 20485 32643 20519
rect 32585 20479 32643 20485
rect 33226 20476 33232 20528
rect 33284 20476 33290 20528
rect 34238 20476 34244 20528
rect 34296 20516 34302 20528
rect 34333 20519 34391 20525
rect 34333 20516 34345 20519
rect 34296 20488 34345 20516
rect 34296 20476 34302 20488
rect 34333 20485 34345 20488
rect 34379 20485 34391 20519
rect 34333 20479 34391 20485
rect 34698 20476 34704 20528
rect 34756 20516 34762 20528
rect 36538 20516 36544 20528
rect 34756 20488 36544 20516
rect 34756 20476 34762 20488
rect 36538 20476 36544 20488
rect 36596 20476 36602 20528
rect 36722 20476 36728 20528
rect 36780 20516 36786 20528
rect 37568 20516 37596 20544
rect 38304 20525 38332 20556
rect 41874 20544 41880 20556
rect 41932 20544 41938 20596
rect 41966 20544 41972 20596
rect 42024 20584 42030 20596
rect 42061 20587 42119 20593
rect 42061 20584 42073 20587
rect 42024 20556 42073 20584
rect 42024 20544 42030 20556
rect 42061 20553 42073 20556
rect 42107 20553 42119 20587
rect 42061 20547 42119 20553
rect 43257 20587 43315 20593
rect 43257 20553 43269 20587
rect 43303 20584 43315 20587
rect 43714 20584 43720 20596
rect 43303 20556 43720 20584
rect 43303 20553 43315 20556
rect 43257 20547 43315 20553
rect 43714 20544 43720 20556
rect 43772 20544 43778 20596
rect 45462 20544 45468 20596
rect 45520 20544 45526 20596
rect 45646 20544 45652 20596
rect 45704 20584 45710 20596
rect 47029 20587 47087 20593
rect 47029 20584 47041 20587
rect 45704 20556 47041 20584
rect 45704 20544 45710 20556
rect 47029 20553 47041 20556
rect 47075 20553 47087 20587
rect 47029 20547 47087 20553
rect 36780 20488 37596 20516
rect 38289 20519 38347 20525
rect 36780 20476 36786 20488
rect 38289 20485 38301 20519
rect 38335 20485 38347 20519
rect 38289 20479 38347 20485
rect 38930 20476 38936 20528
rect 38988 20476 38994 20528
rect 40310 20476 40316 20528
rect 40368 20516 40374 20528
rect 42242 20516 42248 20528
rect 40368 20488 42248 20516
rect 40368 20476 40374 20488
rect 42242 20476 42248 20488
rect 42300 20476 42306 20528
rect 46569 20519 46627 20525
rect 46569 20516 46581 20519
rect 43732 20488 46581 20516
rect 28353 20451 28411 20457
rect 27632 20420 27752 20448
rect 27525 20411 27583 20417
rect 27724 20389 27752 20420
rect 28353 20417 28365 20451
rect 28399 20448 28411 20451
rect 28626 20448 28632 20460
rect 28399 20420 28632 20448
rect 28399 20417 28411 20420
rect 28353 20411 28411 20417
rect 28626 20408 28632 20420
rect 28684 20408 28690 20460
rect 29638 20408 29644 20460
rect 29696 20448 29702 20460
rect 29696 20420 30512 20448
rect 29696 20408 29702 20420
rect 27617 20383 27675 20389
rect 27617 20380 27629 20383
rect 27264 20352 27629 20380
rect 27617 20349 27629 20352
rect 27663 20349 27675 20383
rect 27617 20343 27675 20349
rect 27709 20383 27767 20389
rect 27709 20349 27721 20383
rect 27755 20349 27767 20383
rect 27709 20343 27767 20349
rect 27798 20340 27804 20392
rect 27856 20380 27862 20392
rect 30484 20389 30512 20420
rect 31110 20408 31116 20460
rect 31168 20408 31174 20460
rect 35066 20408 35072 20460
rect 35124 20448 35130 20460
rect 35253 20451 35311 20457
rect 35253 20448 35265 20451
rect 35124 20420 35265 20448
rect 35124 20408 35130 20420
rect 35253 20417 35265 20420
rect 35299 20417 35311 20451
rect 35253 20411 35311 20417
rect 35894 20408 35900 20460
rect 35952 20448 35958 20460
rect 36449 20451 36507 20457
rect 36449 20448 36461 20451
rect 35952 20420 36461 20448
rect 35952 20408 35958 20420
rect 36449 20417 36461 20420
rect 36495 20448 36507 20451
rect 36998 20448 37004 20460
rect 36495 20420 37004 20448
rect 36495 20417 36507 20420
rect 36449 20411 36507 20417
rect 36998 20408 37004 20420
rect 37056 20408 37062 20460
rect 37458 20408 37464 20460
rect 37516 20448 37522 20460
rect 37826 20448 37832 20460
rect 37516 20420 37832 20448
rect 37516 20408 37522 20420
rect 37826 20408 37832 20420
rect 37884 20448 37890 20460
rect 38013 20451 38071 20457
rect 38013 20448 38025 20451
rect 37884 20420 38025 20448
rect 37884 20408 37890 20420
rect 38013 20417 38025 20420
rect 38059 20417 38071 20451
rect 38013 20411 38071 20417
rect 39666 20408 39672 20460
rect 39724 20448 39730 20460
rect 40126 20448 40132 20460
rect 39724 20420 40132 20448
rect 39724 20408 39730 20420
rect 40126 20408 40132 20420
rect 40184 20408 40190 20460
rect 40589 20451 40647 20457
rect 40589 20417 40601 20451
rect 40635 20417 40647 20451
rect 40589 20411 40647 20417
rect 40681 20451 40739 20457
rect 40681 20417 40693 20451
rect 40727 20448 40739 20451
rect 40770 20448 40776 20460
rect 40727 20420 40776 20448
rect 40727 20417 40739 20420
rect 40681 20411 40739 20417
rect 30377 20383 30435 20389
rect 30377 20380 30389 20383
rect 27856 20352 30389 20380
rect 27856 20340 27862 20352
rect 30377 20349 30389 20352
rect 30423 20349 30435 20383
rect 30377 20343 30435 20349
rect 30469 20383 30527 20389
rect 30469 20349 30481 20383
rect 30515 20380 30527 20383
rect 30515 20352 31754 20380
rect 30515 20349 30527 20352
rect 30469 20343 30527 20349
rect 27062 20312 27068 20324
rect 26160 20284 27068 20312
rect 27062 20272 27068 20284
rect 27120 20312 27126 20324
rect 28350 20312 28356 20324
rect 27120 20284 28356 20312
rect 27120 20272 27126 20284
rect 28350 20272 28356 20284
rect 28408 20272 28414 20324
rect 30392 20312 30420 20343
rect 30558 20312 30564 20324
rect 30392 20284 30564 20312
rect 30558 20272 30564 20284
rect 30616 20272 30622 20324
rect 31726 20312 31754 20352
rect 32306 20340 32312 20392
rect 32364 20340 32370 20392
rect 34054 20340 34060 20392
rect 34112 20340 34118 20392
rect 35342 20340 35348 20392
rect 35400 20340 35406 20392
rect 35529 20383 35587 20389
rect 35529 20349 35541 20383
rect 35575 20380 35587 20383
rect 35802 20380 35808 20392
rect 35575 20352 35808 20380
rect 35575 20349 35587 20352
rect 35529 20343 35587 20349
rect 35802 20340 35808 20352
rect 35860 20340 35866 20392
rect 36633 20383 36691 20389
rect 36633 20349 36645 20383
rect 36679 20349 36691 20383
rect 40310 20380 40316 20392
rect 36633 20343 36691 20349
rect 38120 20352 40316 20380
rect 34517 20315 34575 20321
rect 34517 20312 34529 20315
rect 31726 20284 32444 20312
rect 19260 20216 21036 20244
rect 21266 20204 21272 20256
rect 21324 20244 21330 20256
rect 21361 20247 21419 20253
rect 21361 20244 21373 20247
rect 21324 20216 21373 20244
rect 21324 20204 21330 20216
rect 21361 20213 21373 20216
rect 21407 20213 21419 20247
rect 21361 20207 21419 20213
rect 22462 20204 22468 20256
rect 22520 20244 22526 20256
rect 23290 20244 23296 20256
rect 22520 20216 23296 20244
rect 22520 20204 22526 20216
rect 23290 20204 23296 20216
rect 23348 20204 23354 20256
rect 23474 20204 23480 20256
rect 23532 20244 23538 20256
rect 24949 20247 25007 20253
rect 24949 20244 24961 20247
rect 23532 20216 24961 20244
rect 23532 20204 23538 20216
rect 24949 20213 24961 20216
rect 24995 20213 25007 20247
rect 24949 20207 25007 20213
rect 25498 20204 25504 20256
rect 25556 20244 25562 20256
rect 28997 20247 29055 20253
rect 28997 20244 29009 20247
rect 25556 20216 29009 20244
rect 25556 20204 25562 20216
rect 28997 20213 29009 20216
rect 29043 20213 29055 20247
rect 28997 20207 29055 20213
rect 29270 20204 29276 20256
rect 29328 20204 29334 20256
rect 29914 20204 29920 20256
rect 29972 20204 29978 20256
rect 30098 20204 30104 20256
rect 30156 20244 30162 20256
rect 31757 20247 31815 20253
rect 31757 20244 31769 20247
rect 30156 20216 31769 20244
rect 30156 20204 30162 20216
rect 31757 20213 31769 20216
rect 31803 20213 31815 20247
rect 32416 20244 32444 20284
rect 33612 20284 34529 20312
rect 33612 20244 33640 20284
rect 34517 20281 34529 20284
rect 34563 20281 34575 20315
rect 36446 20312 36452 20324
rect 34517 20275 34575 20281
rect 34624 20284 36452 20312
rect 32416 20216 33640 20244
rect 31757 20207 31815 20213
rect 34054 20204 34060 20256
rect 34112 20244 34118 20256
rect 34624 20244 34652 20284
rect 36446 20272 36452 20284
rect 36504 20272 36510 20324
rect 34112 20216 34652 20244
rect 34112 20204 34118 20216
rect 34882 20204 34888 20256
rect 34940 20204 34946 20256
rect 35342 20204 35348 20256
rect 35400 20244 35406 20256
rect 36081 20247 36139 20253
rect 36081 20244 36093 20247
rect 35400 20216 36093 20244
rect 35400 20204 35406 20216
rect 36081 20213 36093 20216
rect 36127 20213 36139 20247
rect 36648 20244 36676 20343
rect 36814 20272 36820 20324
rect 36872 20312 36878 20324
rect 38120 20312 38148 20352
rect 40310 20340 40316 20352
rect 40368 20340 40374 20392
rect 40402 20340 40408 20392
rect 40460 20380 40466 20392
rect 40604 20380 40632 20411
rect 40770 20408 40776 20420
rect 40828 20448 40834 20460
rect 41138 20448 41144 20460
rect 40828 20420 41144 20448
rect 40828 20408 40834 20420
rect 41138 20408 41144 20420
rect 41196 20408 41202 20460
rect 41417 20451 41475 20457
rect 41417 20417 41429 20451
rect 41463 20448 41475 20451
rect 42058 20448 42064 20460
rect 41463 20420 42064 20448
rect 41463 20417 41475 20420
rect 41417 20411 41475 20417
rect 42058 20408 42064 20420
rect 42116 20408 42122 20460
rect 42613 20451 42671 20457
rect 42613 20417 42625 20451
rect 42659 20448 42671 20451
rect 42978 20448 42984 20460
rect 42659 20420 42984 20448
rect 42659 20417 42671 20420
rect 42613 20411 42671 20417
rect 42978 20408 42984 20420
rect 43036 20408 43042 20460
rect 43732 20457 43760 20488
rect 46569 20485 46581 20488
rect 46615 20485 46627 20519
rect 46569 20479 46627 20485
rect 47762 20476 47768 20528
rect 47820 20516 47826 20528
rect 49418 20516 49424 20528
rect 47820 20488 49424 20516
rect 47820 20476 47826 20488
rect 49418 20476 49424 20488
rect 49476 20476 49482 20528
rect 43717 20451 43775 20457
rect 43717 20417 43729 20451
rect 43763 20417 43775 20451
rect 43717 20411 43775 20417
rect 44821 20451 44879 20457
rect 44821 20417 44833 20451
rect 44867 20448 44879 20451
rect 45830 20448 45836 20460
rect 44867 20420 45836 20448
rect 44867 20417 44879 20420
rect 44821 20411 44879 20417
rect 45830 20408 45836 20420
rect 45888 20408 45894 20460
rect 45925 20451 45983 20457
rect 45925 20417 45937 20451
rect 45971 20417 45983 20451
rect 45925 20411 45983 20417
rect 40460 20352 40632 20380
rect 40865 20383 40923 20389
rect 40460 20340 40466 20352
rect 40865 20349 40877 20383
rect 40911 20349 40923 20383
rect 40865 20343 40923 20349
rect 36872 20284 38148 20312
rect 36872 20272 36878 20284
rect 39390 20272 39396 20324
rect 39448 20312 39454 20324
rect 39761 20315 39819 20321
rect 39761 20312 39773 20315
rect 39448 20284 39773 20312
rect 39448 20272 39454 20284
rect 39761 20281 39773 20284
rect 39807 20312 39819 20315
rect 40880 20312 40908 20343
rect 44358 20340 44364 20392
rect 44416 20340 44422 20392
rect 44910 20340 44916 20392
rect 44968 20380 44974 20392
rect 45278 20380 45284 20392
rect 44968 20352 45284 20380
rect 44968 20340 44974 20352
rect 45278 20340 45284 20352
rect 45336 20340 45342 20392
rect 45940 20312 45968 20411
rect 46106 20408 46112 20460
rect 46164 20448 46170 20460
rect 48041 20451 48099 20457
rect 48041 20448 48053 20451
rect 46164 20420 48053 20448
rect 46164 20408 46170 20420
rect 48041 20417 48053 20420
rect 48087 20417 48099 20451
rect 48041 20411 48099 20417
rect 49053 20451 49111 20457
rect 49053 20417 49065 20451
rect 49099 20448 49111 20451
rect 49602 20448 49608 20460
rect 49099 20420 49608 20448
rect 49099 20417 49111 20420
rect 49053 20411 49111 20417
rect 49602 20408 49608 20420
rect 49660 20408 49666 20460
rect 46014 20340 46020 20392
rect 46072 20380 46078 20392
rect 47765 20383 47823 20389
rect 47765 20380 47777 20383
rect 46072 20352 47777 20380
rect 46072 20340 46078 20352
rect 47765 20349 47777 20352
rect 47811 20380 47823 20383
rect 49142 20380 49148 20392
rect 47811 20352 49148 20380
rect 47811 20349 47823 20352
rect 47765 20343 47823 20349
rect 49142 20340 49148 20352
rect 49200 20340 49206 20392
rect 39807 20284 45968 20312
rect 39807 20281 39819 20284
rect 39761 20275 39819 20281
rect 46474 20272 46480 20324
rect 46532 20312 46538 20324
rect 46845 20315 46903 20321
rect 46845 20312 46857 20315
rect 46532 20284 46857 20312
rect 46532 20272 46538 20284
rect 46845 20281 46857 20284
rect 46891 20281 46903 20315
rect 46845 20275 46903 20281
rect 37090 20244 37096 20256
rect 36648 20216 37096 20244
rect 36081 20207 36139 20213
rect 37090 20204 37096 20216
rect 37148 20204 37154 20256
rect 37182 20204 37188 20256
rect 37240 20244 37246 20256
rect 37277 20247 37335 20253
rect 37277 20244 37289 20247
rect 37240 20216 37289 20244
rect 37240 20204 37246 20216
rect 37277 20213 37289 20216
rect 37323 20213 37335 20247
rect 37277 20207 37335 20213
rect 37642 20204 37648 20256
rect 37700 20204 37706 20256
rect 37734 20204 37740 20256
rect 37792 20244 37798 20256
rect 40034 20244 40040 20256
rect 37792 20216 40040 20244
rect 37792 20204 37798 20216
rect 40034 20204 40040 20216
rect 40092 20204 40098 20256
rect 40218 20204 40224 20256
rect 40276 20204 40282 20256
rect 40310 20204 40316 20256
rect 40368 20244 40374 20256
rect 40586 20244 40592 20256
rect 40368 20216 40592 20244
rect 40368 20204 40374 20216
rect 40586 20204 40592 20216
rect 40644 20244 40650 20256
rect 42794 20244 42800 20256
rect 40644 20216 42800 20244
rect 40644 20204 40650 20216
rect 42794 20204 42800 20216
rect 42852 20204 42858 20256
rect 44082 20204 44088 20256
rect 44140 20244 44146 20256
rect 44266 20244 44272 20256
rect 44140 20216 44272 20244
rect 44140 20204 44146 20216
rect 44266 20204 44272 20216
rect 44324 20204 44330 20256
rect 45186 20204 45192 20256
rect 45244 20244 45250 20256
rect 46106 20244 46112 20256
rect 45244 20216 46112 20244
rect 45244 20204 45250 20216
rect 46106 20204 46112 20216
rect 46164 20204 46170 20256
rect 47118 20204 47124 20256
rect 47176 20244 47182 20256
rect 47213 20247 47271 20253
rect 47213 20244 47225 20247
rect 47176 20216 47225 20244
rect 47176 20204 47182 20216
rect 47213 20213 47225 20216
rect 47259 20213 47271 20247
rect 47213 20207 47271 20213
rect 49237 20247 49295 20253
rect 49237 20213 49249 20247
rect 49283 20244 49295 20247
rect 49510 20244 49516 20256
rect 49283 20216 49516 20244
rect 49283 20213 49295 20216
rect 49237 20207 49295 20213
rect 49510 20204 49516 20216
rect 49568 20204 49574 20256
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 3421 20043 3479 20049
rect 3421 20009 3433 20043
rect 3467 20040 3479 20043
rect 3510 20040 3516 20052
rect 3467 20012 3516 20040
rect 3467 20009 3479 20012
rect 3421 20003 3479 20009
rect 3510 20000 3516 20012
rect 3568 20000 3574 20052
rect 3605 20043 3663 20049
rect 3605 20009 3617 20043
rect 3651 20040 3663 20043
rect 3651 20012 11100 20040
rect 3651 20009 3663 20012
rect 3605 20003 3663 20009
rect 10962 19972 10968 19984
rect 2746 19944 10968 19972
rect 2746 19904 2774 19944
rect 10962 19932 10968 19944
rect 11020 19932 11026 19984
rect 11072 19972 11100 20012
rect 11146 20000 11152 20052
rect 11204 20040 11210 20052
rect 14182 20040 14188 20052
rect 11204 20012 14188 20040
rect 11204 20000 11210 20012
rect 14182 20000 14188 20012
rect 14240 20000 14246 20052
rect 17862 20000 17868 20052
rect 17920 20040 17926 20052
rect 21082 20040 21088 20052
rect 17920 20012 21088 20040
rect 17920 20000 17926 20012
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 21174 20000 21180 20052
rect 21232 20040 21238 20052
rect 23201 20043 23259 20049
rect 23201 20040 23213 20043
rect 21232 20012 23213 20040
rect 21232 20000 21238 20012
rect 23201 20009 23213 20012
rect 23247 20009 23259 20043
rect 23201 20003 23259 20009
rect 23290 20000 23296 20052
rect 23348 20040 23354 20052
rect 24762 20040 24768 20052
rect 23348 20012 24768 20040
rect 23348 20000 23354 20012
rect 24762 20000 24768 20012
rect 24820 20000 24826 20052
rect 25590 20000 25596 20052
rect 25648 20040 25654 20052
rect 25648 20012 28488 20040
rect 25648 20000 25654 20012
rect 11422 19972 11428 19984
rect 11072 19944 11428 19972
rect 11422 19932 11428 19944
rect 11480 19932 11486 19984
rect 11514 19932 11520 19984
rect 11572 19932 11578 19984
rect 13630 19932 13636 19984
rect 13688 19972 13694 19984
rect 13688 19944 17172 19972
rect 13688 19932 13694 19944
rect 1780 19876 2774 19904
rect 1780 19845 1808 19876
rect 4890 19864 4896 19916
rect 4948 19864 4954 19916
rect 6178 19864 6184 19916
rect 6236 19904 6242 19916
rect 6273 19907 6331 19913
rect 6273 19904 6285 19907
rect 6236 19876 6285 19904
rect 6236 19864 6242 19876
rect 6273 19873 6285 19876
rect 6319 19873 6331 19907
rect 6273 19867 6331 19873
rect 7282 19864 7288 19916
rect 7340 19904 7346 19916
rect 7834 19904 7840 19916
rect 7340 19876 7840 19904
rect 7340 19864 7346 19876
rect 7834 19864 7840 19876
rect 7892 19864 7898 19916
rect 10134 19904 10140 19916
rect 7944 19876 10140 19904
rect 1765 19839 1823 19845
rect 1765 19805 1777 19839
rect 1811 19805 1823 19839
rect 1765 19799 1823 19805
rect 3326 19796 3332 19848
rect 3384 19836 3390 19848
rect 3973 19839 4031 19845
rect 3973 19836 3985 19839
rect 3384 19808 3985 19836
rect 3384 19796 3390 19808
rect 3973 19805 3985 19808
rect 4019 19805 4031 19839
rect 3973 19799 4031 19805
rect 5997 19839 6055 19845
rect 5997 19805 6009 19839
rect 6043 19805 6055 19839
rect 5997 19799 6055 19805
rect 2777 19771 2835 19777
rect 2777 19737 2789 19771
rect 2823 19768 2835 19771
rect 2866 19768 2872 19780
rect 2823 19740 2872 19768
rect 2823 19737 2835 19740
rect 2777 19731 2835 19737
rect 2866 19728 2872 19740
rect 2924 19728 2930 19780
rect 4890 19728 4896 19780
rect 4948 19768 4954 19780
rect 5718 19768 5724 19780
rect 4948 19740 5724 19768
rect 4948 19728 4954 19740
rect 5718 19728 5724 19740
rect 5776 19728 5782 19780
rect 6012 19768 6040 19799
rect 7190 19796 7196 19848
rect 7248 19836 7254 19848
rect 7944 19845 7972 19876
rect 10134 19864 10140 19876
rect 10192 19864 10198 19916
rect 10413 19907 10471 19913
rect 10413 19873 10425 19907
rect 10459 19904 10471 19907
rect 13722 19904 13728 19916
rect 10459 19876 13728 19904
rect 10459 19873 10471 19876
rect 10413 19867 10471 19873
rect 13722 19864 13728 19876
rect 13780 19864 13786 19916
rect 16298 19904 16304 19916
rect 14476 19876 16304 19904
rect 7929 19839 7987 19845
rect 7929 19836 7941 19839
rect 7248 19808 7941 19836
rect 7248 19796 7254 19808
rect 7929 19805 7941 19808
rect 7975 19805 7987 19839
rect 7929 19799 7987 19805
rect 9766 19796 9772 19848
rect 9824 19796 9830 19848
rect 10873 19839 10931 19845
rect 10873 19836 10885 19839
rect 10704 19808 10885 19836
rect 6270 19768 6276 19780
rect 6012 19740 6276 19768
rect 6270 19728 6276 19740
rect 6328 19728 6334 19780
rect 10704 19777 10732 19808
rect 10873 19805 10885 19808
rect 10919 19805 10931 19839
rect 10873 19799 10931 19805
rect 11974 19796 11980 19848
rect 12032 19796 12038 19848
rect 13538 19796 13544 19848
rect 13596 19836 13602 19848
rect 14476 19836 14504 19876
rect 16298 19864 16304 19876
rect 16356 19864 16362 19916
rect 16485 19907 16543 19913
rect 16485 19873 16497 19907
rect 16531 19904 16543 19907
rect 16850 19904 16856 19916
rect 16531 19876 16856 19904
rect 16531 19873 16543 19876
rect 16485 19867 16543 19873
rect 16850 19864 16856 19876
rect 16908 19904 16914 19916
rect 17037 19907 17095 19913
rect 17037 19904 17049 19907
rect 16908 19876 17049 19904
rect 16908 19864 16914 19876
rect 17037 19873 17049 19876
rect 17083 19873 17095 19907
rect 17144 19904 17172 19944
rect 19242 19932 19248 19984
rect 19300 19972 19306 19984
rect 19521 19975 19579 19981
rect 19521 19972 19533 19975
rect 19300 19944 19533 19972
rect 19300 19932 19306 19944
rect 19521 19941 19533 19944
rect 19567 19941 19579 19975
rect 19521 19935 19579 19941
rect 22465 19975 22523 19981
rect 22465 19941 22477 19975
rect 22511 19972 22523 19975
rect 22554 19972 22560 19984
rect 22511 19944 22560 19972
rect 22511 19941 22523 19944
rect 22465 19935 22523 19941
rect 22554 19932 22560 19944
rect 22612 19932 22618 19984
rect 22925 19975 22983 19981
rect 22925 19972 22937 19975
rect 22664 19944 22937 19972
rect 18785 19907 18843 19913
rect 18785 19904 18797 19907
rect 17144 19876 18797 19904
rect 17037 19867 17095 19873
rect 18785 19873 18797 19876
rect 18831 19904 18843 19907
rect 19978 19904 19984 19916
rect 18831 19876 19984 19904
rect 18831 19873 18843 19876
rect 18785 19867 18843 19873
rect 19978 19864 19984 19876
rect 20036 19864 20042 19916
rect 20162 19864 20168 19916
rect 20220 19864 20226 19916
rect 20714 19864 20720 19916
rect 20772 19864 20778 19916
rect 21634 19864 21640 19916
rect 21692 19904 21698 19916
rect 22664 19904 22692 19944
rect 22925 19941 22937 19944
rect 22971 19972 22983 19975
rect 24302 19972 24308 19984
rect 22971 19944 24308 19972
rect 22971 19941 22983 19944
rect 22925 19935 22983 19941
rect 24302 19932 24308 19944
rect 24360 19932 24366 19984
rect 26234 19932 26240 19984
rect 26292 19972 26298 19984
rect 26970 19972 26976 19984
rect 26292 19944 26976 19972
rect 26292 19932 26298 19944
rect 26970 19932 26976 19944
rect 27028 19932 27034 19984
rect 21692 19876 22692 19904
rect 21692 19864 21698 19876
rect 23750 19864 23756 19916
rect 23808 19864 23814 19916
rect 24854 19864 24860 19916
rect 24912 19904 24918 19916
rect 24949 19907 25007 19913
rect 24949 19904 24961 19907
rect 24912 19876 24961 19904
rect 24912 19864 24918 19876
rect 24949 19873 24961 19876
rect 24995 19873 25007 19907
rect 24949 19867 25007 19873
rect 25222 19864 25228 19916
rect 25280 19864 25286 19916
rect 27430 19864 27436 19916
rect 27488 19864 27494 19916
rect 28460 19904 28488 20012
rect 29730 20000 29736 20052
rect 29788 20000 29794 20052
rect 30852 20012 31064 20040
rect 28905 19975 28963 19981
rect 28905 19941 28917 19975
rect 28951 19972 28963 19975
rect 29270 19972 29276 19984
rect 28951 19944 29276 19972
rect 28951 19941 28963 19944
rect 28905 19935 28963 19941
rect 29270 19932 29276 19944
rect 29328 19932 29334 19984
rect 28460 19876 28672 19904
rect 13596 19808 14504 19836
rect 13596 19796 13602 19808
rect 14550 19796 14556 19848
rect 14608 19796 14614 19848
rect 15194 19796 15200 19848
rect 15252 19836 15258 19848
rect 15252 19808 16620 19836
rect 15252 19796 15258 19808
rect 10689 19771 10747 19777
rect 10689 19768 10701 19771
rect 7484 19740 10701 19768
rect 5442 19660 5448 19712
rect 5500 19700 5506 19712
rect 7484 19700 7512 19740
rect 10689 19737 10701 19740
rect 10735 19737 10747 19771
rect 10689 19731 10747 19737
rect 5500 19672 7512 19700
rect 5500 19660 5506 19672
rect 7650 19660 7656 19712
rect 7708 19660 7714 19712
rect 8570 19660 8576 19712
rect 8628 19660 8634 19712
rect 9122 19660 9128 19712
rect 9180 19660 9186 19712
rect 10704 19700 10732 19731
rect 12250 19728 12256 19780
rect 12308 19728 12314 19780
rect 14090 19768 14096 19780
rect 13478 19740 14096 19768
rect 14090 19728 14096 19740
rect 14148 19728 14154 19780
rect 14182 19728 14188 19780
rect 14240 19768 14246 19780
rect 14277 19771 14335 19777
rect 14277 19768 14289 19771
rect 14240 19740 14289 19768
rect 14240 19728 14246 19740
rect 14277 19737 14289 19740
rect 14323 19768 14335 19771
rect 15657 19771 15715 19777
rect 15657 19768 15669 19771
rect 14323 19740 15669 19768
rect 14323 19737 14335 19740
rect 14277 19731 14335 19737
rect 15657 19737 15669 19740
rect 15703 19768 15715 19771
rect 16482 19768 16488 19780
rect 15703 19740 16488 19768
rect 15703 19737 15715 19740
rect 15657 19731 15715 19737
rect 16482 19728 16488 19740
rect 16540 19728 16546 19780
rect 16592 19768 16620 19808
rect 18414 19796 18420 19848
rect 18472 19796 18478 19848
rect 19518 19796 19524 19848
rect 19576 19836 19582 19848
rect 19889 19839 19947 19845
rect 19889 19836 19901 19839
rect 19576 19808 19901 19836
rect 19576 19796 19582 19808
rect 19889 19805 19901 19808
rect 19935 19805 19947 19839
rect 19889 19799 19947 19805
rect 22554 19796 22560 19848
rect 22612 19836 22618 19848
rect 22738 19836 22744 19848
rect 22612 19808 22744 19836
rect 22612 19796 22618 19808
rect 22738 19796 22744 19808
rect 22796 19796 22802 19848
rect 23566 19796 23572 19848
rect 23624 19836 23630 19848
rect 23661 19839 23719 19845
rect 23661 19836 23673 19839
rect 23624 19808 23673 19836
rect 23624 19796 23630 19808
rect 23661 19805 23673 19808
rect 23707 19805 23719 19839
rect 23661 19799 23719 19805
rect 26326 19796 26332 19848
rect 26384 19796 26390 19848
rect 27154 19796 27160 19848
rect 27212 19796 27218 19848
rect 28534 19796 28540 19848
rect 28592 19796 28598 19848
rect 28644 19836 28672 19876
rect 30190 19864 30196 19916
rect 30248 19904 30254 19916
rect 30377 19907 30435 19913
rect 30377 19904 30389 19907
rect 30248 19876 30389 19904
rect 30248 19864 30254 19876
rect 30377 19873 30389 19876
rect 30423 19904 30435 19907
rect 30852 19904 30880 20012
rect 30929 19975 30987 19981
rect 30929 19941 30941 19975
rect 30975 19941 30987 19975
rect 31036 19972 31064 20012
rect 32766 20000 32772 20052
rect 32824 20040 32830 20052
rect 33778 20040 33784 20052
rect 32824 20012 33784 20040
rect 32824 20000 32830 20012
rect 33778 20000 33784 20012
rect 33836 20000 33842 20052
rect 33962 20000 33968 20052
rect 34020 20040 34026 20052
rect 37734 20040 37740 20052
rect 34020 20012 37740 20040
rect 34020 20000 34026 20012
rect 37734 20000 37740 20012
rect 37792 20000 37798 20052
rect 38562 20000 38568 20052
rect 38620 20040 38626 20052
rect 38620 20012 38976 20040
rect 38620 20000 38626 20012
rect 34146 19972 34152 19984
rect 31036 19944 34152 19972
rect 30929 19935 30987 19941
rect 30423 19876 30880 19904
rect 30423 19873 30435 19876
rect 30377 19867 30435 19873
rect 30944 19836 30972 19935
rect 34146 19932 34152 19944
rect 34204 19932 34210 19984
rect 35158 19932 35164 19984
rect 35216 19972 35222 19984
rect 35526 19972 35532 19984
rect 35216 19944 35532 19972
rect 35216 19932 35222 19944
rect 35526 19932 35532 19944
rect 35584 19932 35590 19984
rect 36081 19975 36139 19981
rect 36081 19941 36093 19975
rect 36127 19972 36139 19975
rect 38948 19972 38976 20012
rect 39850 20000 39856 20052
rect 39908 20040 39914 20052
rect 42058 20040 42064 20052
rect 39908 20012 42064 20040
rect 39908 20000 39914 20012
rect 42058 20000 42064 20012
rect 42116 20000 42122 20052
rect 42242 20000 42248 20052
rect 42300 20040 42306 20052
rect 42981 20043 43039 20049
rect 42981 20040 42993 20043
rect 42300 20012 42993 20040
rect 42300 20000 42306 20012
rect 42981 20009 42993 20012
rect 43027 20009 43039 20043
rect 42981 20003 43039 20009
rect 43438 20000 43444 20052
rect 43496 20040 43502 20052
rect 44085 20043 44143 20049
rect 44085 20040 44097 20043
rect 43496 20012 44097 20040
rect 43496 20000 43502 20012
rect 44085 20009 44097 20012
rect 44131 20009 44143 20043
rect 44085 20003 44143 20009
rect 44266 20000 44272 20052
rect 44324 20040 44330 20052
rect 44729 20043 44787 20049
rect 44729 20040 44741 20043
rect 44324 20012 44741 20040
rect 44324 20000 44330 20012
rect 44729 20009 44741 20012
rect 44775 20040 44787 20043
rect 44775 20012 45784 20040
rect 44775 20009 44787 20012
rect 44729 20003 44787 20009
rect 36127 19944 38884 19972
rect 38948 19944 39804 19972
rect 36127 19941 36139 19944
rect 36081 19935 36139 19941
rect 31294 19904 31300 19916
rect 31128 19876 31300 19904
rect 31128 19845 31156 19876
rect 31294 19864 31300 19876
rect 31352 19864 31358 19916
rect 32398 19864 32404 19916
rect 32456 19864 32462 19916
rect 33134 19864 33140 19916
rect 33192 19904 33198 19916
rect 33505 19907 33563 19913
rect 33505 19904 33517 19907
rect 33192 19876 33517 19904
rect 33192 19864 33198 19876
rect 33505 19873 33517 19876
rect 33551 19904 33563 19907
rect 34238 19904 34244 19916
rect 33551 19876 34244 19904
rect 33551 19873 33563 19876
rect 33505 19867 33563 19873
rect 34238 19864 34244 19876
rect 34296 19864 34302 19916
rect 36262 19864 36268 19916
rect 36320 19904 36326 19916
rect 36446 19904 36452 19916
rect 36320 19876 36452 19904
rect 36320 19864 36326 19876
rect 36446 19864 36452 19876
rect 36504 19904 36510 19916
rect 36541 19907 36599 19913
rect 36541 19904 36553 19907
rect 36504 19876 36553 19904
rect 36504 19864 36510 19876
rect 36541 19873 36553 19876
rect 36587 19873 36599 19907
rect 36541 19867 36599 19873
rect 36725 19907 36783 19913
rect 36725 19873 36737 19907
rect 36771 19904 36783 19907
rect 38470 19904 38476 19916
rect 36771 19876 38476 19904
rect 36771 19873 36783 19876
rect 36725 19867 36783 19873
rect 38470 19864 38476 19876
rect 38528 19864 38534 19916
rect 38856 19904 38884 19944
rect 39209 19907 39267 19913
rect 39209 19904 39221 19907
rect 38856 19876 39221 19904
rect 39209 19873 39221 19876
rect 39255 19873 39267 19907
rect 39209 19867 39267 19873
rect 39301 19907 39359 19913
rect 39301 19873 39313 19907
rect 39347 19904 39359 19907
rect 39666 19904 39672 19916
rect 39347 19876 39672 19904
rect 39347 19873 39359 19876
rect 39301 19867 39359 19873
rect 39666 19864 39672 19876
rect 39724 19864 39730 19916
rect 39776 19904 39804 19944
rect 40770 19932 40776 19984
rect 40828 19972 40834 19984
rect 45756 19972 45784 20012
rect 45830 20000 45836 20052
rect 45888 20000 45894 20052
rect 49050 20000 49056 20052
rect 49108 20040 49114 20052
rect 49145 20043 49203 20049
rect 49145 20040 49157 20043
rect 49108 20012 49157 20040
rect 49108 20000 49114 20012
rect 49145 20009 49157 20012
rect 49191 20009 49203 20043
rect 49145 20003 49203 20009
rect 48314 19972 48320 19984
rect 40828 19944 43668 19972
rect 45756 19944 48320 19972
rect 40828 19932 40834 19944
rect 40681 19907 40739 19913
rect 40681 19904 40693 19907
rect 39776 19876 40693 19904
rect 40681 19873 40693 19876
rect 40727 19904 40739 19907
rect 43640 19904 43668 19944
rect 48314 19932 48320 19944
rect 48372 19932 48378 19984
rect 46937 19907 46995 19913
rect 46937 19904 46949 19907
rect 40727 19876 43484 19904
rect 43640 19876 46949 19904
rect 40727 19873 40739 19876
rect 40681 19867 40739 19873
rect 28644 19808 30972 19836
rect 31113 19839 31171 19845
rect 31113 19805 31125 19839
rect 31159 19805 31171 19839
rect 34149 19839 34207 19845
rect 34149 19836 34161 19839
rect 31113 19799 31171 19805
rect 31726 19808 34161 19836
rect 17313 19771 17371 19777
rect 17313 19768 17325 19771
rect 16592 19740 17325 19768
rect 17313 19737 17325 19740
rect 17359 19737 17371 19771
rect 17313 19731 17371 19737
rect 19306 19740 20852 19768
rect 13538 19700 13544 19712
rect 10704 19672 13544 19700
rect 13538 19660 13544 19672
rect 13596 19660 13602 19712
rect 13630 19660 13636 19712
rect 13688 19700 13694 19712
rect 13725 19703 13783 19709
rect 13725 19700 13737 19703
rect 13688 19672 13737 19700
rect 13688 19660 13694 19672
rect 13725 19669 13737 19672
rect 13771 19669 13783 19703
rect 13725 19663 13783 19669
rect 13814 19660 13820 19712
rect 13872 19700 13878 19712
rect 15197 19703 15255 19709
rect 15197 19700 15209 19703
rect 13872 19672 15209 19700
rect 13872 19660 13878 19672
rect 15197 19669 15209 19672
rect 15243 19669 15255 19703
rect 15197 19663 15255 19669
rect 16298 19660 16304 19712
rect 16356 19700 16362 19712
rect 19306 19700 19334 19740
rect 20824 19712 20852 19740
rect 20990 19728 20996 19780
rect 21048 19728 21054 19780
rect 22830 19768 22836 19780
rect 22218 19740 22836 19768
rect 22830 19728 22836 19740
rect 22888 19728 22894 19780
rect 24578 19728 24584 19780
rect 24636 19768 24642 19780
rect 25130 19768 25136 19780
rect 24636 19740 25136 19768
rect 24636 19728 24642 19740
rect 25130 19728 25136 19740
rect 25188 19728 25194 19780
rect 27706 19768 27712 19780
rect 26528 19740 27712 19768
rect 16356 19672 19334 19700
rect 19981 19703 20039 19709
rect 16356 19660 16362 19672
rect 19981 19669 19993 19703
rect 20027 19700 20039 19703
rect 20438 19700 20444 19712
rect 20027 19672 20444 19700
rect 20027 19669 20039 19672
rect 19981 19663 20039 19669
rect 20438 19660 20444 19672
rect 20496 19660 20502 19712
rect 20806 19660 20812 19712
rect 20864 19660 20870 19712
rect 23569 19703 23627 19709
rect 23569 19669 23581 19703
rect 23615 19700 23627 19703
rect 24302 19700 24308 19712
rect 23615 19672 24308 19700
rect 23615 19669 23627 19672
rect 23569 19663 23627 19669
rect 24302 19660 24308 19672
rect 24360 19660 24366 19712
rect 24489 19703 24547 19709
rect 24489 19669 24501 19703
rect 24535 19700 24547 19703
rect 24854 19700 24860 19712
rect 24535 19672 24860 19700
rect 24535 19669 24547 19672
rect 24489 19663 24547 19669
rect 24854 19660 24860 19672
rect 24912 19700 24918 19712
rect 26528 19700 26556 19740
rect 27706 19728 27712 19740
rect 27764 19728 27770 19780
rect 29454 19768 29460 19780
rect 28966 19740 29460 19768
rect 24912 19672 26556 19700
rect 26697 19703 26755 19709
rect 24912 19660 24918 19672
rect 26697 19669 26709 19703
rect 26743 19700 26755 19703
rect 28966 19700 28994 19740
rect 29454 19728 29460 19740
rect 29512 19728 29518 19780
rect 30101 19771 30159 19777
rect 30101 19737 30113 19771
rect 30147 19768 30159 19771
rect 30147 19740 30880 19768
rect 30147 19737 30159 19740
rect 30101 19731 30159 19737
rect 26743 19672 28994 19700
rect 26743 19669 26755 19672
rect 26697 19663 26755 19669
rect 29270 19660 29276 19712
rect 29328 19660 29334 19712
rect 29822 19660 29828 19712
rect 29880 19700 29886 19712
rect 30193 19703 30251 19709
rect 30193 19700 30205 19703
rect 29880 19672 30205 19700
rect 29880 19660 29886 19672
rect 30193 19669 30205 19672
rect 30239 19669 30251 19703
rect 30852 19700 30880 19740
rect 31570 19728 31576 19780
rect 31628 19728 31634 19780
rect 31726 19700 31754 19808
rect 34149 19805 34161 19808
rect 34195 19805 34207 19839
rect 34977 19839 35035 19845
rect 34977 19836 34989 19839
rect 34149 19799 34207 19805
rect 34440 19808 34989 19836
rect 32030 19728 32036 19780
rect 32088 19768 32094 19780
rect 33134 19768 33140 19780
rect 32088 19740 33140 19768
rect 32088 19728 32094 19740
rect 33134 19728 33140 19740
rect 33192 19728 33198 19780
rect 33321 19771 33379 19777
rect 33321 19737 33333 19771
rect 33367 19768 33379 19771
rect 33594 19768 33600 19780
rect 33367 19740 33600 19768
rect 33367 19737 33379 19740
rect 33321 19731 33379 19737
rect 33594 19728 33600 19740
rect 33652 19728 33658 19780
rect 33778 19728 33784 19780
rect 33836 19768 33842 19780
rect 34440 19768 34468 19808
rect 34977 19805 34989 19808
rect 35023 19836 35035 19839
rect 36630 19836 36636 19848
rect 35023 19808 36636 19836
rect 35023 19805 35035 19808
rect 34977 19799 35035 19805
rect 36630 19796 36636 19808
rect 36688 19796 36694 19848
rect 38654 19836 38660 19848
rect 37384 19808 38660 19836
rect 37384 19780 37412 19808
rect 38654 19796 38660 19808
rect 38712 19796 38718 19848
rect 39117 19839 39175 19845
rect 39117 19805 39129 19839
rect 39163 19836 39175 19839
rect 40218 19836 40224 19848
rect 39163 19808 40224 19836
rect 39163 19805 39175 19808
rect 39117 19799 39175 19805
rect 40218 19796 40224 19808
rect 40276 19796 40282 19848
rect 40310 19796 40316 19848
rect 40368 19836 40374 19848
rect 40405 19839 40463 19845
rect 40405 19836 40417 19839
rect 40368 19808 40417 19836
rect 40368 19796 40374 19808
rect 40405 19805 40417 19808
rect 40451 19805 40463 19839
rect 40405 19799 40463 19805
rect 41233 19839 41291 19845
rect 41233 19805 41245 19839
rect 41279 19805 41291 19839
rect 41233 19799 41291 19805
rect 33836 19740 34468 19768
rect 33836 19728 33842 19740
rect 34514 19728 34520 19780
rect 34572 19768 34578 19780
rect 35345 19771 35403 19777
rect 35345 19768 35357 19771
rect 34572 19740 35357 19768
rect 34572 19728 34578 19740
rect 35345 19737 35357 19740
rect 35391 19737 35403 19771
rect 35345 19731 35403 19737
rect 36354 19728 36360 19780
rect 36412 19768 36418 19780
rect 36449 19771 36507 19777
rect 36449 19768 36461 19771
rect 36412 19740 36461 19768
rect 36412 19728 36418 19740
rect 36449 19737 36461 19740
rect 36495 19768 36507 19771
rect 36998 19768 37004 19780
rect 36495 19740 37004 19768
rect 36495 19737 36507 19740
rect 36449 19731 36507 19737
rect 36998 19728 37004 19740
rect 37056 19728 37062 19780
rect 37366 19728 37372 19780
rect 37424 19728 37430 19780
rect 38197 19771 38255 19777
rect 38197 19737 38209 19771
rect 38243 19768 38255 19771
rect 38286 19768 38292 19780
rect 38243 19740 38292 19768
rect 38243 19737 38255 19740
rect 38197 19731 38255 19737
rect 38286 19728 38292 19740
rect 38344 19728 38350 19780
rect 41248 19768 41276 19799
rect 41874 19796 41880 19848
rect 41932 19796 41938 19848
rect 42337 19839 42395 19845
rect 42337 19805 42349 19839
rect 42383 19836 42395 19839
rect 43254 19836 43260 19848
rect 42383 19808 43260 19836
rect 42383 19805 42395 19808
rect 42337 19799 42395 19805
rect 43254 19796 43260 19808
rect 43312 19796 43318 19848
rect 43456 19845 43484 19876
rect 46937 19873 46949 19876
rect 46983 19873 46995 19907
rect 46937 19867 46995 19873
rect 43441 19839 43499 19845
rect 43441 19805 43453 19839
rect 43487 19805 43499 19839
rect 43441 19799 43499 19805
rect 44174 19796 44180 19848
rect 44232 19836 44238 19848
rect 45189 19839 45247 19845
rect 45189 19836 45201 19839
rect 44232 19808 45201 19836
rect 44232 19796 44238 19808
rect 45189 19805 45201 19808
rect 45235 19805 45247 19839
rect 45189 19799 45247 19805
rect 46290 19796 46296 19848
rect 46348 19796 46354 19848
rect 47397 19839 47455 19845
rect 47397 19805 47409 19839
rect 47443 19836 47455 19839
rect 48406 19836 48412 19848
rect 47443 19808 48412 19836
rect 47443 19805 47455 19808
rect 47397 19799 47455 19805
rect 48406 19796 48412 19808
rect 48464 19796 48470 19848
rect 48498 19796 48504 19848
rect 48556 19796 48562 19848
rect 38672 19740 41276 19768
rect 30852 19672 31754 19700
rect 30193 19663 30251 19669
rect 32766 19660 32772 19712
rect 32824 19700 32830 19712
rect 32953 19703 33011 19709
rect 32953 19700 32965 19703
rect 32824 19672 32965 19700
rect 32824 19660 32830 19672
rect 32953 19669 32965 19672
rect 32999 19669 33011 19703
rect 32953 19663 33011 19669
rect 33226 19660 33232 19712
rect 33284 19700 33290 19712
rect 33413 19703 33471 19709
rect 33413 19700 33425 19703
rect 33284 19672 33425 19700
rect 33284 19660 33290 19672
rect 33413 19669 33425 19672
rect 33459 19669 33471 19703
rect 33413 19663 33471 19669
rect 33502 19660 33508 19712
rect 33560 19700 33566 19712
rect 34790 19700 34796 19712
rect 33560 19672 34796 19700
rect 33560 19660 33566 19672
rect 34790 19660 34796 19672
rect 34848 19660 34854 19712
rect 36630 19660 36636 19712
rect 36688 19700 36694 19712
rect 38672 19700 38700 19740
rect 41322 19728 41328 19780
rect 41380 19728 41386 19780
rect 42058 19728 42064 19780
rect 42116 19768 42122 19780
rect 44361 19771 44419 19777
rect 44361 19768 44373 19771
rect 42116 19740 44373 19768
rect 42116 19728 42122 19740
rect 44361 19737 44373 19740
rect 44407 19768 44419 19771
rect 44450 19768 44456 19780
rect 44407 19740 44456 19768
rect 44407 19737 44419 19740
rect 44361 19731 44419 19737
rect 44450 19728 44456 19740
rect 44508 19728 44514 19780
rect 44637 19771 44695 19777
rect 44637 19737 44649 19771
rect 44683 19768 44695 19771
rect 49694 19768 49700 19780
rect 44683 19740 49700 19768
rect 44683 19737 44695 19740
rect 44637 19731 44695 19737
rect 36688 19672 38700 19700
rect 36688 19660 36694 19672
rect 38746 19660 38752 19712
rect 38804 19660 38810 19712
rect 40037 19703 40095 19709
rect 40037 19669 40049 19703
rect 40083 19700 40095 19703
rect 40310 19700 40316 19712
rect 40083 19672 40316 19700
rect 40083 19669 40095 19672
rect 40037 19663 40095 19669
rect 40310 19660 40316 19672
rect 40368 19660 40374 19712
rect 40402 19660 40408 19712
rect 40460 19700 40466 19712
rect 40497 19703 40555 19709
rect 40497 19700 40509 19703
rect 40460 19672 40509 19700
rect 40460 19660 40466 19672
rect 40497 19669 40509 19672
rect 40543 19669 40555 19703
rect 40497 19663 40555 19669
rect 40586 19660 40592 19712
rect 40644 19700 40650 19712
rect 41340 19700 41368 19728
rect 45204 19712 45232 19740
rect 49694 19728 49700 19740
rect 49752 19728 49758 19780
rect 40644 19672 41368 19700
rect 40644 19660 40650 19672
rect 42794 19660 42800 19712
rect 42852 19700 42858 19712
rect 43346 19700 43352 19712
rect 42852 19672 43352 19700
rect 42852 19660 42858 19672
rect 43346 19660 43352 19672
rect 43404 19660 43410 19712
rect 45186 19660 45192 19712
rect 45244 19660 45250 19712
rect 47026 19660 47032 19712
rect 47084 19700 47090 19712
rect 48041 19703 48099 19709
rect 48041 19700 48053 19703
rect 47084 19672 48053 19700
rect 47084 19660 47090 19672
rect 48041 19669 48053 19672
rect 48087 19669 48099 19703
rect 48041 19663 48099 19669
rect 49513 19703 49571 19709
rect 49513 19669 49525 19703
rect 49559 19700 49571 19703
rect 50614 19700 50620 19712
rect 49559 19672 50620 19700
rect 49559 19669 49571 19672
rect 49513 19663 49571 19669
rect 50614 19660 50620 19672
rect 50672 19660 50678 19712
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 3620 19468 9904 19496
rect 1762 19320 1768 19372
rect 1820 19320 1826 19372
rect 3620 19369 3648 19468
rect 4522 19388 4528 19440
rect 4580 19388 4586 19440
rect 7006 19428 7012 19440
rect 5368 19400 7012 19428
rect 5368 19369 5396 19400
rect 7006 19388 7012 19400
rect 7064 19388 7070 19440
rect 8849 19431 8907 19437
rect 8849 19428 8861 19431
rect 7116 19400 8861 19428
rect 3605 19363 3663 19369
rect 3605 19329 3617 19363
rect 3651 19329 3663 19363
rect 3605 19323 3663 19329
rect 5353 19363 5411 19369
rect 5353 19329 5365 19363
rect 5399 19329 5411 19363
rect 5353 19323 5411 19329
rect 5997 19363 6055 19369
rect 5997 19329 6009 19363
rect 6043 19360 6055 19363
rect 6822 19360 6828 19372
rect 6043 19332 6828 19360
rect 6043 19329 6055 19332
rect 5997 19323 6055 19329
rect 6822 19320 6828 19332
rect 6880 19320 6886 19372
rect 7116 19369 7144 19400
rect 8849 19397 8861 19400
rect 8895 19397 8907 19431
rect 9876 19428 9904 19468
rect 9950 19456 9956 19508
rect 10008 19456 10014 19508
rect 10134 19456 10140 19508
rect 10192 19496 10198 19508
rect 10413 19499 10471 19505
rect 10413 19496 10425 19499
rect 10192 19468 10425 19496
rect 10192 19456 10198 19468
rect 10413 19465 10425 19468
rect 10459 19465 10471 19499
rect 10413 19459 10471 19465
rect 10873 19499 10931 19505
rect 10873 19465 10885 19499
rect 10919 19496 10931 19499
rect 11698 19496 11704 19508
rect 10919 19468 11704 19496
rect 10919 19465 10931 19468
rect 10873 19459 10931 19465
rect 11698 19456 11704 19468
rect 11756 19456 11762 19508
rect 12897 19499 12955 19505
rect 12897 19465 12909 19499
rect 12943 19496 12955 19499
rect 15470 19496 15476 19508
rect 12943 19468 15476 19496
rect 12943 19465 12955 19468
rect 12897 19459 12955 19465
rect 15470 19456 15476 19468
rect 15528 19456 15534 19508
rect 15562 19456 15568 19508
rect 15620 19456 15626 19508
rect 19242 19456 19248 19508
rect 19300 19496 19306 19508
rect 19300 19468 20208 19496
rect 19300 19456 19306 19468
rect 10226 19428 10232 19440
rect 9876 19400 10232 19428
rect 8849 19391 8907 19397
rect 10226 19388 10232 19400
rect 10284 19388 10290 19440
rect 11330 19428 11336 19440
rect 10888 19400 11336 19428
rect 7101 19363 7159 19369
rect 7101 19329 7113 19363
rect 7147 19329 7159 19363
rect 7101 19323 7159 19329
rect 7742 19320 7748 19372
rect 7800 19320 7806 19372
rect 8202 19320 8208 19372
rect 8260 19320 8266 19372
rect 8570 19320 8576 19372
rect 8628 19360 8634 19372
rect 9309 19363 9367 19369
rect 9309 19360 9321 19363
rect 8628 19332 9321 19360
rect 8628 19320 8634 19332
rect 9309 19329 9321 19332
rect 9355 19329 9367 19363
rect 9309 19323 9367 19329
rect 10321 19363 10379 19369
rect 10321 19329 10333 19363
rect 10367 19360 10379 19363
rect 10686 19360 10692 19372
rect 10367 19332 10692 19360
rect 10367 19329 10379 19332
rect 10321 19323 10379 19329
rect 10686 19320 10692 19332
rect 10744 19360 10750 19372
rect 10781 19363 10839 19369
rect 10781 19360 10793 19363
rect 10744 19332 10793 19360
rect 10744 19320 10750 19332
rect 10781 19329 10793 19332
rect 10827 19329 10839 19363
rect 10781 19323 10839 19329
rect 2038 19252 2044 19304
rect 2096 19252 2102 19304
rect 5718 19252 5724 19304
rect 5776 19292 5782 19304
rect 10888 19292 10916 19400
rect 11330 19388 11336 19400
rect 11388 19388 11394 19440
rect 11422 19388 11428 19440
rect 11480 19428 11486 19440
rect 11793 19431 11851 19437
rect 11793 19428 11805 19431
rect 11480 19400 11805 19428
rect 11480 19388 11486 19400
rect 11793 19397 11805 19400
rect 11839 19428 11851 19431
rect 13354 19428 13360 19440
rect 11839 19400 13360 19428
rect 11839 19397 11851 19400
rect 11793 19391 11851 19397
rect 13354 19388 13360 19400
rect 13412 19388 13418 19440
rect 13817 19431 13875 19437
rect 13817 19397 13829 19431
rect 13863 19428 13875 19431
rect 14826 19428 14832 19440
rect 13863 19400 14832 19428
rect 13863 19397 13875 19400
rect 13817 19391 13875 19397
rect 14826 19388 14832 19400
rect 14884 19388 14890 19440
rect 18506 19388 18512 19440
rect 18564 19428 18570 19440
rect 18564 19400 18722 19428
rect 18564 19388 18570 19400
rect 12158 19320 12164 19372
rect 12216 19360 12222 19372
rect 12805 19363 12863 19369
rect 12805 19360 12817 19363
rect 12216 19332 12817 19360
rect 12216 19320 12222 19332
rect 12805 19329 12817 19332
rect 12851 19329 12863 19363
rect 12805 19323 12863 19329
rect 13372 19332 14136 19360
rect 13372 19304 13400 19332
rect 14108 19304 14136 19332
rect 14458 19320 14464 19372
rect 14516 19320 14522 19372
rect 14918 19320 14924 19372
rect 14976 19360 14982 19372
rect 15105 19363 15163 19369
rect 15105 19360 15117 19363
rect 14976 19332 15117 19360
rect 14976 19320 14982 19332
rect 15105 19329 15117 19332
rect 15151 19329 15163 19363
rect 15105 19323 15163 19329
rect 15378 19320 15384 19372
rect 15436 19360 15442 19372
rect 15933 19363 15991 19369
rect 15933 19360 15945 19363
rect 15436 19332 15945 19360
rect 15436 19320 15442 19332
rect 15933 19329 15945 19332
rect 15979 19329 15991 19363
rect 15933 19323 15991 19329
rect 16022 19320 16028 19372
rect 16080 19320 16086 19372
rect 16574 19320 16580 19372
rect 16632 19360 16638 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 16632 19332 16865 19360
rect 16632 19320 16638 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 17862 19320 17868 19372
rect 17920 19360 17926 19372
rect 17957 19363 18015 19369
rect 17957 19360 17969 19363
rect 17920 19332 17969 19360
rect 17920 19320 17926 19332
rect 17957 19329 17969 19332
rect 18003 19329 18015 19363
rect 17957 19323 18015 19329
rect 19702 19320 19708 19372
rect 19760 19360 19766 19372
rect 19981 19363 20039 19369
rect 19981 19360 19993 19363
rect 19760 19332 19993 19360
rect 19760 19320 19766 19332
rect 19981 19329 19993 19332
rect 20027 19329 20039 19363
rect 20180 19360 20208 19468
rect 21266 19456 21272 19508
rect 21324 19496 21330 19508
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 21324 19468 22017 19496
rect 21324 19456 21330 19468
rect 22005 19465 22017 19468
rect 22051 19465 22063 19499
rect 22005 19459 22063 19465
rect 22373 19499 22431 19505
rect 22373 19465 22385 19499
rect 22419 19496 22431 19499
rect 24581 19499 24639 19505
rect 24581 19496 24593 19499
rect 22419 19468 24593 19496
rect 22419 19465 22431 19468
rect 22373 19459 22431 19465
rect 24581 19465 24593 19468
rect 24627 19465 24639 19499
rect 24581 19459 24639 19465
rect 25038 19456 25044 19508
rect 25096 19496 25102 19508
rect 25866 19496 25872 19508
rect 25096 19468 25872 19496
rect 25096 19456 25102 19468
rect 25866 19456 25872 19468
rect 25924 19496 25930 19508
rect 27893 19499 27951 19505
rect 27893 19496 27905 19499
rect 25924 19468 27905 19496
rect 25924 19456 25930 19468
rect 27893 19465 27905 19468
rect 27939 19496 27951 19499
rect 28074 19496 28080 19508
rect 27939 19468 28080 19496
rect 27939 19465 27951 19468
rect 27893 19459 27951 19465
rect 28074 19456 28080 19468
rect 28132 19496 28138 19508
rect 28718 19496 28724 19508
rect 28132 19468 28724 19496
rect 28132 19456 28138 19468
rect 28718 19456 28724 19468
rect 28776 19456 28782 19508
rect 28810 19456 28816 19508
rect 28868 19496 28874 19508
rect 28905 19499 28963 19505
rect 28905 19496 28917 19499
rect 28868 19468 28917 19496
rect 28868 19456 28874 19468
rect 28905 19465 28917 19468
rect 28951 19465 28963 19499
rect 28905 19459 28963 19465
rect 29086 19456 29092 19508
rect 29144 19496 29150 19508
rect 29273 19499 29331 19505
rect 29273 19496 29285 19499
rect 29144 19468 29285 19496
rect 29144 19456 29150 19468
rect 29273 19465 29285 19468
rect 29319 19496 29331 19499
rect 30466 19496 30472 19508
rect 29319 19468 30472 19496
rect 29319 19465 29331 19468
rect 29273 19459 29331 19465
rect 30466 19456 30472 19468
rect 30524 19496 30530 19508
rect 30561 19499 30619 19505
rect 30561 19496 30573 19499
rect 30524 19468 30573 19496
rect 30524 19456 30530 19468
rect 30561 19465 30573 19468
rect 30607 19465 30619 19499
rect 30561 19459 30619 19465
rect 30929 19499 30987 19505
rect 30929 19465 30941 19499
rect 30975 19496 30987 19499
rect 32490 19496 32496 19508
rect 30975 19468 32496 19496
rect 30975 19465 30987 19468
rect 30929 19459 30987 19465
rect 32490 19456 32496 19468
rect 32548 19456 32554 19508
rect 32585 19499 32643 19505
rect 32585 19465 32597 19499
rect 32631 19465 32643 19499
rect 32585 19459 32643 19465
rect 32953 19499 33011 19505
rect 32953 19465 32965 19499
rect 32999 19496 33011 19499
rect 33042 19496 33048 19508
rect 32999 19468 33048 19496
rect 32999 19465 33011 19468
rect 32953 19459 33011 19465
rect 20533 19431 20591 19437
rect 20533 19397 20545 19431
rect 20579 19428 20591 19431
rect 21358 19428 21364 19440
rect 20579 19400 21364 19428
rect 20579 19397 20591 19400
rect 20533 19391 20591 19397
rect 21358 19388 21364 19400
rect 21416 19388 21422 19440
rect 21726 19388 21732 19440
rect 21784 19428 21790 19440
rect 22278 19428 22284 19440
rect 21784 19400 22284 19428
rect 21784 19388 21790 19400
rect 22278 19388 22284 19400
rect 22336 19388 22342 19440
rect 22465 19431 22523 19437
rect 22465 19397 22477 19431
rect 22511 19428 22523 19431
rect 24118 19428 24124 19440
rect 22511 19400 24124 19428
rect 22511 19397 22523 19400
rect 22465 19391 22523 19397
rect 24118 19388 24124 19400
rect 24176 19388 24182 19440
rect 24302 19388 24308 19440
rect 24360 19428 24366 19440
rect 30101 19431 30159 19437
rect 30101 19428 30113 19431
rect 24360 19400 30113 19428
rect 24360 19388 24366 19400
rect 30101 19397 30113 19400
rect 30147 19397 30159 19431
rect 31478 19428 31484 19440
rect 30101 19391 30159 19397
rect 30208 19400 31484 19428
rect 20180 19332 21036 19360
rect 19981 19323 20039 19329
rect 5776 19264 10916 19292
rect 10965 19295 11023 19301
rect 5776 19252 5782 19264
rect 10965 19261 10977 19295
rect 11011 19261 11023 19295
rect 10965 19255 11023 19261
rect 2314 19184 2320 19236
rect 2372 19224 2378 19236
rect 4614 19224 4620 19236
rect 2372 19196 4620 19224
rect 2372 19184 2378 19196
rect 4614 19184 4620 19196
rect 4672 19184 4678 19236
rect 5074 19184 5080 19236
rect 5132 19224 5138 19236
rect 6457 19227 6515 19233
rect 6457 19224 6469 19227
rect 5132 19196 6469 19224
rect 5132 19184 5138 19196
rect 6457 19193 6469 19196
rect 6503 19224 6515 19227
rect 7742 19224 7748 19236
rect 6503 19196 7748 19224
rect 6503 19193 6515 19196
rect 6457 19187 6515 19193
rect 7742 19184 7748 19196
rect 7800 19184 7806 19236
rect 7834 19184 7840 19236
rect 7892 19224 7898 19236
rect 10502 19224 10508 19236
rect 7892 19196 10508 19224
rect 7892 19184 7898 19196
rect 10502 19184 10508 19196
rect 10560 19184 10566 19236
rect 10980 19224 11008 19255
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 11977 19295 12035 19301
rect 11977 19292 11989 19295
rect 11112 19264 11989 19292
rect 11112 19252 11118 19264
rect 11977 19261 11989 19264
rect 12023 19261 12035 19295
rect 11977 19255 12035 19261
rect 12710 19252 12716 19304
rect 12768 19292 12774 19304
rect 12989 19295 13047 19301
rect 12989 19292 13001 19295
rect 12768 19264 13001 19292
rect 12768 19252 12774 19264
rect 12989 19261 13001 19264
rect 13035 19261 13047 19295
rect 12989 19255 13047 19261
rect 13354 19252 13360 19304
rect 13412 19252 13418 19304
rect 13998 19252 14004 19304
rect 14056 19252 14062 19304
rect 14090 19252 14096 19304
rect 14148 19292 14154 19304
rect 14826 19292 14832 19304
rect 14148 19264 14832 19292
rect 14148 19252 14154 19264
rect 14826 19252 14832 19264
rect 14884 19292 14890 19304
rect 15010 19292 15016 19304
rect 14884 19264 15016 19292
rect 14884 19252 14890 19264
rect 15010 19252 15016 19264
rect 15068 19252 15074 19304
rect 15194 19252 15200 19304
rect 15252 19292 15258 19304
rect 16114 19292 16120 19304
rect 15252 19264 16120 19292
rect 15252 19252 15258 19264
rect 16114 19252 16120 19264
rect 16172 19252 16178 19304
rect 18233 19295 18291 19301
rect 18233 19292 18245 19295
rect 16224 19264 18245 19292
rect 10869 19196 11008 19224
rect 6546 19116 6552 19168
rect 6604 19116 6610 19168
rect 6825 19159 6883 19165
rect 6825 19125 6837 19159
rect 6871 19156 6883 19159
rect 7098 19156 7104 19168
rect 6871 19128 7104 19156
rect 6871 19125 6883 19128
rect 6825 19119 6883 19125
rect 7098 19116 7104 19128
rect 7156 19156 7162 19168
rect 7650 19156 7656 19168
rect 7156 19128 7656 19156
rect 7156 19116 7162 19128
rect 7650 19116 7656 19128
rect 7708 19156 7714 19168
rect 7926 19156 7932 19168
rect 7708 19128 7932 19156
rect 7708 19116 7714 19128
rect 7926 19116 7932 19128
rect 7984 19116 7990 19168
rect 8018 19116 8024 19168
rect 8076 19156 8082 19168
rect 9214 19156 9220 19168
rect 8076 19128 9220 19156
rect 8076 19116 8082 19128
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 9582 19116 9588 19168
rect 9640 19156 9646 19168
rect 10869 19156 10897 19196
rect 12066 19184 12072 19236
rect 12124 19224 12130 19236
rect 12124 19196 13676 19224
rect 12124 19184 12130 19196
rect 9640 19128 10897 19156
rect 9640 19116 9646 19128
rect 11054 19116 11060 19168
rect 11112 19156 11118 19168
rect 11241 19159 11299 19165
rect 11241 19156 11253 19159
rect 11112 19128 11253 19156
rect 11112 19116 11118 19128
rect 11241 19125 11253 19128
rect 11287 19125 11299 19159
rect 11241 19119 11299 19125
rect 11330 19116 11336 19168
rect 11388 19156 11394 19168
rect 12158 19156 12164 19168
rect 11388 19128 12164 19156
rect 11388 19116 11394 19128
rect 12158 19116 12164 19128
rect 12216 19156 12222 19168
rect 12253 19159 12311 19165
rect 12253 19156 12265 19159
rect 12216 19128 12265 19156
rect 12216 19116 12222 19128
rect 12253 19125 12265 19128
rect 12299 19125 12311 19159
rect 12253 19119 12311 19125
rect 12434 19116 12440 19168
rect 12492 19116 12498 19168
rect 13648 19156 13676 19196
rect 13722 19184 13728 19236
rect 13780 19224 13786 19236
rect 16224 19224 16252 19264
rect 18233 19261 18245 19264
rect 18279 19261 18291 19295
rect 21008 19292 21036 19332
rect 21082 19320 21088 19372
rect 21140 19360 21146 19372
rect 21269 19363 21327 19369
rect 21269 19360 21281 19363
rect 21140 19332 21281 19360
rect 21140 19320 21146 19332
rect 21269 19329 21281 19332
rect 21315 19329 21327 19363
rect 21450 19360 21456 19372
rect 21269 19323 21327 19329
rect 21376 19332 21456 19360
rect 21376 19292 21404 19332
rect 21450 19320 21456 19332
rect 21508 19320 21514 19372
rect 22002 19320 22008 19372
rect 22060 19360 22066 19372
rect 22060 19332 22416 19360
rect 22060 19320 22066 19332
rect 21008 19264 21404 19292
rect 18233 19255 18291 19261
rect 21910 19252 21916 19304
rect 21968 19292 21974 19304
rect 22388 19292 22416 19332
rect 23474 19320 23480 19372
rect 23532 19334 23538 19372
rect 23753 19363 23811 19369
rect 23532 19320 23612 19334
rect 23753 19329 23765 19363
rect 23799 19360 23811 19363
rect 24854 19360 24860 19372
rect 23799 19332 24860 19360
rect 23799 19329 23811 19332
rect 23753 19323 23811 19329
rect 24854 19320 24860 19332
rect 24912 19320 24918 19372
rect 24949 19363 25007 19369
rect 24949 19329 24961 19363
rect 24995 19329 25007 19363
rect 24949 19323 25007 19329
rect 25041 19363 25099 19369
rect 25041 19329 25053 19363
rect 25087 19360 25099 19363
rect 25590 19360 25596 19372
rect 25087 19332 25596 19360
rect 25087 19329 25099 19332
rect 25041 19323 25099 19329
rect 23492 19306 23612 19320
rect 22462 19292 22468 19304
rect 21968 19264 22324 19292
rect 22388 19264 22468 19292
rect 21968 19252 21974 19264
rect 17954 19224 17960 19236
rect 13780 19196 16252 19224
rect 17420 19196 17960 19224
rect 13780 19184 13786 19196
rect 17420 19156 17448 19196
rect 17954 19184 17960 19196
rect 18012 19184 18018 19236
rect 19426 19184 19432 19236
rect 19484 19224 19490 19236
rect 21726 19224 21732 19236
rect 19484 19196 21732 19224
rect 19484 19184 19490 19196
rect 21726 19184 21732 19196
rect 21784 19184 21790 19236
rect 22296 19224 22324 19264
rect 22462 19252 22468 19264
rect 22520 19252 22526 19304
rect 22557 19295 22615 19301
rect 22557 19261 22569 19295
rect 22603 19261 22615 19295
rect 22557 19255 22615 19261
rect 22572 19224 22600 19255
rect 22296 19196 22600 19224
rect 23385 19227 23443 19233
rect 23385 19193 23397 19227
rect 23431 19224 23443 19227
rect 23584 19224 23612 19306
rect 23842 19292 23848 19304
rect 23431 19196 23612 19224
rect 23676 19264 23848 19292
rect 23431 19193 23443 19196
rect 23385 19187 23443 19193
rect 13648 19128 17448 19156
rect 17497 19159 17555 19165
rect 17497 19125 17509 19159
rect 17543 19156 17555 19159
rect 17862 19156 17868 19168
rect 17543 19128 17868 19156
rect 17543 19125 17555 19128
rect 17497 19119 17555 19125
rect 17862 19116 17868 19128
rect 17920 19116 17926 19168
rect 20806 19116 20812 19168
rect 20864 19156 20870 19168
rect 21450 19156 21456 19168
rect 20864 19128 21456 19156
rect 20864 19116 20870 19128
rect 21450 19116 21456 19128
rect 21508 19156 21514 19168
rect 22002 19156 22008 19168
rect 21508 19128 22008 19156
rect 21508 19116 21514 19128
rect 22002 19116 22008 19128
rect 22060 19116 22066 19168
rect 22278 19116 22284 19168
rect 22336 19156 22342 19168
rect 23109 19159 23167 19165
rect 23109 19156 23121 19159
rect 22336 19128 23121 19156
rect 22336 19116 22342 19128
rect 23109 19125 23121 19128
rect 23155 19125 23167 19159
rect 23109 19119 23167 19125
rect 23474 19116 23480 19168
rect 23532 19156 23538 19168
rect 23676 19156 23704 19264
rect 23842 19252 23848 19264
rect 23900 19252 23906 19304
rect 23934 19252 23940 19304
rect 23992 19292 23998 19304
rect 24029 19295 24087 19301
rect 24029 19292 24041 19295
rect 23992 19264 24041 19292
rect 23992 19252 23998 19264
rect 24029 19261 24041 19264
rect 24075 19292 24087 19295
rect 24578 19292 24584 19304
rect 24075 19264 24584 19292
rect 24075 19261 24087 19264
rect 24029 19255 24087 19261
rect 24578 19252 24584 19264
rect 24636 19252 24642 19304
rect 24964 19292 24992 19323
rect 25590 19320 25596 19332
rect 25648 19320 25654 19372
rect 25961 19363 26019 19369
rect 25961 19329 25973 19363
rect 26007 19360 26019 19363
rect 26007 19332 26188 19360
rect 26007 19329 26019 19332
rect 25961 19323 26019 19329
rect 24780 19264 24992 19292
rect 24780 19224 24808 19264
rect 25130 19252 25136 19304
rect 25188 19292 25194 19304
rect 26160 19292 26188 19332
rect 26234 19320 26240 19372
rect 26292 19360 26298 19372
rect 26605 19363 26663 19369
rect 26605 19360 26617 19363
rect 26292 19332 26617 19360
rect 26292 19320 26298 19332
rect 26605 19329 26617 19332
rect 26651 19329 26663 19363
rect 26605 19323 26663 19329
rect 27065 19363 27123 19369
rect 27065 19329 27077 19363
rect 27111 19360 27123 19363
rect 27111 19332 28120 19360
rect 27111 19329 27123 19332
rect 27065 19323 27123 19329
rect 27246 19292 27252 19304
rect 25188 19264 26004 19292
rect 26160 19264 27252 19292
rect 25188 19252 25194 19264
rect 25976 19236 26004 19264
rect 27246 19252 27252 19264
rect 27304 19252 27310 19304
rect 27982 19292 27988 19304
rect 27356 19264 27988 19292
rect 25222 19224 25228 19236
rect 24780 19196 25228 19224
rect 25222 19184 25228 19196
rect 25280 19224 25286 19236
rect 25593 19227 25651 19233
rect 25593 19224 25605 19227
rect 25280 19196 25605 19224
rect 25280 19184 25286 19196
rect 25593 19193 25605 19196
rect 25639 19193 25651 19227
rect 25593 19187 25651 19193
rect 25958 19184 25964 19236
rect 26016 19184 26022 19236
rect 26878 19184 26884 19236
rect 26936 19224 26942 19236
rect 27157 19227 27215 19233
rect 27157 19224 27169 19227
rect 26936 19196 27169 19224
rect 26936 19184 26942 19196
rect 27157 19193 27169 19196
rect 27203 19224 27215 19227
rect 27356 19224 27384 19264
rect 27982 19252 27988 19264
rect 28040 19252 28046 19304
rect 28092 19292 28120 19332
rect 29270 19320 29276 19372
rect 29328 19360 29334 19372
rect 29365 19363 29423 19369
rect 29365 19360 29377 19363
rect 29328 19332 29377 19360
rect 29328 19320 29334 19332
rect 29365 19329 29377 19332
rect 29411 19329 29423 19363
rect 29365 19323 29423 19329
rect 29454 19320 29460 19372
rect 29512 19360 29518 19372
rect 30208 19360 30236 19400
rect 31478 19388 31484 19400
rect 31536 19388 31542 19440
rect 32600 19428 32628 19459
rect 33042 19456 33048 19468
rect 33100 19456 33106 19508
rect 33318 19456 33324 19508
rect 33376 19496 33382 19508
rect 34241 19499 34299 19505
rect 34241 19496 34253 19499
rect 33376 19468 34253 19496
rect 33376 19456 33382 19468
rect 34241 19465 34253 19468
rect 34287 19465 34299 19499
rect 40494 19496 40500 19508
rect 34241 19459 34299 19465
rect 38856 19468 40500 19496
rect 34054 19428 34060 19440
rect 32600 19400 34060 19428
rect 34054 19388 34060 19400
rect 34112 19388 34118 19440
rect 34422 19388 34428 19440
rect 34480 19428 34486 19440
rect 38856 19437 38884 19468
rect 40494 19456 40500 19468
rect 40552 19456 40558 19508
rect 40773 19499 40831 19505
rect 40773 19465 40785 19499
rect 40819 19496 40831 19499
rect 40954 19496 40960 19508
rect 40819 19468 40960 19496
rect 40819 19465 40831 19468
rect 40773 19459 40831 19465
rect 40954 19456 40960 19468
rect 41012 19456 41018 19508
rect 41874 19456 41880 19508
rect 41932 19496 41938 19508
rect 42610 19496 42616 19508
rect 41932 19468 42616 19496
rect 41932 19456 41938 19468
rect 42610 19456 42616 19468
rect 42668 19456 42674 19508
rect 43254 19456 43260 19508
rect 43312 19456 43318 19508
rect 43438 19456 43444 19508
rect 43496 19496 43502 19508
rect 46569 19499 46627 19505
rect 46569 19496 46581 19499
rect 43496 19468 46581 19496
rect 43496 19456 43502 19468
rect 46569 19465 46581 19468
rect 46615 19465 46627 19499
rect 46569 19459 46627 19465
rect 35989 19431 36047 19437
rect 35989 19428 36001 19431
rect 34480 19400 36001 19428
rect 34480 19388 34486 19400
rect 35989 19397 36001 19400
rect 36035 19428 36047 19431
rect 38841 19431 38899 19437
rect 36035 19400 37228 19428
rect 36035 19397 36047 19400
rect 35989 19391 36047 19397
rect 29512 19332 29592 19360
rect 29512 19320 29518 19332
rect 28169 19295 28227 19301
rect 28169 19292 28181 19295
rect 28092 19264 28181 19292
rect 28169 19261 28181 19264
rect 28215 19292 28227 19295
rect 28534 19292 28540 19304
rect 28215 19264 28540 19292
rect 28215 19261 28227 19264
rect 28169 19255 28227 19261
rect 28534 19252 28540 19264
rect 28592 19292 28598 19304
rect 29564 19301 29592 19332
rect 29840 19332 30236 19360
rect 29549 19295 29607 19301
rect 28592 19264 29408 19292
rect 28592 19252 28598 19264
rect 27203 19196 27384 19224
rect 27203 19193 27215 19196
rect 27157 19187 27215 19193
rect 27430 19184 27436 19236
rect 27488 19224 27494 19236
rect 28629 19227 28687 19233
rect 28629 19224 28641 19227
rect 27488 19196 28641 19224
rect 27488 19184 27494 19196
rect 28629 19193 28641 19196
rect 28675 19224 28687 19227
rect 29270 19224 29276 19236
rect 28675 19196 29276 19224
rect 28675 19193 28687 19196
rect 28629 19187 28687 19193
rect 29270 19184 29276 19196
rect 29328 19184 29334 19236
rect 29380 19224 29408 19264
rect 29549 19261 29561 19295
rect 29595 19292 29607 19295
rect 29595 19264 29629 19292
rect 29595 19261 29607 19264
rect 29549 19255 29607 19261
rect 29840 19224 29868 19332
rect 31294 19320 31300 19372
rect 31352 19320 31358 19372
rect 31386 19320 31392 19372
rect 31444 19320 31450 19372
rect 34146 19320 34152 19372
rect 34204 19320 34210 19372
rect 34238 19320 34244 19372
rect 34296 19360 34302 19372
rect 34296 19332 34468 19360
rect 34296 19320 34302 19332
rect 31573 19295 31631 19301
rect 31573 19261 31585 19295
rect 31619 19292 31631 19295
rect 32122 19292 32128 19304
rect 31619 19264 32128 19292
rect 31619 19261 31631 19264
rect 31573 19255 31631 19261
rect 32122 19252 32128 19264
rect 32180 19252 32186 19304
rect 32950 19252 32956 19304
rect 33008 19292 33014 19304
rect 33045 19295 33103 19301
rect 33045 19292 33057 19295
rect 33008 19264 33057 19292
rect 33008 19252 33014 19264
rect 33045 19261 33057 19264
rect 33091 19261 33103 19295
rect 33045 19255 33103 19261
rect 33229 19295 33287 19301
rect 33229 19261 33241 19295
rect 33275 19292 33287 19295
rect 33275 19264 34008 19292
rect 33275 19261 33287 19264
rect 33229 19255 33287 19261
rect 29380 19196 29868 19224
rect 30006 19184 30012 19236
rect 30064 19224 30070 19236
rect 30064 19196 30696 19224
rect 30064 19184 30070 19196
rect 23532 19128 23704 19156
rect 23532 19116 23538 19128
rect 26510 19116 26516 19168
rect 26568 19156 26574 19168
rect 27525 19159 27583 19165
rect 27525 19156 27537 19159
rect 26568 19128 27537 19156
rect 26568 19116 26574 19128
rect 27525 19125 27537 19128
rect 27571 19125 27583 19159
rect 27525 19119 27583 19125
rect 28166 19116 28172 19168
rect 28224 19156 28230 19168
rect 28994 19156 29000 19168
rect 28224 19128 29000 19156
rect 28224 19116 28230 19128
rect 28994 19116 29000 19128
rect 29052 19156 29058 19168
rect 30558 19156 30564 19168
rect 29052 19128 30564 19156
rect 29052 19116 29058 19128
rect 30558 19116 30564 19128
rect 30616 19116 30622 19168
rect 30668 19156 30696 19196
rect 33778 19184 33784 19236
rect 33836 19184 33842 19236
rect 33980 19224 34008 19264
rect 34330 19252 34336 19304
rect 34388 19252 34394 19304
rect 34440 19292 34468 19332
rect 34790 19320 34796 19372
rect 34848 19320 34854 19372
rect 35253 19363 35311 19369
rect 35253 19329 35265 19363
rect 35299 19360 35311 19363
rect 36078 19360 36084 19372
rect 35299 19332 36084 19360
rect 35299 19329 35311 19332
rect 35253 19323 35311 19329
rect 36078 19320 36084 19332
rect 36136 19320 36142 19372
rect 36170 19320 36176 19372
rect 36228 19360 36234 19372
rect 36725 19363 36783 19369
rect 36725 19360 36737 19363
rect 36228 19332 36737 19360
rect 36228 19320 36234 19332
rect 36725 19329 36737 19332
rect 36771 19329 36783 19363
rect 37200 19360 37228 19400
rect 38841 19397 38853 19431
rect 38887 19397 38899 19431
rect 38841 19391 38899 19397
rect 39114 19388 39120 19440
rect 39172 19428 39178 19440
rect 39172 19400 39330 19428
rect 39172 19388 39178 19400
rect 41138 19388 41144 19440
rect 41196 19388 41202 19440
rect 41322 19388 41328 19440
rect 41380 19428 41386 19440
rect 41380 19400 43852 19428
rect 41380 19388 41386 19400
rect 37353 19360 37359 19372
rect 37200 19332 37359 19360
rect 36725 19323 36783 19329
rect 37353 19320 37359 19332
rect 37411 19320 37417 19372
rect 37458 19369 37464 19372
rect 37449 19363 37464 19369
rect 37449 19329 37461 19363
rect 37449 19323 37464 19329
rect 37458 19320 37464 19323
rect 37516 19320 37522 19372
rect 37826 19320 37832 19372
rect 37884 19360 37890 19372
rect 38565 19363 38623 19369
rect 38565 19360 38577 19363
rect 37884 19332 38577 19360
rect 37884 19320 37890 19332
rect 38565 19329 38577 19332
rect 38611 19329 38623 19363
rect 38565 19323 38623 19329
rect 40218 19320 40224 19372
rect 40276 19360 40282 19372
rect 40402 19360 40408 19372
rect 40276 19332 40408 19360
rect 40276 19320 40282 19332
rect 40402 19320 40408 19332
rect 40460 19320 40466 19372
rect 41233 19363 41291 19369
rect 40604 19332 41000 19360
rect 40126 19292 40132 19304
rect 34440 19264 36584 19292
rect 35158 19224 35164 19236
rect 33980 19196 35164 19224
rect 35158 19184 35164 19196
rect 35216 19184 35222 19236
rect 35437 19227 35495 19233
rect 35437 19193 35449 19227
rect 35483 19224 35495 19227
rect 35618 19224 35624 19236
rect 35483 19196 35624 19224
rect 35483 19193 35495 19196
rect 35437 19187 35495 19193
rect 35618 19184 35624 19196
rect 35676 19184 35682 19236
rect 36446 19224 36452 19236
rect 35728 19196 36452 19224
rect 30834 19156 30840 19168
rect 30668 19128 30840 19156
rect 30834 19116 30840 19128
rect 30892 19156 30898 19168
rect 32214 19156 32220 19168
rect 30892 19128 32220 19156
rect 30892 19116 30898 19128
rect 32214 19116 32220 19128
rect 32272 19116 32278 19168
rect 34054 19116 34060 19168
rect 34112 19156 34118 19168
rect 35728 19156 35756 19196
rect 36446 19184 36452 19196
rect 36504 19184 36510 19236
rect 36556 19224 36584 19264
rect 38626 19264 40132 19292
rect 38626 19224 38654 19264
rect 40126 19252 40132 19264
rect 40184 19252 40190 19304
rect 40310 19252 40316 19304
rect 40368 19292 40374 19304
rect 40494 19292 40500 19304
rect 40368 19264 40500 19292
rect 40368 19252 40374 19264
rect 40494 19252 40500 19264
rect 40552 19252 40558 19304
rect 36556 19196 38654 19224
rect 34112 19128 35756 19156
rect 34112 19116 34118 19128
rect 35894 19116 35900 19168
rect 35952 19156 35958 19168
rect 38105 19159 38163 19165
rect 38105 19156 38117 19159
rect 35952 19128 38117 19156
rect 35952 19116 35958 19128
rect 38105 19125 38117 19128
rect 38151 19125 38163 19159
rect 38105 19119 38163 19125
rect 38194 19116 38200 19168
rect 38252 19156 38258 19168
rect 40034 19156 40040 19168
rect 38252 19128 40040 19156
rect 38252 19116 38258 19128
rect 40034 19116 40040 19128
rect 40092 19116 40098 19168
rect 40218 19116 40224 19168
rect 40276 19156 40282 19168
rect 40313 19159 40371 19165
rect 40313 19156 40325 19159
rect 40276 19128 40325 19156
rect 40276 19116 40282 19128
rect 40313 19125 40325 19128
rect 40359 19156 40371 19159
rect 40604 19156 40632 19332
rect 40972 19224 41000 19332
rect 41233 19329 41245 19363
rect 41279 19360 41291 19363
rect 41279 19332 42104 19360
rect 41279 19329 41291 19332
rect 41233 19323 41291 19329
rect 41340 19304 41368 19332
rect 41322 19252 41328 19304
rect 41380 19252 41386 19304
rect 41417 19295 41475 19301
rect 41417 19261 41429 19295
rect 41463 19292 41475 19295
rect 41463 19264 41736 19292
rect 41463 19261 41475 19264
rect 41417 19255 41475 19261
rect 41230 19224 41236 19236
rect 40972 19196 41236 19224
rect 41230 19184 41236 19196
rect 41288 19184 41294 19236
rect 41708 19168 41736 19264
rect 41966 19252 41972 19304
rect 42024 19252 42030 19304
rect 42076 19292 42104 19332
rect 42610 19320 42616 19372
rect 42668 19320 42674 19372
rect 43705 19363 43763 19369
rect 43705 19329 43717 19363
rect 43751 19329 43763 19363
rect 43824 19360 43852 19400
rect 44082 19388 44088 19440
rect 44140 19428 44146 19440
rect 45465 19431 45523 19437
rect 45465 19428 45477 19431
rect 44140 19400 45477 19428
rect 44140 19388 44146 19400
rect 45465 19397 45477 19400
rect 45511 19397 45523 19431
rect 45465 19391 45523 19397
rect 44821 19363 44879 19369
rect 44821 19360 44833 19363
rect 43824 19332 44833 19360
rect 43705 19323 43763 19329
rect 44821 19329 44833 19332
rect 44867 19329 44879 19363
rect 44821 19323 44879 19329
rect 42794 19292 42800 19304
rect 42076 19264 42800 19292
rect 42794 19252 42800 19264
rect 42852 19252 42858 19304
rect 43732 19292 43760 19323
rect 45922 19320 45928 19372
rect 45980 19320 45986 19372
rect 46934 19320 46940 19372
rect 46992 19360 46998 19372
rect 48041 19363 48099 19369
rect 48041 19360 48053 19363
rect 46992 19332 48053 19360
rect 46992 19320 46998 19332
rect 48041 19329 48053 19332
rect 48087 19329 48099 19363
rect 48041 19323 48099 19329
rect 49142 19320 49148 19372
rect 49200 19320 49206 19372
rect 50062 19320 50068 19372
rect 50120 19360 50126 19372
rect 50798 19360 50804 19372
rect 50120 19332 50804 19360
rect 50120 19320 50126 19332
rect 50798 19320 50804 19332
rect 50856 19320 50862 19372
rect 44082 19292 44088 19304
rect 43732 19264 44088 19292
rect 44082 19252 44088 19264
rect 44140 19252 44146 19304
rect 44450 19252 44456 19304
rect 44508 19292 44514 19304
rect 47213 19295 47271 19301
rect 47213 19292 47225 19295
rect 44508 19264 47225 19292
rect 44508 19252 44514 19264
rect 47213 19261 47225 19264
rect 47259 19261 47271 19295
rect 47213 19255 47271 19261
rect 47765 19295 47823 19301
rect 47765 19261 47777 19295
rect 47811 19261 47823 19295
rect 47765 19255 47823 19261
rect 42610 19184 42616 19236
rect 42668 19224 42674 19236
rect 44361 19227 44419 19233
rect 44361 19224 44373 19227
rect 42668 19196 44373 19224
rect 42668 19184 42674 19196
rect 44361 19193 44373 19196
rect 44407 19193 44419 19227
rect 44361 19187 44419 19193
rect 45646 19184 45652 19236
rect 45704 19224 45710 19236
rect 46845 19227 46903 19233
rect 46845 19224 46857 19227
rect 45704 19196 46857 19224
rect 45704 19184 45710 19196
rect 46845 19193 46857 19196
rect 46891 19224 46903 19227
rect 46891 19196 47256 19224
rect 46891 19193 46903 19196
rect 46845 19187 46903 19193
rect 47228 19168 47256 19196
rect 40359 19128 40632 19156
rect 40359 19125 40371 19128
rect 40313 19119 40371 19125
rect 41690 19116 41696 19168
rect 41748 19116 41754 19168
rect 41877 19159 41935 19165
rect 41877 19125 41889 19159
rect 41923 19156 41935 19159
rect 41966 19156 41972 19168
rect 41923 19128 41972 19156
rect 41923 19125 41935 19128
rect 41877 19119 41935 19125
rect 41966 19116 41972 19128
rect 42024 19116 42030 19168
rect 42242 19116 42248 19168
rect 42300 19116 42306 19168
rect 46934 19116 46940 19168
rect 46992 19156 46998 19168
rect 47029 19159 47087 19165
rect 47029 19156 47041 19159
rect 46992 19128 47041 19156
rect 46992 19116 46998 19128
rect 47029 19125 47041 19128
rect 47075 19125 47087 19159
rect 47029 19119 47087 19125
rect 47210 19116 47216 19168
rect 47268 19116 47274 19168
rect 47673 19159 47731 19165
rect 47673 19125 47685 19159
rect 47719 19156 47731 19159
rect 47780 19156 47808 19255
rect 47854 19184 47860 19236
rect 47912 19224 47918 19236
rect 49329 19227 49387 19233
rect 49329 19224 49341 19227
rect 47912 19196 49341 19224
rect 47912 19184 47918 19196
rect 49329 19193 49341 19196
rect 49375 19193 49387 19227
rect 49329 19187 49387 19193
rect 48222 19156 48228 19168
rect 47719 19128 48228 19156
rect 47719 19125 47731 19128
rect 47673 19119 47731 19125
rect 48222 19116 48228 19128
rect 48280 19156 48286 19168
rect 48685 19159 48743 19165
rect 48685 19156 48697 19159
rect 48280 19128 48697 19156
rect 48280 19116 48286 19128
rect 48685 19125 48697 19128
rect 48731 19125 48743 19159
rect 48685 19119 48743 19125
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 3421 18955 3479 18961
rect 3421 18921 3433 18955
rect 3467 18952 3479 18955
rect 5442 18952 5448 18964
rect 3467 18924 5448 18952
rect 3467 18921 3479 18924
rect 3421 18915 3479 18921
rect 5442 18912 5448 18924
rect 5500 18912 5506 18964
rect 5534 18912 5540 18964
rect 5592 18952 5598 18964
rect 6273 18955 6331 18961
rect 6273 18952 6285 18955
rect 5592 18924 6285 18952
rect 5592 18912 5598 18924
rect 6273 18921 6285 18924
rect 6319 18921 6331 18955
rect 6273 18915 6331 18921
rect 7006 18912 7012 18964
rect 7064 18952 7070 18964
rect 7469 18955 7527 18961
rect 7469 18952 7481 18955
rect 7064 18924 7481 18952
rect 7064 18912 7070 18924
rect 7469 18921 7481 18924
rect 7515 18921 7527 18955
rect 7469 18915 7527 18921
rect 7742 18912 7748 18964
rect 7800 18952 7806 18964
rect 8018 18952 8024 18964
rect 7800 18924 8024 18952
rect 7800 18912 7806 18924
rect 8018 18912 8024 18924
rect 8076 18912 8082 18964
rect 9030 18912 9036 18964
rect 9088 18912 9094 18964
rect 10854 18955 10912 18961
rect 10854 18952 10866 18955
rect 9140 18924 10866 18952
rect 3510 18844 3516 18896
rect 3568 18884 3574 18896
rect 3568 18856 7236 18884
rect 3568 18844 3574 18856
rect 3418 18776 3424 18828
rect 3476 18816 3482 18828
rect 4433 18819 4491 18825
rect 4433 18816 4445 18819
rect 3476 18788 4445 18816
rect 3476 18776 3482 18788
rect 4433 18785 4445 18788
rect 4479 18785 4491 18819
rect 7098 18816 7104 18828
rect 4433 18779 4491 18785
rect 4540 18788 7104 18816
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18748 1823 18751
rect 3878 18748 3884 18760
rect 1811 18720 3884 18748
rect 1811 18717 1823 18720
rect 1765 18711 1823 18717
rect 3878 18708 3884 18720
rect 3936 18708 3942 18760
rect 3973 18751 4031 18757
rect 3973 18717 3985 18751
rect 4019 18717 4031 18751
rect 3973 18711 4031 18717
rect 2774 18640 2780 18692
rect 2832 18640 2838 18692
rect 3418 18640 3424 18692
rect 3476 18680 3482 18692
rect 3988 18680 4016 18711
rect 3476 18652 4016 18680
rect 3476 18640 3482 18652
rect 2866 18572 2872 18624
rect 2924 18612 2930 18624
rect 3605 18615 3663 18621
rect 3605 18612 3617 18615
rect 2924 18584 3617 18612
rect 2924 18572 2930 18584
rect 3605 18581 3617 18584
rect 3651 18612 3663 18615
rect 4540 18612 4568 18788
rect 7098 18776 7104 18788
rect 7156 18776 7162 18828
rect 7208 18816 7236 18856
rect 7650 18844 7656 18896
rect 7708 18884 7714 18896
rect 9140 18884 9168 18924
rect 10854 18921 10866 18924
rect 10900 18921 10912 18955
rect 10854 18915 10912 18921
rect 11054 18912 11060 18964
rect 11112 18952 11118 18964
rect 15102 18952 15108 18964
rect 11112 18924 15108 18952
rect 11112 18912 11118 18924
rect 15102 18912 15108 18924
rect 15160 18912 15166 18964
rect 16666 18912 16672 18964
rect 16724 18952 16730 18964
rect 19613 18955 19671 18961
rect 19613 18952 19625 18955
rect 16724 18924 19625 18952
rect 16724 18912 16730 18924
rect 19613 18921 19625 18924
rect 19659 18921 19671 18955
rect 19613 18915 19671 18921
rect 20162 18912 20168 18964
rect 20220 18912 20226 18964
rect 20990 18952 20996 18964
rect 20272 18924 20996 18952
rect 7708 18856 9168 18884
rect 7708 18844 7714 18856
rect 9214 18844 9220 18896
rect 9272 18884 9278 18896
rect 10318 18884 10324 18896
rect 9272 18856 10324 18884
rect 9272 18844 9278 18856
rect 10318 18844 10324 18856
rect 10376 18844 10382 18896
rect 13722 18844 13728 18896
rect 13780 18844 13786 18896
rect 20272 18884 20300 18924
rect 20990 18912 20996 18924
rect 21048 18912 21054 18964
rect 22278 18912 22284 18964
rect 22336 18952 22342 18964
rect 23474 18952 23480 18964
rect 22336 18924 23480 18952
rect 22336 18912 22342 18924
rect 23474 18912 23480 18924
rect 23532 18912 23538 18964
rect 23658 18912 23664 18964
rect 23716 18952 23722 18964
rect 25501 18955 25559 18961
rect 25501 18952 25513 18955
rect 23716 18924 25513 18952
rect 23716 18912 23722 18924
rect 25501 18921 25513 18924
rect 25547 18921 25559 18955
rect 25501 18915 25559 18921
rect 28994 18912 29000 18964
rect 29052 18912 29058 18964
rect 29733 18955 29791 18961
rect 29733 18921 29745 18955
rect 29779 18952 29791 18955
rect 30098 18952 30104 18964
rect 29779 18924 30104 18952
rect 29779 18921 29791 18924
rect 29733 18915 29791 18921
rect 30098 18912 30104 18924
rect 30156 18912 30162 18964
rect 30374 18952 30380 18964
rect 30208 18924 30380 18952
rect 17328 18856 20300 18884
rect 20640 18856 20944 18884
rect 10042 18816 10048 18828
rect 7208 18788 9168 18816
rect 4982 18708 4988 18760
rect 5040 18748 5046 18760
rect 6546 18748 6552 18760
rect 5040 18720 6552 18748
rect 5040 18708 5046 18720
rect 6546 18708 6552 18720
rect 6604 18708 6610 18760
rect 6825 18751 6883 18757
rect 6825 18717 6837 18751
rect 6871 18748 6883 18751
rect 7834 18748 7840 18760
rect 6871 18720 7840 18748
rect 6871 18717 6883 18720
rect 6825 18711 6883 18717
rect 7834 18708 7840 18720
rect 7892 18708 7898 18760
rect 7929 18751 7987 18757
rect 7929 18717 7941 18751
rect 7975 18717 7987 18751
rect 9140 18748 9168 18788
rect 9324 18788 10048 18816
rect 9324 18748 9352 18788
rect 10042 18776 10048 18788
rect 10100 18776 10106 18828
rect 10137 18819 10195 18825
rect 10137 18785 10149 18819
rect 10183 18816 10195 18819
rect 13740 18816 13768 18844
rect 10183 18788 13032 18816
rect 10183 18785 10195 18788
rect 10137 18779 10195 18785
rect 9140 18720 9352 18748
rect 7929 18711 7987 18717
rect 5534 18640 5540 18692
rect 5592 18680 5598 18692
rect 5718 18680 5724 18692
rect 5592 18652 5724 18680
rect 5592 18640 5598 18652
rect 5718 18640 5724 18652
rect 5776 18640 5782 18692
rect 6178 18640 6184 18692
rect 6236 18640 6242 18692
rect 7742 18640 7748 18692
rect 7800 18680 7806 18692
rect 7944 18680 7972 18711
rect 9490 18708 9496 18760
rect 9548 18708 9554 18760
rect 10597 18751 10655 18757
rect 10597 18717 10609 18751
rect 10643 18717 10655 18751
rect 10597 18711 10655 18717
rect 7800 18652 7972 18680
rect 7800 18640 7806 18652
rect 8478 18640 8484 18692
rect 8536 18680 8542 18692
rect 10612 18680 10640 18711
rect 11146 18680 11152 18692
rect 8536 18652 11152 18680
rect 8536 18640 8542 18652
rect 11146 18640 11152 18652
rect 11204 18640 11210 18692
rect 12158 18680 12164 18692
rect 12098 18652 12164 18680
rect 12158 18640 12164 18652
rect 12216 18640 12222 18692
rect 13004 18680 13032 18788
rect 13096 18788 13768 18816
rect 13096 18757 13124 18788
rect 14274 18776 14280 18828
rect 14332 18776 14338 18828
rect 13081 18751 13139 18757
rect 13081 18717 13093 18751
rect 13127 18717 13139 18751
rect 17328 18748 17356 18856
rect 17954 18776 17960 18828
rect 18012 18816 18018 18828
rect 18417 18819 18475 18825
rect 18417 18816 18429 18819
rect 18012 18788 18429 18816
rect 18012 18776 18018 18788
rect 18417 18785 18429 18788
rect 18463 18816 18475 18819
rect 18874 18816 18880 18828
rect 18463 18788 18880 18816
rect 18463 18785 18475 18788
rect 18417 18779 18475 18785
rect 18874 18776 18880 18788
rect 18932 18776 18938 18828
rect 19978 18776 19984 18828
rect 20036 18816 20042 18828
rect 20640 18825 20668 18856
rect 20625 18819 20683 18825
rect 20036 18788 20484 18816
rect 20036 18776 20042 18788
rect 13081 18711 13139 18717
rect 15856 18720 17356 18748
rect 18325 18751 18383 18757
rect 14182 18680 14188 18692
rect 13004 18652 14188 18680
rect 14182 18640 14188 18652
rect 14240 18640 14246 18692
rect 14550 18640 14556 18692
rect 14608 18640 14614 18692
rect 14826 18640 14832 18692
rect 14884 18680 14890 18692
rect 15010 18680 15016 18692
rect 14884 18652 15016 18680
rect 14884 18640 14890 18652
rect 15010 18640 15016 18652
rect 15068 18640 15074 18692
rect 3651 18584 4568 18612
rect 3651 18581 3663 18584
rect 3605 18575 3663 18581
rect 5810 18572 5816 18624
rect 5868 18572 5874 18624
rect 8570 18572 8576 18624
rect 8628 18572 8634 18624
rect 8938 18572 8944 18624
rect 8996 18612 9002 18624
rect 9125 18615 9183 18621
rect 9125 18612 9137 18615
rect 8996 18584 9137 18612
rect 8996 18572 9002 18584
rect 9125 18581 9137 18584
rect 9171 18581 9183 18615
rect 9125 18575 9183 18581
rect 9582 18572 9588 18624
rect 9640 18612 9646 18624
rect 12345 18615 12403 18621
rect 12345 18612 12357 18615
rect 9640 18584 12357 18612
rect 9640 18572 9646 18584
rect 12345 18581 12357 18584
rect 12391 18581 12403 18615
rect 12345 18575 12403 18581
rect 12802 18572 12808 18624
rect 12860 18572 12866 18624
rect 13725 18615 13783 18621
rect 13725 18581 13737 18615
rect 13771 18612 13783 18615
rect 15856 18612 15884 18720
rect 18325 18717 18337 18751
rect 18371 18748 18383 18751
rect 20346 18748 20352 18760
rect 18371 18720 20352 18748
rect 18371 18717 18383 18720
rect 18325 18711 18383 18717
rect 20346 18708 20352 18720
rect 20404 18708 20410 18760
rect 20456 18748 20484 18788
rect 20625 18785 20637 18819
rect 20671 18785 20683 18819
rect 20625 18779 20683 18785
rect 20809 18819 20867 18825
rect 20809 18785 20821 18819
rect 20855 18785 20867 18819
rect 20916 18816 20944 18856
rect 21726 18844 21732 18896
rect 21784 18884 21790 18896
rect 23109 18887 23167 18893
rect 23109 18884 23121 18887
rect 21784 18856 23121 18884
rect 21784 18844 21790 18856
rect 23109 18853 23121 18856
rect 23155 18853 23167 18887
rect 23109 18847 23167 18853
rect 23216 18856 24072 18884
rect 23216 18816 23244 18856
rect 20916 18788 23244 18816
rect 23753 18819 23811 18825
rect 20809 18779 20867 18785
rect 23753 18785 23765 18819
rect 23799 18816 23811 18819
rect 23934 18816 23940 18828
rect 23799 18788 23940 18816
rect 23799 18785 23811 18788
rect 23753 18779 23811 18785
rect 20824 18748 20852 18779
rect 23934 18776 23940 18788
rect 23992 18776 23998 18828
rect 24044 18816 24072 18856
rect 24854 18844 24860 18896
rect 24912 18844 24918 18896
rect 27062 18884 27068 18896
rect 25516 18856 27068 18884
rect 25314 18816 25320 18828
rect 24044 18788 25320 18816
rect 25314 18776 25320 18788
rect 25372 18776 25378 18828
rect 21174 18748 21180 18760
rect 20456 18720 20852 18748
rect 20916 18720 21180 18748
rect 16482 18640 16488 18692
rect 16540 18640 16546 18692
rect 17313 18683 17371 18689
rect 17313 18649 17325 18683
rect 17359 18680 17371 18683
rect 17494 18680 17500 18692
rect 17359 18652 17500 18680
rect 17359 18649 17371 18652
rect 17313 18643 17371 18649
rect 17494 18640 17500 18652
rect 17552 18640 17558 18692
rect 18233 18683 18291 18689
rect 18233 18649 18245 18683
rect 18279 18649 18291 18683
rect 18233 18643 18291 18649
rect 13771 18584 15884 18612
rect 16025 18615 16083 18621
rect 13771 18581 13783 18584
rect 13725 18575 13783 18581
rect 16025 18581 16037 18615
rect 16071 18612 16083 18615
rect 16114 18612 16120 18624
rect 16071 18584 16120 18612
rect 16071 18581 16083 18584
rect 16025 18575 16083 18581
rect 16114 18572 16120 18584
rect 16172 18572 16178 18624
rect 16942 18572 16948 18624
rect 17000 18612 17006 18624
rect 17865 18615 17923 18621
rect 17865 18612 17877 18615
rect 17000 18584 17877 18612
rect 17000 18572 17006 18584
rect 17865 18581 17877 18584
rect 17911 18581 17923 18615
rect 18248 18612 18276 18643
rect 18874 18640 18880 18692
rect 18932 18680 18938 18692
rect 18932 18652 19104 18680
rect 18932 18640 18938 18652
rect 18322 18612 18328 18624
rect 18248 18584 18328 18612
rect 17865 18575 17923 18581
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 18966 18572 18972 18624
rect 19024 18572 19030 18624
rect 19076 18612 19104 18652
rect 19518 18640 19524 18692
rect 19576 18640 19582 18692
rect 20533 18683 20591 18689
rect 20533 18649 20545 18683
rect 20579 18680 20591 18683
rect 20916 18680 20944 18720
rect 21174 18708 21180 18720
rect 21232 18708 21238 18760
rect 21358 18708 21364 18760
rect 21416 18748 21422 18760
rect 22738 18748 22744 18760
rect 21416 18720 22744 18748
rect 21416 18708 21422 18720
rect 22738 18708 22744 18720
rect 22796 18708 22802 18760
rect 23569 18751 23627 18757
rect 23569 18717 23581 18751
rect 23615 18748 23627 18751
rect 25516 18748 25544 18856
rect 27062 18844 27068 18856
rect 27120 18844 27126 18896
rect 27706 18844 27712 18896
rect 27764 18884 27770 18896
rect 27893 18887 27951 18893
rect 27893 18884 27905 18887
rect 27764 18856 27905 18884
rect 27764 18844 27770 18856
rect 27893 18853 27905 18856
rect 27939 18853 27951 18887
rect 30208 18884 30236 18924
rect 30374 18912 30380 18924
rect 30432 18912 30438 18964
rect 32214 18912 32220 18964
rect 32272 18952 32278 18964
rect 32272 18924 44128 18952
rect 32272 18912 32278 18924
rect 30558 18884 30564 18896
rect 27893 18847 27951 18853
rect 28460 18856 30236 18884
rect 30300 18856 30564 18884
rect 25958 18776 25964 18828
rect 26016 18816 26022 18828
rect 26053 18819 26111 18825
rect 26053 18816 26065 18819
rect 26016 18788 26065 18816
rect 26016 18776 26022 18788
rect 26053 18785 26065 18788
rect 26099 18785 26111 18819
rect 26053 18779 26111 18785
rect 26510 18776 26516 18828
rect 26568 18776 26574 18828
rect 27338 18776 27344 18828
rect 27396 18776 27402 18828
rect 28460 18816 28488 18856
rect 27540 18788 28488 18816
rect 28537 18819 28595 18825
rect 23615 18720 25544 18748
rect 25869 18751 25927 18757
rect 23615 18717 23627 18720
rect 23569 18711 23627 18717
rect 25869 18717 25881 18751
rect 25915 18748 25927 18751
rect 26528 18748 26556 18776
rect 25915 18720 26556 18748
rect 27157 18751 27215 18757
rect 25915 18717 25927 18720
rect 25869 18711 25927 18717
rect 27157 18717 27169 18751
rect 27203 18748 27215 18751
rect 27430 18748 27436 18760
rect 27203 18720 27436 18748
rect 27203 18717 27215 18720
rect 27157 18711 27215 18717
rect 27430 18708 27436 18720
rect 27488 18708 27494 18760
rect 20579 18652 20944 18680
rect 22189 18683 22247 18689
rect 20579 18649 20591 18652
rect 20533 18643 20591 18649
rect 22189 18649 22201 18683
rect 22235 18680 22247 18683
rect 22830 18680 22836 18692
rect 22235 18652 22836 18680
rect 22235 18649 22247 18652
rect 22189 18643 22247 18649
rect 22830 18640 22836 18652
rect 22888 18640 22894 18692
rect 24673 18683 24731 18689
rect 24673 18649 24685 18683
rect 24719 18649 24731 18683
rect 24673 18643 24731 18649
rect 25961 18683 26019 18689
rect 25961 18649 25973 18683
rect 26007 18680 26019 18683
rect 27540 18680 27568 18788
rect 28537 18785 28549 18819
rect 28583 18816 28595 18819
rect 28718 18816 28724 18828
rect 28583 18788 28724 18816
rect 28583 18785 28595 18788
rect 28537 18779 28595 18785
rect 28718 18776 28724 18788
rect 28776 18776 28782 18828
rect 29362 18776 29368 18828
rect 29420 18816 29426 18828
rect 30300 18825 30328 18856
rect 30558 18844 30564 18856
rect 30616 18844 30622 18896
rect 32582 18844 32588 18896
rect 32640 18884 32646 18896
rect 32769 18887 32827 18893
rect 32769 18884 32781 18887
rect 32640 18856 32781 18884
rect 32640 18844 32646 18856
rect 32769 18853 32781 18856
rect 32815 18853 32827 18887
rect 38013 18887 38071 18893
rect 32769 18847 32827 18853
rect 33244 18856 36400 18884
rect 30193 18819 30251 18825
rect 30193 18816 30205 18819
rect 29420 18788 30205 18816
rect 29420 18776 29426 18788
rect 30193 18785 30205 18788
rect 30239 18785 30251 18819
rect 30193 18779 30251 18785
rect 30285 18819 30343 18825
rect 30285 18785 30297 18819
rect 30331 18785 30343 18819
rect 30285 18779 30343 18785
rect 32217 18819 32275 18825
rect 32217 18785 32229 18819
rect 32263 18816 32275 18819
rect 32306 18816 32312 18828
rect 32263 18788 32312 18816
rect 32263 18785 32275 18788
rect 32217 18779 32275 18785
rect 28261 18751 28319 18757
rect 28261 18717 28273 18751
rect 28307 18748 28319 18751
rect 28902 18748 28908 18760
rect 28307 18720 28908 18748
rect 28307 18717 28319 18720
rect 28261 18711 28319 18717
rect 28902 18708 28908 18720
rect 28960 18708 28966 18760
rect 29270 18708 29276 18760
rect 29328 18708 29334 18760
rect 29730 18708 29736 18760
rect 29788 18748 29794 18760
rect 30101 18751 30159 18757
rect 30101 18748 30113 18751
rect 29788 18720 30113 18748
rect 29788 18708 29794 18720
rect 30101 18717 30113 18720
rect 30147 18717 30159 18751
rect 30208 18748 30236 18779
rect 32306 18776 32312 18788
rect 32364 18776 32370 18828
rect 33244 18825 33272 18856
rect 33229 18819 33287 18825
rect 33229 18785 33241 18819
rect 33275 18785 33287 18819
rect 33229 18779 33287 18785
rect 33413 18819 33471 18825
rect 33413 18785 33425 18819
rect 33459 18785 33471 18819
rect 33413 18779 33471 18785
rect 31389 18751 31447 18757
rect 30208 18720 31340 18748
rect 30101 18711 30159 18717
rect 28166 18680 28172 18692
rect 26007 18652 27568 18680
rect 27816 18652 28172 18680
rect 26007 18649 26019 18652
rect 25961 18643 26019 18649
rect 22278 18612 22284 18624
rect 19076 18584 22284 18612
rect 22278 18572 22284 18584
rect 22336 18612 22342 18624
rect 22557 18615 22615 18621
rect 22557 18612 22569 18615
rect 22336 18584 22569 18612
rect 22336 18572 22342 18584
rect 22557 18581 22569 18584
rect 22603 18581 22615 18615
rect 22557 18575 22615 18581
rect 22738 18572 22744 18624
rect 22796 18572 22802 18624
rect 23474 18572 23480 18624
rect 23532 18572 23538 18624
rect 23750 18572 23756 18624
rect 23808 18612 23814 18624
rect 24121 18615 24179 18621
rect 24121 18612 24133 18615
rect 23808 18584 24133 18612
rect 23808 18572 23814 18584
rect 24121 18581 24133 18584
rect 24167 18581 24179 18615
rect 24121 18575 24179 18581
rect 24302 18572 24308 18624
rect 24360 18612 24366 18624
rect 24688 18612 24716 18643
rect 25225 18615 25283 18621
rect 25225 18612 25237 18615
rect 24360 18584 25237 18612
rect 24360 18572 24366 18584
rect 25225 18581 25237 18584
rect 25271 18612 25283 18615
rect 25866 18612 25872 18624
rect 25271 18584 25872 18612
rect 25271 18581 25283 18584
rect 25225 18575 25283 18581
rect 25866 18572 25872 18584
rect 25924 18572 25930 18624
rect 26326 18572 26332 18624
rect 26384 18612 26390 18624
rect 26697 18615 26755 18621
rect 26697 18612 26709 18615
rect 26384 18584 26709 18612
rect 26384 18572 26390 18584
rect 26697 18581 26709 18584
rect 26743 18581 26755 18615
rect 26697 18575 26755 18581
rect 27065 18615 27123 18621
rect 27065 18581 27077 18615
rect 27111 18612 27123 18615
rect 27816 18612 27844 18652
rect 28166 18640 28172 18652
rect 28224 18640 28230 18692
rect 28353 18683 28411 18689
rect 28353 18649 28365 18683
rect 28399 18680 28411 18683
rect 29822 18680 29828 18692
rect 28399 18652 29828 18680
rect 28399 18649 28411 18652
rect 28353 18643 28411 18649
rect 29822 18640 29828 18652
rect 29880 18640 29886 18692
rect 30116 18680 30144 18711
rect 30929 18683 30987 18689
rect 30929 18680 30941 18683
rect 30116 18652 30941 18680
rect 30929 18649 30941 18652
rect 30975 18680 30987 18683
rect 31110 18680 31116 18692
rect 30975 18652 31116 18680
rect 30975 18649 30987 18652
rect 30929 18643 30987 18649
rect 31110 18640 31116 18652
rect 31168 18640 31174 18692
rect 31312 18680 31340 18720
rect 31389 18717 31401 18751
rect 31435 18748 31447 18751
rect 31570 18748 31576 18760
rect 31435 18720 31576 18748
rect 31435 18717 31447 18720
rect 31389 18711 31447 18717
rect 31570 18708 31576 18720
rect 31628 18708 31634 18760
rect 32122 18708 32128 18760
rect 32180 18748 32186 18760
rect 33428 18748 33456 18779
rect 33594 18776 33600 18828
rect 33652 18816 33658 18828
rect 33870 18816 33876 18828
rect 33652 18788 33876 18816
rect 33652 18776 33658 18788
rect 33870 18776 33876 18788
rect 33928 18776 33934 18828
rect 34238 18776 34244 18828
rect 34296 18816 34302 18828
rect 34333 18819 34391 18825
rect 34333 18816 34345 18819
rect 34296 18788 34345 18816
rect 34296 18776 34302 18788
rect 34333 18785 34345 18788
rect 34379 18785 34391 18819
rect 34333 18779 34391 18785
rect 34606 18776 34612 18828
rect 34664 18816 34670 18828
rect 35437 18819 35495 18825
rect 35437 18816 35449 18819
rect 34664 18788 35449 18816
rect 34664 18776 34670 18788
rect 35437 18785 35449 18788
rect 35483 18785 35495 18819
rect 35437 18779 35495 18785
rect 35989 18819 36047 18825
rect 35989 18785 36001 18819
rect 36035 18816 36047 18819
rect 36078 18816 36084 18828
rect 36035 18788 36084 18816
rect 36035 18785 36047 18788
rect 35989 18779 36047 18785
rect 36078 18776 36084 18788
rect 36136 18776 36142 18828
rect 36262 18776 36268 18828
rect 36320 18776 36326 18828
rect 36372 18816 36400 18856
rect 38013 18853 38025 18887
rect 38059 18884 38071 18887
rect 38562 18884 38568 18896
rect 38059 18856 38568 18884
rect 38059 18853 38071 18856
rect 38013 18847 38071 18853
rect 38562 18844 38568 18856
rect 38620 18844 38626 18896
rect 39574 18844 39580 18896
rect 39632 18844 39638 18896
rect 39666 18844 39672 18896
rect 39724 18884 39730 18896
rect 44100 18884 44128 18924
rect 44174 18912 44180 18964
rect 44232 18952 44238 18964
rect 44453 18955 44511 18961
rect 44453 18952 44465 18955
rect 44232 18924 44465 18952
rect 44232 18912 44238 18924
rect 44453 18921 44465 18924
rect 44499 18921 44511 18955
rect 44453 18915 44511 18921
rect 45833 18955 45891 18961
rect 45833 18921 45845 18955
rect 45879 18952 45891 18955
rect 46290 18952 46296 18964
rect 45879 18924 46296 18952
rect 45879 18921 45891 18924
rect 45833 18915 45891 18921
rect 46290 18912 46296 18924
rect 46348 18912 46354 18964
rect 47394 18912 47400 18964
rect 47452 18912 47458 18964
rect 48406 18912 48412 18964
rect 48464 18912 48470 18964
rect 48958 18912 48964 18964
rect 49016 18952 49022 18964
rect 49053 18955 49111 18961
rect 49053 18952 49065 18955
rect 49016 18924 49065 18952
rect 49016 18912 49022 18924
rect 49053 18921 49065 18924
rect 49099 18921 49111 18955
rect 49053 18915 49111 18921
rect 47118 18884 47124 18896
rect 39724 18856 40172 18884
rect 39724 18844 39730 18856
rect 38746 18816 38752 18828
rect 36372 18788 38752 18816
rect 38746 18776 38752 18788
rect 38804 18776 38810 18828
rect 39117 18819 39175 18825
rect 39117 18785 39129 18819
rect 39163 18816 39175 18819
rect 39850 18816 39856 18828
rect 39163 18788 39856 18816
rect 39163 18785 39175 18788
rect 39117 18779 39175 18785
rect 39850 18776 39856 18788
rect 39908 18776 39914 18828
rect 40144 18816 40172 18856
rect 41340 18856 43392 18884
rect 44100 18856 47124 18884
rect 41340 18816 41368 18856
rect 40144 18788 41368 18816
rect 41598 18776 41604 18828
rect 41656 18816 41662 18828
rect 42610 18816 42616 18828
rect 41656 18788 42616 18816
rect 41656 18776 41662 18788
rect 42610 18776 42616 18788
rect 42668 18776 42674 18828
rect 36170 18748 36176 18760
rect 32180 18720 33272 18748
rect 33428 18720 36176 18748
rect 32180 18708 32186 18720
rect 32214 18680 32220 18692
rect 31312 18652 32220 18680
rect 32214 18640 32220 18652
rect 32272 18640 32278 18692
rect 32398 18640 32404 18692
rect 32456 18680 32462 18692
rect 33137 18683 33195 18689
rect 33137 18680 33149 18683
rect 32456 18652 33149 18680
rect 32456 18640 32462 18652
rect 33137 18649 33149 18652
rect 33183 18649 33195 18683
rect 33244 18680 33272 18720
rect 36170 18708 36176 18720
rect 36228 18708 36234 18760
rect 38654 18708 38660 18760
rect 38712 18748 38718 18760
rect 39758 18748 39764 18760
rect 38712 18720 39764 18748
rect 38712 18708 38718 18720
rect 39758 18708 39764 18720
rect 39816 18708 39822 18760
rect 40034 18708 40040 18760
rect 40092 18708 40098 18760
rect 42150 18748 42156 18760
rect 41708 18744 42156 18748
rect 41616 18720 42156 18744
rect 41616 18716 41736 18720
rect 34054 18680 34060 18692
rect 33244 18652 34060 18680
rect 33137 18643 33195 18649
rect 34054 18640 34060 18652
rect 34112 18640 34118 18692
rect 34149 18683 34207 18689
rect 34149 18649 34161 18683
rect 34195 18680 34207 18683
rect 34330 18680 34336 18692
rect 34195 18652 34336 18680
rect 34195 18649 34207 18652
rect 34149 18643 34207 18649
rect 34330 18640 34336 18652
rect 34388 18640 34394 18692
rect 34440 18652 35204 18680
rect 27111 18584 27844 18612
rect 27111 18581 27123 18584
rect 27065 18575 27123 18581
rect 28074 18572 28080 18624
rect 28132 18612 28138 18624
rect 29181 18615 29239 18621
rect 29181 18612 29193 18615
rect 28132 18584 29193 18612
rect 28132 18572 28138 18584
rect 29181 18581 29193 18584
rect 29227 18612 29239 18615
rect 29362 18612 29368 18624
rect 29227 18584 29368 18612
rect 29227 18581 29239 18584
rect 29181 18575 29239 18581
rect 29362 18572 29368 18584
rect 29420 18572 29426 18624
rect 29454 18572 29460 18624
rect 29512 18612 29518 18624
rect 29638 18612 29644 18624
rect 29512 18584 29644 18612
rect 29512 18572 29518 18584
rect 29638 18572 29644 18584
rect 29696 18612 29702 18624
rect 30745 18615 30803 18621
rect 30745 18612 30757 18615
rect 29696 18584 30757 18612
rect 29696 18572 29702 18584
rect 30745 18581 30757 18584
rect 30791 18581 30803 18615
rect 30745 18575 30803 18581
rect 33318 18572 33324 18624
rect 33376 18612 33382 18624
rect 34440 18612 34468 18652
rect 33376 18584 34468 18612
rect 33376 18572 33382 18584
rect 34790 18572 34796 18624
rect 34848 18612 34854 18624
rect 34885 18615 34943 18621
rect 34885 18612 34897 18615
rect 34848 18584 34897 18612
rect 34848 18572 34854 18584
rect 34885 18581 34897 18584
rect 34931 18581 34943 18615
rect 35176 18612 35204 18652
rect 35250 18640 35256 18692
rect 35308 18640 35314 18692
rect 35345 18683 35403 18689
rect 35345 18649 35357 18683
rect 35391 18680 35403 18683
rect 35434 18680 35440 18692
rect 35391 18652 35440 18680
rect 35391 18649 35403 18652
rect 35345 18643 35403 18649
rect 35434 18640 35440 18652
rect 35492 18640 35498 18692
rect 36541 18683 36599 18689
rect 35544 18652 36032 18680
rect 35544 18612 35572 18652
rect 35176 18584 35572 18612
rect 36004 18612 36032 18652
rect 36541 18649 36553 18683
rect 36587 18680 36599 18683
rect 36814 18680 36820 18692
rect 36587 18652 36820 18680
rect 36587 18649 36599 18652
rect 36541 18643 36599 18649
rect 36814 18640 36820 18652
rect 36872 18640 36878 18692
rect 37826 18680 37832 18692
rect 37766 18652 37832 18680
rect 37826 18640 37832 18652
rect 37884 18680 37890 18692
rect 39942 18680 39948 18692
rect 37884 18652 39948 18680
rect 37884 18640 37890 18652
rect 39942 18640 39948 18652
rect 40000 18640 40006 18692
rect 40310 18689 40316 18692
rect 40300 18683 40316 18689
rect 40300 18649 40312 18683
rect 40300 18643 40316 18649
rect 40310 18640 40316 18643
rect 40368 18640 40374 18692
rect 41616 18680 41644 18716
rect 42150 18708 42156 18720
rect 42208 18708 42214 18760
rect 42242 18708 42248 18760
rect 42300 18708 42306 18760
rect 43364 18757 43392 18856
rect 47118 18844 47124 18856
rect 47176 18844 47182 18896
rect 47412 18884 47440 18912
rect 49421 18887 49479 18893
rect 49421 18884 49433 18887
rect 47412 18856 49433 18884
rect 49421 18853 49433 18856
rect 49467 18853 49479 18887
rect 49421 18847 49479 18853
rect 43714 18776 43720 18828
rect 43772 18816 43778 18828
rect 44818 18816 44824 18828
rect 43772 18788 44824 18816
rect 43772 18776 43778 18788
rect 44818 18776 44824 18788
rect 44876 18776 44882 18828
rect 46937 18819 46995 18825
rect 46937 18816 46949 18819
rect 45204 18788 46949 18816
rect 43349 18751 43407 18757
rect 43349 18717 43361 18751
rect 43395 18717 43407 18751
rect 43349 18711 43407 18717
rect 43898 18708 43904 18760
rect 43956 18748 43962 18760
rect 45204 18757 45232 18788
rect 46937 18785 46949 18788
rect 46983 18785 46995 18819
rect 46937 18779 46995 18785
rect 44637 18751 44695 18757
rect 44637 18748 44649 18751
rect 43956 18720 44649 18748
rect 43956 18708 43962 18720
rect 44637 18717 44649 18720
rect 44683 18717 44695 18751
rect 44637 18711 44695 18717
rect 45189 18751 45247 18757
rect 45189 18717 45201 18751
rect 45235 18717 45247 18751
rect 45189 18711 45247 18717
rect 46290 18708 46296 18760
rect 46348 18708 46354 18760
rect 47765 18751 47823 18757
rect 47765 18717 47777 18751
rect 47811 18717 47823 18751
rect 47765 18711 47823 18717
rect 47780 18680 47808 18711
rect 41538 18652 41644 18680
rect 41800 18652 47808 18680
rect 48961 18683 49019 18689
rect 36722 18612 36728 18624
rect 36004 18584 36728 18612
rect 34885 18575 34943 18581
rect 36722 18572 36728 18584
rect 36780 18572 36786 18624
rect 38473 18615 38531 18621
rect 38473 18581 38485 18615
rect 38519 18612 38531 18615
rect 38746 18612 38752 18624
rect 38519 18584 38752 18612
rect 38519 18581 38531 18584
rect 38473 18575 38531 18581
rect 38746 18572 38752 18584
rect 38804 18572 38810 18624
rect 38838 18572 38844 18624
rect 38896 18572 38902 18624
rect 38930 18572 38936 18624
rect 38988 18572 38994 18624
rect 40586 18572 40592 18624
rect 40644 18612 40650 18624
rect 41598 18612 41604 18624
rect 40644 18584 41604 18612
rect 40644 18572 40650 18584
rect 41598 18572 41604 18584
rect 41656 18572 41662 18624
rect 41690 18572 41696 18624
rect 41748 18612 41754 18624
rect 41800 18621 41828 18652
rect 48961 18649 48973 18683
rect 49007 18680 49019 18683
rect 49694 18680 49700 18692
rect 49007 18652 49700 18680
rect 49007 18649 49019 18652
rect 48961 18643 49019 18649
rect 49694 18640 49700 18652
rect 49752 18640 49758 18692
rect 41785 18615 41843 18621
rect 41785 18612 41797 18615
rect 41748 18584 41797 18612
rect 41748 18572 41754 18584
rect 41785 18581 41797 18584
rect 41831 18581 41843 18615
rect 41785 18575 41843 18581
rect 42610 18572 42616 18624
rect 42668 18612 42674 18624
rect 42889 18615 42947 18621
rect 42889 18612 42901 18615
rect 42668 18584 42901 18612
rect 42668 18572 42674 18584
rect 42889 18581 42901 18584
rect 42935 18581 42947 18615
rect 42889 18575 42947 18581
rect 43714 18572 43720 18624
rect 43772 18612 43778 18624
rect 43993 18615 44051 18621
rect 43993 18612 44005 18615
rect 43772 18584 44005 18612
rect 43772 18572 43778 18584
rect 43993 18581 44005 18584
rect 44039 18581 44051 18615
rect 43993 18575 44051 18581
rect 44266 18572 44272 18624
rect 44324 18612 44330 18624
rect 47213 18615 47271 18621
rect 47213 18612 47225 18615
rect 44324 18584 47225 18612
rect 44324 18572 44330 18584
rect 47213 18581 47225 18584
rect 47259 18581 47271 18615
rect 47213 18575 47271 18581
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 3329 18411 3387 18417
rect 3329 18377 3341 18411
rect 3375 18408 3387 18411
rect 3510 18408 3516 18420
rect 3375 18380 3516 18408
rect 3375 18377 3387 18380
rect 3329 18371 3387 18377
rect 3510 18368 3516 18380
rect 3568 18368 3574 18420
rect 3602 18368 3608 18420
rect 3660 18368 3666 18420
rect 10965 18411 11023 18417
rect 10965 18408 10977 18411
rect 6104 18380 10977 18408
rect 6104 18340 6132 18380
rect 10965 18377 10977 18380
rect 11011 18377 11023 18411
rect 10965 18371 11023 18377
rect 12158 18368 12164 18420
rect 12216 18408 12222 18420
rect 12618 18408 12624 18420
rect 12216 18380 12624 18408
rect 12216 18368 12222 18380
rect 12618 18368 12624 18380
rect 12676 18408 12682 18420
rect 12676 18380 13032 18408
rect 12676 18368 12682 18380
rect 2746 18312 6132 18340
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18272 1823 18275
rect 2746 18272 2774 18312
rect 6546 18300 6552 18352
rect 6604 18340 6610 18352
rect 8757 18343 8815 18349
rect 8757 18340 8769 18343
rect 6604 18312 8769 18340
rect 6604 18300 6610 18312
rect 8757 18309 8769 18312
rect 8803 18309 8815 18343
rect 8757 18303 8815 18309
rect 8846 18300 8852 18352
rect 8904 18340 8910 18352
rect 8904 18312 9246 18340
rect 8904 18300 8910 18312
rect 10042 18300 10048 18352
rect 10100 18340 10106 18352
rect 10870 18340 10876 18352
rect 10100 18312 10876 18340
rect 10100 18300 10106 18312
rect 10870 18300 10876 18312
rect 10928 18300 10934 18352
rect 11054 18300 11060 18352
rect 11112 18340 11118 18352
rect 12897 18343 12955 18349
rect 12897 18340 12909 18343
rect 11112 18312 12909 18340
rect 11112 18300 11118 18312
rect 12897 18309 12909 18312
rect 12943 18309 12955 18343
rect 13004 18340 13032 18380
rect 14642 18368 14648 18420
rect 14700 18408 14706 18420
rect 16853 18411 16911 18417
rect 16853 18408 16865 18411
rect 14700 18380 16865 18408
rect 14700 18368 14706 18380
rect 16853 18377 16865 18380
rect 16899 18377 16911 18411
rect 16853 18371 16911 18377
rect 17310 18368 17316 18420
rect 17368 18368 17374 18420
rect 18233 18411 18291 18417
rect 18233 18377 18245 18411
rect 18279 18408 18291 18411
rect 18690 18408 18696 18420
rect 18279 18380 18696 18408
rect 18279 18377 18291 18380
rect 18233 18371 18291 18377
rect 18690 18368 18696 18380
rect 18748 18368 18754 18420
rect 19153 18411 19211 18417
rect 19153 18377 19165 18411
rect 19199 18408 19211 18411
rect 19199 18380 22094 18408
rect 19199 18377 19211 18380
rect 19153 18371 19211 18377
rect 13354 18340 13360 18352
rect 13004 18312 13360 18340
rect 12897 18303 12955 18309
rect 13354 18300 13360 18312
rect 13412 18300 13418 18352
rect 14182 18300 14188 18352
rect 14240 18340 14246 18352
rect 19889 18343 19947 18349
rect 19889 18340 19901 18343
rect 14240 18312 19901 18340
rect 14240 18300 14246 18312
rect 19889 18309 19901 18312
rect 19935 18309 19947 18343
rect 22066 18340 22094 18380
rect 22186 18368 22192 18420
rect 22244 18368 22250 18420
rect 23474 18368 23480 18420
rect 23532 18408 23538 18420
rect 25501 18411 25559 18417
rect 25501 18408 25513 18411
rect 23532 18380 25513 18408
rect 23532 18368 23538 18380
rect 25501 18377 25513 18380
rect 25547 18377 25559 18411
rect 25501 18371 25559 18377
rect 25774 18368 25780 18420
rect 25832 18408 25838 18420
rect 25869 18411 25927 18417
rect 25869 18408 25881 18411
rect 25832 18380 25881 18408
rect 25832 18368 25838 18380
rect 25869 18377 25881 18380
rect 25915 18408 25927 18411
rect 25915 18380 26372 18408
rect 25915 18377 25927 18380
rect 25869 18371 25927 18377
rect 23109 18343 23167 18349
rect 23109 18340 23121 18343
rect 22066 18312 23121 18340
rect 19889 18303 19947 18309
rect 23109 18309 23121 18312
rect 23155 18309 23167 18343
rect 24762 18340 24768 18352
rect 24334 18312 24768 18340
rect 23109 18303 23167 18309
rect 24762 18300 24768 18312
rect 24820 18300 24826 18352
rect 1811 18244 2774 18272
rect 1811 18241 1823 18244
rect 1765 18235 1823 18241
rect 3602 18232 3608 18284
rect 3660 18272 3666 18284
rect 3789 18275 3847 18281
rect 3789 18272 3801 18275
rect 3660 18244 3801 18272
rect 3660 18232 3666 18244
rect 3789 18241 3801 18244
rect 3835 18241 3847 18275
rect 3789 18235 3847 18241
rect 4249 18275 4307 18281
rect 4249 18241 4261 18275
rect 4295 18241 4307 18275
rect 4249 18235 4307 18241
rect 5353 18275 5411 18281
rect 5353 18241 5365 18275
rect 5399 18272 5411 18275
rect 5994 18272 6000 18284
rect 5399 18244 6000 18272
rect 5399 18241 5411 18244
rect 5353 18235 5411 18241
rect 2038 18164 2044 18216
rect 2096 18164 2102 18216
rect 4264 18204 4292 18235
rect 5994 18232 6000 18244
rect 6052 18232 6058 18284
rect 6917 18275 6975 18281
rect 6917 18241 6929 18275
rect 6963 18272 6975 18275
rect 7006 18272 7012 18284
rect 6963 18244 7012 18272
rect 6963 18241 6975 18244
rect 6917 18235 6975 18241
rect 7006 18232 7012 18244
rect 7064 18232 7070 18284
rect 7374 18232 7380 18284
rect 7432 18232 7438 18284
rect 8478 18232 8484 18284
rect 8536 18232 8542 18284
rect 11790 18232 11796 18284
rect 11848 18232 11854 18284
rect 15197 18275 15255 18281
rect 15197 18241 15209 18275
rect 15243 18272 15255 18275
rect 15562 18272 15568 18284
rect 15243 18244 15568 18272
rect 15243 18241 15255 18244
rect 15197 18235 15255 18241
rect 15562 18232 15568 18244
rect 15620 18232 15626 18284
rect 16117 18275 16175 18281
rect 16117 18241 16129 18275
rect 16163 18241 16175 18275
rect 16117 18235 16175 18241
rect 7098 18204 7104 18216
rect 4264 18176 7104 18204
rect 7098 18164 7104 18176
rect 7156 18164 7162 18216
rect 8846 18164 8852 18216
rect 8904 18204 8910 18216
rect 8904 18176 10180 18204
rect 8904 18164 8910 18176
rect 3878 18096 3884 18148
rect 3936 18136 3942 18148
rect 6733 18139 6791 18145
rect 6733 18136 6745 18139
rect 3936 18108 6745 18136
rect 3936 18096 3942 18108
rect 6733 18105 6745 18108
rect 6779 18105 6791 18139
rect 7834 18136 7840 18148
rect 6733 18099 6791 18105
rect 7576 18108 7840 18136
rect 4893 18071 4951 18077
rect 4893 18037 4905 18071
rect 4939 18068 4951 18071
rect 5718 18068 5724 18080
rect 4939 18040 5724 18068
rect 4939 18037 4951 18040
rect 4893 18031 4951 18037
rect 5718 18028 5724 18040
rect 5776 18028 5782 18080
rect 5902 18028 5908 18080
rect 5960 18068 5966 18080
rect 5997 18071 6055 18077
rect 5997 18068 6009 18071
rect 5960 18040 6009 18068
rect 5960 18028 5966 18040
rect 5997 18037 6009 18040
rect 6043 18037 6055 18071
rect 5997 18031 6055 18037
rect 6457 18071 6515 18077
rect 6457 18037 6469 18071
rect 6503 18068 6515 18071
rect 7576 18068 7604 18108
rect 7834 18096 7840 18108
rect 7892 18136 7898 18148
rect 8294 18136 8300 18148
rect 7892 18108 8300 18136
rect 7892 18096 7898 18108
rect 8294 18096 8300 18108
rect 8352 18096 8358 18148
rect 10152 18136 10180 18176
rect 10226 18164 10232 18216
rect 10284 18164 10290 18216
rect 11974 18164 11980 18216
rect 12032 18204 12038 18216
rect 12621 18207 12679 18213
rect 12621 18204 12633 18207
rect 12032 18176 12633 18204
rect 12032 18164 12038 18176
rect 12621 18173 12633 18176
rect 12667 18173 12679 18207
rect 12621 18167 12679 18173
rect 12158 18136 12164 18148
rect 10152 18108 12164 18136
rect 12158 18096 12164 18108
rect 12216 18096 12222 18148
rect 12345 18139 12403 18145
rect 12345 18105 12357 18139
rect 12391 18136 12403 18139
rect 12526 18136 12532 18148
rect 12391 18108 12532 18136
rect 12391 18105 12403 18108
rect 12345 18099 12403 18105
rect 12526 18096 12532 18108
rect 12584 18096 12590 18148
rect 6503 18040 7604 18068
rect 8021 18071 8079 18077
rect 6503 18037 6515 18040
rect 6457 18031 6515 18037
rect 8021 18037 8033 18071
rect 8067 18068 8079 18071
rect 9398 18068 9404 18080
rect 8067 18040 9404 18068
rect 8067 18037 8079 18040
rect 8021 18031 8079 18037
rect 9398 18028 9404 18040
rect 9456 18028 9462 18080
rect 11238 18028 11244 18080
rect 11296 18068 11302 18080
rect 11885 18071 11943 18077
rect 11885 18068 11897 18071
rect 11296 18040 11897 18068
rect 11296 18028 11302 18040
rect 11885 18037 11897 18040
rect 11931 18037 11943 18071
rect 12636 18068 12664 18167
rect 12894 18164 12900 18216
rect 12952 18204 12958 18216
rect 14369 18207 14427 18213
rect 14369 18204 14381 18207
rect 12952 18176 14381 18204
rect 12952 18164 12958 18176
rect 14369 18173 14381 18176
rect 14415 18173 14427 18207
rect 14369 18167 14427 18173
rect 15286 18164 15292 18216
rect 15344 18164 15350 18216
rect 15473 18207 15531 18213
rect 15473 18173 15485 18207
rect 15519 18204 15531 18207
rect 15838 18204 15844 18216
rect 15519 18176 15844 18204
rect 15519 18173 15531 18176
rect 15473 18167 15531 18173
rect 15838 18164 15844 18176
rect 15896 18164 15902 18216
rect 14642 18096 14648 18148
rect 14700 18136 14706 18148
rect 16132 18136 16160 18235
rect 16298 18232 16304 18284
rect 16356 18272 16362 18284
rect 17221 18275 17279 18281
rect 17221 18272 17233 18275
rect 16356 18244 17233 18272
rect 16356 18232 16362 18244
rect 17221 18241 17233 18244
rect 17267 18241 17279 18275
rect 17221 18235 17279 18241
rect 17862 18232 17868 18284
rect 17920 18272 17926 18284
rect 18509 18275 18567 18281
rect 18509 18272 18521 18275
rect 17920 18244 18521 18272
rect 17920 18232 17926 18244
rect 18509 18241 18521 18244
rect 18555 18241 18567 18275
rect 18509 18235 18567 18241
rect 19150 18232 19156 18284
rect 19208 18272 19214 18284
rect 19426 18272 19432 18284
rect 19208 18244 19432 18272
rect 19208 18232 19214 18244
rect 19426 18232 19432 18244
rect 19484 18232 19490 18284
rect 19613 18275 19671 18281
rect 19613 18272 19625 18275
rect 19536 18244 19625 18272
rect 16206 18164 16212 18216
rect 16264 18204 16270 18216
rect 17405 18207 17463 18213
rect 17405 18204 17417 18207
rect 16264 18176 17417 18204
rect 16264 18164 16270 18176
rect 17405 18173 17417 18176
rect 17451 18173 17463 18207
rect 17405 18167 17463 18173
rect 17494 18164 17500 18216
rect 17552 18204 17558 18216
rect 19536 18204 19564 18244
rect 19613 18241 19625 18244
rect 19659 18241 19671 18275
rect 19613 18235 19671 18241
rect 20990 18232 20996 18284
rect 21048 18272 21054 18284
rect 22002 18272 22008 18284
rect 21048 18244 22008 18272
rect 21048 18232 21054 18244
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 22097 18275 22155 18281
rect 22097 18241 22109 18275
rect 22143 18272 22155 18275
rect 22278 18272 22284 18284
rect 22143 18244 22284 18272
rect 22143 18241 22155 18244
rect 22097 18235 22155 18241
rect 22278 18232 22284 18244
rect 22336 18232 22342 18284
rect 25130 18232 25136 18284
rect 25188 18272 25194 18284
rect 25225 18275 25283 18281
rect 25225 18272 25237 18275
rect 25188 18244 25237 18272
rect 25188 18232 25194 18244
rect 25225 18241 25237 18244
rect 25271 18272 25283 18275
rect 26344 18272 26372 18380
rect 26602 18368 26608 18420
rect 26660 18408 26666 18420
rect 26789 18411 26847 18417
rect 26789 18408 26801 18411
rect 26660 18380 26801 18408
rect 26660 18368 26666 18380
rect 26789 18377 26801 18380
rect 26835 18408 26847 18411
rect 27062 18408 27068 18420
rect 26835 18380 27068 18408
rect 26835 18377 26847 18380
rect 26789 18371 26847 18377
rect 27062 18368 27068 18380
rect 27120 18368 27126 18420
rect 27246 18368 27252 18420
rect 27304 18408 27310 18420
rect 30009 18411 30067 18417
rect 30009 18408 30021 18411
rect 27304 18380 30021 18408
rect 27304 18368 27310 18380
rect 30009 18377 30021 18380
rect 30055 18377 30067 18411
rect 30009 18371 30067 18377
rect 30834 18368 30840 18420
rect 30892 18408 30898 18420
rect 31021 18411 31079 18417
rect 31021 18408 31033 18411
rect 30892 18380 31033 18408
rect 30892 18368 30898 18380
rect 31021 18377 31033 18380
rect 31067 18377 31079 18411
rect 31021 18371 31079 18377
rect 31570 18368 31576 18420
rect 31628 18408 31634 18420
rect 31754 18408 31760 18420
rect 31628 18380 31760 18408
rect 31628 18368 31634 18380
rect 31754 18368 31760 18380
rect 31812 18408 31818 18420
rect 33781 18411 33839 18417
rect 33781 18408 33793 18411
rect 31812 18380 33793 18408
rect 31812 18368 31818 18380
rect 33781 18377 33793 18380
rect 33827 18408 33839 18411
rect 34422 18408 34428 18420
rect 33827 18380 34428 18408
rect 33827 18377 33839 18380
rect 33781 18371 33839 18377
rect 34422 18368 34428 18380
rect 34480 18368 34486 18420
rect 36170 18368 36176 18420
rect 36228 18408 36234 18420
rect 36630 18408 36636 18420
rect 36228 18380 36636 18408
rect 36228 18368 36234 18380
rect 36630 18368 36636 18380
rect 36688 18368 36694 18420
rect 36722 18368 36728 18420
rect 36780 18408 36786 18420
rect 36817 18411 36875 18417
rect 36817 18408 36829 18411
rect 36780 18380 36829 18408
rect 36780 18368 36786 18380
rect 36817 18377 36829 18380
rect 36863 18408 36875 18411
rect 38654 18408 38660 18420
rect 36863 18380 38660 18408
rect 36863 18377 36875 18380
rect 36817 18371 36875 18377
rect 38654 18368 38660 18380
rect 38712 18368 38718 18420
rect 38930 18368 38936 18420
rect 38988 18408 38994 18420
rect 40586 18408 40592 18420
rect 38988 18380 40172 18408
rect 38988 18368 38994 18380
rect 40144 18352 40172 18380
rect 40236 18380 40592 18408
rect 26418 18300 26424 18352
rect 26476 18340 26482 18352
rect 26476 18312 27922 18340
rect 26476 18300 26482 18312
rect 28810 18300 28816 18352
rect 28868 18340 28874 18352
rect 33318 18340 33324 18352
rect 28868 18312 33324 18340
rect 28868 18300 28874 18312
rect 33318 18300 33324 18312
rect 33376 18300 33382 18352
rect 33594 18300 33600 18352
rect 33652 18340 33658 18352
rect 33873 18343 33931 18349
rect 33873 18340 33885 18343
rect 33652 18312 33885 18340
rect 33652 18300 33658 18312
rect 33873 18309 33885 18312
rect 33919 18309 33931 18343
rect 34330 18340 34336 18352
rect 33873 18303 33931 18309
rect 34072 18312 34336 18340
rect 26605 18275 26663 18281
rect 26605 18272 26617 18275
rect 25271 18244 26188 18272
rect 26344 18244 26617 18272
rect 25271 18241 25283 18244
rect 25225 18235 25283 18241
rect 26160 18216 26188 18244
rect 26605 18241 26617 18244
rect 26651 18272 26663 18275
rect 27062 18272 27068 18284
rect 26651 18244 27068 18272
rect 26651 18241 26663 18244
rect 26605 18235 26663 18241
rect 27062 18232 27068 18244
rect 27120 18232 27126 18284
rect 27154 18232 27160 18284
rect 27212 18232 27218 18284
rect 28718 18232 28724 18284
rect 28776 18272 28782 18284
rect 29365 18275 29423 18281
rect 29365 18272 29377 18275
rect 28776 18244 29377 18272
rect 28776 18232 28782 18244
rect 17552 18176 19564 18204
rect 17552 18164 17558 18176
rect 22830 18164 22836 18216
rect 22888 18164 22894 18216
rect 24578 18164 24584 18216
rect 24636 18164 24642 18216
rect 25961 18207 26019 18213
rect 25961 18204 25973 18207
rect 24964 18176 25973 18204
rect 14700 18108 14964 18136
rect 16132 18108 19748 18136
rect 14700 18096 14706 18108
rect 14274 18068 14280 18080
rect 12636 18040 14280 18068
rect 11885 18031 11943 18037
rect 14274 18028 14280 18040
rect 14332 18028 14338 18080
rect 14826 18028 14832 18080
rect 14884 18028 14890 18080
rect 14936 18068 14964 18108
rect 16209 18071 16267 18077
rect 16209 18068 16221 18071
rect 14936 18040 16221 18068
rect 16209 18037 16221 18040
rect 16255 18037 16267 18071
rect 16209 18031 16267 18037
rect 16390 18028 16396 18080
rect 16448 18068 16454 18080
rect 17954 18068 17960 18080
rect 16448 18040 17960 18068
rect 16448 18028 16454 18040
rect 17954 18028 17960 18040
rect 18012 18028 18018 18080
rect 18049 18071 18107 18077
rect 18049 18037 18061 18071
rect 18095 18068 18107 18071
rect 19150 18068 19156 18080
rect 18095 18040 19156 18068
rect 18095 18037 18107 18040
rect 18049 18031 18107 18037
rect 19150 18028 19156 18040
rect 19208 18028 19214 18080
rect 19720 18068 19748 18108
rect 24964 18080 24992 18176
rect 25961 18173 25973 18176
rect 26007 18173 26019 18207
rect 25961 18167 26019 18173
rect 26142 18164 26148 18216
rect 26200 18164 26206 18216
rect 27433 18207 27491 18213
rect 27433 18173 27445 18207
rect 27479 18204 27491 18207
rect 27522 18204 27528 18216
rect 27479 18176 27528 18204
rect 27479 18173 27491 18176
rect 27433 18167 27491 18173
rect 27522 18164 27528 18176
rect 27580 18164 27586 18216
rect 25038 18096 25044 18148
rect 25096 18136 25102 18148
rect 26602 18136 26608 18148
rect 25096 18108 26608 18136
rect 25096 18096 25102 18108
rect 26602 18096 26608 18108
rect 26660 18096 26666 18148
rect 20898 18068 20904 18080
rect 19720 18040 20904 18068
rect 20898 18028 20904 18040
rect 20956 18028 20962 18080
rect 21361 18071 21419 18077
rect 21361 18037 21373 18071
rect 21407 18068 21419 18071
rect 21450 18068 21456 18080
rect 21407 18040 21456 18068
rect 21407 18037 21419 18040
rect 21361 18031 21419 18037
rect 21450 18028 21456 18040
rect 21508 18028 21514 18080
rect 24946 18028 24952 18080
rect 25004 18028 25010 18080
rect 25958 18028 25964 18080
rect 26016 18068 26022 18080
rect 28920 18077 28948 18244
rect 29365 18241 29377 18244
rect 29411 18241 29423 18275
rect 29365 18235 29423 18241
rect 30558 18232 30564 18284
rect 30616 18272 30622 18284
rect 30834 18272 30840 18284
rect 30616 18244 30840 18272
rect 30616 18232 30622 18244
rect 30834 18232 30840 18244
rect 30892 18232 30898 18284
rect 30926 18232 30932 18284
rect 30984 18272 30990 18284
rect 30984 18244 31524 18272
rect 30984 18232 30990 18244
rect 31205 18207 31263 18213
rect 31205 18173 31217 18207
rect 31251 18204 31263 18207
rect 31386 18204 31392 18216
rect 31251 18176 31392 18204
rect 31251 18173 31263 18176
rect 31205 18167 31263 18173
rect 31386 18164 31392 18176
rect 31444 18164 31450 18216
rect 31496 18204 31524 18244
rect 32214 18232 32220 18284
rect 32272 18232 32278 18284
rect 33045 18275 33103 18281
rect 33045 18241 33057 18275
rect 33091 18272 33103 18275
rect 34072 18272 34100 18312
rect 34330 18300 34336 18312
rect 34388 18300 34394 18352
rect 34698 18300 34704 18352
rect 34756 18300 34762 18352
rect 37826 18340 37832 18352
rect 35926 18312 37832 18340
rect 37826 18300 37832 18312
rect 37884 18300 37890 18352
rect 39114 18340 39120 18352
rect 38028 18312 39120 18340
rect 33091 18244 34100 18272
rect 34164 18244 34376 18272
rect 33091 18241 33103 18244
rect 33045 18235 33103 18241
rect 33336 18216 33364 18244
rect 32122 18204 32128 18216
rect 31496 18176 32128 18204
rect 32122 18164 32128 18176
rect 32180 18204 32186 18216
rect 32309 18207 32367 18213
rect 32309 18204 32321 18207
rect 32180 18176 32321 18204
rect 32180 18164 32186 18176
rect 32309 18173 32321 18176
rect 32355 18173 32367 18207
rect 32309 18167 32367 18173
rect 32674 18164 32680 18216
rect 32732 18204 32738 18216
rect 33137 18207 33195 18213
rect 33137 18204 33149 18207
rect 32732 18176 33149 18204
rect 32732 18164 32738 18176
rect 33137 18173 33149 18176
rect 33183 18173 33195 18207
rect 33137 18167 33195 18173
rect 30374 18096 30380 18148
rect 30432 18136 30438 18148
rect 33152 18136 33180 18167
rect 33226 18164 33232 18216
rect 33284 18164 33290 18216
rect 33318 18164 33324 18216
rect 33376 18164 33382 18216
rect 33410 18164 33416 18216
rect 33468 18204 33474 18216
rect 34054 18204 34060 18216
rect 33468 18176 34060 18204
rect 33468 18164 33474 18176
rect 34054 18164 34060 18176
rect 34112 18204 34118 18216
rect 34164 18213 34192 18244
rect 34149 18207 34207 18213
rect 34149 18204 34161 18207
rect 34112 18176 34161 18204
rect 34112 18164 34118 18176
rect 34149 18173 34161 18176
rect 34195 18173 34207 18207
rect 34149 18167 34207 18173
rect 34348 18136 34376 18244
rect 36722 18232 36728 18284
rect 36780 18232 36786 18284
rect 37274 18232 37280 18284
rect 37332 18272 37338 18284
rect 37461 18275 37519 18281
rect 37461 18272 37473 18275
rect 37332 18244 37473 18272
rect 37332 18232 37338 18244
rect 37461 18241 37473 18244
rect 37507 18241 37519 18275
rect 37461 18235 37519 18241
rect 34422 18164 34428 18216
rect 34480 18164 34486 18216
rect 38028 18204 38056 18312
rect 39114 18300 39120 18312
rect 39172 18300 39178 18352
rect 40126 18300 40132 18352
rect 40184 18300 40190 18352
rect 39942 18232 39948 18284
rect 40000 18232 40006 18284
rect 40236 18272 40264 18380
rect 40586 18368 40592 18380
rect 40644 18368 40650 18420
rect 41156 18380 41368 18408
rect 40052 18244 40264 18272
rect 34532 18176 38056 18204
rect 34532 18136 34560 18176
rect 38286 18164 38292 18216
rect 38344 18204 38350 18216
rect 38565 18207 38623 18213
rect 38565 18204 38577 18207
rect 38344 18176 38577 18204
rect 38344 18164 38350 18176
rect 38565 18173 38577 18176
rect 38611 18173 38623 18207
rect 38565 18167 38623 18173
rect 38841 18207 38899 18213
rect 38841 18173 38853 18207
rect 38887 18204 38899 18207
rect 40052 18204 40080 18244
rect 40310 18232 40316 18284
rect 40368 18232 40374 18284
rect 40586 18232 40592 18284
rect 40644 18272 40650 18284
rect 40644 18244 40908 18272
rect 40644 18232 40650 18244
rect 38887 18176 40080 18204
rect 40328 18204 40356 18232
rect 40770 18204 40776 18216
rect 40328 18176 40776 18204
rect 38887 18173 38899 18176
rect 38841 18167 38899 18173
rect 30432 18108 33088 18136
rect 33152 18108 34192 18136
rect 34348 18108 34560 18136
rect 30432 18096 30438 18108
rect 28905 18071 28963 18077
rect 28905 18068 28917 18071
rect 26016 18040 28917 18068
rect 26016 18028 26022 18040
rect 28905 18037 28917 18040
rect 28951 18037 28963 18071
rect 28905 18031 28963 18037
rect 30558 18028 30564 18080
rect 30616 18028 30622 18080
rect 30742 18028 30748 18080
rect 30800 18068 30806 18080
rect 31573 18071 31631 18077
rect 31573 18068 31585 18071
rect 30800 18040 31585 18068
rect 30800 18028 30806 18040
rect 31573 18037 31585 18040
rect 31619 18037 31631 18071
rect 31573 18031 31631 18037
rect 31662 18028 31668 18080
rect 31720 18068 31726 18080
rect 31757 18071 31815 18077
rect 31757 18068 31769 18071
rect 31720 18040 31769 18068
rect 31720 18028 31726 18040
rect 31757 18037 31769 18040
rect 31803 18037 31815 18071
rect 31757 18031 31815 18037
rect 32674 18028 32680 18080
rect 32732 18028 32738 18080
rect 33060 18068 33088 18108
rect 33962 18068 33968 18080
rect 33060 18040 33968 18068
rect 33962 18028 33968 18040
rect 34020 18028 34026 18080
rect 34164 18068 34192 18108
rect 36170 18096 36176 18148
rect 36228 18136 36234 18148
rect 36814 18136 36820 18148
rect 36228 18108 36820 18136
rect 36228 18096 36234 18108
rect 36814 18096 36820 18108
rect 36872 18096 36878 18148
rect 35986 18068 35992 18080
rect 34164 18040 35992 18068
rect 35986 18028 35992 18040
rect 36044 18028 36050 18080
rect 37458 18028 37464 18080
rect 37516 18068 37522 18080
rect 38105 18071 38163 18077
rect 38105 18068 38117 18071
rect 37516 18040 38117 18068
rect 37516 18028 37522 18040
rect 38105 18037 38117 18040
rect 38151 18037 38163 18071
rect 38580 18068 38608 18167
rect 40770 18164 40776 18176
rect 40828 18164 40834 18216
rect 40880 18204 40908 18244
rect 41156 18204 41184 18380
rect 41230 18300 41236 18352
rect 41288 18300 41294 18352
rect 41340 18340 41368 18380
rect 42794 18368 42800 18420
rect 42852 18408 42858 18420
rect 44910 18408 44916 18420
rect 42852 18380 44916 18408
rect 42852 18368 42858 18380
rect 44910 18368 44916 18380
rect 44968 18408 44974 18420
rect 47213 18411 47271 18417
rect 47213 18408 47225 18411
rect 44968 18380 47225 18408
rect 44968 18368 44974 18380
rect 47213 18377 47225 18380
rect 47259 18377 47271 18411
rect 47213 18371 47271 18377
rect 49234 18368 49240 18420
rect 49292 18368 49298 18420
rect 42150 18340 42156 18352
rect 41340 18312 42156 18340
rect 42150 18300 42156 18312
rect 42208 18300 42214 18352
rect 42702 18300 42708 18352
rect 42760 18340 42766 18352
rect 46474 18340 46480 18352
rect 42760 18312 46480 18340
rect 42760 18300 42766 18312
rect 46474 18300 46480 18312
rect 46532 18300 46538 18352
rect 46934 18300 46940 18352
rect 46992 18340 46998 18352
rect 47854 18340 47860 18352
rect 46992 18312 47860 18340
rect 46992 18300 46998 18312
rect 47854 18300 47860 18312
rect 47912 18300 47918 18352
rect 41325 18275 41383 18281
rect 41325 18241 41337 18275
rect 41371 18272 41383 18275
rect 41371 18244 41552 18272
rect 41371 18241 41383 18244
rect 41325 18235 41383 18241
rect 41524 18216 41552 18244
rect 42610 18232 42616 18284
rect 42668 18232 42674 18284
rect 43714 18232 43720 18284
rect 43772 18232 43778 18284
rect 44358 18232 44364 18284
rect 44416 18232 44422 18284
rect 44542 18232 44548 18284
rect 44600 18272 44606 18284
rect 44821 18275 44879 18281
rect 44821 18272 44833 18275
rect 44600 18244 44833 18272
rect 44600 18232 44606 18244
rect 44821 18241 44833 18244
rect 44867 18241 44879 18275
rect 44821 18235 44879 18241
rect 45925 18275 45983 18281
rect 45925 18241 45937 18275
rect 45971 18272 45983 18275
rect 47026 18272 47032 18284
rect 45971 18244 47032 18272
rect 45971 18241 45983 18244
rect 45925 18235 45983 18241
rect 47026 18232 47032 18244
rect 47084 18232 47090 18284
rect 47118 18232 47124 18284
rect 47176 18272 47182 18284
rect 48041 18275 48099 18281
rect 48041 18272 48053 18275
rect 47176 18244 48053 18272
rect 47176 18232 47182 18244
rect 48041 18241 48053 18244
rect 48087 18241 48099 18275
rect 48041 18235 48099 18241
rect 49053 18275 49111 18281
rect 49053 18241 49065 18275
rect 49099 18272 49111 18275
rect 50062 18272 50068 18284
rect 49099 18244 50068 18272
rect 49099 18241 49111 18244
rect 49053 18235 49111 18241
rect 50062 18232 50068 18244
rect 50120 18232 50126 18284
rect 40880 18176 41184 18204
rect 41414 18164 41420 18216
rect 41472 18164 41478 18216
rect 41506 18164 41512 18216
rect 41564 18164 41570 18216
rect 41598 18164 41604 18216
rect 41656 18204 41662 18216
rect 42061 18207 42119 18213
rect 42061 18204 42073 18207
rect 41656 18176 42073 18204
rect 41656 18164 41662 18176
rect 42061 18173 42073 18176
rect 42107 18173 42119 18207
rect 46290 18204 46296 18216
rect 42061 18167 42119 18173
rect 42168 18176 46296 18204
rect 40310 18096 40316 18148
rect 40368 18136 40374 18148
rect 42168 18136 42196 18176
rect 46290 18164 46296 18176
rect 46348 18164 46354 18216
rect 47578 18164 47584 18216
rect 47636 18204 47642 18216
rect 47673 18207 47731 18213
rect 47673 18204 47685 18207
rect 47636 18176 47685 18204
rect 47636 18164 47642 18176
rect 47673 18173 47685 18176
rect 47719 18204 47731 18207
rect 47765 18207 47823 18213
rect 47765 18204 47777 18207
rect 47719 18176 47777 18204
rect 47719 18173 47731 18176
rect 47673 18167 47731 18173
rect 47765 18173 47777 18176
rect 47811 18204 47823 18207
rect 48866 18204 48872 18216
rect 47811 18176 48872 18204
rect 47811 18173 47823 18176
rect 47765 18167 47823 18173
rect 48866 18164 48872 18176
rect 48924 18164 48930 18216
rect 40368 18108 42196 18136
rect 40368 18096 40374 18108
rect 43990 18096 43996 18148
rect 44048 18136 44054 18148
rect 46569 18139 46627 18145
rect 46569 18136 46581 18139
rect 44048 18108 46581 18136
rect 44048 18096 44054 18108
rect 46569 18105 46581 18108
rect 46615 18105 46627 18139
rect 46569 18099 46627 18105
rect 46937 18139 46995 18145
rect 46937 18105 46949 18139
rect 46983 18136 46995 18139
rect 47118 18136 47124 18148
rect 46983 18108 47124 18136
rect 46983 18105 46995 18108
rect 46937 18099 46995 18105
rect 47118 18096 47124 18108
rect 47176 18096 47182 18148
rect 40034 18068 40040 18080
rect 38580 18040 40040 18068
rect 38105 18031 38163 18037
rect 40034 18028 40040 18040
rect 40092 18028 40098 18080
rect 40126 18028 40132 18080
rect 40184 18068 40190 18080
rect 40865 18071 40923 18077
rect 40865 18068 40877 18071
rect 40184 18040 40877 18068
rect 40184 18028 40190 18040
rect 40865 18037 40877 18040
rect 40911 18037 40923 18071
rect 40865 18031 40923 18037
rect 40954 18028 40960 18080
rect 41012 18068 41018 18080
rect 41138 18068 41144 18080
rect 41012 18040 41144 18068
rect 41012 18028 41018 18040
rect 41138 18028 41144 18040
rect 41196 18028 41202 18080
rect 41969 18071 42027 18077
rect 41969 18037 41981 18071
rect 42015 18068 42027 18071
rect 42334 18068 42340 18080
rect 42015 18040 42340 18068
rect 42015 18037 42027 18040
rect 41969 18031 42027 18037
rect 42334 18028 42340 18040
rect 42392 18028 42398 18080
rect 42794 18028 42800 18080
rect 42852 18068 42858 18080
rect 43257 18071 43315 18077
rect 43257 18068 43269 18071
rect 42852 18040 43269 18068
rect 42852 18028 42858 18040
rect 43257 18037 43269 18040
rect 43303 18037 43315 18071
rect 43257 18031 43315 18037
rect 45370 18028 45376 18080
rect 45428 18068 45434 18080
rect 45465 18071 45523 18077
rect 45465 18068 45477 18071
rect 45428 18040 45477 18068
rect 45428 18028 45434 18040
rect 45465 18037 45477 18040
rect 45511 18037 45523 18071
rect 45465 18031 45523 18037
rect 46658 18028 46664 18080
rect 46716 18068 46722 18080
rect 47029 18071 47087 18077
rect 47029 18068 47041 18071
rect 46716 18040 47041 18068
rect 46716 18028 46722 18040
rect 47029 18037 47041 18040
rect 47075 18037 47087 18071
rect 47029 18031 47087 18037
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 2866 17824 2872 17876
rect 2924 17864 2930 17876
rect 3513 17867 3571 17873
rect 3513 17864 3525 17867
rect 2924 17836 3525 17864
rect 2924 17824 2930 17836
rect 3513 17833 3525 17836
rect 3559 17833 3571 17867
rect 3513 17827 3571 17833
rect 6365 17867 6423 17873
rect 6365 17833 6377 17867
rect 6411 17864 6423 17867
rect 6638 17864 6644 17876
rect 6411 17836 6644 17864
rect 6411 17833 6423 17836
rect 6365 17827 6423 17833
rect 6638 17824 6644 17836
rect 6696 17824 6702 17876
rect 8573 17867 8631 17873
rect 8573 17833 8585 17867
rect 8619 17864 8631 17867
rect 9490 17864 9496 17876
rect 8619 17836 9496 17864
rect 8619 17833 8631 17836
rect 8573 17827 8631 17833
rect 9490 17824 9496 17836
rect 9548 17824 9554 17876
rect 14734 17864 14740 17876
rect 11072 17836 14740 17864
rect 10962 17796 10968 17808
rect 7392 17768 10968 17796
rect 1210 17688 1216 17740
rect 1268 17728 1274 17740
rect 2041 17731 2099 17737
rect 2041 17728 2053 17731
rect 1268 17700 2053 17728
rect 1268 17688 1274 17700
rect 2041 17697 2053 17700
rect 2087 17697 2099 17731
rect 2041 17691 2099 17697
rect 3973 17731 4031 17737
rect 3973 17697 3985 17731
rect 4019 17728 4031 17731
rect 4154 17728 4160 17740
rect 4019 17700 4160 17728
rect 4019 17697 4031 17700
rect 3973 17691 4031 17697
rect 4154 17688 4160 17700
rect 4212 17688 4218 17740
rect 5261 17731 5319 17737
rect 5261 17697 5273 17731
rect 5307 17728 5319 17731
rect 7392 17728 7420 17768
rect 10962 17756 10968 17768
rect 11020 17756 11026 17808
rect 5307 17700 7420 17728
rect 7469 17731 7527 17737
rect 5307 17697 5319 17700
rect 5261 17691 5319 17697
rect 7469 17697 7481 17731
rect 7515 17728 7527 17731
rect 9766 17728 9772 17740
rect 7515 17700 9772 17728
rect 7515 17697 7527 17700
rect 7469 17691 7527 17697
rect 9766 17688 9772 17700
rect 9824 17688 9830 17740
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17629 1823 17663
rect 1765 17623 1823 17629
rect 1780 17592 1808 17623
rect 3418 17620 3424 17672
rect 3476 17620 3482 17672
rect 4614 17620 4620 17672
rect 4672 17620 4678 17672
rect 5718 17620 5724 17672
rect 5776 17620 5782 17672
rect 6822 17620 6828 17672
rect 6880 17620 6886 17672
rect 7929 17663 7987 17669
rect 7929 17629 7941 17663
rect 7975 17660 7987 17663
rect 9950 17660 9956 17672
rect 7975 17632 9956 17660
rect 7975 17629 7987 17632
rect 7929 17623 7987 17629
rect 9950 17620 9956 17632
rect 10008 17620 10014 17672
rect 10045 17663 10103 17669
rect 10045 17629 10057 17663
rect 10091 17660 10103 17663
rect 11072 17660 11100 17836
rect 14734 17824 14740 17836
rect 14792 17824 14798 17876
rect 14918 17824 14924 17876
rect 14976 17864 14982 17876
rect 19610 17864 19616 17876
rect 14976 17836 19616 17864
rect 14976 17824 14982 17836
rect 19610 17824 19616 17836
rect 19668 17824 19674 17876
rect 20514 17867 20572 17873
rect 20514 17864 20526 17867
rect 19720 17836 20526 17864
rect 13262 17796 13268 17808
rect 12728 17768 13268 17796
rect 11146 17688 11152 17740
rect 11204 17728 11210 17740
rect 11974 17728 11980 17740
rect 11204 17700 11980 17728
rect 11204 17688 11210 17700
rect 11974 17688 11980 17700
rect 12032 17688 12038 17740
rect 12158 17688 12164 17740
rect 12216 17728 12222 17740
rect 12728 17728 12756 17768
rect 13262 17756 13268 17768
rect 13320 17756 13326 17808
rect 13446 17756 13452 17808
rect 13504 17796 13510 17808
rect 19720 17796 19748 17836
rect 20514 17833 20526 17836
rect 20560 17833 20572 17867
rect 20514 17827 20572 17833
rect 20898 17824 20904 17876
rect 20956 17864 20962 17876
rect 22465 17867 22523 17873
rect 22465 17864 22477 17867
rect 20956 17836 22477 17864
rect 20956 17824 20962 17836
rect 22465 17833 22477 17836
rect 22511 17833 22523 17867
rect 22465 17827 22523 17833
rect 24210 17824 24216 17876
rect 24268 17864 24274 17876
rect 24268 17836 26924 17864
rect 24268 17824 24274 17836
rect 13504 17768 14412 17796
rect 13504 17756 13510 17768
rect 12216 17700 12756 17728
rect 12216 17688 12222 17700
rect 12802 17688 12808 17740
rect 12860 17728 12866 17740
rect 13725 17731 13783 17737
rect 13725 17728 13737 17731
rect 12860 17700 13737 17728
rect 12860 17688 12866 17700
rect 13725 17697 13737 17700
rect 13771 17697 13783 17731
rect 14384 17728 14412 17768
rect 16868 17768 19748 17796
rect 16868 17728 16896 17768
rect 22646 17756 22652 17808
rect 22704 17796 22710 17808
rect 22704 17768 24624 17796
rect 22704 17756 22710 17768
rect 14384 17700 16896 17728
rect 13725 17691 13783 17697
rect 17034 17688 17040 17740
rect 17092 17728 17098 17740
rect 17865 17731 17923 17737
rect 17865 17728 17877 17731
rect 17092 17700 17877 17728
rect 17092 17688 17098 17700
rect 17865 17697 17877 17700
rect 17911 17697 17923 17731
rect 17865 17691 17923 17697
rect 17954 17688 17960 17740
rect 18012 17728 18018 17740
rect 18785 17731 18843 17737
rect 18785 17728 18797 17731
rect 18012 17700 18797 17728
rect 18012 17688 18018 17700
rect 18785 17697 18797 17700
rect 18831 17697 18843 17731
rect 18785 17691 18843 17697
rect 19242 17688 19248 17740
rect 19300 17728 19306 17740
rect 19300 17700 20300 17728
rect 19300 17688 19306 17700
rect 10091 17632 11100 17660
rect 10091 17629 10103 17632
rect 10045 17623 10103 17629
rect 12526 17620 12532 17672
rect 12584 17620 12590 17672
rect 12820 17632 13676 17660
rect 1780 17564 9076 17592
rect 8938 17484 8944 17536
rect 8996 17484 9002 17536
rect 9048 17524 9076 17564
rect 9214 17552 9220 17604
rect 9272 17592 9278 17604
rect 9401 17595 9459 17601
rect 9401 17592 9413 17595
rect 9272 17564 9413 17592
rect 9272 17552 9278 17564
rect 9401 17561 9413 17564
rect 9447 17561 9459 17595
rect 9401 17555 9459 17561
rect 9582 17552 9588 17604
rect 9640 17592 9646 17604
rect 9640 17564 10824 17592
rect 9640 17552 9646 17564
rect 9493 17527 9551 17533
rect 9493 17524 9505 17527
rect 9048 17496 9505 17524
rect 9493 17493 9505 17496
rect 9539 17493 9551 17527
rect 9493 17487 9551 17493
rect 10502 17484 10508 17536
rect 10560 17524 10566 17536
rect 10689 17527 10747 17533
rect 10689 17524 10701 17527
rect 10560 17496 10701 17524
rect 10560 17484 10566 17496
rect 10689 17493 10701 17496
rect 10735 17493 10747 17527
rect 10796 17524 10824 17564
rect 10870 17552 10876 17604
rect 10928 17592 10934 17604
rect 11425 17595 11483 17601
rect 11425 17592 11437 17595
rect 10928 17564 11437 17592
rect 10928 17552 10934 17564
rect 11425 17561 11437 17564
rect 11471 17561 11483 17595
rect 11425 17555 11483 17561
rect 12820 17524 12848 17632
rect 13538 17552 13544 17604
rect 13596 17552 13602 17604
rect 13648 17592 13676 17632
rect 14274 17620 14280 17672
rect 14332 17620 14338 17672
rect 17773 17663 17831 17669
rect 15856 17632 17724 17660
rect 14553 17595 14611 17601
rect 14553 17592 14565 17595
rect 13648 17564 14565 17592
rect 14553 17561 14565 17564
rect 14599 17561 14611 17595
rect 14553 17555 14611 17561
rect 15010 17552 15016 17604
rect 15068 17552 15074 17604
rect 10796 17496 12848 17524
rect 12897 17527 12955 17533
rect 10689 17487 10747 17493
rect 12897 17493 12909 17527
rect 12943 17524 12955 17527
rect 13354 17524 13360 17536
rect 12943 17496 13360 17524
rect 12943 17493 12955 17496
rect 12897 17487 12955 17493
rect 13354 17484 13360 17496
rect 13412 17484 13418 17536
rect 14734 17484 14740 17536
rect 14792 17524 14798 17536
rect 15856 17524 15884 17632
rect 16577 17595 16635 17601
rect 16577 17561 16589 17595
rect 16623 17592 16635 17595
rect 17126 17592 17132 17604
rect 16623 17564 17132 17592
rect 16623 17561 16635 17564
rect 16577 17555 16635 17561
rect 17126 17552 17132 17564
rect 17184 17552 17190 17604
rect 17696 17592 17724 17632
rect 17773 17629 17785 17663
rect 17819 17660 17831 17663
rect 19426 17660 19432 17672
rect 17819 17632 19432 17660
rect 17819 17629 17831 17632
rect 17773 17623 17831 17629
rect 19426 17620 19432 17632
rect 19484 17620 19490 17672
rect 20272 17669 20300 17700
rect 22002 17688 22008 17740
rect 22060 17728 22066 17740
rect 24596 17737 24624 17768
rect 23017 17731 23075 17737
rect 23017 17728 23029 17731
rect 22060 17700 23029 17728
rect 22060 17688 22066 17700
rect 23017 17697 23029 17700
rect 23063 17697 23075 17731
rect 23017 17691 23075 17697
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17697 24639 17731
rect 24581 17691 24639 17697
rect 25685 17731 25743 17737
rect 25685 17697 25697 17731
rect 25731 17728 25743 17731
rect 26234 17728 26240 17740
rect 25731 17700 26240 17728
rect 25731 17697 25743 17700
rect 25685 17691 25743 17697
rect 26234 17688 26240 17700
rect 26292 17688 26298 17740
rect 26896 17728 26924 17836
rect 26970 17824 26976 17876
rect 27028 17864 27034 17876
rect 27430 17864 27436 17876
rect 27028 17836 27436 17864
rect 27028 17824 27034 17836
rect 27430 17824 27436 17836
rect 27488 17824 27494 17876
rect 27614 17824 27620 17876
rect 27672 17824 27678 17876
rect 28074 17824 28080 17876
rect 28132 17864 28138 17876
rect 30190 17864 30196 17876
rect 28132 17836 30196 17864
rect 28132 17824 28138 17836
rect 30190 17824 30196 17836
rect 30248 17824 30254 17876
rect 30650 17824 30656 17876
rect 30708 17864 30714 17876
rect 33597 17867 33655 17873
rect 30708 17836 33548 17864
rect 30708 17824 30714 17836
rect 27246 17756 27252 17808
rect 27304 17796 27310 17808
rect 27304 17768 31340 17796
rect 27304 17756 27310 17768
rect 28074 17728 28080 17740
rect 26896 17700 28080 17728
rect 28074 17688 28080 17700
rect 28132 17688 28138 17740
rect 28626 17688 28632 17740
rect 28684 17728 28690 17740
rect 28997 17731 29055 17737
rect 28997 17728 29009 17731
rect 28684 17700 29009 17728
rect 28684 17688 28690 17700
rect 28997 17697 29009 17700
rect 29043 17697 29055 17731
rect 28997 17691 29055 17697
rect 29454 17688 29460 17740
rect 29512 17728 29518 17740
rect 31312 17737 31340 17768
rect 32582 17756 32588 17808
rect 32640 17796 32646 17808
rect 33045 17799 33103 17805
rect 33045 17796 33057 17799
rect 32640 17768 33057 17796
rect 32640 17756 32646 17768
rect 33045 17765 33057 17768
rect 33091 17796 33103 17799
rect 33410 17796 33416 17808
rect 33091 17768 33416 17796
rect 33091 17765 33103 17768
rect 33045 17759 33103 17765
rect 33410 17756 33416 17768
rect 33468 17756 33474 17808
rect 33520 17796 33548 17836
rect 33597 17833 33609 17867
rect 33643 17864 33655 17867
rect 34146 17864 34152 17876
rect 33643 17836 34152 17864
rect 33643 17833 33655 17836
rect 33597 17827 33655 17833
rect 34146 17824 34152 17836
rect 34204 17824 34210 17876
rect 34885 17867 34943 17873
rect 34885 17833 34897 17867
rect 34931 17864 34943 17867
rect 34974 17864 34980 17876
rect 34931 17836 34980 17864
rect 34931 17833 34943 17836
rect 34885 17827 34943 17833
rect 34974 17824 34980 17836
rect 35032 17824 35038 17876
rect 35986 17824 35992 17876
rect 36044 17824 36050 17876
rect 36712 17867 36770 17873
rect 36712 17833 36724 17867
rect 36758 17864 36770 17867
rect 36758 17836 37872 17864
rect 36758 17833 36770 17836
rect 36712 17827 36770 17833
rect 35894 17796 35900 17808
rect 33520 17768 35900 17796
rect 35894 17756 35900 17768
rect 35952 17756 35958 17808
rect 36173 17799 36231 17805
rect 36173 17765 36185 17799
rect 36219 17796 36231 17799
rect 36446 17796 36452 17808
rect 36219 17768 36452 17796
rect 36219 17765 36231 17768
rect 36173 17759 36231 17765
rect 36446 17756 36452 17768
rect 36504 17756 36510 17808
rect 37844 17796 37872 17836
rect 37918 17824 37924 17876
rect 37976 17864 37982 17876
rect 44269 17867 44327 17873
rect 44269 17864 44281 17867
rect 37976 17836 44281 17864
rect 37976 17824 37982 17836
rect 44269 17833 44281 17836
rect 44315 17864 44327 17867
rect 44450 17864 44456 17876
rect 44315 17836 44456 17864
rect 44315 17833 44327 17836
rect 44269 17827 44327 17833
rect 44450 17824 44456 17836
rect 44508 17824 44514 17876
rect 46474 17824 46480 17876
rect 46532 17864 46538 17876
rect 48041 17867 48099 17873
rect 48041 17864 48053 17867
rect 46532 17836 48053 17864
rect 46532 17824 46538 17836
rect 48041 17833 48053 17836
rect 48087 17833 48099 17867
rect 48041 17827 48099 17833
rect 38470 17796 38476 17808
rect 37844 17768 38476 17796
rect 38470 17756 38476 17768
rect 38528 17756 38534 17808
rect 38562 17756 38568 17808
rect 38620 17796 38626 17808
rect 39666 17796 39672 17808
rect 38620 17768 39672 17796
rect 38620 17756 38626 17768
rect 39666 17756 39672 17768
rect 39724 17756 39730 17808
rect 41506 17756 41512 17808
rect 41564 17796 41570 17808
rect 41785 17799 41843 17805
rect 41785 17796 41797 17799
rect 41564 17768 41797 17796
rect 41564 17756 41570 17768
rect 41785 17765 41797 17768
rect 41831 17796 41843 17799
rect 46014 17796 46020 17808
rect 41831 17768 46020 17796
rect 41831 17765 41843 17768
rect 41785 17759 41843 17765
rect 46014 17756 46020 17768
rect 46072 17756 46078 17808
rect 30285 17731 30343 17737
rect 30285 17728 30297 17731
rect 29512 17700 30297 17728
rect 29512 17688 29518 17700
rect 30285 17697 30297 17700
rect 30331 17697 30343 17731
rect 30285 17691 30343 17697
rect 31297 17731 31355 17737
rect 31297 17697 31309 17731
rect 31343 17728 31355 17731
rect 32306 17728 32312 17740
rect 31343 17700 32312 17728
rect 31343 17697 31355 17700
rect 31297 17691 31355 17697
rect 32306 17688 32312 17700
rect 32364 17688 32370 17740
rect 33594 17688 33600 17740
rect 33652 17728 33658 17740
rect 34057 17731 34115 17737
rect 34057 17728 34069 17731
rect 33652 17700 34069 17728
rect 33652 17688 33658 17700
rect 34057 17697 34069 17700
rect 34103 17697 34115 17731
rect 34057 17691 34115 17697
rect 34146 17688 34152 17740
rect 34204 17688 34210 17740
rect 34514 17728 34520 17740
rect 34256 17700 34520 17728
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17660 19763 17663
rect 20257 17663 20315 17669
rect 19751 17648 19840 17660
rect 19751 17632 19800 17648
rect 19751 17629 19763 17632
rect 19705 17623 19763 17629
rect 17696 17564 18276 17592
rect 14792 17496 15884 17524
rect 14792 17484 14798 17496
rect 15930 17484 15936 17536
rect 15988 17524 15994 17536
rect 16025 17527 16083 17533
rect 16025 17524 16037 17527
rect 15988 17496 16037 17524
rect 15988 17484 15994 17496
rect 16025 17493 16037 17496
rect 16071 17493 16083 17527
rect 16025 17487 16083 17493
rect 16666 17484 16672 17536
rect 16724 17484 16730 17536
rect 17310 17484 17316 17536
rect 17368 17484 17374 17536
rect 17678 17484 17684 17536
rect 17736 17484 17742 17536
rect 18248 17524 18276 17564
rect 18322 17552 18328 17604
rect 18380 17592 18386 17604
rect 18601 17595 18659 17601
rect 18601 17592 18613 17595
rect 18380 17564 18613 17592
rect 18380 17552 18386 17564
rect 18601 17561 18613 17564
rect 18647 17561 18659 17595
rect 18601 17555 18659 17561
rect 18782 17552 18788 17604
rect 18840 17592 18846 17604
rect 19150 17592 19156 17604
rect 18840 17564 19156 17592
rect 18840 17552 18846 17564
rect 19150 17552 19156 17564
rect 19208 17592 19214 17604
rect 19521 17595 19579 17601
rect 19794 17596 19800 17632
rect 19852 17596 19858 17648
rect 20257 17629 20269 17663
rect 20303 17629 20315 17663
rect 20257 17623 20315 17629
rect 19521 17592 19533 17595
rect 19208 17564 19533 17592
rect 19208 17552 19214 17564
rect 19521 17561 19533 17564
rect 19567 17561 19579 17595
rect 20272 17592 20300 17623
rect 22830 17620 22836 17672
rect 22888 17660 22894 17672
rect 23106 17660 23112 17672
rect 22888 17632 23112 17660
rect 22888 17620 22894 17632
rect 23106 17620 23112 17632
rect 23164 17660 23170 17672
rect 25409 17663 25467 17669
rect 25409 17660 25421 17663
rect 23164 17632 25421 17660
rect 23164 17620 23170 17632
rect 25409 17629 25421 17632
rect 25455 17629 25467 17663
rect 25409 17623 25467 17629
rect 27801 17663 27859 17669
rect 27801 17629 27813 17663
rect 27847 17629 27859 17663
rect 27801 17623 27859 17629
rect 20806 17592 20812 17604
rect 20272 17564 20812 17592
rect 19521 17555 19579 17561
rect 20806 17552 20812 17564
rect 20864 17552 20870 17604
rect 21266 17552 21272 17604
rect 21324 17552 21330 17604
rect 22925 17595 22983 17601
rect 22925 17561 22937 17595
rect 22971 17592 22983 17595
rect 23658 17592 23664 17604
rect 22971 17564 23664 17592
rect 22971 17561 22983 17564
rect 22925 17555 22983 17561
rect 23658 17552 23664 17564
rect 23716 17552 23722 17604
rect 23750 17552 23756 17604
rect 23808 17552 23814 17604
rect 24762 17552 24768 17604
rect 24820 17592 24826 17604
rect 24820 17564 26096 17592
rect 24820 17552 24826 17564
rect 19794 17524 19800 17536
rect 18248 17496 19800 17524
rect 19794 17484 19800 17496
rect 19852 17484 19858 17536
rect 21358 17484 21364 17536
rect 21416 17524 21422 17536
rect 21910 17524 21916 17536
rect 21416 17496 21916 17524
rect 21416 17484 21422 17496
rect 21910 17484 21916 17496
rect 21968 17524 21974 17536
rect 22005 17527 22063 17533
rect 22005 17524 22017 17527
rect 21968 17496 22017 17524
rect 21968 17484 21974 17496
rect 22005 17493 22017 17496
rect 22051 17493 22063 17527
rect 22005 17487 22063 17493
rect 22833 17527 22891 17533
rect 22833 17493 22845 17527
rect 22879 17524 22891 17527
rect 23474 17524 23480 17536
rect 22879 17496 23480 17524
rect 22879 17493 22891 17496
rect 22833 17487 22891 17493
rect 23474 17484 23480 17496
rect 23532 17484 23538 17536
rect 23842 17484 23848 17536
rect 23900 17484 23906 17536
rect 24118 17484 24124 17536
rect 24176 17524 24182 17536
rect 25041 17527 25099 17533
rect 25041 17524 25053 17527
rect 24176 17496 25053 17524
rect 24176 17484 24182 17496
rect 25041 17493 25053 17496
rect 25087 17493 25099 17527
rect 26068 17524 26096 17564
rect 26418 17552 26424 17604
rect 26476 17552 26482 17604
rect 27816 17592 27844 17623
rect 28350 17620 28356 17672
rect 28408 17660 28414 17672
rect 28813 17663 28871 17669
rect 28813 17660 28825 17663
rect 28408 17632 28825 17660
rect 28408 17620 28414 17632
rect 28813 17629 28825 17632
rect 28859 17660 28871 17663
rect 30929 17663 30987 17669
rect 30929 17660 30941 17663
rect 28859 17632 30941 17660
rect 28859 17629 28871 17632
rect 28813 17623 28871 17629
rect 30929 17629 30941 17632
rect 30975 17629 30987 17663
rect 30929 17623 30987 17629
rect 32582 17620 32588 17672
rect 32640 17660 32646 17672
rect 34256 17660 34284 17700
rect 34514 17688 34520 17700
rect 34572 17688 34578 17740
rect 34698 17688 34704 17740
rect 34756 17728 34762 17740
rect 35345 17731 35403 17737
rect 35345 17728 35357 17731
rect 34756 17700 35357 17728
rect 34756 17688 34762 17700
rect 35345 17697 35357 17700
rect 35391 17697 35403 17731
rect 35345 17691 35403 17697
rect 35526 17688 35532 17740
rect 35584 17688 35590 17740
rect 35802 17688 35808 17740
rect 35860 17728 35866 17740
rect 35986 17728 35992 17740
rect 35860 17700 35992 17728
rect 35860 17688 35866 17700
rect 35986 17688 35992 17700
rect 36044 17688 36050 17740
rect 38286 17728 38292 17740
rect 36464 17700 38292 17728
rect 32640 17632 34284 17660
rect 32640 17620 32646 17632
rect 34422 17620 34428 17672
rect 34480 17660 34486 17672
rect 36464 17669 36492 17700
rect 38286 17688 38292 17700
rect 38344 17688 38350 17740
rect 38378 17688 38384 17740
rect 38436 17728 38442 17740
rect 39301 17731 39359 17737
rect 38436 17700 39252 17728
rect 38436 17688 38442 17700
rect 36449 17663 36507 17669
rect 36449 17660 36461 17663
rect 34480 17632 36461 17660
rect 34480 17620 34486 17632
rect 36449 17629 36461 17632
rect 36495 17629 36507 17663
rect 38010 17660 38016 17672
rect 37858 17632 38016 17660
rect 36449 17623 36507 17629
rect 38010 17620 38016 17632
rect 38068 17620 38074 17672
rect 39224 17660 39252 17700
rect 39301 17697 39313 17731
rect 39347 17728 39359 17731
rect 39850 17728 39856 17740
rect 39347 17700 39856 17728
rect 39347 17697 39359 17700
rect 39301 17691 39359 17697
rect 39850 17688 39856 17700
rect 39908 17688 39914 17740
rect 40034 17688 40040 17740
rect 40092 17688 40098 17740
rect 40313 17731 40371 17737
rect 40313 17697 40325 17731
rect 40359 17728 40371 17731
rect 43990 17728 43996 17740
rect 40359 17700 43996 17728
rect 40359 17697 40371 17700
rect 40313 17691 40371 17697
rect 43990 17688 43996 17700
rect 44048 17688 44054 17740
rect 44450 17688 44456 17740
rect 44508 17688 44514 17740
rect 39224 17632 39620 17660
rect 27890 17592 27896 17604
rect 27816 17564 27896 17592
rect 27890 17552 27896 17564
rect 27948 17552 27954 17604
rect 28905 17595 28963 17601
rect 28905 17592 28917 17595
rect 28092 17564 28917 17592
rect 27062 17524 27068 17536
rect 26068 17496 27068 17524
rect 25041 17487 25099 17493
rect 27062 17484 27068 17496
rect 27120 17524 27126 17536
rect 27157 17527 27215 17533
rect 27157 17524 27169 17527
rect 27120 17496 27169 17524
rect 27120 17484 27126 17496
rect 27157 17493 27169 17496
rect 27203 17493 27215 17527
rect 27157 17487 27215 17493
rect 27430 17484 27436 17536
rect 27488 17524 27494 17536
rect 28092 17524 28120 17564
rect 28905 17561 28917 17564
rect 28951 17592 28963 17595
rect 31573 17595 31631 17601
rect 28951 17564 30880 17592
rect 28951 17561 28963 17564
rect 28905 17555 28963 17561
rect 27488 17496 28120 17524
rect 27488 17484 27494 17496
rect 28442 17484 28448 17536
rect 28500 17484 28506 17536
rect 28534 17484 28540 17536
rect 28592 17524 28598 17536
rect 28994 17524 29000 17536
rect 28592 17496 29000 17524
rect 28592 17484 28598 17496
rect 28994 17484 29000 17496
rect 29052 17484 29058 17536
rect 29730 17484 29736 17536
rect 29788 17484 29794 17536
rect 30098 17484 30104 17536
rect 30156 17484 30162 17536
rect 30190 17484 30196 17536
rect 30248 17484 30254 17536
rect 30852 17533 30880 17564
rect 31573 17561 31585 17595
rect 31619 17592 31631 17595
rect 35802 17592 35808 17604
rect 31619 17564 31754 17592
rect 31619 17561 31631 17564
rect 31573 17555 31631 17561
rect 30837 17527 30895 17533
rect 30837 17493 30849 17527
rect 30883 17524 30895 17527
rect 30926 17524 30932 17536
rect 30883 17496 30932 17524
rect 30883 17493 30895 17496
rect 30837 17487 30895 17493
rect 30926 17484 30932 17496
rect 30984 17484 30990 17536
rect 31726 17524 31754 17564
rect 32968 17564 35808 17592
rect 32968 17524 32996 17564
rect 35802 17552 35808 17564
rect 35860 17552 35866 17604
rect 36814 17592 36820 17604
rect 36096 17564 36820 17592
rect 31726 17496 32996 17524
rect 33965 17527 34023 17533
rect 33965 17493 33977 17527
rect 34011 17524 34023 17527
rect 34054 17524 34060 17536
rect 34011 17496 34060 17524
rect 34011 17493 34023 17496
rect 33965 17487 34023 17493
rect 34054 17484 34060 17496
rect 34112 17484 34118 17536
rect 35253 17527 35311 17533
rect 35253 17493 35265 17527
rect 35299 17524 35311 17527
rect 36096 17524 36124 17564
rect 36814 17552 36820 17564
rect 36872 17552 36878 17604
rect 39025 17595 39083 17601
rect 38028 17564 38700 17592
rect 35299 17496 36124 17524
rect 35299 17493 35311 17496
rect 35253 17487 35311 17493
rect 36170 17484 36176 17536
rect 36228 17524 36234 17536
rect 38028 17524 38056 17564
rect 36228 17496 38056 17524
rect 38197 17527 38255 17533
rect 36228 17484 36234 17496
rect 38197 17493 38209 17527
rect 38243 17524 38255 17527
rect 38470 17524 38476 17536
rect 38243 17496 38476 17524
rect 38243 17493 38255 17496
rect 38197 17487 38255 17493
rect 38470 17484 38476 17496
rect 38528 17484 38534 17536
rect 38672 17533 38700 17564
rect 39025 17561 39037 17595
rect 39071 17592 39083 17595
rect 39390 17592 39396 17604
rect 39071 17564 39396 17592
rect 39071 17561 39083 17564
rect 39025 17555 39083 17561
rect 39390 17552 39396 17564
rect 39448 17552 39454 17604
rect 38657 17527 38715 17533
rect 38657 17493 38669 17527
rect 38703 17493 38715 17527
rect 38657 17487 38715 17493
rect 39114 17484 39120 17536
rect 39172 17484 39178 17536
rect 39206 17484 39212 17536
rect 39264 17524 39270 17536
rect 39482 17524 39488 17536
rect 39264 17496 39488 17524
rect 39264 17484 39270 17496
rect 39482 17484 39488 17496
rect 39540 17484 39546 17536
rect 39592 17524 39620 17632
rect 42242 17620 42248 17672
rect 42300 17620 42306 17672
rect 43383 17663 43441 17669
rect 43383 17660 43395 17663
rect 42352 17632 43395 17660
rect 40770 17552 40776 17604
rect 40828 17552 40834 17604
rect 42352 17524 42380 17632
rect 43383 17629 43395 17632
rect 43429 17629 43441 17663
rect 43383 17623 43441 17629
rect 45189 17663 45247 17669
rect 45189 17629 45201 17663
rect 45235 17629 45247 17663
rect 45189 17623 45247 17629
rect 44726 17552 44732 17604
rect 44784 17592 44790 17604
rect 45204 17592 45232 17623
rect 46014 17620 46020 17672
rect 46072 17660 46078 17672
rect 46293 17663 46351 17669
rect 46293 17660 46305 17663
rect 46072 17632 46305 17660
rect 46072 17620 46078 17632
rect 46293 17629 46305 17632
rect 46339 17629 46351 17663
rect 46293 17623 46351 17629
rect 47397 17663 47455 17669
rect 47397 17629 47409 17663
rect 47443 17660 47455 17663
rect 48406 17660 48412 17672
rect 47443 17632 48412 17660
rect 47443 17629 47455 17632
rect 47397 17623 47455 17629
rect 48406 17620 48412 17632
rect 48464 17620 48470 17672
rect 48498 17620 48504 17672
rect 48556 17620 48562 17672
rect 44784 17564 45232 17592
rect 44784 17552 44790 17564
rect 47578 17552 47584 17604
rect 47636 17592 47642 17604
rect 49421 17595 49479 17601
rect 49421 17592 49433 17595
rect 47636 17564 49433 17592
rect 47636 17552 47642 17564
rect 49421 17561 49433 17564
rect 49467 17561 49479 17595
rect 49421 17555 49479 17561
rect 39592 17496 42380 17524
rect 42610 17484 42616 17536
rect 42668 17524 42674 17536
rect 42889 17527 42947 17533
rect 42889 17524 42901 17527
rect 42668 17496 42901 17524
rect 42668 17484 42674 17496
rect 42889 17493 42901 17496
rect 42935 17493 42947 17527
rect 42889 17487 42947 17493
rect 43346 17484 43352 17536
rect 43404 17524 43410 17536
rect 43993 17527 44051 17533
rect 43993 17524 44005 17527
rect 43404 17496 44005 17524
rect 43404 17484 43410 17496
rect 43993 17493 44005 17496
rect 44039 17493 44051 17527
rect 43993 17487 44051 17493
rect 45830 17484 45836 17536
rect 45888 17484 45894 17536
rect 45922 17484 45928 17536
rect 45980 17524 45986 17536
rect 46937 17527 46995 17533
rect 46937 17524 46949 17527
rect 45980 17496 46949 17524
rect 45980 17484 45986 17496
rect 46937 17493 46949 17496
rect 46983 17493 46995 17527
rect 46937 17487 46995 17493
rect 47118 17484 47124 17536
rect 47176 17524 47182 17536
rect 49145 17527 49203 17533
rect 49145 17524 49157 17527
rect 47176 17496 49157 17524
rect 47176 17484 47182 17496
rect 49145 17493 49157 17496
rect 49191 17493 49203 17527
rect 49145 17487 49203 17493
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 49970 17348 49976 17400
rect 50028 17388 50034 17400
rect 50706 17388 50712 17400
rect 50028 17360 50712 17388
rect 50028 17348 50034 17360
rect 50706 17348 50712 17360
rect 50764 17348 50770 17400
rect 1762 17280 1768 17332
rect 1820 17320 1826 17332
rect 3605 17323 3663 17329
rect 3605 17320 3617 17323
rect 1820 17292 3617 17320
rect 1820 17280 1826 17292
rect 3605 17289 3617 17292
rect 3651 17289 3663 17323
rect 3605 17283 3663 17289
rect 4614 17280 4620 17332
rect 4672 17320 4678 17332
rect 5997 17323 6055 17329
rect 5997 17320 6009 17323
rect 4672 17292 6009 17320
rect 4672 17280 4678 17292
rect 5997 17289 6009 17292
rect 6043 17289 6055 17323
rect 5997 17283 6055 17289
rect 6362 17280 6368 17332
rect 6420 17320 6426 17332
rect 6733 17323 6791 17329
rect 6733 17320 6745 17323
rect 6420 17292 6745 17320
rect 6420 17280 6426 17292
rect 6733 17289 6745 17292
rect 6779 17289 6791 17323
rect 6733 17283 6791 17289
rect 7374 17280 7380 17332
rect 7432 17320 7438 17332
rect 7745 17323 7803 17329
rect 7745 17320 7757 17323
rect 7432 17292 7757 17320
rect 7432 17280 7438 17292
rect 7745 17289 7757 17292
rect 7791 17289 7803 17323
rect 12066 17320 12072 17332
rect 7745 17283 7803 17289
rect 8220 17292 12072 17320
rect 4798 17212 4804 17264
rect 4856 17252 4862 17264
rect 4893 17255 4951 17261
rect 4893 17252 4905 17255
rect 4856 17224 4905 17252
rect 4856 17212 4862 17224
rect 4893 17221 4905 17224
rect 4939 17221 4951 17255
rect 6457 17255 6515 17261
rect 4893 17215 4951 17221
rect 5276 17224 6408 17252
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17184 1823 17187
rect 1854 17184 1860 17196
rect 1811 17156 1860 17184
rect 1811 17153 1823 17156
rect 1765 17147 1823 17153
rect 1854 17144 1860 17156
rect 1912 17144 1918 17196
rect 2774 17144 2780 17196
rect 2832 17184 2838 17196
rect 3789 17187 3847 17193
rect 3789 17184 3801 17187
rect 2832 17156 3801 17184
rect 2832 17144 2838 17156
rect 3789 17153 3801 17156
rect 3835 17153 3847 17187
rect 3789 17147 3847 17153
rect 4249 17187 4307 17193
rect 4249 17153 4261 17187
rect 4295 17153 4307 17187
rect 4249 17147 4307 17153
rect 1302 17076 1308 17128
rect 1360 17116 1366 17128
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 1360 17088 2053 17116
rect 1360 17076 1366 17088
rect 2041 17085 2053 17088
rect 2087 17085 2099 17119
rect 4264 17116 4292 17147
rect 4338 17144 4344 17196
rect 4396 17184 4402 17196
rect 5276 17184 5304 17224
rect 4396 17156 5304 17184
rect 5353 17187 5411 17193
rect 4396 17144 4402 17156
rect 5353 17153 5365 17187
rect 5399 17184 5411 17187
rect 5442 17184 5448 17196
rect 5399 17156 5448 17184
rect 5399 17153 5411 17156
rect 5353 17147 5411 17153
rect 5442 17144 5448 17156
rect 5500 17144 5506 17196
rect 6380 17184 6408 17224
rect 6457 17221 6469 17255
rect 6503 17252 6515 17255
rect 8110 17252 8116 17264
rect 6503 17224 8116 17252
rect 6503 17221 6515 17224
rect 6457 17215 6515 17221
rect 8110 17212 8116 17224
rect 8168 17212 8174 17264
rect 6549 17187 6607 17193
rect 6549 17184 6561 17187
rect 6380 17156 6561 17184
rect 6549 17153 6561 17156
rect 6595 17184 6607 17187
rect 6730 17184 6736 17196
rect 6595 17156 6736 17184
rect 6595 17153 6607 17156
rect 6549 17147 6607 17153
rect 6730 17144 6736 17156
rect 6788 17144 6794 17196
rect 8220 17193 8248 17292
rect 12066 17280 12072 17292
rect 12124 17280 12130 17332
rect 12434 17280 12440 17332
rect 12492 17280 12498 17332
rect 13814 17320 13820 17332
rect 13188 17292 13820 17320
rect 8680 17224 9536 17252
rect 7101 17187 7159 17193
rect 7101 17153 7113 17187
rect 7147 17153 7159 17187
rect 7101 17147 7159 17153
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17153 8263 17187
rect 8205 17147 8263 17153
rect 7006 17116 7012 17128
rect 4264 17088 7012 17116
rect 2041 17079 2099 17085
rect 7006 17076 7012 17088
rect 7064 17076 7070 17128
rect 7116 17116 7144 17147
rect 8478 17116 8484 17128
rect 7116 17088 8484 17116
rect 8478 17076 8484 17088
rect 8536 17076 8542 17128
rect 3329 17051 3387 17057
rect 3329 17017 3341 17051
rect 3375 17048 3387 17051
rect 7742 17048 7748 17060
rect 3375 17020 7748 17048
rect 3375 17017 3387 17020
rect 3329 17011 3387 17017
rect 7742 17008 7748 17020
rect 7800 17048 7806 17060
rect 8680 17048 8708 17224
rect 9309 17187 9367 17193
rect 9309 17153 9321 17187
rect 9355 17184 9367 17187
rect 9508 17184 9536 17224
rect 9950 17212 9956 17264
rect 10008 17212 10014 17264
rect 11517 17255 11575 17261
rect 11517 17252 11529 17255
rect 10152 17224 11529 17252
rect 10152 17184 10180 17224
rect 11517 17221 11529 17224
rect 11563 17252 11575 17255
rect 13188 17252 13216 17292
rect 13814 17280 13820 17292
rect 13872 17280 13878 17332
rect 14001 17323 14059 17329
rect 14001 17289 14013 17323
rect 14047 17320 14059 17323
rect 14458 17320 14464 17332
rect 14047 17292 14464 17320
rect 14047 17289 14059 17292
rect 14001 17283 14059 17289
rect 14458 17280 14464 17292
rect 14516 17280 14522 17332
rect 15470 17280 15476 17332
rect 15528 17320 15534 17332
rect 15565 17323 15623 17329
rect 15565 17320 15577 17323
rect 15528 17292 15577 17320
rect 15528 17280 15534 17292
rect 15565 17289 15577 17292
rect 15611 17289 15623 17323
rect 18877 17323 18935 17329
rect 18877 17320 18889 17323
rect 15565 17283 15623 17289
rect 17052 17292 18889 17320
rect 17052 17264 17080 17292
rect 18877 17289 18889 17292
rect 18923 17289 18935 17323
rect 24854 17320 24860 17332
rect 18877 17283 18935 17289
rect 22940 17292 24860 17320
rect 11563 17224 13216 17252
rect 11563 17221 11575 17224
rect 11517 17215 11575 17221
rect 13262 17212 13268 17264
rect 13320 17252 13326 17264
rect 13320 17224 13860 17252
rect 13320 17212 13326 17224
rect 9355 17156 9444 17184
rect 9508 17156 10180 17184
rect 9355 17153 9367 17156
rect 9309 17147 9367 17153
rect 9416 17048 9444 17156
rect 10226 17144 10232 17196
rect 10284 17184 10290 17196
rect 10781 17187 10839 17193
rect 10781 17184 10793 17187
rect 10284 17156 10793 17184
rect 10284 17144 10290 17156
rect 10781 17153 10793 17156
rect 10827 17153 10839 17187
rect 10781 17147 10839 17153
rect 10962 17144 10968 17196
rect 11020 17184 11026 17196
rect 12529 17187 12587 17193
rect 12529 17184 12541 17187
rect 11020 17156 12541 17184
rect 11020 17144 11026 17156
rect 12529 17153 12541 17156
rect 12575 17153 12587 17187
rect 12529 17147 12587 17153
rect 13357 17187 13415 17193
rect 13357 17153 13369 17187
rect 13403 17153 13415 17187
rect 13832 17184 13860 17224
rect 13906 17212 13912 17264
rect 13964 17252 13970 17264
rect 17034 17252 17040 17264
rect 13964 17224 17040 17252
rect 13964 17212 13970 17224
rect 17034 17212 17040 17224
rect 17092 17212 17098 17264
rect 17494 17252 17500 17264
rect 17144 17224 17500 17252
rect 14461 17187 14519 17193
rect 14461 17184 14473 17187
rect 13832 17156 14473 17184
rect 13357 17147 13415 17153
rect 14461 17153 14473 17156
rect 14507 17184 14519 17187
rect 15010 17184 15016 17196
rect 14507 17156 15016 17184
rect 14507 17153 14519 17156
rect 14461 17147 14519 17153
rect 10042 17076 10048 17128
rect 10100 17116 10106 17128
rect 10594 17116 10600 17128
rect 10100 17088 10600 17116
rect 10100 17076 10106 17088
rect 10594 17076 10600 17088
rect 10652 17116 10658 17128
rect 10873 17119 10931 17125
rect 10873 17116 10885 17119
rect 10652 17088 10885 17116
rect 10652 17076 10658 17088
rect 10873 17085 10885 17088
rect 10919 17085 10931 17119
rect 10873 17079 10931 17085
rect 11057 17119 11115 17125
rect 11057 17085 11069 17119
rect 11103 17116 11115 17119
rect 12618 17116 12624 17128
rect 11103 17088 12624 17116
rect 11103 17085 11115 17088
rect 11057 17079 11115 17085
rect 12618 17076 12624 17088
rect 12676 17076 12682 17128
rect 13372 17116 13400 17147
rect 15010 17144 15016 17156
rect 15068 17144 15074 17196
rect 15470 17144 15476 17196
rect 15528 17184 15534 17196
rect 17144 17193 17172 17224
rect 17494 17212 17500 17224
rect 17552 17212 17558 17264
rect 17954 17212 17960 17264
rect 18012 17212 18018 17264
rect 19610 17212 19616 17264
rect 19668 17212 19674 17264
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 15528 17156 15945 17184
rect 15528 17144 15534 17156
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 17129 17187 17187 17193
rect 17129 17153 17141 17187
rect 17175 17153 17187 17187
rect 17129 17147 17187 17153
rect 18690 17144 18696 17196
rect 18748 17184 18754 17196
rect 18748 17156 19196 17184
rect 18748 17144 18754 17156
rect 15746 17116 15752 17128
rect 13372 17088 15752 17116
rect 15746 17076 15752 17088
rect 15804 17076 15810 17128
rect 16022 17076 16028 17128
rect 16080 17076 16086 17128
rect 16114 17076 16120 17128
rect 16172 17076 16178 17128
rect 16298 17076 16304 17128
rect 16356 17116 16362 17128
rect 17405 17119 17463 17125
rect 17405 17116 17417 17119
rect 16356 17088 17417 17116
rect 16356 17076 16362 17088
rect 17405 17085 17417 17088
rect 17451 17085 17463 17119
rect 19168 17116 19196 17156
rect 19242 17144 19248 17196
rect 19300 17184 19306 17196
rect 19337 17187 19395 17193
rect 19337 17184 19349 17187
rect 19300 17156 19349 17184
rect 19300 17144 19306 17156
rect 19337 17153 19349 17156
rect 19383 17153 19395 17187
rect 20990 17184 20996 17196
rect 20746 17156 20996 17184
rect 19337 17147 19395 17153
rect 20990 17144 20996 17156
rect 21048 17184 21054 17196
rect 22005 17187 22063 17193
rect 21048 17156 21312 17184
rect 21048 17144 21054 17156
rect 21284 17128 21312 17156
rect 22005 17153 22017 17187
rect 22051 17184 22063 17187
rect 22940 17184 22968 17292
rect 24854 17280 24860 17292
rect 24912 17280 24918 17332
rect 25317 17323 25375 17329
rect 25317 17289 25329 17323
rect 25363 17320 25375 17323
rect 25406 17320 25412 17332
rect 25363 17292 25412 17320
rect 25363 17289 25375 17292
rect 25317 17283 25375 17289
rect 25406 17280 25412 17292
rect 25464 17280 25470 17332
rect 26605 17323 26663 17329
rect 26605 17289 26617 17323
rect 26651 17320 26663 17323
rect 26786 17320 26792 17332
rect 26651 17292 26792 17320
rect 26651 17289 26663 17292
rect 26605 17283 26663 17289
rect 26786 17280 26792 17292
rect 26844 17280 26850 17332
rect 30098 17280 30104 17332
rect 30156 17320 30162 17332
rect 31573 17323 31631 17329
rect 31573 17320 31585 17323
rect 30156 17292 31585 17320
rect 30156 17280 30162 17292
rect 31573 17289 31585 17292
rect 31619 17320 31631 17323
rect 31938 17320 31944 17332
rect 31619 17292 31944 17320
rect 31619 17289 31631 17292
rect 31573 17283 31631 17289
rect 31938 17280 31944 17292
rect 31996 17280 32002 17332
rect 32030 17280 32036 17332
rect 32088 17280 32094 17332
rect 32674 17280 32680 17332
rect 32732 17320 32738 17332
rect 32732 17292 34192 17320
rect 32732 17280 32738 17292
rect 24118 17212 24124 17264
rect 24176 17212 24182 17264
rect 26418 17212 26424 17264
rect 26476 17252 26482 17264
rect 27430 17252 27436 17264
rect 26476 17224 27436 17252
rect 26476 17212 26482 17224
rect 27430 17212 27436 17224
rect 27488 17252 27494 17264
rect 28810 17252 28816 17264
rect 27488 17224 28816 17252
rect 27488 17212 27494 17224
rect 28810 17212 28816 17224
rect 28868 17252 28874 17264
rect 28868 17224 29026 17252
rect 28868 17212 28874 17224
rect 30466 17212 30472 17264
rect 30524 17252 30530 17264
rect 31202 17252 31208 17264
rect 30524 17224 31208 17252
rect 30524 17212 30530 17224
rect 31202 17212 31208 17224
rect 31260 17212 31266 17264
rect 22051 17156 22968 17184
rect 22051 17153 22063 17156
rect 22005 17147 22063 17153
rect 23106 17144 23112 17196
rect 23164 17144 23170 17196
rect 25406 17144 25412 17196
rect 25464 17184 25470 17196
rect 25685 17187 25743 17193
rect 25685 17184 25697 17187
rect 25464 17156 25697 17184
rect 25464 17144 25470 17156
rect 25685 17153 25697 17156
rect 25731 17153 25743 17187
rect 25685 17147 25743 17153
rect 25777 17187 25835 17193
rect 25777 17153 25789 17187
rect 25823 17184 25835 17187
rect 26142 17184 26148 17196
rect 25823 17156 26148 17184
rect 25823 17153 25835 17156
rect 25777 17147 25835 17153
rect 26142 17144 26148 17156
rect 26200 17144 26206 17196
rect 26234 17144 26240 17196
rect 26292 17184 26298 17196
rect 27157 17187 27215 17193
rect 27157 17184 27169 17187
rect 26292 17156 27169 17184
rect 26292 17144 26298 17156
rect 27157 17153 27169 17156
rect 27203 17153 27215 17187
rect 27157 17147 27215 17153
rect 27246 17144 27252 17196
rect 27304 17184 27310 17196
rect 28261 17187 28319 17193
rect 28261 17184 28273 17187
rect 27304 17156 28273 17184
rect 27304 17144 27310 17156
rect 28261 17153 28273 17156
rect 28307 17153 28319 17187
rect 28261 17147 28319 17153
rect 30742 17144 30748 17196
rect 30800 17184 30806 17196
rect 30837 17187 30895 17193
rect 30837 17184 30849 17187
rect 30800 17156 30849 17184
rect 30800 17144 30806 17156
rect 30837 17153 30849 17156
rect 30883 17153 30895 17187
rect 30837 17147 30895 17153
rect 30929 17187 30987 17193
rect 30929 17153 30941 17187
rect 30975 17184 30987 17187
rect 30975 17156 31524 17184
rect 30975 17153 30987 17156
rect 30929 17147 30987 17153
rect 19168 17088 20760 17116
rect 17405 17079 17463 17085
rect 20732 17060 20760 17088
rect 21266 17076 21272 17128
rect 21324 17116 21330 17128
rect 21453 17119 21511 17125
rect 21453 17116 21465 17119
rect 21324 17088 21465 17116
rect 21324 17076 21330 17088
rect 21453 17085 21465 17088
rect 21499 17116 21511 17119
rect 21637 17119 21695 17125
rect 21637 17116 21649 17119
rect 21499 17088 21649 17116
rect 21499 17085 21511 17088
rect 21453 17079 21511 17085
rect 21637 17085 21649 17088
rect 21683 17116 21695 17119
rect 22370 17116 22376 17128
rect 21683 17088 22376 17116
rect 21683 17085 21695 17088
rect 21637 17079 21695 17085
rect 22370 17076 22376 17088
rect 22428 17076 22434 17128
rect 23385 17119 23443 17125
rect 23385 17085 23397 17119
rect 23431 17116 23443 17119
rect 25498 17116 25504 17128
rect 23431 17088 25504 17116
rect 23431 17085 23443 17088
rect 23385 17079 23443 17085
rect 25498 17076 25504 17088
rect 25556 17076 25562 17128
rect 25590 17076 25596 17128
rect 25648 17116 25654 17128
rect 25869 17119 25927 17125
rect 25869 17116 25881 17119
rect 25648 17088 25881 17116
rect 25648 17076 25654 17088
rect 25869 17085 25881 17088
rect 25915 17085 25927 17119
rect 25869 17079 25927 17085
rect 26421 17119 26479 17125
rect 26421 17085 26433 17119
rect 26467 17116 26479 17119
rect 26602 17116 26608 17128
rect 26467 17088 26608 17116
rect 26467 17085 26479 17088
rect 26421 17079 26479 17085
rect 26602 17076 26608 17088
rect 26660 17076 26666 17128
rect 26694 17076 26700 17128
rect 26752 17076 26758 17128
rect 28537 17119 28595 17125
rect 28537 17085 28549 17119
rect 28583 17116 28595 17119
rect 30006 17116 30012 17128
rect 28583 17088 30012 17116
rect 28583 17085 28595 17088
rect 28537 17079 28595 17085
rect 30006 17076 30012 17088
rect 30064 17076 30070 17128
rect 31021 17119 31079 17125
rect 31021 17085 31033 17119
rect 31067 17085 31079 17119
rect 31496 17116 31524 17156
rect 31570 17144 31576 17196
rect 31628 17184 31634 17196
rect 31846 17184 31852 17196
rect 31628 17156 31852 17184
rect 31628 17144 31634 17156
rect 31846 17144 31852 17156
rect 31904 17144 31910 17196
rect 31662 17116 31668 17128
rect 31496 17088 31668 17116
rect 31021 17079 31079 17085
rect 7800 17020 8708 17048
rect 8772 17020 9352 17048
rect 9416 17020 11744 17048
rect 7800 17008 7806 17020
rect 2038 16940 2044 16992
rect 2096 16980 2102 16992
rect 3602 16980 3608 16992
rect 2096 16952 3608 16980
rect 2096 16940 2102 16952
rect 3602 16940 3608 16952
rect 3660 16980 3666 16992
rect 8772 16980 8800 17020
rect 3660 16952 8800 16980
rect 8849 16983 8907 16989
rect 3660 16940 3666 16952
rect 8849 16949 8861 16983
rect 8895 16980 8907 16983
rect 9122 16980 9128 16992
rect 8895 16952 9128 16980
rect 8895 16949 8907 16952
rect 8849 16943 8907 16949
rect 9122 16940 9128 16952
rect 9180 16940 9186 16992
rect 9324 16980 9352 17020
rect 10042 16980 10048 16992
rect 9324 16952 10048 16980
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 10410 16940 10416 16992
rect 10468 16940 10474 16992
rect 11716 16980 11744 17020
rect 11790 17008 11796 17060
rect 11848 17008 11854 17060
rect 16206 17048 16212 17060
rect 11900 17020 16212 17048
rect 11900 16980 11928 17020
rect 16206 17008 16212 17020
rect 16264 17008 16270 17060
rect 18506 17008 18512 17060
rect 18564 17048 18570 17060
rect 18690 17048 18696 17060
rect 18564 17020 18696 17048
rect 18564 17008 18570 17020
rect 18690 17008 18696 17020
rect 18748 17008 18754 17060
rect 20714 17008 20720 17060
rect 20772 17008 20778 17060
rect 20898 17008 20904 17060
rect 20956 17048 20962 17060
rect 22002 17048 22008 17060
rect 20956 17020 22008 17048
rect 20956 17008 20962 17020
rect 22002 17008 22008 17020
rect 22060 17048 22066 17060
rect 22060 17020 23244 17048
rect 22060 17008 22066 17020
rect 11716 16952 11928 16980
rect 12066 16940 12072 16992
rect 12124 16940 12130 16992
rect 15102 16940 15108 16992
rect 15160 16940 15166 16992
rect 16853 16983 16911 16989
rect 16853 16949 16865 16983
rect 16899 16980 16911 16983
rect 17954 16980 17960 16992
rect 16899 16952 17960 16980
rect 16899 16949 16911 16952
rect 16853 16943 16911 16949
rect 17954 16940 17960 16952
rect 18012 16940 18018 16992
rect 18046 16940 18052 16992
rect 18104 16980 18110 16992
rect 19150 16980 19156 16992
rect 18104 16952 19156 16980
rect 18104 16940 18110 16952
rect 19150 16940 19156 16952
rect 19208 16940 19214 16992
rect 20346 16940 20352 16992
rect 20404 16980 20410 16992
rect 21085 16983 21143 16989
rect 21085 16980 21097 16983
rect 20404 16952 21097 16980
rect 20404 16940 20410 16952
rect 21085 16949 21097 16952
rect 21131 16949 21143 16983
rect 21085 16943 21143 16949
rect 22186 16940 22192 16992
rect 22244 16980 22250 16992
rect 22649 16983 22707 16989
rect 22649 16980 22661 16983
rect 22244 16952 22661 16980
rect 22244 16940 22250 16952
rect 22649 16949 22661 16952
rect 22695 16949 22707 16983
rect 23216 16980 23244 17020
rect 24486 17008 24492 17060
rect 24544 17048 24550 17060
rect 27706 17048 27712 17060
rect 24544 17020 27712 17048
rect 24544 17008 24550 17020
rect 27706 17008 27712 17020
rect 27764 17008 27770 17060
rect 29546 17008 29552 17060
rect 29604 17048 29610 17060
rect 30374 17048 30380 17060
rect 29604 17020 30380 17048
rect 29604 17008 29610 17020
rect 30374 17008 30380 17020
rect 30432 17008 30438 17060
rect 30742 17008 30748 17060
rect 30800 17048 30806 17060
rect 31036 17048 31064 17079
rect 31662 17076 31668 17088
rect 31720 17076 31726 17128
rect 31757 17119 31815 17125
rect 31757 17085 31769 17119
rect 31803 17116 31815 17119
rect 32048 17116 32076 17280
rect 32858 17212 32864 17264
rect 32916 17212 32922 17264
rect 34164 17252 34192 17292
rect 34882 17280 34888 17332
rect 34940 17320 34946 17332
rect 35253 17323 35311 17329
rect 35253 17320 35265 17323
rect 34940 17292 35265 17320
rect 34940 17280 34946 17292
rect 35253 17289 35265 17292
rect 35299 17289 35311 17323
rect 35253 17283 35311 17289
rect 35526 17280 35532 17332
rect 35584 17320 35590 17332
rect 35584 17292 37412 17320
rect 35584 17280 35590 17292
rect 35161 17255 35219 17261
rect 35161 17252 35173 17255
rect 34164 17224 35173 17252
rect 35161 17221 35173 17224
rect 35207 17221 35219 17255
rect 37274 17252 37280 17264
rect 35161 17215 35219 17221
rect 35268 17224 37280 17252
rect 32306 17144 32312 17196
rect 32364 17184 32370 17196
rect 32585 17187 32643 17193
rect 32585 17184 32597 17187
rect 32364 17156 32597 17184
rect 32364 17144 32370 17156
rect 32585 17153 32597 17156
rect 32631 17153 32643 17187
rect 34514 17184 34520 17196
rect 33994 17156 34520 17184
rect 32585 17147 32643 17153
rect 34514 17144 34520 17156
rect 34572 17144 34578 17196
rect 32122 17116 32128 17128
rect 31803 17088 32128 17116
rect 31803 17085 31815 17088
rect 31757 17079 31815 17085
rect 32122 17076 32128 17088
rect 32180 17076 32186 17128
rect 33318 17076 33324 17128
rect 33376 17116 33382 17128
rect 35268 17116 35296 17224
rect 37274 17212 37280 17224
rect 37332 17212 37338 17264
rect 37384 17252 37412 17292
rect 37550 17280 37556 17332
rect 37608 17320 37614 17332
rect 38105 17323 38163 17329
rect 38105 17320 38117 17323
rect 37608 17292 38117 17320
rect 37608 17280 37614 17292
rect 38105 17289 38117 17292
rect 38151 17289 38163 17323
rect 38105 17283 38163 17289
rect 38194 17280 38200 17332
rect 38252 17320 38258 17332
rect 38838 17320 38844 17332
rect 38252 17292 38844 17320
rect 38252 17280 38258 17292
rect 38838 17280 38844 17292
rect 38896 17280 38902 17332
rect 39022 17280 39028 17332
rect 39080 17280 39086 17332
rect 39114 17280 39120 17332
rect 39172 17320 39178 17332
rect 40865 17323 40923 17329
rect 40865 17320 40877 17323
rect 39172 17292 40877 17320
rect 39172 17280 39178 17292
rect 40865 17289 40877 17292
rect 40911 17289 40923 17323
rect 40865 17283 40923 17289
rect 40954 17280 40960 17332
rect 41012 17320 41018 17332
rect 46569 17323 46627 17329
rect 46569 17320 46581 17323
rect 41012 17292 46581 17320
rect 41012 17280 41018 17292
rect 46569 17289 46581 17292
rect 46615 17289 46627 17323
rect 46569 17283 46627 17289
rect 48406 17280 48412 17332
rect 48464 17280 48470 17332
rect 49050 17280 49056 17332
rect 49108 17320 49114 17332
rect 49108 17292 49924 17320
rect 49108 17280 49114 17292
rect 39040 17252 39068 17280
rect 40770 17252 40776 17264
rect 37384 17224 39068 17252
rect 40066 17224 40776 17252
rect 40770 17212 40776 17224
rect 40828 17212 40834 17264
rect 41138 17212 41144 17264
rect 41196 17252 41202 17264
rect 41325 17255 41383 17261
rect 41325 17252 41337 17255
rect 41196 17224 41337 17252
rect 41196 17212 41202 17224
rect 41325 17221 41337 17224
rect 41371 17221 41383 17255
rect 45830 17252 45836 17264
rect 41325 17215 41383 17221
rect 41432 17224 45836 17252
rect 35526 17144 35532 17196
rect 35584 17184 35590 17196
rect 36357 17187 36415 17193
rect 36357 17184 36369 17187
rect 35584 17156 36369 17184
rect 35584 17144 35590 17156
rect 36357 17153 36369 17156
rect 36403 17153 36415 17187
rect 36357 17147 36415 17153
rect 36538 17144 36544 17196
rect 36596 17184 36602 17196
rect 36596 17156 37136 17184
rect 36596 17144 36602 17156
rect 33376 17088 35296 17116
rect 35437 17119 35495 17125
rect 33376 17076 33382 17088
rect 35437 17085 35449 17119
rect 35483 17116 35495 17119
rect 35710 17116 35716 17128
rect 35483 17088 35716 17116
rect 35483 17085 35495 17088
rect 35437 17079 35495 17085
rect 35710 17076 35716 17088
rect 35768 17076 35774 17128
rect 36449 17119 36507 17125
rect 36449 17085 36461 17119
rect 36495 17085 36507 17119
rect 36449 17079 36507 17085
rect 30800 17020 31064 17048
rect 30800 17008 30806 17020
rect 31478 17008 31484 17060
rect 31536 17048 31542 17060
rect 32582 17048 32588 17060
rect 31536 17020 32588 17048
rect 31536 17008 31542 17020
rect 32582 17008 32588 17020
rect 32640 17008 32646 17060
rect 33870 17008 33876 17060
rect 33928 17048 33934 17060
rect 36464 17048 36492 17079
rect 36630 17076 36636 17128
rect 36688 17076 36694 17128
rect 36814 17076 36820 17128
rect 36872 17116 36878 17128
rect 37001 17119 37059 17125
rect 37001 17116 37013 17119
rect 36872 17088 37013 17116
rect 36872 17076 36878 17088
rect 37001 17085 37013 17088
rect 37047 17085 37059 17119
rect 37108 17116 37136 17156
rect 37458 17144 37464 17196
rect 37516 17144 37522 17196
rect 38286 17144 38292 17196
rect 38344 17184 38350 17196
rect 38565 17187 38623 17193
rect 38565 17184 38577 17187
rect 38344 17156 38577 17184
rect 38344 17144 38350 17156
rect 38565 17153 38577 17156
rect 38611 17153 38623 17187
rect 38565 17147 38623 17153
rect 41230 17144 41236 17196
rect 41288 17144 41294 17196
rect 41432 17184 41460 17224
rect 45830 17212 45836 17224
rect 45888 17212 45894 17264
rect 47118 17212 47124 17264
rect 47176 17252 47182 17264
rect 48961 17255 49019 17261
rect 48961 17252 48973 17255
rect 47176 17224 47808 17252
rect 47176 17212 47182 17224
rect 41386 17156 41460 17184
rect 38378 17116 38384 17128
rect 37108 17088 38384 17116
rect 37001 17079 37059 17085
rect 38378 17076 38384 17088
rect 38436 17076 38442 17128
rect 38841 17119 38899 17125
rect 38841 17085 38853 17119
rect 38887 17116 38899 17119
rect 41386 17116 41414 17156
rect 42150 17144 42156 17196
rect 42208 17144 42214 17196
rect 42610 17144 42616 17196
rect 42668 17144 42674 17196
rect 43714 17144 43720 17196
rect 43772 17144 43778 17196
rect 44821 17187 44879 17193
rect 44821 17153 44833 17187
rect 44867 17184 44879 17187
rect 45462 17184 45468 17196
rect 44867 17156 45468 17184
rect 44867 17153 44879 17156
rect 44821 17147 44879 17153
rect 45462 17144 45468 17156
rect 45520 17144 45526 17196
rect 45922 17144 45928 17196
rect 45980 17144 45986 17196
rect 47780 17193 47808 17224
rect 48700 17224 48973 17252
rect 47765 17187 47823 17193
rect 47765 17153 47777 17187
rect 47811 17153 47823 17187
rect 47765 17147 47823 17153
rect 38887 17088 41414 17116
rect 38887 17085 38899 17088
rect 38841 17079 38899 17085
rect 41506 17076 41512 17128
rect 41564 17076 41570 17128
rect 43254 17076 43260 17128
rect 43312 17076 43318 17128
rect 44082 17076 44088 17128
rect 44140 17116 44146 17128
rect 46937 17119 46995 17125
rect 46937 17116 46949 17119
rect 44140 17088 46949 17116
rect 44140 17076 44146 17088
rect 46937 17085 46949 17088
rect 46983 17116 46995 17119
rect 47029 17119 47087 17125
rect 47029 17116 47041 17119
rect 46983 17088 47041 17116
rect 46983 17085 46995 17088
rect 46937 17079 46995 17085
rect 47029 17085 47041 17088
rect 47075 17085 47087 17119
rect 47029 17079 47087 17085
rect 47118 17076 47124 17128
rect 47176 17116 47182 17128
rect 48700 17116 48728 17224
rect 48961 17221 48973 17224
rect 49007 17252 49019 17255
rect 49142 17252 49148 17264
rect 49007 17224 49148 17252
rect 49007 17221 49019 17224
rect 48961 17215 49019 17221
rect 49142 17212 49148 17224
rect 49200 17212 49206 17264
rect 48774 17144 48780 17196
rect 48832 17184 48838 17196
rect 49050 17184 49056 17196
rect 48832 17156 49056 17184
rect 48832 17144 48838 17156
rect 49050 17144 49056 17156
rect 49108 17144 49114 17196
rect 49896 17128 49924 17292
rect 47176 17088 48728 17116
rect 47176 17076 47182 17088
rect 49878 17076 49884 17128
rect 49936 17076 49942 17128
rect 37642 17048 37648 17060
rect 33928 17020 36492 17048
rect 36924 17020 37648 17048
rect 33928 17008 33934 17020
rect 24857 16983 24915 16989
rect 24857 16980 24869 16983
rect 23216 16952 24869 16980
rect 22649 16943 22707 16949
rect 24857 16949 24869 16952
rect 24903 16949 24915 16983
rect 24857 16943 24915 16949
rect 27801 16983 27859 16989
rect 27801 16949 27813 16983
rect 27847 16980 27859 16983
rect 28350 16980 28356 16992
rect 27847 16952 28356 16980
rect 27847 16949 27859 16952
rect 27801 16943 27859 16949
rect 28350 16940 28356 16952
rect 28408 16940 28414 16992
rect 29178 16940 29184 16992
rect 29236 16980 29242 16992
rect 29638 16980 29644 16992
rect 29236 16952 29644 16980
rect 29236 16940 29242 16952
rect 29638 16940 29644 16952
rect 29696 16940 29702 16992
rect 30006 16940 30012 16992
rect 30064 16940 30070 16992
rect 30469 16983 30527 16989
rect 30469 16949 30481 16983
rect 30515 16980 30527 16983
rect 31202 16980 31208 16992
rect 30515 16952 31208 16980
rect 30515 16949 30527 16952
rect 30469 16943 30527 16949
rect 31202 16940 31208 16952
rect 31260 16940 31266 16992
rect 31846 16940 31852 16992
rect 31904 16940 31910 16992
rect 32217 16983 32275 16989
rect 32217 16949 32229 16983
rect 32263 16980 32275 16983
rect 32858 16980 32864 16992
rect 32263 16952 32864 16980
rect 32263 16949 32275 16952
rect 32217 16943 32275 16949
rect 32858 16940 32864 16952
rect 32916 16940 32922 16992
rect 34330 16940 34336 16992
rect 34388 16940 34394 16992
rect 34793 16983 34851 16989
rect 34793 16949 34805 16983
rect 34839 16980 34851 16983
rect 35894 16980 35900 16992
rect 34839 16952 35900 16980
rect 34839 16949 34851 16952
rect 34793 16943 34851 16949
rect 35894 16940 35900 16952
rect 35952 16940 35958 16992
rect 35989 16983 36047 16989
rect 35989 16949 36001 16983
rect 36035 16980 36047 16983
rect 36924 16980 36952 17020
rect 37642 17008 37648 17020
rect 37700 17008 37706 17060
rect 44361 17051 44419 17057
rect 44361 17048 44373 17051
rect 39868 17020 44373 17048
rect 36035 16952 36952 16980
rect 36035 16949 36047 16952
rect 35989 16943 36047 16949
rect 38194 16940 38200 16992
rect 38252 16980 38258 16992
rect 39868 16980 39896 17020
rect 44361 17017 44373 17020
rect 44407 17017 44419 17051
rect 44361 17011 44419 17017
rect 44726 17008 44732 17060
rect 44784 17048 44790 17060
rect 45465 17051 45523 17057
rect 45465 17048 45477 17051
rect 44784 17020 45477 17048
rect 44784 17008 44790 17020
rect 45465 17017 45477 17020
rect 45511 17017 45523 17051
rect 45465 17011 45523 17017
rect 46474 17008 46480 17060
rect 46532 17048 46538 17060
rect 46750 17048 46756 17060
rect 46532 17020 46756 17048
rect 46532 17008 46538 17020
rect 46750 17008 46756 17020
rect 46808 17008 46814 17060
rect 47762 17008 47768 17060
rect 47820 17048 47826 17060
rect 49421 17051 49479 17057
rect 49421 17048 49433 17051
rect 47820 17020 49433 17048
rect 47820 17008 47826 17020
rect 49421 17017 49433 17020
rect 49467 17017 49479 17051
rect 49421 17011 49479 17017
rect 38252 16952 39896 16980
rect 40313 16983 40371 16989
rect 38252 16940 38258 16952
rect 40313 16949 40325 16983
rect 40359 16980 40371 16983
rect 40954 16980 40960 16992
rect 40359 16952 40960 16980
rect 40359 16949 40371 16952
rect 40313 16943 40371 16949
rect 40954 16940 40960 16952
rect 41012 16940 41018 16992
rect 41414 16940 41420 16992
rect 41472 16980 41478 16992
rect 41877 16983 41935 16989
rect 41877 16980 41889 16983
rect 41472 16952 41889 16980
rect 41472 16940 41478 16952
rect 41877 16949 41889 16952
rect 41923 16949 41935 16983
rect 41877 16943 41935 16949
rect 44082 16940 44088 16992
rect 44140 16980 44146 16992
rect 44266 16980 44272 16992
rect 44140 16952 44272 16980
rect 44140 16940 44146 16952
rect 44266 16940 44272 16952
rect 44324 16940 44330 16992
rect 45554 16940 45560 16992
rect 45612 16980 45618 16992
rect 49053 16983 49111 16989
rect 49053 16980 49065 16983
rect 45612 16952 49065 16980
rect 45612 16940 45618 16952
rect 49053 16949 49065 16952
rect 49099 16949 49111 16983
rect 49053 16943 49111 16949
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 2924 16748 8064 16776
rect 2924 16736 2930 16748
rect 3605 16711 3663 16717
rect 3605 16677 3617 16711
rect 3651 16708 3663 16711
rect 5350 16708 5356 16720
rect 3651 16680 5356 16708
rect 3651 16677 3663 16680
rect 3605 16671 3663 16677
rect 5350 16668 5356 16680
rect 5408 16668 5414 16720
rect 7190 16708 7196 16720
rect 6288 16680 7196 16708
rect 3421 16643 3479 16649
rect 3421 16609 3433 16643
rect 3467 16640 3479 16643
rect 6288 16640 6316 16680
rect 7190 16668 7196 16680
rect 7248 16668 7254 16720
rect 7561 16711 7619 16717
rect 7561 16677 7573 16711
rect 7607 16677 7619 16711
rect 7561 16671 7619 16677
rect 3467 16612 6316 16640
rect 6380 16612 6592 16640
rect 3467 16609 3479 16612
rect 3421 16603 3479 16609
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16572 1823 16575
rect 3878 16572 3884 16584
rect 1811 16544 3884 16572
rect 1811 16541 1823 16544
rect 1765 16535 1823 16541
rect 3878 16532 3884 16544
rect 3936 16532 3942 16584
rect 4249 16575 4307 16581
rect 4249 16541 4261 16575
rect 4295 16572 4307 16575
rect 5258 16572 5264 16584
rect 4295 16544 5264 16572
rect 4295 16541 4307 16544
rect 4249 16535 4307 16541
rect 5258 16532 5264 16544
rect 5316 16532 5322 16584
rect 5353 16575 5411 16581
rect 5353 16541 5365 16575
rect 5399 16541 5411 16575
rect 5353 16535 5411 16541
rect 1302 16464 1308 16516
rect 1360 16504 1366 16516
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1360 16476 2513 16504
rect 1360 16464 1366 16476
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 5368 16504 5396 16535
rect 5442 16532 5448 16584
rect 5500 16572 5506 16584
rect 6380 16572 6408 16612
rect 5500 16544 6408 16572
rect 6457 16575 6515 16581
rect 5500 16532 5506 16544
rect 6457 16541 6469 16575
rect 6503 16541 6515 16575
rect 6564 16572 6592 16612
rect 7101 16575 7159 16581
rect 7101 16572 7113 16575
rect 6564 16544 7113 16572
rect 6457 16535 6515 16541
rect 7101 16541 7113 16544
rect 7147 16541 7159 16575
rect 7576 16572 7604 16671
rect 8036 16649 8064 16748
rect 8294 16736 8300 16788
rect 8352 16776 8358 16788
rect 8938 16776 8944 16788
rect 8352 16748 8944 16776
rect 8352 16736 8358 16748
rect 8938 16736 8944 16748
rect 8996 16736 9002 16788
rect 10042 16736 10048 16788
rect 10100 16776 10106 16788
rect 10962 16776 10968 16788
rect 10100 16748 10968 16776
rect 10100 16736 10106 16748
rect 10962 16736 10968 16748
rect 11020 16736 11026 16788
rect 11054 16736 11060 16788
rect 11112 16776 11118 16788
rect 11112 16748 12434 16776
rect 11112 16736 11118 16748
rect 8757 16711 8815 16717
rect 8757 16677 8769 16711
rect 8803 16708 8815 16711
rect 12158 16708 12164 16720
rect 8803 16680 12164 16708
rect 8803 16677 8815 16680
rect 8757 16671 8815 16677
rect 12158 16668 12164 16680
rect 12216 16668 12222 16720
rect 12406 16708 12434 16748
rect 12618 16736 12624 16788
rect 12676 16776 12682 16788
rect 13630 16776 13636 16788
rect 12676 16748 13636 16776
rect 12676 16736 12682 16748
rect 13630 16736 13636 16748
rect 13688 16736 13694 16788
rect 13814 16736 13820 16788
rect 13872 16736 13878 16788
rect 15381 16779 15439 16785
rect 15381 16745 15393 16779
rect 15427 16776 15439 16779
rect 16022 16776 16028 16788
rect 15427 16748 16028 16776
rect 15427 16745 15439 16748
rect 15381 16739 15439 16745
rect 16022 16736 16028 16748
rect 16080 16776 16086 16788
rect 17770 16776 17776 16788
rect 16080 16748 17776 16776
rect 16080 16736 16086 16748
rect 17770 16736 17776 16748
rect 17828 16736 17834 16788
rect 17862 16736 17868 16788
rect 17920 16736 17926 16788
rect 17954 16736 17960 16788
rect 18012 16776 18018 16788
rect 18966 16776 18972 16788
rect 18012 16748 18972 16776
rect 18012 16736 18018 16748
rect 18966 16736 18972 16748
rect 19024 16776 19030 16788
rect 20533 16779 20591 16785
rect 20533 16776 20545 16779
rect 19024 16748 20545 16776
rect 19024 16736 19030 16748
rect 20533 16745 20545 16748
rect 20579 16776 20591 16779
rect 20990 16776 20996 16788
rect 20579 16748 20996 16776
rect 20579 16745 20591 16748
rect 20533 16739 20591 16745
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 21726 16776 21732 16788
rect 21100 16748 21732 16776
rect 16114 16708 16120 16720
rect 12406 16680 16120 16708
rect 16114 16668 16120 16680
rect 16172 16668 16178 16720
rect 16206 16668 16212 16720
rect 16264 16708 16270 16720
rect 18046 16708 18052 16720
rect 16264 16680 18052 16708
rect 16264 16668 16270 16680
rect 18046 16668 18052 16680
rect 18104 16668 18110 16720
rect 18340 16680 18552 16708
rect 8021 16643 8079 16649
rect 8021 16609 8033 16643
rect 8067 16609 8079 16643
rect 8021 16603 8079 16609
rect 8110 16600 8116 16652
rect 8168 16600 8174 16652
rect 8938 16600 8944 16652
rect 8996 16640 9002 16652
rect 8996 16612 11560 16640
rect 8996 16600 9002 16612
rect 9122 16572 9128 16584
rect 7576 16544 9128 16572
rect 7101 16535 7159 16541
rect 6362 16504 6368 16516
rect 5368 16476 6368 16504
rect 2501 16467 2559 16473
rect 6362 16464 6368 16476
rect 6420 16464 6426 16516
rect 6472 16504 6500 16535
rect 9122 16532 9128 16544
rect 9180 16532 9186 16584
rect 9214 16532 9220 16584
rect 9272 16532 9278 16584
rect 9861 16575 9919 16581
rect 9861 16541 9873 16575
rect 9907 16572 9919 16575
rect 10321 16575 10379 16581
rect 10321 16572 10333 16575
rect 9907 16544 10333 16572
rect 9907 16541 9919 16544
rect 9861 16535 9919 16541
rect 10321 16541 10333 16544
rect 10367 16541 10379 16575
rect 10321 16535 10379 16541
rect 10962 16532 10968 16584
rect 11020 16532 11026 16584
rect 11532 16572 11560 16612
rect 11606 16600 11612 16652
rect 11664 16640 11670 16652
rect 11977 16643 12035 16649
rect 11977 16640 11989 16643
rect 11664 16612 11989 16640
rect 11664 16600 11670 16612
rect 11977 16609 11989 16612
rect 12023 16609 12035 16643
rect 11977 16603 12035 16609
rect 13081 16643 13139 16649
rect 13081 16609 13093 16643
rect 13127 16609 13139 16643
rect 13081 16603 13139 16609
rect 13096 16572 13124 16603
rect 13262 16600 13268 16652
rect 13320 16600 13326 16652
rect 13814 16600 13820 16652
rect 13872 16640 13878 16652
rect 14829 16643 14887 16649
rect 14829 16640 14841 16643
rect 13872 16612 14841 16640
rect 13872 16600 13878 16612
rect 14829 16609 14841 16612
rect 14875 16609 14887 16643
rect 14829 16603 14887 16609
rect 11532 16544 13492 16572
rect 11054 16504 11060 16516
rect 6472 16476 11060 16504
rect 11054 16464 11060 16476
rect 11112 16464 11118 16516
rect 11146 16464 11152 16516
rect 11204 16504 11210 16516
rect 13464 16504 13492 16544
rect 13538 16532 13544 16584
rect 13596 16572 13602 16584
rect 14642 16572 14648 16584
rect 13596 16544 14648 16572
rect 13596 16532 13602 16544
rect 14642 16532 14648 16544
rect 14700 16532 14706 16584
rect 14734 16532 14740 16584
rect 14792 16532 14798 16584
rect 14844 16572 14872 16603
rect 15746 16600 15752 16652
rect 15804 16640 15810 16652
rect 17954 16640 17960 16652
rect 15804 16612 17960 16640
rect 15804 16600 15810 16612
rect 17954 16600 17960 16612
rect 18012 16600 18018 16652
rect 18340 16640 18368 16680
rect 18156 16612 18368 16640
rect 18417 16643 18475 16649
rect 15102 16572 15108 16584
rect 14844 16544 15108 16572
rect 15102 16532 15108 16544
rect 15160 16532 15166 16584
rect 15645 16575 15703 16581
rect 15645 16572 15657 16575
rect 15580 16544 15657 16572
rect 13725 16507 13783 16513
rect 11204 16476 12112 16504
rect 13464 16476 13676 16504
rect 11204 16464 11210 16476
rect 3602 16396 3608 16448
rect 3660 16436 3666 16448
rect 3881 16439 3939 16445
rect 3881 16436 3893 16439
rect 3660 16408 3893 16436
rect 3660 16396 3666 16408
rect 3881 16405 3893 16408
rect 3927 16405 3939 16439
rect 3881 16399 3939 16405
rect 4893 16439 4951 16445
rect 4893 16405 4905 16439
rect 4939 16436 4951 16439
rect 5902 16436 5908 16448
rect 4939 16408 5908 16436
rect 4939 16405 4951 16408
rect 4893 16399 4951 16405
rect 5902 16396 5908 16408
rect 5960 16396 5966 16448
rect 5997 16439 6055 16445
rect 5997 16405 6009 16439
rect 6043 16436 6055 16439
rect 6822 16436 6828 16448
rect 6043 16408 6828 16436
rect 6043 16405 6055 16408
rect 5997 16399 6055 16405
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 7190 16396 7196 16448
rect 7248 16436 7254 16448
rect 7929 16439 7987 16445
rect 7929 16436 7941 16439
rect 7248 16408 7941 16436
rect 7248 16396 7254 16408
rect 7929 16405 7941 16408
rect 7975 16405 7987 16439
rect 7929 16399 7987 16405
rect 9030 16396 9036 16448
rect 9088 16436 9094 16448
rect 9214 16436 9220 16448
rect 9088 16408 9220 16436
rect 9088 16396 9094 16408
rect 9214 16396 9220 16408
rect 9272 16396 9278 16448
rect 10870 16396 10876 16448
rect 10928 16436 10934 16448
rect 11425 16439 11483 16445
rect 11425 16436 11437 16439
rect 10928 16408 11437 16436
rect 10928 16396 10934 16408
rect 11425 16405 11437 16408
rect 11471 16405 11483 16439
rect 11425 16399 11483 16405
rect 11790 16396 11796 16448
rect 11848 16396 11854 16448
rect 11882 16396 11888 16448
rect 11940 16396 11946 16448
rect 12084 16436 12112 16476
rect 12342 16436 12348 16448
rect 12084 16408 12348 16436
rect 12342 16396 12348 16408
rect 12400 16396 12406 16448
rect 12434 16396 12440 16448
rect 12492 16436 12498 16448
rect 12621 16439 12679 16445
rect 12621 16436 12633 16439
rect 12492 16408 12633 16436
rect 12492 16396 12498 16408
rect 12621 16405 12633 16408
rect 12667 16405 12679 16439
rect 12621 16399 12679 16405
rect 12986 16396 12992 16448
rect 13044 16436 13050 16448
rect 13538 16436 13544 16448
rect 13044 16408 13544 16436
rect 13044 16396 13050 16408
rect 13538 16396 13544 16408
rect 13596 16396 13602 16448
rect 13648 16436 13676 16476
rect 13725 16473 13737 16507
rect 13771 16504 13783 16507
rect 13814 16504 13820 16516
rect 13771 16476 13820 16504
rect 13771 16473 13783 16476
rect 13725 16467 13783 16473
rect 13814 16464 13820 16476
rect 13872 16464 13878 16516
rect 14752 16504 14780 16532
rect 14200 16476 14780 16504
rect 15580 16504 15608 16544
rect 15645 16541 15657 16544
rect 15691 16541 15703 16575
rect 15645 16535 15703 16541
rect 16301 16575 16359 16581
rect 16301 16541 16313 16575
rect 16347 16572 16359 16575
rect 16574 16572 16580 16584
rect 16347 16544 16580 16572
rect 16347 16541 16359 16544
rect 16301 16535 16359 16541
rect 16574 16532 16580 16544
rect 16632 16532 16638 16584
rect 16758 16532 16764 16584
rect 16816 16532 16822 16584
rect 17405 16575 17463 16581
rect 17405 16541 17417 16575
rect 17451 16572 17463 16575
rect 18156 16572 18184 16612
rect 18417 16609 18429 16643
rect 18463 16609 18475 16643
rect 18417 16603 18475 16609
rect 18432 16572 18460 16603
rect 17451 16544 18184 16572
rect 18248 16544 18460 16572
rect 18524 16572 18552 16680
rect 19150 16668 19156 16720
rect 19208 16708 19214 16720
rect 21100 16708 21128 16748
rect 21726 16736 21732 16748
rect 21784 16736 21790 16788
rect 21910 16736 21916 16788
rect 21968 16776 21974 16788
rect 23750 16776 23756 16788
rect 21968 16748 23756 16776
rect 21968 16736 21974 16748
rect 23750 16736 23756 16748
rect 23808 16736 23814 16788
rect 24302 16736 24308 16788
rect 24360 16776 24366 16788
rect 24581 16779 24639 16785
rect 24581 16776 24593 16779
rect 24360 16748 24593 16776
rect 24360 16736 24366 16748
rect 24581 16745 24593 16748
rect 24627 16745 24639 16779
rect 24581 16739 24639 16745
rect 25212 16779 25270 16785
rect 25212 16745 25224 16779
rect 25258 16776 25270 16779
rect 26602 16776 26608 16788
rect 25258 16748 26608 16776
rect 25258 16745 25270 16748
rect 25212 16739 25270 16745
rect 26602 16736 26608 16748
rect 26660 16736 26666 16788
rect 26694 16736 26700 16788
rect 26752 16776 26758 16788
rect 27157 16779 27215 16785
rect 27157 16776 27169 16779
rect 26752 16748 27169 16776
rect 26752 16736 26758 16748
rect 27157 16745 27169 16748
rect 27203 16776 27215 16779
rect 27982 16776 27988 16788
rect 27203 16748 27988 16776
rect 27203 16745 27215 16748
rect 27157 16739 27215 16745
rect 27982 16736 27988 16748
rect 28040 16736 28046 16788
rect 29546 16776 29552 16788
rect 28644 16748 29552 16776
rect 19208 16680 20116 16708
rect 19208 16668 19214 16680
rect 18966 16600 18972 16652
rect 19024 16640 19030 16652
rect 19702 16640 19708 16652
rect 19024 16612 19708 16640
rect 19024 16600 19030 16612
rect 19702 16600 19708 16612
rect 19760 16600 19766 16652
rect 20088 16649 20116 16680
rect 20640 16680 21128 16708
rect 27065 16711 27123 16717
rect 20073 16643 20131 16649
rect 20073 16609 20085 16643
rect 20119 16640 20131 16643
rect 20346 16640 20352 16652
rect 20119 16612 20352 16640
rect 20119 16609 20131 16612
rect 20073 16603 20131 16609
rect 20346 16600 20352 16612
rect 20404 16600 20410 16652
rect 19889 16575 19947 16581
rect 18524 16544 19380 16572
rect 17451 16541 17463 16544
rect 17405 16535 17463 16541
rect 16390 16504 16396 16516
rect 15580 16476 16396 16504
rect 14200 16436 14228 16476
rect 16390 16464 16396 16476
rect 16448 16464 16454 16516
rect 17862 16504 17868 16516
rect 16776 16476 17868 16504
rect 13648 16408 14228 16436
rect 14277 16439 14335 16445
rect 14277 16405 14289 16439
rect 14323 16436 14335 16439
rect 14458 16436 14464 16448
rect 14323 16408 14464 16436
rect 14323 16405 14335 16408
rect 14277 16399 14335 16405
rect 14458 16396 14464 16408
rect 14516 16396 14522 16448
rect 15010 16396 15016 16448
rect 15068 16436 15074 16448
rect 16776 16436 16804 16476
rect 17862 16464 17868 16476
rect 17920 16464 17926 16516
rect 18248 16504 18276 16544
rect 18156 16476 18276 16504
rect 18325 16507 18383 16513
rect 15068 16408 16804 16436
rect 15068 16396 15074 16408
rect 16850 16396 16856 16448
rect 16908 16436 16914 16448
rect 18156 16436 18184 16476
rect 18325 16473 18337 16507
rect 18371 16504 18383 16507
rect 19352 16504 19380 16544
rect 19889 16541 19901 16575
rect 19935 16572 19947 16575
rect 20640 16572 20668 16680
rect 27065 16677 27077 16711
rect 27111 16708 27123 16711
rect 27522 16708 27528 16720
rect 27111 16680 27528 16708
rect 27111 16677 27123 16680
rect 27065 16671 27123 16677
rect 27522 16668 27528 16680
rect 27580 16668 27586 16720
rect 28644 16708 28672 16748
rect 29546 16736 29552 16748
rect 29604 16736 29610 16788
rect 29638 16736 29644 16788
rect 29696 16776 29702 16788
rect 29733 16779 29791 16785
rect 29733 16776 29745 16779
rect 29696 16748 29745 16776
rect 29696 16736 29702 16748
rect 29733 16745 29745 16748
rect 29779 16745 29791 16779
rect 29733 16739 29791 16745
rect 30006 16736 30012 16788
rect 30064 16776 30070 16788
rect 30190 16776 30196 16788
rect 30064 16748 30196 16776
rect 30064 16736 30070 16748
rect 30190 16736 30196 16748
rect 30248 16776 30254 16788
rect 33318 16776 33324 16788
rect 30248 16748 33324 16776
rect 30248 16736 30254 16748
rect 33318 16736 33324 16748
rect 33376 16736 33382 16788
rect 33686 16736 33692 16788
rect 33744 16776 33750 16788
rect 34238 16776 34244 16788
rect 33744 16748 34244 16776
rect 33744 16736 33750 16748
rect 34238 16736 34244 16748
rect 34296 16736 34302 16788
rect 34698 16736 34704 16788
rect 34756 16776 34762 16788
rect 35526 16776 35532 16788
rect 34756 16748 35532 16776
rect 34756 16736 34762 16748
rect 35526 16736 35532 16748
rect 35584 16736 35590 16788
rect 37093 16779 37151 16785
rect 36188 16748 37044 16776
rect 27724 16680 28672 16708
rect 20714 16600 20720 16652
rect 20772 16600 20778 16652
rect 20806 16600 20812 16652
rect 20864 16640 20870 16652
rect 20993 16643 21051 16649
rect 20993 16640 21005 16643
rect 20864 16612 21005 16640
rect 20864 16600 20870 16612
rect 20993 16609 21005 16612
rect 21039 16640 21051 16643
rect 22830 16640 22836 16652
rect 21039 16612 22836 16640
rect 21039 16609 21051 16612
rect 20993 16603 21051 16609
rect 22830 16600 22836 16612
rect 22888 16600 22894 16652
rect 23937 16643 23995 16649
rect 23937 16609 23949 16643
rect 23983 16640 23995 16643
rect 24762 16640 24768 16652
rect 23983 16612 24768 16640
rect 23983 16609 23995 16612
rect 23937 16603 23995 16609
rect 24762 16600 24768 16612
rect 24820 16600 24826 16652
rect 24949 16643 25007 16649
rect 24949 16609 24961 16643
rect 24995 16640 25007 16643
rect 25958 16640 25964 16652
rect 24995 16612 25964 16640
rect 24995 16609 25007 16612
rect 24949 16603 25007 16609
rect 25958 16600 25964 16612
rect 26016 16600 26022 16652
rect 27338 16600 27344 16652
rect 27396 16640 27402 16652
rect 27724 16640 27752 16680
rect 29822 16668 29828 16720
rect 29880 16708 29886 16720
rect 32309 16711 32367 16717
rect 29880 16680 30236 16708
rect 29880 16668 29886 16680
rect 27396 16612 27752 16640
rect 27396 16600 27402 16612
rect 27982 16600 27988 16652
rect 28040 16600 28046 16652
rect 28169 16643 28227 16649
rect 28169 16609 28181 16643
rect 28215 16640 28227 16643
rect 28534 16640 28540 16652
rect 28215 16612 28540 16640
rect 28215 16609 28227 16612
rect 28169 16603 28227 16609
rect 28534 16600 28540 16612
rect 28592 16600 28598 16652
rect 28810 16600 28816 16652
rect 28868 16640 28874 16652
rect 30006 16640 30012 16652
rect 28868 16612 30012 16640
rect 28868 16600 28874 16612
rect 30006 16600 30012 16612
rect 30064 16600 30070 16652
rect 30098 16600 30104 16652
rect 30156 16600 30162 16652
rect 30208 16640 30236 16680
rect 31680 16680 31892 16708
rect 31680 16640 31708 16680
rect 30208 16612 31708 16640
rect 31864 16640 31892 16680
rect 32309 16677 32321 16711
rect 32355 16708 32367 16711
rect 32355 16680 34008 16708
rect 32355 16677 32367 16680
rect 32309 16671 32367 16677
rect 32769 16643 32827 16649
rect 32769 16640 32781 16643
rect 31864 16612 32781 16640
rect 32769 16609 32781 16612
rect 32815 16609 32827 16643
rect 32769 16603 32827 16609
rect 32953 16643 33011 16649
rect 32953 16609 32965 16643
rect 32999 16640 33011 16643
rect 33318 16640 33324 16652
rect 32999 16612 33324 16640
rect 32999 16609 33011 16612
rect 32953 16603 33011 16609
rect 33318 16600 33324 16612
rect 33376 16600 33382 16652
rect 33410 16600 33416 16652
rect 33468 16600 33474 16652
rect 33980 16649 34008 16680
rect 33965 16643 34023 16649
rect 33965 16609 33977 16643
rect 34011 16609 34023 16643
rect 33965 16603 34023 16609
rect 34149 16643 34207 16649
rect 34149 16609 34161 16643
rect 34195 16640 34207 16643
rect 34195 16612 34376 16640
rect 34195 16609 34207 16612
rect 34149 16603 34207 16609
rect 19935 16544 20668 16572
rect 19935 16541 19947 16544
rect 19889 16535 19947 16541
rect 22370 16532 22376 16584
rect 22428 16572 22434 16584
rect 23382 16572 23388 16584
rect 22428 16544 23388 16572
rect 22428 16532 22434 16544
rect 23382 16532 23388 16544
rect 23440 16572 23446 16584
rect 24118 16572 24124 16584
rect 23440 16544 24124 16572
rect 23440 16532 23446 16544
rect 24118 16532 24124 16544
rect 24176 16572 24182 16584
rect 24397 16575 24455 16581
rect 24397 16572 24409 16575
rect 24176 16544 24409 16572
rect 24176 16532 24182 16544
rect 24397 16541 24409 16544
rect 24443 16541 24455 16575
rect 24397 16535 24455 16541
rect 21269 16507 21327 16513
rect 21269 16504 21281 16507
rect 18371 16476 18644 16504
rect 19352 16476 21281 16504
rect 18371 16473 18383 16476
rect 18325 16467 18383 16473
rect 18616 16448 18644 16476
rect 21269 16473 21281 16476
rect 21315 16473 21327 16507
rect 23842 16504 23848 16516
rect 21269 16467 21327 16473
rect 22756 16476 23848 16504
rect 16908 16408 18184 16436
rect 16908 16396 16914 16408
rect 18230 16396 18236 16448
rect 18288 16396 18294 16448
rect 18598 16396 18604 16448
rect 18656 16396 18662 16448
rect 19426 16396 19432 16448
rect 19484 16396 19490 16448
rect 19794 16396 19800 16448
rect 19852 16396 19858 16448
rect 19886 16396 19892 16448
rect 19944 16436 19950 16448
rect 22756 16445 22784 16476
rect 23842 16464 23848 16476
rect 23900 16464 23906 16516
rect 24412 16504 24440 16535
rect 27890 16532 27896 16584
rect 27948 16532 27954 16584
rect 29270 16532 29276 16584
rect 29328 16572 29334 16584
rect 29546 16572 29552 16584
rect 29328 16544 29552 16572
rect 29328 16532 29334 16544
rect 29546 16532 29552 16544
rect 29604 16532 29610 16584
rect 31478 16532 31484 16584
rect 31536 16532 31542 16584
rect 31938 16532 31944 16584
rect 31996 16572 32002 16584
rect 33428 16572 33456 16600
rect 31996 16544 33456 16572
rect 31996 16532 32002 16544
rect 24412 16476 25714 16504
rect 26620 16476 27568 16504
rect 22741 16439 22799 16445
rect 22741 16436 22753 16439
rect 19944 16408 22753 16436
rect 19944 16396 19950 16408
rect 22741 16405 22753 16408
rect 22787 16405 22799 16439
rect 22741 16399 22799 16405
rect 23290 16396 23296 16448
rect 23348 16396 23354 16448
rect 23658 16396 23664 16448
rect 23716 16396 23722 16448
rect 23753 16439 23811 16445
rect 23753 16405 23765 16439
rect 23799 16436 23811 16439
rect 24486 16436 24492 16448
rect 23799 16408 24492 16436
rect 23799 16405 23811 16408
rect 23753 16399 23811 16405
rect 24486 16396 24492 16408
rect 24544 16396 24550 16448
rect 26142 16396 26148 16448
rect 26200 16436 26206 16448
rect 26620 16436 26648 16476
rect 26200 16408 26648 16436
rect 26200 16396 26206 16408
rect 26694 16396 26700 16448
rect 26752 16396 26758 16448
rect 27540 16445 27568 16476
rect 27614 16464 27620 16516
rect 27672 16504 27678 16516
rect 28718 16504 28724 16516
rect 27672 16476 28724 16504
rect 27672 16464 27678 16476
rect 28718 16464 28724 16476
rect 28776 16464 28782 16516
rect 30377 16507 30435 16513
rect 30377 16473 30389 16507
rect 30423 16504 30435 16507
rect 30650 16504 30656 16516
rect 30423 16476 30656 16504
rect 30423 16473 30435 16476
rect 30377 16467 30435 16473
rect 30650 16464 30656 16476
rect 30708 16464 30714 16516
rect 34348 16504 34376 16612
rect 34422 16600 34428 16652
rect 34480 16640 34486 16652
rect 35161 16643 35219 16649
rect 34480 16612 34928 16640
rect 34480 16600 34486 16612
rect 34900 16584 34928 16612
rect 35161 16609 35173 16643
rect 35207 16640 35219 16643
rect 36188 16640 36216 16748
rect 37016 16708 37044 16748
rect 37093 16745 37105 16779
rect 37139 16776 37151 16779
rect 38102 16776 38108 16788
rect 37139 16748 38108 16776
rect 37139 16745 37151 16748
rect 37093 16739 37151 16745
rect 38102 16736 38108 16748
rect 38160 16736 38166 16788
rect 38746 16736 38752 16788
rect 38804 16736 38810 16788
rect 41322 16776 41328 16788
rect 40696 16748 41328 16776
rect 38194 16708 38200 16720
rect 37016 16680 38200 16708
rect 38194 16668 38200 16680
rect 38252 16668 38258 16720
rect 38562 16668 38568 16720
rect 38620 16708 38626 16720
rect 38764 16708 38792 16736
rect 40696 16708 40724 16748
rect 41322 16736 41328 16748
rect 41380 16736 41386 16788
rect 41877 16779 41935 16785
rect 41877 16745 41889 16779
rect 41923 16776 41935 16779
rect 42242 16776 42248 16788
rect 41923 16748 42248 16776
rect 41923 16745 41935 16748
rect 41877 16739 41935 16745
rect 42242 16736 42248 16748
rect 42300 16736 42306 16788
rect 42981 16779 43039 16785
rect 42981 16745 42993 16779
rect 43027 16776 43039 16779
rect 43714 16776 43720 16788
rect 43027 16748 43720 16776
rect 43027 16745 43039 16748
rect 42981 16739 43039 16745
rect 43714 16736 43720 16748
rect 43772 16736 43778 16788
rect 44818 16736 44824 16788
rect 44876 16776 44882 16788
rect 49421 16779 49479 16785
rect 49421 16776 49433 16779
rect 44876 16748 49433 16776
rect 44876 16736 44882 16748
rect 47228 16720 47256 16748
rect 49421 16745 49433 16748
rect 49467 16745 49479 16779
rect 49421 16739 49479 16745
rect 44542 16708 44548 16720
rect 38620 16680 38792 16708
rect 40236 16680 40724 16708
rect 41616 16680 44548 16708
rect 38620 16668 38626 16680
rect 40236 16652 40264 16680
rect 35207 16612 36216 16640
rect 37737 16643 37795 16649
rect 35207 16609 35219 16612
rect 35161 16603 35219 16609
rect 37737 16609 37749 16643
rect 37783 16640 37795 16643
rect 38838 16640 38844 16652
rect 37783 16612 38844 16640
rect 37783 16609 37795 16612
rect 37737 16603 37795 16609
rect 38838 16600 38844 16612
rect 38896 16600 38902 16652
rect 38933 16643 38991 16649
rect 38933 16609 38945 16643
rect 38979 16640 38991 16643
rect 39298 16640 39304 16652
rect 38979 16612 39304 16640
rect 38979 16609 38991 16612
rect 38933 16603 38991 16609
rect 39298 16600 39304 16612
rect 39356 16600 39362 16652
rect 39482 16600 39488 16652
rect 39540 16600 39546 16652
rect 40218 16600 40224 16652
rect 40276 16600 40282 16652
rect 40494 16600 40500 16652
rect 40552 16600 40558 16652
rect 40681 16643 40739 16649
rect 40681 16609 40693 16643
rect 40727 16640 40739 16643
rect 40954 16640 40960 16652
rect 40727 16612 40960 16640
rect 40727 16609 40739 16612
rect 40681 16603 40739 16609
rect 40954 16600 40960 16612
rect 41012 16640 41018 16652
rect 41616 16640 41644 16680
rect 44542 16668 44548 16680
rect 44600 16668 44606 16720
rect 45186 16668 45192 16720
rect 45244 16708 45250 16720
rect 45830 16708 45836 16720
rect 45244 16680 45836 16708
rect 45244 16668 45250 16680
rect 45830 16668 45836 16680
rect 45888 16668 45894 16720
rect 47210 16668 47216 16720
rect 47268 16668 47274 16720
rect 41012 16612 41644 16640
rect 41012 16600 41018 16612
rect 41966 16600 41972 16652
rect 42024 16640 42030 16652
rect 44266 16640 44272 16652
rect 42024 16612 44272 16640
rect 42024 16600 42030 16612
rect 44266 16600 44272 16612
rect 44324 16600 44330 16652
rect 48406 16600 48412 16652
rect 48464 16640 48470 16652
rect 48958 16640 48964 16652
rect 48464 16612 48964 16640
rect 48464 16600 48470 16612
rect 48958 16600 48964 16612
rect 49016 16600 49022 16652
rect 34882 16532 34888 16584
rect 34940 16532 34946 16584
rect 41233 16575 41291 16581
rect 41233 16572 41245 16575
rect 36464 16544 41245 16572
rect 31864 16476 34376 16504
rect 27525 16439 27583 16445
rect 27525 16405 27537 16439
rect 27571 16405 27583 16439
rect 27525 16399 27583 16405
rect 27706 16396 27712 16448
rect 27764 16436 27770 16448
rect 28537 16439 28595 16445
rect 28537 16436 28549 16439
rect 27764 16408 28549 16436
rect 27764 16396 27770 16408
rect 28537 16405 28549 16408
rect 28583 16405 28595 16439
rect 28537 16399 28595 16405
rect 28902 16396 28908 16448
rect 28960 16396 28966 16448
rect 31864 16445 31892 16476
rect 31849 16439 31907 16445
rect 31849 16405 31861 16439
rect 31895 16405 31907 16439
rect 31849 16399 31907 16405
rect 32677 16439 32735 16445
rect 32677 16405 32689 16439
rect 32723 16436 32735 16439
rect 33318 16436 33324 16448
rect 32723 16408 33324 16436
rect 32723 16405 32735 16408
rect 32677 16399 32735 16405
rect 33318 16396 33324 16408
rect 33376 16396 33382 16448
rect 33505 16439 33563 16445
rect 33505 16405 33517 16439
rect 33551 16436 33563 16439
rect 33594 16436 33600 16448
rect 33551 16408 33600 16436
rect 33551 16405 33563 16408
rect 33505 16399 33563 16405
rect 33594 16396 33600 16408
rect 33652 16396 33658 16448
rect 33686 16396 33692 16448
rect 33744 16436 33750 16448
rect 33873 16439 33931 16445
rect 33873 16436 33885 16439
rect 33744 16408 33885 16436
rect 33744 16396 33750 16408
rect 33873 16405 33885 16408
rect 33919 16405 33931 16439
rect 34348 16436 34376 16476
rect 35802 16464 35808 16516
rect 35860 16464 35866 16516
rect 36464 16436 36492 16544
rect 41233 16541 41245 16544
rect 41279 16541 41291 16575
rect 41233 16535 41291 16541
rect 42337 16575 42395 16581
rect 42337 16541 42349 16575
rect 42383 16572 42395 16575
rect 43346 16572 43352 16584
rect 42383 16544 43352 16572
rect 42383 16541 42395 16544
rect 42337 16535 42395 16541
rect 43346 16532 43352 16544
rect 43404 16532 43410 16584
rect 43441 16575 43499 16581
rect 43441 16541 43453 16575
rect 43487 16572 43499 16575
rect 44358 16572 44364 16584
rect 43487 16544 44364 16572
rect 43487 16541 43499 16544
rect 43441 16535 43499 16541
rect 44358 16532 44364 16544
rect 44416 16532 44422 16584
rect 44450 16532 44456 16584
rect 44508 16572 44514 16584
rect 44729 16575 44787 16581
rect 44729 16572 44741 16575
rect 44508 16544 44741 16572
rect 44508 16532 44514 16544
rect 44729 16541 44741 16544
rect 44775 16541 44787 16575
rect 44729 16535 44787 16541
rect 45186 16532 45192 16584
rect 45244 16532 45250 16584
rect 45462 16532 45468 16584
rect 45520 16572 45526 16584
rect 45833 16575 45891 16581
rect 45833 16572 45845 16575
rect 45520 16544 45845 16572
rect 45520 16532 45526 16544
rect 45833 16541 45845 16544
rect 45879 16541 45891 16575
rect 45833 16535 45891 16541
rect 46293 16575 46351 16581
rect 46293 16541 46305 16575
rect 46339 16541 46351 16575
rect 46293 16535 46351 16541
rect 37001 16507 37059 16513
rect 37001 16473 37013 16507
rect 37047 16504 37059 16507
rect 37461 16507 37519 16513
rect 37461 16504 37473 16507
rect 37047 16476 37473 16504
rect 37047 16473 37059 16476
rect 37001 16467 37059 16473
rect 37461 16473 37473 16476
rect 37507 16504 37519 16507
rect 37734 16504 37740 16516
rect 37507 16476 37740 16504
rect 37507 16473 37519 16476
rect 37461 16467 37519 16473
rect 37734 16464 37740 16476
rect 37792 16464 37798 16516
rect 39482 16504 39488 16516
rect 38212 16476 39488 16504
rect 34348 16408 36492 16436
rect 33873 16399 33931 16405
rect 36630 16396 36636 16448
rect 36688 16396 36694 16448
rect 37553 16439 37611 16445
rect 37553 16405 37565 16439
rect 37599 16436 37611 16439
rect 38212 16436 38240 16476
rect 39482 16464 39488 16476
rect 39540 16464 39546 16516
rect 40405 16507 40463 16513
rect 40405 16473 40417 16507
rect 40451 16504 40463 16507
rect 41874 16504 41880 16516
rect 40451 16476 41880 16504
rect 40451 16473 40463 16476
rect 40405 16467 40463 16473
rect 41874 16464 41880 16476
rect 41932 16504 41938 16516
rect 44545 16507 44603 16513
rect 44545 16504 44557 16507
rect 41932 16476 44557 16504
rect 41932 16464 41938 16476
rect 44545 16473 44557 16476
rect 44591 16473 44603 16507
rect 44545 16467 44603 16473
rect 45370 16464 45376 16516
rect 45428 16504 45434 16516
rect 46308 16504 46336 16535
rect 47210 16532 47216 16584
rect 47268 16572 47274 16584
rect 47397 16575 47455 16581
rect 47397 16572 47409 16575
rect 47268 16544 47409 16572
rect 47268 16532 47274 16544
rect 47397 16541 47409 16544
rect 47443 16541 47455 16575
rect 47397 16535 47455 16541
rect 48501 16575 48559 16581
rect 48501 16541 48513 16575
rect 48547 16572 48559 16575
rect 48774 16572 48780 16584
rect 48547 16544 48780 16572
rect 48547 16541 48559 16544
rect 48501 16535 48559 16541
rect 48774 16532 48780 16544
rect 48832 16532 48838 16584
rect 45428 16476 46336 16504
rect 45428 16464 45434 16476
rect 49234 16464 49240 16516
rect 49292 16504 49298 16516
rect 49292 16476 49924 16504
rect 49292 16464 49298 16476
rect 37599 16408 38240 16436
rect 38289 16439 38347 16445
rect 37599 16405 37611 16408
rect 37553 16399 37611 16405
rect 38289 16405 38301 16439
rect 38335 16436 38347 16439
rect 38378 16436 38384 16448
rect 38335 16408 38384 16436
rect 38335 16405 38347 16408
rect 38289 16399 38347 16405
rect 38378 16396 38384 16408
rect 38436 16396 38442 16448
rect 38654 16396 38660 16448
rect 38712 16396 38718 16448
rect 38746 16396 38752 16448
rect 38804 16396 38810 16448
rect 39393 16439 39451 16445
rect 39393 16405 39405 16439
rect 39439 16436 39451 16439
rect 39666 16436 39672 16448
rect 39439 16408 39672 16436
rect 39439 16405 39451 16408
rect 39393 16399 39451 16405
rect 39666 16396 39672 16408
rect 39724 16396 39730 16448
rect 40034 16396 40040 16448
rect 40092 16396 40098 16448
rect 42242 16396 42248 16448
rect 42300 16436 42306 16448
rect 44085 16439 44143 16445
rect 44085 16436 44097 16439
rect 42300 16408 44097 16436
rect 42300 16396 42306 16408
rect 44085 16405 44097 16408
rect 44131 16405 44143 16439
rect 44085 16399 44143 16405
rect 44453 16439 44511 16445
rect 44453 16405 44465 16439
rect 44499 16436 44511 16439
rect 45462 16436 45468 16448
rect 44499 16408 45468 16436
rect 44499 16405 44511 16408
rect 44453 16399 44511 16405
rect 45462 16396 45468 16408
rect 45520 16396 45526 16448
rect 45922 16396 45928 16448
rect 45980 16436 45986 16448
rect 46937 16439 46995 16445
rect 46937 16436 46949 16439
rect 45980 16408 46949 16436
rect 45980 16396 45986 16408
rect 46937 16405 46949 16408
rect 46983 16405 46995 16439
rect 46937 16399 46995 16405
rect 47026 16396 47032 16448
rect 47084 16436 47090 16448
rect 47394 16436 47400 16448
rect 47084 16408 47400 16436
rect 47084 16396 47090 16408
rect 47394 16396 47400 16408
rect 47452 16396 47458 16448
rect 48041 16439 48099 16445
rect 48041 16405 48053 16439
rect 48087 16436 48099 16439
rect 48498 16436 48504 16448
rect 48087 16408 48504 16436
rect 48087 16405 48099 16408
rect 48041 16399 48099 16405
rect 48498 16396 48504 16408
rect 48556 16396 48562 16448
rect 48958 16396 48964 16448
rect 49016 16436 49022 16448
rect 49145 16439 49203 16445
rect 49145 16436 49157 16439
rect 49016 16408 49157 16436
rect 49016 16396 49022 16408
rect 49145 16405 49157 16408
rect 49191 16405 49203 16439
rect 49145 16399 49203 16405
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 5994 16192 6000 16244
rect 6052 16192 6058 16244
rect 6362 16192 6368 16244
rect 6420 16232 6426 16244
rect 7742 16232 7748 16244
rect 6420 16204 7748 16232
rect 6420 16192 6426 16204
rect 7742 16192 7748 16204
rect 7800 16192 7806 16244
rect 7834 16192 7840 16244
rect 7892 16232 7898 16244
rect 7892 16204 8248 16232
rect 7892 16192 7898 16204
rect 3789 16167 3847 16173
rect 3789 16133 3801 16167
rect 3835 16164 3847 16167
rect 3970 16164 3976 16176
rect 3835 16136 3976 16164
rect 3835 16133 3847 16136
rect 3789 16127 3847 16133
rect 3970 16124 3976 16136
rect 4028 16124 4034 16176
rect 7098 16124 7104 16176
rect 7156 16164 7162 16176
rect 7285 16167 7343 16173
rect 7285 16164 7297 16167
rect 7156 16136 7297 16164
rect 7156 16124 7162 16136
rect 7285 16133 7297 16136
rect 7331 16133 7343 16167
rect 7285 16127 7343 16133
rect 1762 16056 1768 16108
rect 1820 16056 1826 16108
rect 3602 16056 3608 16108
rect 3660 16056 3666 16108
rect 4249 16099 4307 16105
rect 4249 16065 4261 16099
rect 4295 16096 4307 16099
rect 5258 16096 5264 16108
rect 4295 16068 5264 16096
rect 4295 16065 4307 16068
rect 4249 16059 4307 16065
rect 5258 16056 5264 16068
rect 5316 16056 5322 16108
rect 5353 16099 5411 16105
rect 5353 16065 5365 16099
rect 5399 16065 5411 16099
rect 5353 16059 5411 16065
rect 1302 15988 1308 16040
rect 1360 16028 1366 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1360 16000 2053 16028
rect 1360 15988 1366 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 3878 15988 3884 16040
rect 3936 16028 3942 16040
rect 5368 16028 5396 16059
rect 6454 16056 6460 16108
rect 6512 16096 6518 16108
rect 6641 16099 6699 16105
rect 6641 16096 6653 16099
rect 6512 16068 6653 16096
rect 6512 16056 6518 16068
rect 6641 16065 6653 16068
rect 6687 16065 6699 16099
rect 6641 16059 6699 16065
rect 8110 16056 8116 16108
rect 8168 16056 8174 16108
rect 8220 16096 8248 16204
rect 8846 16192 8852 16244
rect 8904 16232 8910 16244
rect 8904 16204 11836 16232
rect 8904 16192 8910 16204
rect 8662 16124 8668 16176
rect 8720 16164 8726 16176
rect 10778 16164 10784 16176
rect 8720 16136 10784 16164
rect 8720 16124 8726 16136
rect 10778 16124 10784 16136
rect 10836 16124 10842 16176
rect 11808 16164 11836 16204
rect 11882 16192 11888 16244
rect 11940 16232 11946 16244
rect 11977 16235 12035 16241
rect 11977 16232 11989 16235
rect 11940 16204 11989 16232
rect 11940 16192 11946 16204
rect 11977 16201 11989 16204
rect 12023 16201 12035 16235
rect 11977 16195 12035 16201
rect 12434 16192 12440 16244
rect 12492 16192 12498 16244
rect 13173 16235 13231 16241
rect 13173 16232 13185 16235
rect 12636 16204 13185 16232
rect 12158 16164 12164 16176
rect 11808 16136 12164 16164
rect 12158 16124 12164 16136
rect 12216 16124 12222 16176
rect 12345 16167 12403 16173
rect 12345 16133 12357 16167
rect 12391 16164 12403 16167
rect 12636 16164 12664 16204
rect 13173 16201 13185 16204
rect 13219 16201 13231 16235
rect 13173 16195 13231 16201
rect 13446 16192 13452 16244
rect 13504 16232 13510 16244
rect 13541 16235 13599 16241
rect 13541 16232 13553 16235
rect 13504 16204 13553 16232
rect 13504 16192 13510 16204
rect 13541 16201 13553 16204
rect 13587 16201 13599 16235
rect 13541 16195 13599 16201
rect 14826 16192 14832 16244
rect 14884 16232 14890 16244
rect 15378 16232 15384 16244
rect 14884 16204 15384 16232
rect 14884 16192 14890 16204
rect 15378 16192 15384 16204
rect 15436 16192 15442 16244
rect 15562 16192 15568 16244
rect 15620 16232 15626 16244
rect 15933 16235 15991 16241
rect 15933 16232 15945 16235
rect 15620 16204 15945 16232
rect 15620 16192 15626 16204
rect 15933 16201 15945 16204
rect 15979 16201 15991 16235
rect 15933 16195 15991 16201
rect 16022 16192 16028 16244
rect 16080 16192 16086 16244
rect 16390 16192 16396 16244
rect 16448 16232 16454 16244
rect 20898 16232 20904 16244
rect 16448 16204 20904 16232
rect 16448 16192 16454 16204
rect 20898 16192 20904 16204
rect 20956 16192 20962 16244
rect 21174 16192 21180 16244
rect 21232 16232 21238 16244
rect 23290 16232 23296 16244
rect 21232 16204 23296 16232
rect 21232 16192 21238 16204
rect 23290 16192 23296 16204
rect 23348 16192 23354 16244
rect 24302 16192 24308 16244
rect 24360 16232 24366 16244
rect 24765 16235 24823 16241
rect 24765 16232 24777 16235
rect 24360 16204 24777 16232
rect 24360 16192 24366 16204
rect 24765 16201 24777 16204
rect 24811 16201 24823 16235
rect 24765 16195 24823 16201
rect 24854 16192 24860 16244
rect 24912 16232 24918 16244
rect 25866 16232 25872 16244
rect 24912 16204 25872 16232
rect 24912 16192 24918 16204
rect 25866 16192 25872 16204
rect 25924 16232 25930 16244
rect 26694 16232 26700 16244
rect 25924 16204 26700 16232
rect 25924 16192 25930 16204
rect 26694 16192 26700 16204
rect 26752 16192 26758 16244
rect 27338 16192 27344 16244
rect 27396 16232 27402 16244
rect 27617 16235 27675 16241
rect 27617 16232 27629 16235
rect 27396 16204 27629 16232
rect 27396 16192 27402 16204
rect 27617 16201 27629 16204
rect 27663 16201 27675 16235
rect 27617 16195 27675 16201
rect 28902 16192 28908 16244
rect 28960 16232 28966 16244
rect 29917 16235 29975 16241
rect 29917 16232 29929 16235
rect 28960 16204 29929 16232
rect 28960 16192 28966 16204
rect 29917 16201 29929 16204
rect 29963 16201 29975 16235
rect 29917 16195 29975 16201
rect 30650 16192 30656 16244
rect 30708 16232 30714 16244
rect 30834 16232 30840 16244
rect 30708 16204 30840 16232
rect 30708 16192 30714 16204
rect 30834 16192 30840 16204
rect 30892 16192 30898 16244
rect 31205 16235 31263 16241
rect 31205 16201 31217 16235
rect 31251 16232 31263 16235
rect 31570 16232 31576 16244
rect 31251 16204 31576 16232
rect 31251 16201 31263 16204
rect 31205 16195 31263 16201
rect 31570 16192 31576 16204
rect 31628 16232 31634 16244
rect 31846 16232 31852 16244
rect 31628 16204 31852 16232
rect 31628 16192 31634 16204
rect 31846 16192 31852 16204
rect 31904 16192 31910 16244
rect 31938 16192 31944 16244
rect 31996 16232 32002 16244
rect 32214 16232 32220 16244
rect 31996 16204 32220 16232
rect 31996 16192 32002 16204
rect 32214 16192 32220 16204
rect 32272 16192 32278 16244
rect 32309 16235 32367 16241
rect 32309 16201 32321 16235
rect 32355 16232 32367 16235
rect 32398 16232 32404 16244
rect 32355 16204 32404 16232
rect 32355 16201 32367 16204
rect 32309 16195 32367 16201
rect 32398 16192 32404 16204
rect 32456 16192 32462 16244
rect 32769 16235 32827 16241
rect 32769 16201 32781 16235
rect 32815 16232 32827 16235
rect 32858 16232 32864 16244
rect 32815 16204 32864 16232
rect 32815 16201 32827 16204
rect 32769 16195 32827 16201
rect 32858 16192 32864 16204
rect 32916 16192 32922 16244
rect 33505 16235 33563 16241
rect 33505 16201 33517 16235
rect 33551 16232 33563 16235
rect 34698 16232 34704 16244
rect 33551 16204 34704 16232
rect 33551 16201 33563 16204
rect 33505 16195 33563 16201
rect 34698 16192 34704 16204
rect 34756 16192 34762 16244
rect 35268 16204 39896 16232
rect 14550 16164 14556 16176
rect 12391 16136 12664 16164
rect 12728 16136 14556 16164
rect 12391 16133 12403 16136
rect 12345 16127 12403 16133
rect 8220 16068 8432 16096
rect 3936 16000 5396 16028
rect 3936 15988 3942 16000
rect 4798 15852 4804 15904
rect 4856 15892 4862 15904
rect 4893 15895 4951 15901
rect 4893 15892 4905 15895
rect 4856 15864 4905 15892
rect 4856 15852 4862 15864
rect 4893 15861 4905 15864
rect 4939 15861 4951 15895
rect 5368 15892 5396 16000
rect 5810 15988 5816 16040
rect 5868 16028 5874 16040
rect 8404 16037 8432 16068
rect 8570 16056 8576 16108
rect 8628 16096 8634 16108
rect 9401 16099 9459 16105
rect 9401 16096 9413 16099
rect 8628 16068 9413 16096
rect 8628 16056 8634 16068
rect 9401 16065 9413 16068
rect 9447 16065 9459 16099
rect 9401 16059 9459 16065
rect 10502 16056 10508 16108
rect 10560 16056 10566 16108
rect 12728 16096 12756 16136
rect 14550 16124 14556 16136
rect 14608 16124 14614 16176
rect 14936 16136 16712 16164
rect 13538 16096 13544 16108
rect 12084 16068 12756 16096
rect 13004 16068 13544 16096
rect 8205 16031 8263 16037
rect 8205 16028 8217 16031
rect 5868 16000 8217 16028
rect 5868 15988 5874 16000
rect 8205 15997 8217 16000
rect 8251 15997 8263 16031
rect 8205 15991 8263 15997
rect 8389 16031 8447 16037
rect 8389 15997 8401 16031
rect 8435 16028 8447 16031
rect 9030 16028 9036 16040
rect 8435 16000 9036 16028
rect 8435 15997 8447 16000
rect 8389 15991 8447 15997
rect 9030 15988 9036 16000
rect 9088 15988 9094 16040
rect 12084 16028 12112 16068
rect 9140 16000 12112 16028
rect 12621 16031 12679 16037
rect 7742 15920 7748 15972
rect 7800 15920 7806 15972
rect 7926 15920 7932 15972
rect 7984 15960 7990 15972
rect 9140 15960 9168 16000
rect 12621 15997 12633 16031
rect 12667 16028 12679 16031
rect 13004 16028 13032 16068
rect 13538 16056 13544 16068
rect 13596 16056 13602 16108
rect 13633 16099 13691 16105
rect 13633 16065 13645 16099
rect 13679 16096 13691 16099
rect 13906 16096 13912 16108
rect 13679 16068 13912 16096
rect 13679 16065 13691 16068
rect 13633 16059 13691 16065
rect 13906 16056 13912 16068
rect 13964 16056 13970 16108
rect 14734 16056 14740 16108
rect 14792 16056 14798 16108
rect 12667 16000 13032 16028
rect 12667 15997 12679 16000
rect 12621 15991 12679 15997
rect 13262 15988 13268 16040
rect 13320 16028 13326 16040
rect 13722 16028 13728 16040
rect 13320 16000 13728 16028
rect 13320 15988 13326 16000
rect 13722 15988 13728 16000
rect 13780 16028 13786 16040
rect 14936 16037 14964 16136
rect 14921 16031 14979 16037
rect 14921 16028 14933 16031
rect 13780 16000 14933 16028
rect 13780 15988 13786 16000
rect 14921 15997 14933 16000
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 15102 15988 15108 16040
rect 15160 16028 15166 16040
rect 16114 16028 16120 16040
rect 15160 16000 16120 16028
rect 15160 15988 15166 16000
rect 16114 15988 16120 16000
rect 16172 15988 16178 16040
rect 16298 15988 16304 16040
rect 16356 15988 16362 16040
rect 16684 16028 16712 16136
rect 16850 16124 16856 16176
rect 16908 16124 16914 16176
rect 17681 16167 17739 16173
rect 17681 16133 17693 16167
rect 17727 16164 17739 16167
rect 17770 16164 17776 16176
rect 17727 16136 17776 16164
rect 17727 16133 17739 16136
rect 17681 16127 17739 16133
rect 17770 16124 17776 16136
rect 17828 16124 17834 16176
rect 17954 16124 17960 16176
rect 18012 16164 18018 16176
rect 19429 16167 19487 16173
rect 19429 16164 19441 16167
rect 18012 16136 19441 16164
rect 18012 16124 18018 16136
rect 19429 16133 19441 16136
rect 19475 16133 19487 16167
rect 19429 16127 19487 16133
rect 20714 16124 20720 16176
rect 20772 16164 20778 16176
rect 20772 16136 26832 16164
rect 20772 16124 20778 16136
rect 16761 16099 16819 16105
rect 16761 16065 16773 16099
rect 16807 16096 16819 16099
rect 17589 16099 17647 16105
rect 17589 16096 17601 16099
rect 16807 16068 17601 16096
rect 16807 16065 16819 16068
rect 16761 16059 16819 16065
rect 17589 16065 17601 16068
rect 17635 16096 17647 16099
rect 18509 16099 18567 16105
rect 17635 16068 18460 16096
rect 17635 16065 17647 16068
rect 17589 16059 17647 16065
rect 17402 16028 17408 16040
rect 16684 16000 17408 16028
rect 17402 15988 17408 16000
rect 17460 15988 17466 16040
rect 17773 16031 17831 16037
rect 17773 15997 17785 16031
rect 17819 15997 17831 16031
rect 18432 16028 18460 16068
rect 18509 16065 18521 16099
rect 18555 16096 18567 16099
rect 18598 16096 18604 16108
rect 18555 16068 18604 16096
rect 18555 16065 18567 16068
rect 18509 16059 18567 16065
rect 18598 16056 18604 16068
rect 18656 16056 18662 16108
rect 18690 16056 18696 16108
rect 18748 16056 18754 16108
rect 19150 16056 19156 16108
rect 19208 16056 19214 16108
rect 20990 16096 20996 16108
rect 20562 16068 20996 16096
rect 20990 16056 20996 16068
rect 21048 16056 21054 16108
rect 21082 16056 21088 16108
rect 21140 16096 21146 16108
rect 21361 16099 21419 16105
rect 21361 16096 21373 16099
rect 21140 16068 21373 16096
rect 21140 16056 21146 16068
rect 21361 16065 21373 16068
rect 21407 16096 21419 16099
rect 21634 16096 21640 16108
rect 21407 16068 21640 16096
rect 21407 16065 21419 16068
rect 21361 16059 21419 16065
rect 21634 16056 21640 16068
rect 21692 16056 21698 16108
rect 22373 16099 22431 16105
rect 22373 16096 22385 16099
rect 21744 16068 22385 16096
rect 18782 16028 18788 16040
rect 18432 16000 18788 16028
rect 17773 15991 17831 15997
rect 7984 15932 9168 15960
rect 7984 15920 7990 15932
rect 9306 15920 9312 15972
rect 9364 15960 9370 15972
rect 11054 15960 11060 15972
rect 9364 15932 11060 15960
rect 9364 15920 9370 15932
rect 11054 15920 11060 15932
rect 11112 15920 11118 15972
rect 11149 15963 11207 15969
rect 11149 15929 11161 15963
rect 11195 15960 11207 15963
rect 16316 15960 16344 15988
rect 11195 15932 16344 15960
rect 11195 15929 11207 15932
rect 11149 15923 11207 15929
rect 16574 15920 16580 15972
rect 16632 15960 16638 15972
rect 17788 15960 17816 15991
rect 18782 15988 18788 16000
rect 18840 15988 18846 16040
rect 18892 16000 20576 16028
rect 16632 15932 17816 15960
rect 16632 15920 16638 15932
rect 17862 15920 17868 15972
rect 17920 15960 17926 15972
rect 18506 15960 18512 15972
rect 17920 15932 18512 15960
rect 17920 15920 17926 15932
rect 18506 15920 18512 15932
rect 18564 15960 18570 15972
rect 18892 15960 18920 16000
rect 18564 15932 18920 15960
rect 18564 15920 18570 15932
rect 8294 15892 8300 15904
rect 5368 15864 8300 15892
rect 4893 15855 4951 15861
rect 8294 15852 8300 15864
rect 8352 15852 8358 15904
rect 8846 15852 8852 15904
rect 8904 15852 8910 15904
rect 8938 15852 8944 15904
rect 8996 15892 9002 15904
rect 9033 15895 9091 15901
rect 9033 15892 9045 15895
rect 8996 15864 9045 15892
rect 8996 15852 9002 15864
rect 9033 15861 9045 15864
rect 9079 15861 9091 15895
rect 9033 15855 9091 15861
rect 10045 15895 10103 15901
rect 10045 15861 10057 15895
rect 10091 15892 10103 15895
rect 10594 15892 10600 15904
rect 10091 15864 10600 15892
rect 10091 15861 10103 15864
rect 10045 15855 10103 15861
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 11701 15895 11759 15901
rect 11701 15861 11713 15895
rect 11747 15892 11759 15895
rect 11882 15892 11888 15904
rect 11747 15864 11888 15892
rect 11747 15861 11759 15864
rect 11701 15855 11759 15861
rect 11882 15852 11888 15864
rect 11940 15852 11946 15904
rect 12158 15852 12164 15904
rect 12216 15892 12222 15904
rect 13906 15892 13912 15904
rect 12216 15864 13912 15892
rect 12216 15852 12222 15864
rect 13906 15852 13912 15864
rect 13964 15852 13970 15904
rect 14369 15895 14427 15901
rect 14369 15861 14381 15895
rect 14415 15892 14427 15895
rect 14734 15892 14740 15904
rect 14415 15864 14740 15892
rect 14415 15861 14427 15864
rect 14369 15855 14427 15861
rect 14734 15852 14740 15864
rect 14792 15852 14798 15904
rect 15565 15895 15623 15901
rect 15565 15861 15577 15895
rect 15611 15892 15623 15895
rect 16298 15892 16304 15904
rect 15611 15864 16304 15892
rect 15611 15861 15623 15864
rect 15565 15855 15623 15861
rect 16298 15852 16304 15864
rect 16356 15852 16362 15904
rect 17218 15852 17224 15904
rect 17276 15852 17282 15904
rect 17586 15852 17592 15904
rect 17644 15892 17650 15904
rect 17954 15892 17960 15904
rect 17644 15864 17960 15892
rect 17644 15852 17650 15864
rect 17954 15852 17960 15864
rect 18012 15852 18018 15904
rect 18782 15852 18788 15904
rect 18840 15892 18846 15904
rect 19610 15892 19616 15904
rect 18840 15864 19616 15892
rect 18840 15852 18846 15864
rect 19610 15852 19616 15864
rect 19668 15852 19674 15904
rect 20548 15892 20576 16000
rect 20898 15988 20904 16040
rect 20956 16028 20962 16040
rect 21744 16028 21772 16068
rect 22373 16065 22385 16068
rect 22419 16065 22431 16099
rect 22373 16059 22431 16065
rect 23569 16099 23627 16105
rect 23569 16065 23581 16099
rect 23615 16096 23627 16099
rect 23842 16096 23848 16108
rect 23615 16068 23848 16096
rect 23615 16065 23627 16068
rect 23569 16059 23627 16065
rect 23842 16056 23848 16068
rect 23900 16056 23906 16108
rect 24762 16056 24768 16108
rect 24820 16096 24826 16108
rect 24857 16099 24915 16105
rect 24857 16096 24869 16099
rect 24820 16068 24869 16096
rect 24820 16056 24826 16068
rect 24857 16065 24869 16068
rect 24903 16065 24915 16099
rect 24857 16059 24915 16065
rect 25314 16056 25320 16108
rect 25372 16096 25378 16108
rect 25774 16096 25780 16108
rect 25372 16068 25780 16096
rect 25372 16056 25378 16068
rect 25774 16056 25780 16068
rect 25832 16096 25838 16108
rect 25961 16099 26019 16105
rect 25961 16096 25973 16099
rect 25832 16068 25973 16096
rect 25832 16056 25838 16068
rect 25961 16065 25973 16068
rect 26007 16065 26019 16099
rect 25961 16059 26019 16065
rect 26053 16099 26111 16105
rect 26053 16065 26065 16099
rect 26099 16096 26111 16099
rect 26694 16096 26700 16108
rect 26099 16068 26700 16096
rect 26099 16065 26111 16068
rect 26053 16059 26111 16065
rect 20956 16000 21772 16028
rect 20956 15988 20962 16000
rect 22462 15988 22468 16040
rect 22520 15988 22526 16040
rect 22557 16031 22615 16037
rect 22557 15997 22569 16031
rect 22603 15997 22615 16031
rect 22557 15991 22615 15997
rect 20622 15920 20628 15972
rect 20680 15960 20686 15972
rect 22005 15963 22063 15969
rect 22005 15960 22017 15963
rect 20680 15932 22017 15960
rect 20680 15920 20686 15932
rect 22005 15929 22017 15932
rect 22051 15929 22063 15963
rect 22005 15923 22063 15929
rect 20901 15895 20959 15901
rect 20901 15892 20913 15895
rect 20548 15864 20913 15892
rect 20901 15861 20913 15864
rect 20947 15892 20959 15895
rect 20990 15892 20996 15904
rect 20947 15864 20996 15892
rect 20947 15861 20959 15864
rect 20901 15855 20959 15861
rect 20990 15852 20996 15864
rect 21048 15852 21054 15904
rect 21358 15852 21364 15904
rect 21416 15892 21422 15904
rect 21545 15895 21603 15901
rect 21545 15892 21557 15895
rect 21416 15864 21557 15892
rect 21416 15852 21422 15864
rect 21545 15861 21557 15864
rect 21591 15861 21603 15895
rect 21545 15855 21603 15861
rect 21634 15852 21640 15904
rect 21692 15892 21698 15904
rect 22572 15892 22600 15991
rect 22830 15988 22836 16040
rect 22888 16028 22894 16040
rect 23661 16031 23719 16037
rect 23661 16028 23673 16031
rect 22888 16000 23673 16028
rect 22888 15988 22894 16000
rect 23661 15997 23673 16000
rect 23707 15997 23719 16031
rect 23661 15991 23719 15997
rect 23753 16031 23811 16037
rect 23753 15997 23765 16031
rect 23799 16028 23811 16031
rect 24394 16028 24400 16040
rect 23799 16000 24400 16028
rect 23799 15997 23811 16000
rect 23753 15991 23811 15997
rect 24394 15988 24400 16000
rect 24452 15988 24458 16040
rect 25038 15988 25044 16040
rect 25096 15988 25102 16040
rect 25866 15988 25872 16040
rect 25924 16028 25930 16040
rect 26068 16028 26096 16059
rect 26694 16056 26700 16068
rect 26752 16056 26758 16108
rect 25924 16000 26096 16028
rect 26145 16031 26203 16037
rect 25924 15988 25930 16000
rect 26145 15997 26157 16031
rect 26191 15997 26203 16031
rect 26804 16028 26832 16136
rect 26878 16124 26884 16176
rect 26936 16164 26942 16176
rect 33686 16164 33692 16176
rect 26936 16136 27752 16164
rect 26936 16124 26942 16136
rect 27338 16056 27344 16108
rect 27396 16096 27402 16108
rect 27525 16099 27583 16105
rect 27525 16096 27537 16099
rect 27396 16068 27537 16096
rect 27396 16056 27402 16068
rect 27525 16065 27537 16068
rect 27571 16065 27583 16099
rect 27525 16059 27583 16065
rect 27614 16028 27620 16040
rect 26804 16000 27620 16028
rect 26145 15991 26203 15997
rect 23201 15963 23259 15969
rect 23201 15929 23213 15963
rect 23247 15960 23259 15963
rect 23566 15960 23572 15972
rect 23247 15932 23572 15960
rect 23247 15929 23259 15932
rect 23201 15923 23259 15929
rect 23566 15920 23572 15932
rect 23624 15920 23630 15972
rect 25774 15920 25780 15972
rect 25832 15960 25838 15972
rect 26160 15960 26188 15991
rect 27614 15988 27620 16000
rect 27672 15988 27678 16040
rect 27724 16037 27752 16136
rect 29564 16136 33692 16164
rect 28350 16056 28356 16108
rect 28408 16056 28414 16108
rect 27709 16031 27767 16037
rect 27709 15997 27721 16031
rect 27755 15997 27767 16031
rect 27709 15991 27767 15997
rect 28997 16031 29055 16037
rect 28997 15997 29009 16031
rect 29043 16028 29055 16031
rect 29270 16028 29276 16040
rect 29043 16000 29276 16028
rect 29043 15997 29055 16000
rect 28997 15991 29055 15997
rect 29270 15988 29276 16000
rect 29328 15988 29334 16040
rect 25832 15932 26188 15960
rect 25832 15920 25838 15932
rect 27246 15920 27252 15972
rect 27304 15960 27310 15972
rect 29564 15969 29592 16136
rect 33686 16124 33692 16136
rect 33744 16124 33750 16176
rect 34790 16124 34796 16176
rect 34848 16164 34854 16176
rect 35158 16164 35164 16176
rect 34848 16136 35164 16164
rect 34848 16124 34854 16136
rect 35158 16124 35164 16136
rect 35216 16124 35222 16176
rect 35268 16173 35296 16204
rect 35253 16167 35311 16173
rect 35253 16133 35265 16167
rect 35299 16133 35311 16167
rect 35253 16127 35311 16133
rect 35802 16124 35808 16176
rect 35860 16124 35866 16176
rect 38470 16164 38476 16176
rect 36556 16136 38476 16164
rect 29638 16056 29644 16108
rect 29696 16096 29702 16108
rect 29696 16068 30328 16096
rect 29696 16056 29702 16068
rect 30009 16031 30067 16037
rect 30009 15997 30021 16031
rect 30055 15997 30067 16031
rect 30009 15991 30067 15997
rect 29549 15963 29607 15969
rect 27304 15932 29132 15960
rect 27304 15920 27310 15932
rect 21692 15864 22600 15892
rect 21692 15852 21698 15864
rect 23290 15852 23296 15904
rect 23348 15892 23354 15904
rect 24397 15895 24455 15901
rect 24397 15892 24409 15895
rect 23348 15864 24409 15892
rect 23348 15852 23354 15864
rect 24397 15861 24409 15864
rect 24443 15861 24455 15895
rect 24397 15855 24455 15861
rect 24486 15852 24492 15904
rect 24544 15892 24550 15904
rect 25593 15895 25651 15901
rect 25593 15892 25605 15895
rect 24544 15864 25605 15892
rect 24544 15852 24550 15864
rect 25593 15861 25605 15864
rect 25639 15861 25651 15895
rect 25593 15855 25651 15861
rect 26786 15852 26792 15904
rect 26844 15892 26850 15904
rect 27157 15895 27215 15901
rect 27157 15892 27169 15895
rect 26844 15864 27169 15892
rect 26844 15852 26850 15864
rect 27157 15861 27169 15864
rect 27203 15861 27215 15895
rect 27157 15855 27215 15861
rect 27338 15852 27344 15904
rect 27396 15892 27402 15904
rect 27706 15892 27712 15904
rect 27396 15864 27712 15892
rect 27396 15852 27402 15864
rect 27706 15852 27712 15864
rect 27764 15852 27770 15904
rect 29104 15892 29132 15932
rect 29549 15929 29561 15963
rect 29595 15929 29607 15963
rect 29549 15923 29607 15929
rect 30024 15892 30052 15991
rect 30190 15988 30196 16040
rect 30248 15988 30254 16040
rect 30300 16028 30328 16068
rect 30558 16056 30564 16108
rect 30616 16096 30622 16108
rect 30616 16068 32168 16096
rect 30616 16056 30622 16068
rect 32140 16040 32168 16068
rect 32398 16056 32404 16108
rect 32456 16096 32462 16108
rect 32677 16099 32735 16105
rect 32677 16096 32689 16099
rect 32456 16068 32689 16096
rect 32456 16056 32462 16068
rect 32677 16065 32689 16068
rect 32723 16065 32735 16099
rect 32677 16059 32735 16065
rect 33873 16099 33931 16105
rect 33873 16065 33885 16099
rect 33919 16096 33931 16099
rect 34146 16096 34152 16108
rect 33919 16068 34152 16096
rect 33919 16065 33931 16068
rect 33873 16059 33931 16065
rect 34146 16056 34152 16068
rect 34204 16056 34210 16108
rect 34882 16056 34888 16108
rect 34940 16096 34946 16108
rect 34977 16099 35035 16105
rect 34977 16096 34989 16099
rect 34940 16068 34989 16096
rect 34940 16056 34946 16068
rect 34977 16065 34989 16068
rect 35023 16065 35035 16099
rect 34977 16059 35035 16065
rect 31297 16031 31355 16037
rect 31297 16028 31309 16031
rect 30300 16000 31309 16028
rect 31297 15997 31309 16000
rect 31343 15997 31355 16031
rect 31297 15991 31355 15997
rect 31389 16031 31447 16037
rect 31389 15997 31401 16031
rect 31435 15997 31447 16031
rect 31389 15991 31447 15997
rect 30374 15920 30380 15972
rect 30432 15960 30438 15972
rect 31404 15960 31432 15991
rect 32122 15988 32128 16040
rect 32180 15988 32186 16040
rect 32953 16031 33011 16037
rect 32953 15997 32965 16031
rect 32999 15997 33011 16031
rect 32953 15991 33011 15997
rect 32306 15960 32312 15972
rect 30432 15932 32312 15960
rect 30432 15920 30438 15932
rect 32306 15920 32312 15932
rect 32364 15920 32370 15972
rect 32968 15960 32996 15991
rect 33962 15988 33968 16040
rect 34020 15988 34026 16040
rect 34057 16031 34115 16037
rect 34057 15997 34069 16031
rect 34103 16028 34115 16031
rect 34330 16028 34336 16040
rect 34103 16000 34336 16028
rect 34103 15997 34115 16000
rect 34057 15991 34115 15997
rect 34330 15988 34336 16000
rect 34388 15988 34394 16040
rect 36556 16028 36584 16136
rect 38470 16124 38476 16136
rect 38528 16124 38534 16176
rect 38562 16124 38568 16176
rect 38620 16124 38626 16176
rect 39868 16164 39896 16204
rect 40034 16192 40040 16244
rect 40092 16232 40098 16244
rect 41233 16235 41291 16241
rect 41233 16232 41245 16235
rect 40092 16204 41245 16232
rect 40092 16192 40098 16204
rect 41233 16201 41245 16204
rect 41279 16201 41291 16235
rect 41233 16195 41291 16201
rect 41322 16192 41328 16244
rect 41380 16232 41386 16244
rect 42245 16235 42303 16241
rect 42245 16232 42257 16235
rect 41380 16204 42257 16232
rect 41380 16192 41386 16204
rect 42245 16201 42257 16204
rect 42291 16232 42303 16235
rect 42291 16204 42840 16232
rect 42291 16201 42303 16204
rect 42245 16195 42303 16201
rect 42702 16164 42708 16176
rect 39868 16136 42708 16164
rect 42702 16124 42708 16136
rect 42760 16124 42766 16176
rect 42812 16164 42840 16204
rect 44358 16192 44364 16244
rect 44416 16192 44422 16244
rect 44542 16192 44548 16244
rect 44600 16232 44606 16244
rect 47765 16235 47823 16241
rect 47765 16232 47777 16235
rect 44600 16204 47777 16232
rect 44600 16192 44606 16204
rect 47765 16201 47777 16204
rect 47811 16201 47823 16235
rect 47765 16195 47823 16201
rect 48774 16192 48780 16244
rect 48832 16192 48838 16244
rect 49513 16235 49571 16241
rect 49513 16201 49525 16235
rect 49559 16232 49571 16235
rect 49896 16232 49924 16476
rect 49559 16204 49924 16232
rect 49559 16201 49571 16204
rect 49513 16195 49571 16201
rect 45554 16164 45560 16176
rect 42812 16136 45560 16164
rect 45554 16124 45560 16136
rect 45612 16124 45618 16176
rect 46566 16164 46572 16176
rect 45664 16136 46572 16164
rect 36814 16056 36820 16108
rect 36872 16096 36878 16108
rect 37645 16099 37703 16105
rect 37645 16096 37657 16099
rect 36872 16068 37657 16096
rect 36872 16056 36878 16068
rect 37645 16065 37657 16068
rect 37691 16065 37703 16099
rect 37645 16059 37703 16065
rect 38286 16056 38292 16108
rect 38344 16056 38350 16108
rect 39666 16056 39672 16108
rect 39724 16056 39730 16108
rect 40402 16056 40408 16108
rect 40460 16056 40466 16108
rect 41138 16056 41144 16108
rect 41196 16056 41202 16108
rect 41248 16068 42564 16096
rect 35084 16000 36584 16028
rect 35084 15960 35112 16000
rect 36630 15988 36636 16040
rect 36688 16028 36694 16040
rect 41248 16028 41276 16068
rect 36688 16000 41276 16028
rect 36688 15988 36694 16000
rect 41322 15988 41328 16040
rect 41380 15988 41386 16040
rect 41877 16031 41935 16037
rect 41877 15997 41889 16031
rect 41923 16028 41935 16031
rect 42058 16028 42064 16040
rect 41923 16000 42064 16028
rect 41923 15997 41935 16000
rect 41877 15991 41935 15997
rect 42058 15988 42064 16000
rect 42116 16028 42122 16040
rect 42334 16028 42340 16040
rect 42116 16000 42340 16028
rect 42116 15988 42122 16000
rect 42334 15988 42340 16000
rect 42392 15988 42398 16040
rect 42536 16028 42564 16068
rect 42610 16056 42616 16108
rect 42668 16056 42674 16108
rect 43717 16099 43775 16105
rect 43717 16065 43729 16099
rect 43763 16065 43775 16099
rect 43717 16059 43775 16065
rect 43732 16028 43760 16059
rect 44818 16056 44824 16108
rect 44876 16056 44882 16108
rect 45664 16096 45692 16136
rect 46566 16124 46572 16136
rect 46624 16164 46630 16176
rect 46624 16136 47256 16164
rect 46624 16124 46630 16136
rect 45388 16068 45692 16096
rect 42536 16000 43760 16028
rect 44358 15988 44364 16040
rect 44416 16028 44422 16040
rect 45388 16028 45416 16068
rect 45922 16056 45928 16108
rect 45980 16056 45986 16108
rect 47228 16096 47256 16136
rect 47394 16124 47400 16176
rect 47452 16164 47458 16176
rect 48314 16164 48320 16176
rect 47452 16136 48320 16164
rect 47452 16124 47458 16136
rect 48314 16124 48320 16136
rect 48372 16164 48378 16176
rect 49329 16167 49387 16173
rect 49329 16164 49341 16167
rect 48372 16136 49341 16164
rect 48372 16124 48378 16136
rect 49329 16133 49341 16136
rect 49375 16133 49387 16167
rect 49329 16127 49387 16133
rect 47581 16099 47639 16105
rect 47581 16096 47593 16099
rect 46032 16068 47164 16096
rect 47228 16068 47593 16096
rect 44416 16000 45416 16028
rect 44416 15988 44422 16000
rect 45462 15988 45468 16040
rect 45520 16028 45526 16040
rect 46032 16028 46060 16068
rect 45520 16000 46060 16028
rect 47029 16031 47087 16037
rect 45520 15988 45526 16000
rect 47029 15997 47041 16031
rect 47075 15997 47087 16031
rect 47136 16028 47164 16068
rect 47581 16065 47593 16068
rect 47627 16065 47639 16099
rect 47581 16059 47639 16065
rect 48133 16099 48191 16105
rect 48133 16065 48145 16099
rect 48179 16096 48191 16099
rect 49234 16096 49240 16108
rect 48179 16068 49240 16096
rect 48179 16065 48191 16068
rect 48133 16059 48191 16065
rect 49234 16056 49240 16068
rect 49292 16056 49298 16108
rect 47136 16000 48820 16028
rect 47029 15991 47087 15997
rect 32968 15932 35112 15960
rect 36725 15963 36783 15969
rect 36725 15929 36737 15963
rect 36771 15960 36783 15963
rect 36814 15960 36820 15972
rect 36771 15932 36820 15960
rect 36771 15929 36783 15932
rect 36725 15923 36783 15929
rect 36814 15920 36820 15932
rect 36872 15920 36878 15972
rect 36998 15920 37004 15972
rect 37056 15960 37062 15972
rect 40773 15963 40831 15969
rect 40773 15960 40785 15963
rect 37056 15932 37872 15960
rect 37056 15920 37062 15932
rect 29104 15864 30052 15892
rect 30282 15852 30288 15904
rect 30340 15892 30346 15904
rect 30558 15892 30564 15904
rect 30340 15864 30564 15892
rect 30340 15852 30346 15864
rect 30558 15852 30564 15864
rect 30616 15852 30622 15904
rect 30834 15852 30840 15904
rect 30892 15852 30898 15904
rect 31938 15852 31944 15904
rect 31996 15892 32002 15904
rect 33502 15892 33508 15904
rect 31996 15864 33508 15892
rect 31996 15852 32002 15864
rect 33502 15852 33508 15864
rect 33560 15852 33566 15904
rect 34609 15895 34667 15901
rect 34609 15861 34621 15895
rect 34655 15892 34667 15895
rect 34698 15892 34704 15904
rect 34655 15864 34704 15892
rect 34655 15861 34667 15864
rect 34609 15855 34667 15861
rect 34698 15852 34704 15864
rect 34756 15852 34762 15904
rect 35618 15852 35624 15904
rect 35676 15892 35682 15904
rect 35802 15892 35808 15904
rect 35676 15864 35808 15892
rect 35676 15852 35682 15864
rect 35802 15852 35808 15864
rect 35860 15852 35866 15904
rect 37734 15852 37740 15904
rect 37792 15852 37798 15904
rect 37844 15892 37872 15932
rect 39592 15932 40785 15960
rect 39592 15892 39620 15932
rect 40773 15929 40785 15932
rect 40819 15929 40831 15963
rect 45186 15960 45192 15972
rect 40773 15923 40831 15929
rect 40880 15932 45192 15960
rect 37844 15864 39620 15892
rect 39850 15852 39856 15904
rect 39908 15892 39914 15904
rect 40037 15895 40095 15901
rect 40037 15892 40049 15895
rect 39908 15864 40049 15892
rect 39908 15852 39914 15864
rect 40037 15861 40049 15864
rect 40083 15892 40095 15895
rect 40880 15892 40908 15932
rect 45186 15920 45192 15932
rect 45244 15920 45250 15972
rect 47044 15904 47072 15991
rect 48792 15904 48820 16000
rect 40083 15864 40908 15892
rect 40083 15861 40095 15864
rect 40037 15855 40095 15861
rect 40954 15852 40960 15904
rect 41012 15892 41018 15904
rect 41414 15892 41420 15904
rect 41012 15864 41420 15892
rect 41012 15852 41018 15864
rect 41414 15852 41420 15864
rect 41472 15852 41478 15904
rect 41874 15852 41880 15904
rect 41932 15892 41938 15904
rect 42061 15895 42119 15901
rect 42061 15892 42073 15895
rect 41932 15864 42073 15892
rect 41932 15852 41938 15864
rect 42061 15861 42073 15864
rect 42107 15892 42119 15895
rect 42518 15892 42524 15904
rect 42107 15864 42524 15892
rect 42107 15861 42119 15864
rect 42061 15855 42119 15861
rect 42518 15852 42524 15864
rect 42576 15852 42582 15904
rect 42794 15852 42800 15904
rect 42852 15892 42858 15904
rect 43257 15895 43315 15901
rect 43257 15892 43269 15895
rect 42852 15864 43269 15892
rect 42852 15852 42858 15864
rect 43257 15861 43269 15864
rect 43303 15861 43315 15895
rect 43257 15855 43315 15861
rect 45462 15852 45468 15904
rect 45520 15852 45526 15904
rect 46566 15852 46572 15904
rect 46624 15852 46630 15904
rect 47026 15852 47032 15904
rect 47084 15852 47090 15904
rect 48774 15852 48780 15904
rect 48832 15892 48838 15904
rect 49053 15895 49111 15901
rect 49053 15892 49065 15895
rect 48832 15864 49065 15892
rect 48832 15852 48838 15864
rect 49053 15861 49065 15864
rect 49099 15861 49111 15895
rect 49053 15855 49111 15861
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 3605 15691 3663 15697
rect 3605 15657 3617 15691
rect 3651 15688 3663 15691
rect 3878 15688 3884 15700
rect 3651 15660 3884 15688
rect 3651 15657 3663 15660
rect 3605 15651 3663 15657
rect 3878 15648 3884 15660
rect 3936 15648 3942 15700
rect 3973 15691 4031 15697
rect 3973 15657 3985 15691
rect 4019 15688 4031 15691
rect 4062 15688 4068 15700
rect 4019 15660 4068 15688
rect 4019 15657 4031 15660
rect 3973 15651 4031 15657
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 5261 15691 5319 15697
rect 5261 15657 5273 15691
rect 5307 15688 5319 15691
rect 5350 15688 5356 15700
rect 5307 15660 5356 15688
rect 5307 15657 5319 15660
rect 5261 15651 5319 15657
rect 5350 15648 5356 15660
rect 5408 15648 5414 15700
rect 7374 15648 7380 15700
rect 7432 15648 7438 15700
rect 7469 15691 7527 15697
rect 7469 15657 7481 15691
rect 7515 15688 7527 15691
rect 7926 15688 7932 15700
rect 7515 15660 7932 15688
rect 7515 15657 7527 15660
rect 7469 15651 7527 15657
rect 7926 15648 7932 15660
rect 7984 15648 7990 15700
rect 8220 15660 11652 15688
rect 3421 15623 3479 15629
rect 3421 15589 3433 15623
rect 3467 15620 3479 15623
rect 7392 15620 7420 15648
rect 3467 15592 7420 15620
rect 3467 15589 3479 15592
rect 3421 15583 3479 15589
rect 1302 15512 1308 15564
rect 1360 15552 1366 15564
rect 2041 15555 2099 15561
rect 2041 15552 2053 15555
rect 1360 15524 2053 15552
rect 1360 15512 1366 15524
rect 2041 15521 2053 15524
rect 2087 15521 2099 15555
rect 2041 15515 2099 15521
rect 7374 15512 7380 15564
rect 7432 15552 7438 15564
rect 8110 15552 8116 15564
rect 7432 15524 8116 15552
rect 7432 15512 7438 15524
rect 8110 15512 8116 15524
rect 8168 15512 8174 15564
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15484 1823 15487
rect 3602 15484 3608 15496
rect 1811 15456 3608 15484
rect 1811 15453 1823 15456
rect 1765 15447 1823 15453
rect 3602 15444 3608 15456
rect 3660 15444 3666 15496
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15453 4215 15487
rect 4157 15447 4215 15453
rect 3418 15376 3424 15428
rect 3476 15416 3482 15428
rect 4172 15416 4200 15447
rect 4614 15444 4620 15496
rect 4672 15444 4678 15496
rect 5718 15444 5724 15496
rect 5776 15444 5782 15496
rect 6822 15444 6828 15496
rect 6880 15444 6886 15496
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15484 7987 15487
rect 8220 15484 8248 15660
rect 8478 15580 8484 15632
rect 8536 15620 8542 15632
rect 8573 15623 8631 15629
rect 8573 15620 8585 15623
rect 8536 15592 8585 15620
rect 8536 15580 8542 15592
rect 8573 15589 8585 15592
rect 8619 15589 8631 15623
rect 9214 15620 9220 15632
rect 8573 15583 8631 15589
rect 8956 15592 9220 15620
rect 8294 15512 8300 15564
rect 8352 15552 8358 15564
rect 8956 15552 8984 15592
rect 9214 15580 9220 15592
rect 9272 15580 9278 15632
rect 8352 15524 8984 15552
rect 9125 15555 9183 15561
rect 8352 15512 8358 15524
rect 9125 15521 9137 15555
rect 9171 15552 9183 15555
rect 10042 15552 10048 15564
rect 9171 15524 10048 15552
rect 9171 15521 9183 15524
rect 9125 15515 9183 15521
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 10137 15555 10195 15561
rect 10137 15521 10149 15555
rect 10183 15552 10195 15555
rect 10778 15552 10784 15564
rect 10183 15524 10784 15552
rect 10183 15521 10195 15524
rect 10137 15515 10195 15521
rect 10778 15512 10784 15524
rect 10836 15512 10842 15564
rect 11624 15484 11652 15660
rect 11698 15648 11704 15700
rect 11756 15688 11762 15700
rect 12345 15691 12403 15697
rect 12345 15688 12357 15691
rect 11756 15660 12357 15688
rect 11756 15648 11762 15660
rect 12345 15657 12357 15660
rect 12391 15657 12403 15691
rect 12345 15651 12403 15657
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 13446 15688 13452 15700
rect 12492 15660 13452 15688
rect 12492 15648 12498 15660
rect 13446 15648 13452 15660
rect 13504 15688 13510 15700
rect 13504 15660 15240 15688
rect 13504 15648 13510 15660
rect 11790 15580 11796 15632
rect 11848 15620 11854 15632
rect 14277 15623 14335 15629
rect 14277 15620 14289 15623
rect 11848 15592 14289 15620
rect 11848 15580 11854 15592
rect 14277 15589 14289 15592
rect 14323 15589 14335 15623
rect 15212 15620 15240 15660
rect 15286 15648 15292 15700
rect 15344 15688 15350 15700
rect 16761 15691 16819 15697
rect 16761 15688 16773 15691
rect 15344 15660 16773 15688
rect 15344 15648 15350 15660
rect 16761 15657 16773 15660
rect 16807 15657 16819 15691
rect 19337 15691 19395 15697
rect 19337 15688 19349 15691
rect 16761 15651 16819 15657
rect 16868 15660 19349 15688
rect 15746 15620 15752 15632
rect 14277 15583 14335 15589
rect 14660 15592 15056 15620
rect 15212 15592 15752 15620
rect 12802 15512 12808 15564
rect 12860 15512 12866 15564
rect 12986 15512 12992 15564
rect 13044 15552 13050 15564
rect 13354 15552 13360 15564
rect 13044 15524 13360 15552
rect 13044 15512 13050 15524
rect 13354 15512 13360 15524
rect 13412 15512 13418 15564
rect 13906 15512 13912 15564
rect 13964 15552 13970 15564
rect 14660 15552 14688 15592
rect 13964 15524 14688 15552
rect 13964 15512 13970 15524
rect 14734 15512 14740 15564
rect 14792 15512 14798 15564
rect 14918 15512 14924 15564
rect 14976 15512 14982 15564
rect 15028 15552 15056 15592
rect 15746 15580 15752 15592
rect 15804 15580 15810 15632
rect 16114 15620 16120 15632
rect 15856 15592 16120 15620
rect 15856 15552 15884 15592
rect 15948 15561 15976 15592
rect 16114 15580 16120 15592
rect 16172 15580 16178 15632
rect 16868 15620 16896 15660
rect 19337 15657 19349 15660
rect 19383 15688 19395 15691
rect 19518 15688 19524 15700
rect 19383 15660 19524 15688
rect 19383 15657 19395 15660
rect 19337 15651 19395 15657
rect 19518 15648 19524 15660
rect 19576 15688 19582 15700
rect 19886 15688 19892 15700
rect 19576 15660 19892 15688
rect 19576 15648 19582 15660
rect 19886 15648 19892 15660
rect 19944 15648 19950 15700
rect 20438 15648 20444 15700
rect 20496 15688 20502 15700
rect 20901 15691 20959 15697
rect 20901 15688 20913 15691
rect 20496 15660 20913 15688
rect 20496 15648 20502 15660
rect 20901 15657 20913 15660
rect 20947 15657 20959 15691
rect 20901 15651 20959 15657
rect 20990 15648 20996 15700
rect 21048 15688 21054 15700
rect 24118 15688 24124 15700
rect 21048 15660 24124 15688
rect 21048 15648 21054 15660
rect 24118 15648 24124 15660
rect 24176 15648 24182 15700
rect 24581 15691 24639 15697
rect 24581 15657 24593 15691
rect 24627 15688 24639 15691
rect 24762 15688 24768 15700
rect 24627 15660 24768 15688
rect 24627 15657 24639 15660
rect 24581 15651 24639 15657
rect 24762 15648 24768 15660
rect 24820 15648 24826 15700
rect 25501 15691 25559 15697
rect 25501 15657 25513 15691
rect 25547 15688 25559 15691
rect 26234 15688 26240 15700
rect 25547 15660 26240 15688
rect 25547 15657 25559 15660
rect 25501 15651 25559 15657
rect 26234 15648 26240 15660
rect 26292 15648 26298 15700
rect 26602 15648 26608 15700
rect 26660 15648 26666 15700
rect 29273 15691 29331 15697
rect 29273 15688 29285 15691
rect 27448 15660 29285 15688
rect 18690 15620 18696 15632
rect 16776 15592 16896 15620
rect 17236 15592 18696 15620
rect 15028 15524 15884 15552
rect 15933 15555 15991 15561
rect 15933 15521 15945 15555
rect 15979 15521 15991 15555
rect 15933 15515 15991 15521
rect 16022 15512 16028 15564
rect 16080 15552 16086 15564
rect 16776 15552 16804 15592
rect 16080 15524 16804 15552
rect 16080 15512 16086 15524
rect 16850 15512 16856 15564
rect 16908 15552 16914 15564
rect 17236 15561 17264 15592
rect 18690 15580 18696 15592
rect 18748 15580 18754 15632
rect 21818 15620 21824 15632
rect 21376 15592 21824 15620
rect 17221 15555 17279 15561
rect 17221 15552 17233 15555
rect 16908 15524 17233 15552
rect 16908 15512 16914 15524
rect 17221 15521 17233 15524
rect 17267 15521 17279 15555
rect 17221 15515 17279 15521
rect 17313 15555 17371 15561
rect 17313 15521 17325 15555
rect 17359 15521 17371 15555
rect 17313 15515 17371 15521
rect 16390 15484 16396 15496
rect 7975 15456 8248 15484
rect 8404 15456 9628 15484
rect 11624 15456 16396 15484
rect 7975 15453 7987 15456
rect 7929 15447 7987 15453
rect 5350 15416 5356 15428
rect 3476 15388 5356 15416
rect 3476 15376 3482 15388
rect 5350 15376 5356 15388
rect 5408 15376 5414 15428
rect 6365 15419 6423 15425
rect 6365 15385 6377 15419
rect 6411 15416 6423 15419
rect 8404 15416 8432 15456
rect 6411 15388 8432 15416
rect 6411 15385 6423 15388
rect 6365 15379 6423 15385
rect 9490 15376 9496 15428
rect 9548 15376 9554 15428
rect 9600 15416 9628 15456
rect 16390 15444 16396 15456
rect 16448 15484 16454 15496
rect 17328 15484 17356 15515
rect 17402 15512 17408 15564
rect 17460 15552 17466 15564
rect 18509 15555 18567 15561
rect 18509 15552 18521 15555
rect 17460 15524 18521 15552
rect 17460 15512 17466 15524
rect 18509 15521 18521 15524
rect 18555 15521 18567 15555
rect 18509 15515 18567 15521
rect 20441 15555 20499 15561
rect 20441 15521 20453 15555
rect 20487 15552 20499 15555
rect 20714 15552 20720 15564
rect 20487 15524 20720 15552
rect 20487 15521 20499 15524
rect 20441 15515 20499 15521
rect 20714 15512 20720 15524
rect 20772 15512 20778 15564
rect 20806 15512 20812 15564
rect 20864 15552 20870 15564
rect 21376 15561 21404 15592
rect 21818 15580 21824 15592
rect 21876 15580 21882 15632
rect 22278 15580 22284 15632
rect 22336 15620 22342 15632
rect 27065 15623 27123 15629
rect 27065 15620 27077 15623
rect 22336 15592 27077 15620
rect 22336 15580 22342 15592
rect 27065 15589 27077 15592
rect 27111 15589 27123 15623
rect 27065 15583 27123 15589
rect 21361 15555 21419 15561
rect 21361 15552 21373 15555
rect 20864 15524 21373 15552
rect 20864 15512 20870 15524
rect 21361 15521 21373 15524
rect 21407 15521 21419 15555
rect 21361 15515 21419 15521
rect 21450 15512 21456 15564
rect 21508 15512 21514 15564
rect 23477 15555 23535 15561
rect 23477 15552 23489 15555
rect 22756 15524 23489 15552
rect 16448 15456 17356 15484
rect 18325 15487 18383 15493
rect 16448 15444 16454 15456
rect 18325 15453 18337 15487
rect 18371 15484 18383 15487
rect 18414 15484 18420 15496
rect 18371 15456 18420 15484
rect 18371 15453 18383 15456
rect 18325 15447 18383 15453
rect 18414 15444 18420 15456
rect 18472 15484 18478 15496
rect 18969 15487 19027 15493
rect 18969 15484 18981 15487
rect 18472 15456 18981 15484
rect 18472 15444 18478 15456
rect 18969 15453 18981 15456
rect 19015 15453 19027 15487
rect 18969 15447 19027 15453
rect 19797 15487 19855 15493
rect 19797 15453 19809 15487
rect 19843 15484 19855 15487
rect 22186 15484 22192 15496
rect 19843 15456 22192 15484
rect 19843 15453 19855 15456
rect 19797 15447 19855 15453
rect 22186 15444 22192 15456
rect 22244 15444 22250 15496
rect 22281 15487 22339 15493
rect 22281 15453 22293 15487
rect 22327 15484 22339 15487
rect 22646 15484 22652 15496
rect 22327 15456 22652 15484
rect 22327 15453 22339 15456
rect 22281 15447 22339 15453
rect 22646 15444 22652 15456
rect 22704 15444 22710 15496
rect 10413 15419 10471 15425
rect 10413 15416 10425 15419
rect 9600 15388 10425 15416
rect 10413 15385 10425 15388
rect 10459 15385 10471 15419
rect 12434 15416 12440 15428
rect 11638 15388 12440 15416
rect 10413 15379 10471 15385
rect 12434 15376 12440 15388
rect 12492 15376 12498 15428
rect 14645 15419 14703 15425
rect 14645 15385 14657 15419
rect 14691 15416 14703 15419
rect 14691 15388 18000 15416
rect 14691 15385 14703 15388
rect 14645 15379 14703 15385
rect 6638 15308 6644 15360
rect 6696 15348 6702 15360
rect 9306 15348 9312 15360
rect 6696 15320 9312 15348
rect 6696 15308 6702 15320
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 9582 15308 9588 15360
rect 9640 15308 9646 15360
rect 11698 15308 11704 15360
rect 11756 15348 11762 15360
rect 11885 15351 11943 15357
rect 11885 15348 11897 15351
rect 11756 15320 11897 15348
rect 11756 15308 11762 15320
rect 11885 15317 11897 15320
rect 11931 15348 11943 15351
rect 12158 15348 12164 15360
rect 11931 15320 12164 15348
rect 11931 15317 11943 15320
rect 11885 15311 11943 15317
rect 12158 15308 12164 15320
rect 12216 15308 12222 15360
rect 12710 15308 12716 15360
rect 12768 15308 12774 15360
rect 13541 15351 13599 15357
rect 13541 15317 13553 15351
rect 13587 15348 13599 15351
rect 13630 15348 13636 15360
rect 13587 15320 13636 15348
rect 13587 15317 13599 15320
rect 13541 15311 13599 15317
rect 13630 15308 13636 15320
rect 13688 15308 13694 15360
rect 15194 15308 15200 15360
rect 15252 15348 15258 15360
rect 15473 15351 15531 15357
rect 15473 15348 15485 15351
rect 15252 15320 15485 15348
rect 15252 15308 15258 15320
rect 15473 15317 15485 15320
rect 15519 15317 15531 15351
rect 15473 15311 15531 15317
rect 15746 15308 15752 15360
rect 15804 15348 15810 15360
rect 15841 15351 15899 15357
rect 15841 15348 15853 15351
rect 15804 15320 15853 15348
rect 15804 15308 15810 15320
rect 15841 15317 15853 15320
rect 15887 15348 15899 15351
rect 16666 15348 16672 15360
rect 15887 15320 16672 15348
rect 15887 15317 15899 15320
rect 15841 15311 15899 15317
rect 16666 15308 16672 15320
rect 16724 15308 16730 15360
rect 17126 15308 17132 15360
rect 17184 15308 17190 15360
rect 17218 15308 17224 15360
rect 17276 15348 17282 15360
rect 17402 15348 17408 15360
rect 17276 15320 17408 15348
rect 17276 15308 17282 15320
rect 17402 15308 17408 15320
rect 17460 15308 17466 15360
rect 17972 15357 18000 15388
rect 21266 15376 21272 15428
rect 21324 15416 21330 15428
rect 21324 15388 21496 15416
rect 21324 15376 21330 15388
rect 17957 15351 18015 15357
rect 17957 15317 17969 15351
rect 18003 15317 18015 15351
rect 17957 15311 18015 15317
rect 18414 15308 18420 15360
rect 18472 15308 18478 15360
rect 19521 15351 19579 15357
rect 19521 15317 19533 15351
rect 19567 15348 19579 15351
rect 19610 15348 19616 15360
rect 19567 15320 19616 15348
rect 19567 15317 19579 15320
rect 19521 15311 19579 15317
rect 19610 15308 19616 15320
rect 19668 15348 19674 15360
rect 20254 15348 20260 15360
rect 19668 15320 20260 15348
rect 19668 15308 19674 15320
rect 20254 15308 20260 15320
rect 20312 15308 20318 15360
rect 21468 15348 21496 15388
rect 21634 15376 21640 15428
rect 21692 15416 21698 15428
rect 22756 15416 22784 15524
rect 23477 15521 23489 15524
rect 23523 15521 23535 15555
rect 23477 15515 23535 15521
rect 23566 15512 23572 15564
rect 23624 15552 23630 15564
rect 24394 15552 24400 15564
rect 23624 15524 24400 15552
rect 23624 15512 23630 15524
rect 24394 15512 24400 15524
rect 24452 15512 24458 15564
rect 26326 15552 26332 15564
rect 24780 15524 26332 15552
rect 23290 15444 23296 15496
rect 23348 15444 23354 15496
rect 23385 15487 23443 15493
rect 23385 15453 23397 15487
rect 23431 15484 23443 15487
rect 24780 15484 24808 15524
rect 26326 15512 26332 15524
rect 26384 15512 26390 15564
rect 23431 15456 24808 15484
rect 24857 15487 24915 15493
rect 23431 15453 23443 15456
rect 23385 15447 23443 15453
rect 24857 15453 24869 15487
rect 24903 15484 24915 15487
rect 24946 15484 24952 15496
rect 24903 15456 24952 15484
rect 24903 15453 24915 15456
rect 24857 15447 24915 15453
rect 24946 15444 24952 15456
rect 25004 15484 25010 15496
rect 25590 15484 25596 15496
rect 25004 15456 25596 15484
rect 25004 15444 25010 15456
rect 25590 15444 25596 15456
rect 25648 15444 25654 15496
rect 25961 15487 26019 15493
rect 25961 15453 25973 15487
rect 26007 15484 26019 15487
rect 26142 15484 26148 15496
rect 26007 15456 26148 15484
rect 26007 15453 26019 15456
rect 25961 15447 26019 15453
rect 26142 15444 26148 15456
rect 26200 15444 26206 15496
rect 21692 15388 22784 15416
rect 21692 15376 21698 15388
rect 24394 15376 24400 15428
rect 24452 15416 24458 15428
rect 24670 15416 24676 15428
rect 24452 15388 24676 15416
rect 24452 15376 24458 15388
rect 24670 15376 24676 15388
rect 24728 15376 24734 15428
rect 25222 15376 25228 15428
rect 25280 15416 25286 15428
rect 27448 15425 27476 15660
rect 29273 15657 29285 15660
rect 29319 15688 29331 15691
rect 31757 15691 31815 15697
rect 29319 15660 30420 15688
rect 29319 15657 29331 15660
rect 29273 15651 29331 15657
rect 27522 15580 27528 15632
rect 27580 15620 27586 15632
rect 29638 15620 29644 15632
rect 27580 15592 29644 15620
rect 27580 15580 27586 15592
rect 29638 15580 29644 15592
rect 29696 15580 29702 15632
rect 29733 15623 29791 15629
rect 29733 15589 29745 15623
rect 29779 15620 29791 15623
rect 30190 15620 30196 15632
rect 29779 15592 30196 15620
rect 29779 15589 29791 15592
rect 29733 15583 29791 15589
rect 30190 15580 30196 15592
rect 30248 15580 30254 15632
rect 27614 15512 27620 15564
rect 27672 15512 27678 15564
rect 27706 15512 27712 15564
rect 27764 15552 27770 15564
rect 27764 15524 28304 15552
rect 27764 15512 27770 15524
rect 28276 15493 28304 15524
rect 28350 15512 28356 15564
rect 28408 15552 28414 15564
rect 28902 15552 28908 15564
rect 28408 15524 28908 15552
rect 28408 15512 28414 15524
rect 28902 15512 28908 15524
rect 28960 15512 28966 15564
rect 29914 15512 29920 15564
rect 29972 15552 29978 15564
rect 29972 15524 30236 15552
rect 29972 15512 29978 15524
rect 28261 15487 28319 15493
rect 28261 15453 28273 15487
rect 28307 15453 28319 15487
rect 28261 15447 28319 15453
rect 29730 15444 29736 15496
rect 29788 15484 29794 15496
rect 30208 15493 30236 15524
rect 30282 15512 30288 15564
rect 30340 15512 30346 15564
rect 30392 15552 30420 15660
rect 31757 15657 31769 15691
rect 31803 15688 31815 15691
rect 34698 15688 34704 15700
rect 31803 15660 33364 15688
rect 31803 15657 31815 15660
rect 31757 15651 31815 15657
rect 30558 15580 30564 15632
rect 30616 15620 30622 15632
rect 32306 15620 32312 15632
rect 30616 15592 32312 15620
rect 30616 15580 30622 15592
rect 32306 15580 32312 15592
rect 32364 15580 32370 15632
rect 31938 15552 31944 15564
rect 30392 15524 31944 15552
rect 31938 15512 31944 15524
rect 31996 15512 32002 15564
rect 32401 15555 32459 15561
rect 32401 15521 32413 15555
rect 32447 15552 32459 15555
rect 32582 15552 32588 15564
rect 32447 15524 32588 15552
rect 32447 15521 32459 15524
rect 32401 15515 32459 15521
rect 32582 15512 32588 15524
rect 32640 15512 32646 15564
rect 30101 15487 30159 15493
rect 30101 15484 30113 15487
rect 29788 15456 30113 15484
rect 29788 15444 29794 15456
rect 30101 15453 30113 15456
rect 30147 15453 30159 15487
rect 30101 15447 30159 15453
rect 30193 15487 30251 15493
rect 30193 15453 30205 15487
rect 30239 15453 30251 15487
rect 30193 15447 30251 15453
rect 30374 15444 30380 15496
rect 30432 15484 30438 15496
rect 30558 15484 30564 15496
rect 30432 15456 30564 15484
rect 30432 15444 30438 15456
rect 30558 15444 30564 15456
rect 30616 15444 30622 15496
rect 30834 15444 30840 15496
rect 30892 15484 30898 15496
rect 32125 15487 32183 15493
rect 32125 15484 32137 15487
rect 30892 15456 32137 15484
rect 30892 15444 30898 15456
rect 32125 15453 32137 15456
rect 32171 15453 32183 15487
rect 32125 15447 32183 15453
rect 32217 15487 32275 15493
rect 32217 15453 32229 15487
rect 32263 15484 32275 15487
rect 32766 15484 32772 15496
rect 32263 15456 32772 15484
rect 32263 15453 32275 15456
rect 32217 15447 32275 15453
rect 32766 15444 32772 15456
rect 32824 15444 32830 15496
rect 27433 15419 27491 15425
rect 27433 15416 27445 15419
rect 25280 15388 27445 15416
rect 25280 15376 25286 15388
rect 27433 15385 27445 15388
rect 27479 15385 27491 15419
rect 27433 15379 27491 15385
rect 27522 15376 27528 15428
rect 27580 15416 27586 15428
rect 27580 15388 27752 15416
rect 27580 15376 27586 15388
rect 21913 15351 21971 15357
rect 21913 15348 21925 15351
rect 21468 15320 21925 15348
rect 21913 15317 21925 15320
rect 21959 15317 21971 15351
rect 21913 15311 21971 15317
rect 22554 15308 22560 15360
rect 22612 15348 22618 15360
rect 22925 15351 22983 15357
rect 22925 15348 22937 15351
rect 22612 15320 22937 15348
rect 22612 15308 22618 15320
rect 22925 15317 22937 15320
rect 22971 15317 22983 15351
rect 22925 15311 22983 15317
rect 23474 15308 23480 15360
rect 23532 15348 23538 15360
rect 23750 15348 23756 15360
rect 23532 15320 23756 15348
rect 23532 15308 23538 15320
rect 23750 15308 23756 15320
rect 23808 15308 23814 15360
rect 23842 15308 23848 15360
rect 23900 15348 23906 15360
rect 23937 15351 23995 15357
rect 23937 15348 23949 15351
rect 23900 15320 23949 15348
rect 23900 15308 23906 15320
rect 23937 15317 23949 15320
rect 23983 15317 23995 15351
rect 23937 15311 23995 15317
rect 24118 15308 24124 15360
rect 24176 15348 24182 15360
rect 24213 15351 24271 15357
rect 24213 15348 24225 15351
rect 24176 15320 24225 15348
rect 24176 15308 24182 15320
rect 24213 15317 24225 15320
rect 24259 15348 24271 15351
rect 25038 15348 25044 15360
rect 24259 15320 25044 15348
rect 24259 15317 24271 15320
rect 24213 15311 24271 15317
rect 25038 15308 25044 15320
rect 25096 15308 25102 15360
rect 27724 15348 27752 15388
rect 27890 15376 27896 15428
rect 27948 15416 27954 15428
rect 28905 15419 28963 15425
rect 28905 15416 28917 15419
rect 27948 15388 28917 15416
rect 27948 15376 27954 15388
rect 28905 15385 28917 15388
rect 28951 15385 28963 15419
rect 32490 15416 32496 15428
rect 28905 15379 28963 15385
rect 32416 15388 32496 15416
rect 30834 15348 30840 15360
rect 27724 15320 30840 15348
rect 30834 15308 30840 15320
rect 30892 15308 30898 15360
rect 31113 15351 31171 15357
rect 31113 15317 31125 15351
rect 31159 15348 31171 15351
rect 32416 15348 32444 15388
rect 32490 15376 32496 15388
rect 32548 15376 32554 15428
rect 33336 15416 33364 15660
rect 33612 15660 34704 15688
rect 33410 15512 33416 15564
rect 33468 15512 33474 15564
rect 33612 15561 33640 15660
rect 34698 15648 34704 15660
rect 34756 15648 34762 15700
rect 35161 15691 35219 15697
rect 35161 15657 35173 15691
rect 35207 15688 35219 15691
rect 37724 15691 37782 15697
rect 35207 15660 37412 15688
rect 35207 15657 35219 15660
rect 35161 15651 35219 15657
rect 37090 15620 37096 15632
rect 35544 15592 37096 15620
rect 33597 15555 33655 15561
rect 33597 15521 33609 15555
rect 33643 15521 33655 15555
rect 33597 15515 33655 15521
rect 34146 15512 34152 15564
rect 34204 15512 34210 15564
rect 34330 15512 34336 15564
rect 34388 15552 34394 15564
rect 35544 15552 35572 15592
rect 37090 15580 37096 15592
rect 37148 15580 37154 15632
rect 34388 15524 35572 15552
rect 34388 15512 34394 15524
rect 35802 15512 35808 15564
rect 35860 15512 35866 15564
rect 33428 15484 33456 15512
rect 34701 15487 34759 15493
rect 34701 15484 34713 15487
rect 33428 15456 34713 15484
rect 34701 15453 34713 15456
rect 34747 15453 34759 15487
rect 34701 15447 34759 15453
rect 36354 15444 36360 15496
rect 36412 15444 36418 15496
rect 37274 15416 37280 15428
rect 33336 15388 37280 15416
rect 37274 15376 37280 15388
rect 37332 15376 37338 15428
rect 31159 15320 32444 15348
rect 31159 15317 31171 15320
rect 31113 15311 31171 15317
rect 32950 15308 32956 15360
rect 33008 15308 33014 15360
rect 33321 15351 33379 15357
rect 33321 15317 33333 15351
rect 33367 15348 33379 15351
rect 34054 15348 34060 15360
rect 33367 15320 34060 15348
rect 33367 15317 33379 15320
rect 33321 15311 33379 15317
rect 34054 15308 34060 15320
rect 34112 15348 34118 15360
rect 34606 15348 34612 15360
rect 34112 15320 34612 15348
rect 34112 15308 34118 15320
rect 34606 15308 34612 15320
rect 34664 15308 34670 15360
rect 35069 15351 35127 15357
rect 35069 15317 35081 15351
rect 35115 15348 35127 15351
rect 35526 15348 35532 15360
rect 35115 15320 35532 15348
rect 35115 15317 35127 15320
rect 35069 15311 35127 15317
rect 35526 15308 35532 15320
rect 35584 15308 35590 15360
rect 35621 15351 35679 15357
rect 35621 15317 35633 15351
rect 35667 15348 35679 15351
rect 36814 15348 36820 15360
rect 35667 15320 36820 15348
rect 35667 15317 35679 15320
rect 35621 15311 35679 15317
rect 36814 15308 36820 15320
rect 36872 15308 36878 15360
rect 36998 15308 37004 15360
rect 37056 15308 37062 15360
rect 37384 15348 37412 15660
rect 37724 15657 37736 15691
rect 37770 15688 37782 15691
rect 45462 15688 45468 15700
rect 37770 15660 45468 15688
rect 37770 15657 37782 15660
rect 37724 15651 37782 15657
rect 45462 15648 45468 15660
rect 45520 15648 45526 15700
rect 39482 15580 39488 15632
rect 39540 15580 39546 15632
rect 41322 15580 41328 15632
rect 41380 15620 41386 15632
rect 41785 15623 41843 15629
rect 41785 15620 41797 15623
rect 41380 15592 41797 15620
rect 41380 15580 41386 15592
rect 41785 15589 41797 15592
rect 41831 15589 41843 15623
rect 41785 15583 41843 15589
rect 42702 15580 42708 15632
rect 42760 15620 42766 15632
rect 42889 15623 42947 15629
rect 42889 15620 42901 15623
rect 42760 15592 42901 15620
rect 42760 15580 42766 15592
rect 42889 15589 42901 15592
rect 42935 15589 42947 15623
rect 46566 15620 46572 15632
rect 42889 15583 42947 15589
rect 44008 15592 46572 15620
rect 40037 15555 40095 15561
rect 40037 15552 40049 15555
rect 37476 15524 40049 15552
rect 37476 15496 37504 15524
rect 40037 15521 40049 15524
rect 40083 15521 40095 15555
rect 40037 15515 40095 15521
rect 40313 15555 40371 15561
rect 40313 15521 40325 15555
rect 40359 15552 40371 15555
rect 44008 15552 44036 15592
rect 46566 15580 46572 15592
rect 46624 15580 46630 15632
rect 40359 15524 44036 15552
rect 40359 15521 40371 15524
rect 40313 15515 40371 15521
rect 44266 15512 44272 15564
rect 44324 15552 44330 15564
rect 45002 15552 45008 15564
rect 44324 15524 45008 15552
rect 44324 15512 44330 15524
rect 45002 15512 45008 15524
rect 45060 15552 45066 15564
rect 45189 15555 45247 15561
rect 45189 15552 45201 15555
rect 45060 15524 45201 15552
rect 45060 15512 45066 15524
rect 45189 15521 45201 15524
rect 45235 15521 45247 15555
rect 45189 15515 45247 15521
rect 45462 15512 45468 15564
rect 45520 15512 45526 15564
rect 49878 15512 49884 15564
rect 49936 15552 49942 15564
rect 49936 15524 50936 15552
rect 49936 15512 49942 15524
rect 37458 15444 37464 15496
rect 37516 15444 37522 15496
rect 38838 15444 38844 15496
rect 38896 15444 38902 15496
rect 39114 15444 39120 15496
rect 39172 15484 39178 15496
rect 39390 15484 39396 15496
rect 39172 15456 39396 15484
rect 39172 15444 39178 15456
rect 39390 15444 39396 15456
rect 39448 15444 39454 15496
rect 42242 15444 42248 15496
rect 42300 15444 42306 15496
rect 43349 15487 43407 15493
rect 43349 15453 43361 15487
rect 43395 15453 43407 15487
rect 43349 15447 43407 15453
rect 41690 15416 41696 15428
rect 41538 15388 41696 15416
rect 41690 15376 41696 15388
rect 41748 15376 41754 15428
rect 43364 15416 43392 15447
rect 44634 15444 44640 15496
rect 44692 15444 44698 15496
rect 46661 15487 46719 15493
rect 46661 15453 46673 15487
rect 46707 15453 46719 15487
rect 46661 15447 46719 15453
rect 47121 15487 47179 15493
rect 47121 15453 47133 15487
rect 47167 15453 47179 15487
rect 47121 15447 47179 15453
rect 48225 15487 48283 15493
rect 48225 15453 48237 15487
rect 48271 15484 48283 15487
rect 49326 15484 49332 15496
rect 48271 15456 49332 15484
rect 48271 15453 48283 15456
rect 48225 15447 48283 15453
rect 42352 15388 43392 15416
rect 39114 15348 39120 15360
rect 37384 15320 39120 15348
rect 39114 15308 39120 15320
rect 39172 15308 39178 15360
rect 39209 15351 39267 15357
rect 39209 15317 39221 15351
rect 39255 15348 39267 15351
rect 39298 15348 39304 15360
rect 39255 15320 39304 15348
rect 39255 15317 39267 15320
rect 39209 15311 39267 15317
rect 39298 15308 39304 15320
rect 39356 15308 39362 15360
rect 39758 15308 39764 15360
rect 39816 15348 39822 15360
rect 42352 15348 42380 15388
rect 43438 15376 43444 15428
rect 43496 15416 43502 15428
rect 46676 15416 46704 15447
rect 43496 15388 46704 15416
rect 47136 15416 47164 15447
rect 49326 15444 49332 15456
rect 49384 15444 49390 15496
rect 48314 15416 48320 15428
rect 47136 15388 48320 15416
rect 43496 15376 43502 15388
rect 48314 15376 48320 15388
rect 48372 15376 48378 15428
rect 49237 15419 49295 15425
rect 49237 15385 49249 15419
rect 49283 15416 49295 15419
rect 49421 15419 49479 15425
rect 49421 15416 49433 15419
rect 49283 15388 49433 15416
rect 49283 15385 49295 15388
rect 49237 15379 49295 15385
rect 49421 15385 49433 15388
rect 49467 15416 49479 15419
rect 50430 15416 50436 15428
rect 49467 15388 50436 15416
rect 49467 15385 49479 15388
rect 49421 15379 49479 15385
rect 50430 15376 50436 15388
rect 50488 15376 50494 15428
rect 39816 15320 42380 15348
rect 39816 15308 39822 15320
rect 43990 15308 43996 15360
rect 44048 15308 44054 15360
rect 44450 15308 44456 15360
rect 44508 15308 44514 15360
rect 46477 15351 46535 15357
rect 46477 15317 46489 15351
rect 46523 15348 46535 15351
rect 46842 15348 46848 15360
rect 46523 15320 46848 15348
rect 46523 15317 46535 15320
rect 46477 15311 46535 15317
rect 46842 15308 46848 15320
rect 46900 15308 46906 15360
rect 47762 15308 47768 15360
rect 47820 15308 47826 15360
rect 48590 15308 48596 15360
rect 48648 15348 48654 15360
rect 48869 15351 48927 15357
rect 48869 15348 48881 15351
rect 48648 15320 48881 15348
rect 48648 15308 48654 15320
rect 48869 15317 48881 15320
rect 48915 15317 48927 15351
rect 48869 15311 48927 15317
rect 49602 15308 49608 15360
rect 49660 15348 49666 15360
rect 49786 15348 49792 15360
rect 49660 15320 49792 15348
rect 49660 15308 49666 15320
rect 49786 15308 49792 15320
rect 49844 15308 49850 15360
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 3605 15147 3663 15153
rect 3605 15144 3617 15147
rect 2746 15116 3617 15144
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 2746 15008 2774 15116
rect 3605 15113 3617 15116
rect 3651 15113 3663 15147
rect 3605 15107 3663 15113
rect 7006 15104 7012 15156
rect 7064 15144 7070 15156
rect 7561 15147 7619 15153
rect 7561 15144 7573 15147
rect 7064 15116 7573 15144
rect 7064 15104 7070 15116
rect 7561 15113 7573 15116
rect 7607 15113 7619 15147
rect 7561 15107 7619 15113
rect 7742 15104 7748 15156
rect 7800 15144 7806 15156
rect 9493 15147 9551 15153
rect 9493 15144 9505 15147
rect 7800 15116 9505 15144
rect 7800 15104 7806 15116
rect 9493 15113 9505 15116
rect 9539 15113 9551 15147
rect 9493 15107 9551 15113
rect 9674 15104 9680 15156
rect 9732 15144 9738 15156
rect 10413 15147 10471 15153
rect 10413 15144 10425 15147
rect 9732 15116 10425 15144
rect 9732 15104 9738 15116
rect 10413 15113 10425 15116
rect 10459 15113 10471 15147
rect 10413 15107 10471 15113
rect 10781 15147 10839 15153
rect 10781 15113 10793 15147
rect 10827 15144 10839 15147
rect 11885 15147 11943 15153
rect 11885 15144 11897 15147
rect 10827 15116 11897 15144
rect 10827 15113 10839 15116
rect 10781 15107 10839 15113
rect 11885 15113 11897 15116
rect 11931 15113 11943 15147
rect 12894 15144 12900 15156
rect 11885 15107 11943 15113
rect 12084 15116 12900 15144
rect 3329 15079 3387 15085
rect 3329 15045 3341 15079
rect 3375 15076 3387 15079
rect 3418 15076 3424 15088
rect 3375 15048 3424 15076
rect 3375 15045 3387 15048
rect 3329 15039 3387 15045
rect 3418 15036 3424 15048
rect 3476 15036 3482 15088
rect 6730 15076 6736 15088
rect 3804 15048 6736 15076
rect 3804 15017 3832 15048
rect 6730 15036 6736 15048
rect 6788 15036 6794 15088
rect 7834 15036 7840 15088
rect 7892 15076 7898 15088
rect 8665 15079 8723 15085
rect 8665 15076 8677 15079
rect 7892 15048 8677 15076
rect 7892 15036 7898 15048
rect 8665 15045 8677 15048
rect 8711 15045 8723 15079
rect 8665 15039 8723 15045
rect 9122 15036 9128 15088
rect 9180 15076 9186 15088
rect 9585 15079 9643 15085
rect 9585 15076 9597 15079
rect 9180 15048 9597 15076
rect 9180 15036 9186 15048
rect 9585 15045 9597 15048
rect 9631 15045 9643 15079
rect 9585 15039 9643 15045
rect 10870 15036 10876 15088
rect 10928 15036 10934 15088
rect 1811 14980 2774 15008
rect 3789 15011 3847 15017
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 3789 14977 3801 15011
rect 3835 14977 3847 15011
rect 3789 14971 3847 14977
rect 4249 15011 4307 15017
rect 4249 14977 4261 15011
rect 4295 14977 4307 15011
rect 4249 14971 4307 14977
rect 5353 15011 5411 15017
rect 5353 14977 5365 15011
rect 5399 15008 5411 15011
rect 6822 15008 6828 15020
rect 5399 14980 6828 15008
rect 5399 14977 5411 14980
rect 5353 14971 5411 14977
rect 1302 14900 1308 14952
rect 1360 14940 1366 14952
rect 2041 14943 2099 14949
rect 2041 14940 2053 14943
rect 1360 14912 2053 14940
rect 1360 14900 1366 14912
rect 2041 14909 2053 14912
rect 2087 14909 2099 14943
rect 4264 14940 4292 14971
rect 6822 14968 6828 14980
rect 6880 14968 6886 15020
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 15008 6975 15011
rect 7926 15008 7932 15020
rect 6963 14980 7932 15008
rect 6963 14977 6975 14980
rect 6917 14971 6975 14977
rect 7926 14968 7932 14980
rect 7984 14968 7990 15020
rect 8018 14968 8024 15020
rect 8076 14968 8082 15020
rect 8478 14968 8484 15020
rect 8536 15008 8542 15020
rect 11698 15008 11704 15020
rect 8536 14980 11704 15008
rect 8536 14968 8542 14980
rect 11698 14968 11704 14980
rect 11756 14968 11762 15020
rect 6178 14940 6184 14952
rect 4264 14912 6184 14940
rect 2041 14903 2099 14909
rect 6178 14900 6184 14912
rect 6236 14900 6242 14952
rect 6457 14943 6515 14949
rect 6457 14909 6469 14943
rect 6503 14940 6515 14943
rect 9490 14940 9496 14952
rect 6503 14912 9496 14940
rect 6503 14909 6515 14912
rect 6457 14903 6515 14909
rect 9490 14900 9496 14912
rect 9548 14900 9554 14952
rect 9769 14943 9827 14949
rect 9769 14909 9781 14943
rect 9815 14940 9827 14943
rect 9858 14940 9864 14952
rect 9815 14912 9864 14940
rect 9815 14909 9827 14912
rect 9769 14903 9827 14909
rect 9858 14900 9864 14912
rect 9916 14900 9922 14952
rect 10318 14900 10324 14952
rect 10376 14940 10382 14952
rect 10965 14943 11023 14949
rect 10965 14940 10977 14943
rect 10376 14912 10977 14940
rect 10376 14900 10382 14912
rect 10965 14909 10977 14912
rect 11011 14909 11023 14943
rect 10965 14903 11023 14909
rect 4893 14875 4951 14881
rect 4893 14841 4905 14875
rect 4939 14872 4951 14875
rect 7098 14872 7104 14884
rect 4939 14844 7104 14872
rect 4939 14841 4951 14844
rect 4893 14835 4951 14841
rect 7098 14832 7104 14844
rect 7156 14832 7162 14884
rect 7558 14832 7564 14884
rect 7616 14872 7622 14884
rect 7742 14872 7748 14884
rect 7616 14844 7748 14872
rect 7616 14832 7622 14844
rect 7742 14832 7748 14844
rect 7800 14832 7806 14884
rect 7834 14832 7840 14884
rect 7892 14872 7898 14884
rect 12084 14872 12112 15116
rect 12894 15104 12900 15116
rect 12952 15104 12958 15156
rect 13262 15104 13268 15156
rect 13320 15144 13326 15156
rect 14734 15144 14740 15156
rect 13320 15116 14740 15144
rect 13320 15104 13326 15116
rect 14734 15104 14740 15116
rect 14792 15104 14798 15156
rect 16025 15147 16083 15153
rect 16025 15113 16037 15147
rect 16071 15144 16083 15147
rect 16390 15144 16396 15156
rect 16071 15116 16396 15144
rect 16071 15113 16083 15116
rect 16025 15107 16083 15113
rect 16390 15104 16396 15116
rect 16448 15104 16454 15156
rect 18233 15147 18291 15153
rect 18233 15113 18245 15147
rect 18279 15144 18291 15147
rect 18322 15144 18328 15156
rect 18279 15116 18328 15144
rect 18279 15113 18291 15116
rect 18233 15107 18291 15113
rect 18322 15104 18328 15116
rect 18380 15144 18386 15156
rect 18874 15144 18880 15156
rect 18380 15116 18880 15144
rect 18380 15104 18386 15116
rect 18874 15104 18880 15116
rect 18932 15104 18938 15156
rect 19429 15147 19487 15153
rect 19429 15113 19441 15147
rect 19475 15144 19487 15147
rect 19610 15144 19616 15156
rect 19475 15116 19616 15144
rect 19475 15113 19487 15116
rect 19429 15107 19487 15113
rect 19610 15104 19616 15116
rect 19668 15104 19674 15156
rect 19794 15104 19800 15156
rect 19852 15144 19858 15156
rect 20257 15147 20315 15153
rect 20257 15144 20269 15147
rect 19852 15116 20269 15144
rect 19852 15104 19858 15116
rect 20257 15113 20269 15116
rect 20303 15113 20315 15147
rect 20257 15107 20315 15113
rect 21450 15104 21456 15156
rect 21508 15104 21514 15156
rect 21637 15147 21695 15153
rect 21637 15113 21649 15147
rect 21683 15144 21695 15147
rect 21818 15144 21824 15156
rect 21683 15116 21824 15144
rect 21683 15113 21695 15116
rect 21637 15107 21695 15113
rect 21818 15104 21824 15116
rect 21876 15104 21882 15156
rect 22002 15104 22008 15156
rect 22060 15144 22066 15156
rect 23569 15147 23627 15153
rect 23569 15144 23581 15147
rect 22060 15116 23581 15144
rect 22060 15104 22066 15116
rect 23569 15113 23581 15116
rect 23615 15113 23627 15147
rect 23569 15107 23627 15113
rect 23750 15104 23756 15156
rect 23808 15144 23814 15156
rect 24121 15147 24179 15153
rect 24121 15144 24133 15147
rect 23808 15116 24133 15144
rect 23808 15104 23814 15116
rect 24121 15113 24133 15116
rect 24167 15113 24179 15147
rect 24121 15107 24179 15113
rect 25406 15104 25412 15156
rect 25464 15104 25470 15156
rect 27157 15147 27215 15153
rect 27157 15113 27169 15147
rect 27203 15144 27215 15147
rect 27246 15144 27252 15156
rect 27203 15116 27252 15144
rect 27203 15113 27215 15116
rect 27157 15107 27215 15113
rect 27246 15104 27252 15116
rect 27304 15104 27310 15156
rect 27525 15147 27583 15153
rect 27525 15144 27537 15147
rect 27356 15116 27537 15144
rect 12253 15079 12311 15085
rect 12253 15045 12265 15079
rect 12299 15076 12311 15079
rect 13998 15076 14004 15088
rect 12299 15048 14004 15076
rect 12299 15045 12311 15048
rect 12253 15039 12311 15045
rect 13998 15036 14004 15048
rect 14056 15036 14062 15088
rect 14553 15079 14611 15085
rect 14553 15076 14565 15079
rect 14108 15048 14565 15076
rect 12158 14968 12164 15020
rect 12216 15008 12222 15020
rect 12216 14980 12480 15008
rect 12216 14968 12222 14980
rect 12250 14900 12256 14952
rect 12308 14940 12314 14952
rect 12452 14949 12480 14980
rect 12526 14968 12532 15020
rect 12584 15008 12590 15020
rect 13449 15011 13507 15017
rect 13449 15008 13461 15011
rect 12584 14980 13461 15008
rect 12584 14968 12590 14980
rect 13449 14977 13461 14980
rect 13495 14977 13507 15011
rect 13449 14971 13507 14977
rect 13538 14968 13544 15020
rect 13596 14968 13602 15020
rect 12345 14943 12403 14949
rect 12345 14940 12357 14943
rect 12308 14912 12357 14940
rect 12308 14900 12314 14912
rect 12345 14909 12357 14912
rect 12391 14909 12403 14943
rect 12345 14903 12403 14909
rect 12437 14943 12495 14949
rect 12437 14909 12449 14943
rect 12483 14909 12495 14943
rect 13262 14940 13268 14952
rect 12437 14903 12495 14909
rect 12544 14912 13268 14940
rect 7892 14844 12112 14872
rect 7892 14832 7898 14844
rect 5994 14764 6000 14816
rect 6052 14764 6058 14816
rect 6641 14807 6699 14813
rect 6641 14773 6653 14807
rect 6687 14804 6699 14807
rect 8294 14804 8300 14816
rect 6687 14776 8300 14804
rect 6687 14773 6699 14776
rect 6641 14767 6699 14773
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 9125 14807 9183 14813
rect 9125 14773 9137 14807
rect 9171 14804 9183 14807
rect 9766 14804 9772 14816
rect 9171 14776 9772 14804
rect 9171 14773 9183 14776
rect 9125 14767 9183 14773
rect 9766 14764 9772 14776
rect 9824 14764 9830 14816
rect 9950 14764 9956 14816
rect 10008 14804 10014 14816
rect 11517 14807 11575 14813
rect 11517 14804 11529 14807
rect 10008 14776 11529 14804
rect 10008 14764 10014 14776
rect 11517 14773 11529 14776
rect 11563 14804 11575 14807
rect 12544 14804 12572 14912
rect 13262 14900 13268 14912
rect 13320 14900 13326 14952
rect 13725 14943 13783 14949
rect 13725 14909 13737 14943
rect 13771 14909 13783 14943
rect 13725 14903 13783 14909
rect 12802 14832 12808 14884
rect 12860 14872 12866 14884
rect 13740 14872 13768 14903
rect 13814 14900 13820 14952
rect 13872 14940 13878 14952
rect 14108 14940 14136 15048
rect 14553 15045 14565 15048
rect 14599 15045 14611 15079
rect 14553 15039 14611 15045
rect 16206 15036 16212 15088
rect 16264 15076 16270 15088
rect 17589 15079 17647 15085
rect 16264 15048 17540 15076
rect 16264 15036 16270 15048
rect 16022 15008 16028 15020
rect 15686 14980 16028 15008
rect 16022 14968 16028 14980
rect 16080 14968 16086 15020
rect 16390 14968 16396 15020
rect 16448 14968 16454 15020
rect 16666 14968 16672 15020
rect 16724 15008 16730 15020
rect 16945 15011 17003 15017
rect 16945 15008 16957 15011
rect 16724 14980 16957 15008
rect 16724 14968 16730 14980
rect 16945 14977 16957 14980
rect 16991 14977 17003 15011
rect 16945 14971 17003 14977
rect 17034 14968 17040 15020
rect 17092 15008 17098 15020
rect 17129 15011 17187 15017
rect 17129 15008 17141 15011
rect 17092 14980 17141 15008
rect 17092 14968 17098 14980
rect 17129 14977 17141 14980
rect 17175 14977 17187 15011
rect 17512 15008 17540 15048
rect 17589 15045 17601 15079
rect 17635 15076 17647 15079
rect 17770 15076 17776 15088
rect 17635 15048 17776 15076
rect 17635 15045 17647 15048
rect 17589 15039 17647 15045
rect 17770 15036 17776 15048
rect 17828 15076 17834 15088
rect 19518 15076 19524 15088
rect 17828 15048 19524 15076
rect 17828 15036 17834 15048
rect 19518 15036 19524 15048
rect 19576 15036 19582 15088
rect 20806 15076 20812 15088
rect 19628 15048 20812 15076
rect 18325 15011 18383 15017
rect 17512 14980 18092 15008
rect 17129 14971 17187 14977
rect 13872 14912 14136 14940
rect 13872 14900 13878 14912
rect 14274 14900 14280 14952
rect 14332 14900 14338 14952
rect 15838 14940 15844 14952
rect 14384 14912 15844 14940
rect 14384 14872 14412 14912
rect 15838 14900 15844 14912
rect 15896 14900 15902 14952
rect 16114 14900 16120 14952
rect 16172 14940 16178 14952
rect 18064 14940 18092 14980
rect 18325 14977 18337 15011
rect 18371 15008 18383 15011
rect 18506 15008 18512 15020
rect 18371 14980 18512 15008
rect 18371 14977 18383 14980
rect 18325 14971 18383 14977
rect 18506 14968 18512 14980
rect 18564 14968 18570 15020
rect 18690 14968 18696 15020
rect 18748 15008 18754 15020
rect 19628 15008 19656 15048
rect 20806 15036 20812 15048
rect 20864 15036 20870 15088
rect 22830 15036 22836 15088
rect 22888 15076 22894 15088
rect 25777 15079 25835 15085
rect 22888 15048 24808 15076
rect 22888 15036 22894 15048
rect 18748 14980 19656 15008
rect 18748 14968 18754 14980
rect 19794 14968 19800 15020
rect 19852 15008 19858 15020
rect 20162 15008 20168 15020
rect 19852 14980 20168 15008
rect 19852 14968 19858 14980
rect 20162 14968 20168 14980
rect 20220 14968 20226 15020
rect 20622 14968 20628 15020
rect 20680 14968 20686 15020
rect 21542 14968 21548 15020
rect 21600 15008 21606 15020
rect 22002 15008 22008 15020
rect 21600 14980 22008 15008
rect 21600 14968 21606 14980
rect 22002 14968 22008 14980
rect 22060 14968 22066 15020
rect 23293 15011 23351 15017
rect 23293 14977 23305 15011
rect 23339 15008 23351 15011
rect 23566 15008 23572 15020
rect 23339 14980 23572 15008
rect 23339 14977 23351 14980
rect 23293 14971 23351 14977
rect 23566 14968 23572 14980
rect 23624 14968 23630 15020
rect 23845 15011 23903 15017
rect 23845 15008 23857 15011
rect 23676 14980 23857 15008
rect 18417 14943 18475 14949
rect 18417 14940 18429 14943
rect 16172 14912 18000 14940
rect 18064 14912 18429 14940
rect 16172 14900 16178 14912
rect 17865 14875 17923 14881
rect 17865 14872 17877 14875
rect 12860 14844 14412 14872
rect 15580 14844 17877 14872
rect 12860 14832 12866 14844
rect 11563 14776 12572 14804
rect 11563 14773 11575 14776
rect 11517 14767 11575 14773
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 13081 14807 13139 14813
rect 13081 14804 13093 14807
rect 12676 14776 13093 14804
rect 12676 14764 12682 14776
rect 13081 14773 13093 14776
rect 13127 14773 13139 14807
rect 13081 14767 13139 14773
rect 13538 14764 13544 14816
rect 13596 14804 13602 14816
rect 15580 14804 15608 14844
rect 17865 14841 17877 14844
rect 17911 14841 17923 14875
rect 17972 14872 18000 14912
rect 18417 14909 18429 14912
rect 18463 14909 18475 14943
rect 18417 14903 18475 14909
rect 19518 14900 19524 14952
rect 19576 14900 19582 14952
rect 19613 14943 19671 14949
rect 19613 14909 19625 14943
rect 19659 14940 19671 14943
rect 19886 14940 19892 14952
rect 19659 14912 19892 14940
rect 19659 14909 19671 14912
rect 19613 14903 19671 14909
rect 19886 14900 19892 14912
rect 19944 14900 19950 14952
rect 20714 14900 20720 14952
rect 20772 14900 20778 14952
rect 20809 14943 20867 14949
rect 20809 14909 20821 14943
rect 20855 14909 20867 14943
rect 20809 14903 20867 14909
rect 17972 14844 19334 14872
rect 17865 14835 17923 14841
rect 13596 14776 15608 14804
rect 13596 14764 13602 14776
rect 15654 14764 15660 14816
rect 15712 14804 15718 14816
rect 18690 14804 18696 14816
rect 15712 14776 18696 14804
rect 15712 14764 15718 14776
rect 18690 14764 18696 14776
rect 18748 14764 18754 14816
rect 19058 14764 19064 14816
rect 19116 14764 19122 14816
rect 19306 14804 19334 14844
rect 19702 14832 19708 14884
rect 19760 14872 19766 14884
rect 20824 14872 20852 14903
rect 22462 14900 22468 14952
rect 22520 14940 22526 14952
rect 22741 14943 22799 14949
rect 22741 14940 22753 14943
rect 22520 14912 22753 14940
rect 22520 14900 22526 14912
rect 22741 14909 22753 14912
rect 22787 14909 22799 14943
rect 22741 14903 22799 14909
rect 23106 14900 23112 14952
rect 23164 14940 23170 14952
rect 23676 14940 23704 14980
rect 23845 14977 23857 14980
rect 23891 14977 23903 15011
rect 23845 14971 23903 14977
rect 24026 14968 24032 15020
rect 24084 15008 24090 15020
rect 24489 15011 24547 15017
rect 24489 15008 24501 15011
rect 24084 14980 24501 15008
rect 24084 14968 24090 14980
rect 24489 14977 24501 14980
rect 24535 14977 24547 15011
rect 24489 14971 24547 14977
rect 23164 14912 23704 14940
rect 23164 14900 23170 14912
rect 19760 14844 20852 14872
rect 19760 14832 19766 14844
rect 22186 14832 22192 14884
rect 22244 14872 22250 14884
rect 22244 14844 23520 14872
rect 22244 14832 22250 14844
rect 23492 14816 23520 14844
rect 23198 14804 23204 14816
rect 19306 14776 23204 14804
rect 23198 14764 23204 14776
rect 23256 14764 23262 14816
rect 23474 14764 23480 14816
rect 23532 14764 23538 14816
rect 23676 14804 23704 14912
rect 23750 14900 23756 14952
rect 23808 14940 23814 14952
rect 24581 14943 24639 14949
rect 24581 14940 24593 14943
rect 23808 14912 24593 14940
rect 23808 14900 23814 14912
rect 24581 14909 24593 14912
rect 24627 14909 24639 14943
rect 24581 14903 24639 14909
rect 24670 14900 24676 14952
rect 24728 14900 24734 14952
rect 24780 14872 24808 15048
rect 25777 15045 25789 15079
rect 25823 15076 25835 15079
rect 25866 15076 25872 15088
rect 25823 15048 25872 15076
rect 25823 15045 25835 15048
rect 25777 15039 25835 15045
rect 25866 15036 25872 15048
rect 25924 15036 25930 15088
rect 26970 15076 26976 15088
rect 25976 15048 26976 15076
rect 25976 15008 26004 15048
rect 26970 15036 26976 15048
rect 27028 15036 27034 15088
rect 27356 15076 27384 15116
rect 27525 15113 27537 15116
rect 27571 15113 27583 15147
rect 27525 15107 27583 15113
rect 27617 15147 27675 15153
rect 27617 15113 27629 15147
rect 27663 15144 27675 15147
rect 27982 15144 27988 15156
rect 27663 15116 27988 15144
rect 27663 15113 27675 15116
rect 27617 15107 27675 15113
rect 27982 15104 27988 15116
rect 28040 15104 28046 15156
rect 28442 15104 28448 15156
rect 28500 15144 28506 15156
rect 28718 15144 28724 15156
rect 28500 15116 28724 15144
rect 28500 15104 28506 15116
rect 28718 15104 28724 15116
rect 28776 15104 28782 15156
rect 28810 15104 28816 15156
rect 28868 15104 28874 15156
rect 28902 15104 28908 15156
rect 28960 15144 28966 15156
rect 29822 15144 29828 15156
rect 28960 15116 29828 15144
rect 28960 15104 28966 15116
rect 29822 15104 29828 15116
rect 29880 15104 29886 15156
rect 29917 15147 29975 15153
rect 29917 15113 29929 15147
rect 29963 15144 29975 15147
rect 32214 15144 32220 15156
rect 29963 15116 32220 15144
rect 29963 15113 29975 15116
rect 29917 15107 29975 15113
rect 32214 15104 32220 15116
rect 32272 15104 32278 15156
rect 32309 15147 32367 15153
rect 32309 15113 32321 15147
rect 32355 15113 32367 15147
rect 33226 15144 33232 15156
rect 32309 15107 32367 15113
rect 32416 15116 33232 15144
rect 27264 15048 27384 15076
rect 27264 15008 27292 15048
rect 27798 15036 27804 15088
rect 27856 15076 27862 15088
rect 27856 15048 29224 15076
rect 27856 15036 27862 15048
rect 28258 15008 28264 15020
rect 25884 14980 26004 15008
rect 26436 14980 27292 15008
rect 27356 14980 28264 15008
rect 24854 14900 24860 14952
rect 24912 14940 24918 14952
rect 25884 14949 25912 14980
rect 26436 14952 26464 14980
rect 25869 14943 25927 14949
rect 25869 14940 25881 14943
rect 24912 14912 25881 14940
rect 24912 14900 24918 14912
rect 25869 14909 25881 14912
rect 25915 14909 25927 14943
rect 25869 14903 25927 14909
rect 26053 14943 26111 14949
rect 26053 14909 26065 14943
rect 26099 14940 26111 14943
rect 26234 14940 26240 14952
rect 26099 14912 26240 14940
rect 26099 14909 26111 14912
rect 26053 14903 26111 14909
rect 26234 14900 26240 14912
rect 26292 14900 26298 14952
rect 26418 14900 26424 14952
rect 26476 14900 26482 14952
rect 26602 14900 26608 14952
rect 26660 14900 26666 14952
rect 27154 14900 27160 14952
rect 27212 14940 27218 14952
rect 27356 14940 27384 14980
rect 28258 14968 28264 14980
rect 28316 14968 28322 15020
rect 28718 14968 28724 15020
rect 28776 15008 28782 15020
rect 29086 15008 29092 15020
rect 28776 14980 29092 15008
rect 28776 14968 28782 14980
rect 29086 14968 29092 14980
rect 29144 14968 29150 15020
rect 27212 14912 27384 14940
rect 27801 14943 27859 14949
rect 27212 14900 27218 14912
rect 27801 14909 27813 14943
rect 27847 14940 27859 14943
rect 27890 14940 27896 14952
rect 27847 14912 27896 14940
rect 27847 14909 27859 14912
rect 27801 14903 27859 14909
rect 27890 14900 27896 14912
rect 27948 14900 27954 14952
rect 28905 14943 28963 14949
rect 28905 14940 28917 14943
rect 28828 14912 28917 14940
rect 28353 14875 28411 14881
rect 28353 14872 28365 14875
rect 24780 14844 28365 14872
rect 28353 14841 28365 14844
rect 28399 14841 28411 14875
rect 28353 14835 28411 14841
rect 28718 14832 28724 14884
rect 28776 14872 28782 14884
rect 28828 14872 28856 14912
rect 28905 14909 28917 14912
rect 28951 14909 28963 14943
rect 29196 14940 29224 15048
rect 29270 15036 29276 15088
rect 29328 15076 29334 15088
rect 29730 15076 29736 15088
rect 29328 15048 29736 15076
rect 29328 15036 29334 15048
rect 29730 15036 29736 15048
rect 29788 15036 29794 15088
rect 32324 15076 32352 15107
rect 29840 15048 32352 15076
rect 29840 14940 29868 15048
rect 30650 15008 30656 15020
rect 30208 14980 30656 15008
rect 30208 14949 30236 14980
rect 30650 14968 30656 14980
rect 30708 15008 30714 15020
rect 30834 15008 30840 15020
rect 30708 14980 30840 15008
rect 30708 14968 30714 14980
rect 30834 14968 30840 14980
rect 30892 14968 30898 15020
rect 31205 15011 31263 15017
rect 31205 14977 31217 15011
rect 31251 15008 31263 15011
rect 32416 15008 32444 15116
rect 33226 15104 33232 15116
rect 33284 15104 33290 15156
rect 33505 15147 33563 15153
rect 33505 15113 33517 15147
rect 33551 15144 33563 15147
rect 35253 15147 35311 15153
rect 35253 15144 35265 15147
rect 33551 15116 35265 15144
rect 33551 15113 33563 15116
rect 33505 15107 33563 15113
rect 35253 15113 35265 15116
rect 35299 15113 35311 15147
rect 35253 15107 35311 15113
rect 35342 15104 35348 15156
rect 35400 15104 35406 15156
rect 35986 15104 35992 15156
rect 36044 15144 36050 15156
rect 37366 15144 37372 15156
rect 36044 15116 37372 15144
rect 36044 15104 36050 15116
rect 37366 15104 37372 15116
rect 37424 15144 37430 15156
rect 37645 15147 37703 15153
rect 37645 15144 37657 15147
rect 37424 15116 37657 15144
rect 37424 15104 37430 15116
rect 37645 15113 37657 15116
rect 37691 15113 37703 15147
rect 40221 15147 40279 15153
rect 40221 15144 40233 15147
rect 37645 15107 37703 15113
rect 37752 15116 40233 15144
rect 32769 15079 32827 15085
rect 32769 15045 32781 15079
rect 32815 15076 32827 15079
rect 37752 15076 37780 15116
rect 40221 15113 40233 15116
rect 40267 15113 40279 15147
rect 40221 15107 40279 15113
rect 40862 15104 40868 15156
rect 40920 15144 40926 15156
rect 40920 15116 43944 15144
rect 40920 15104 40926 15116
rect 32815 15048 37780 15076
rect 32815 15045 32827 15048
rect 32769 15039 32827 15045
rect 37826 15036 37832 15088
rect 37884 15076 37890 15088
rect 38746 15076 38752 15088
rect 37884 15048 38752 15076
rect 37884 15036 37890 15048
rect 38746 15036 38752 15048
rect 38804 15036 38810 15088
rect 40589 15079 40647 15085
rect 40589 15045 40601 15079
rect 40635 15076 40647 15079
rect 40770 15076 40776 15088
rect 40635 15048 40776 15076
rect 40635 15045 40647 15048
rect 40589 15039 40647 15045
rect 40770 15036 40776 15048
rect 40828 15036 40834 15088
rect 42794 15076 42800 15088
rect 41432 15048 42800 15076
rect 31251 14980 32444 15008
rect 31251 14977 31263 14980
rect 31205 14971 31263 14977
rect 32490 14968 32496 15020
rect 32548 15008 32554 15020
rect 32677 15011 32735 15017
rect 32677 15008 32689 15011
rect 32548 14980 32689 15008
rect 32548 14968 32554 14980
rect 32677 14977 32689 14980
rect 32723 14977 32735 15011
rect 33410 15008 33416 15020
rect 32677 14971 32735 14977
rect 32784 14980 33416 15008
rect 29196 14912 29868 14940
rect 30009 14943 30067 14949
rect 28905 14903 28963 14909
rect 30009 14909 30021 14943
rect 30055 14909 30067 14943
rect 30009 14903 30067 14909
rect 30193 14943 30251 14949
rect 30193 14909 30205 14943
rect 30239 14909 30251 14943
rect 30193 14903 30251 14909
rect 30024 14872 30052 14903
rect 30374 14900 30380 14952
rect 30432 14940 30438 14952
rect 31297 14943 31355 14949
rect 31297 14940 31309 14943
rect 30432 14912 31309 14940
rect 30432 14900 30438 14912
rect 31297 14909 31309 14912
rect 31343 14909 31355 14943
rect 31297 14903 31355 14909
rect 31386 14900 31392 14952
rect 31444 14900 31450 14952
rect 32784 14940 32812 14980
rect 33410 14968 33416 14980
rect 33468 14968 33474 15020
rect 33686 14968 33692 15020
rect 33744 15008 33750 15020
rect 33873 15011 33931 15017
rect 33873 15008 33885 15011
rect 33744 14980 33885 15008
rect 33744 14968 33750 14980
rect 33873 14977 33885 14980
rect 33919 14977 33931 15011
rect 33873 14971 33931 14977
rect 33965 15011 34023 15017
rect 33965 14977 33977 15011
rect 34011 15008 34023 15011
rect 34882 15008 34888 15020
rect 34011 14980 34888 15008
rect 34011 14977 34023 14980
rect 33965 14971 34023 14977
rect 34882 14968 34888 14980
rect 34940 14968 34946 15020
rect 36446 14968 36452 15020
rect 36504 14968 36510 15020
rect 36541 15011 36599 15017
rect 36541 14977 36553 15011
rect 36587 15008 36599 15011
rect 37090 15008 37096 15020
rect 36587 14980 37096 15008
rect 36587 14977 36599 14980
rect 36541 14971 36599 14977
rect 37090 14968 37096 14980
rect 37148 14968 37154 15020
rect 37458 14968 37464 15020
rect 37516 15008 37522 15020
rect 38013 15011 38071 15017
rect 38013 15008 38025 15011
rect 37516 14980 38025 15008
rect 37516 14968 37522 14980
rect 38013 14977 38025 14980
rect 38059 14977 38071 15011
rect 38013 14971 38071 14977
rect 39942 14968 39948 15020
rect 40000 15008 40006 15020
rect 41432 15017 41460 15048
rect 42794 15036 42800 15048
rect 42852 15036 42858 15088
rect 41417 15011 41475 15017
rect 40000 14980 40816 15008
rect 40000 14968 40006 14980
rect 31726 14912 32812 14940
rect 32953 14943 33011 14949
rect 28776 14844 28856 14872
rect 29380 14844 30052 14872
rect 30837 14875 30895 14881
rect 28776 14832 28782 14844
rect 29380 14816 29408 14844
rect 30837 14841 30849 14875
rect 30883 14872 30895 14875
rect 31726 14872 31754 14912
rect 32953 14909 32965 14943
rect 32999 14940 33011 14943
rect 33502 14940 33508 14952
rect 32999 14912 33508 14940
rect 32999 14909 33011 14912
rect 32953 14903 33011 14909
rect 33502 14900 33508 14912
rect 33560 14900 33566 14952
rect 34149 14943 34207 14949
rect 34149 14909 34161 14943
rect 34195 14940 34207 14943
rect 34330 14940 34336 14952
rect 34195 14912 34336 14940
rect 34195 14909 34207 14912
rect 34149 14903 34207 14909
rect 34330 14900 34336 14912
rect 34388 14900 34394 14952
rect 35526 14900 35532 14952
rect 35584 14900 35590 14952
rect 35618 14900 35624 14952
rect 35676 14940 35682 14952
rect 36725 14943 36783 14949
rect 35676 14912 36676 14940
rect 35676 14900 35682 14912
rect 30883 14844 31754 14872
rect 30883 14841 30895 14844
rect 30837 14835 30895 14841
rect 32214 14832 32220 14884
rect 32272 14872 32278 14884
rect 36354 14872 36360 14884
rect 32272 14844 36360 14872
rect 32272 14832 32278 14844
rect 36354 14832 36360 14844
rect 36412 14832 36418 14884
rect 28442 14804 28448 14816
rect 23676 14776 28448 14804
rect 28442 14764 28448 14776
rect 28500 14764 28506 14816
rect 28534 14764 28540 14816
rect 28592 14804 28598 14816
rect 29086 14804 29092 14816
rect 28592 14776 29092 14804
rect 28592 14764 28598 14776
rect 29086 14764 29092 14776
rect 29144 14764 29150 14816
rect 29362 14764 29368 14816
rect 29420 14764 29426 14816
rect 29549 14807 29607 14813
rect 29549 14773 29561 14807
rect 29595 14804 29607 14807
rect 30650 14804 30656 14816
rect 29595 14776 30656 14804
rect 29595 14773 29607 14776
rect 29549 14767 29607 14773
rect 30650 14764 30656 14776
rect 30708 14764 30714 14816
rect 31570 14764 31576 14816
rect 31628 14804 31634 14816
rect 31941 14807 31999 14813
rect 31941 14804 31953 14807
rect 31628 14776 31953 14804
rect 31628 14764 31634 14776
rect 31941 14773 31953 14776
rect 31987 14804 31999 14807
rect 32858 14804 32864 14816
rect 31987 14776 32864 14804
rect 31987 14773 31999 14776
rect 31941 14767 31999 14773
rect 32858 14764 32864 14776
rect 32916 14764 32922 14816
rect 33226 14764 33232 14816
rect 33284 14804 33290 14816
rect 34330 14804 34336 14816
rect 33284 14776 34336 14804
rect 33284 14764 33290 14776
rect 34330 14764 34336 14776
rect 34388 14804 34394 14816
rect 34517 14807 34575 14813
rect 34517 14804 34529 14807
rect 34388 14776 34529 14804
rect 34388 14764 34394 14776
rect 34517 14773 34529 14776
rect 34563 14773 34575 14807
rect 34517 14767 34575 14773
rect 34885 14807 34943 14813
rect 34885 14773 34897 14807
rect 34931 14804 34943 14807
rect 35894 14804 35900 14816
rect 34931 14776 35900 14804
rect 34931 14773 34943 14776
rect 34885 14767 34943 14773
rect 35894 14764 35900 14776
rect 35952 14764 35958 14816
rect 36081 14807 36139 14813
rect 36081 14773 36093 14807
rect 36127 14804 36139 14807
rect 36262 14804 36268 14816
rect 36127 14776 36268 14804
rect 36127 14773 36139 14776
rect 36081 14767 36139 14773
rect 36262 14764 36268 14776
rect 36320 14764 36326 14816
rect 36648 14804 36676 14912
rect 36725 14909 36737 14943
rect 36771 14909 36783 14943
rect 36725 14903 36783 14909
rect 36740 14872 36768 14903
rect 36814 14900 36820 14952
rect 36872 14940 36878 14952
rect 37369 14943 37427 14949
rect 37369 14940 37381 14943
rect 36872 14912 37381 14940
rect 36872 14900 36878 14912
rect 37369 14909 37381 14912
rect 37415 14940 37427 14943
rect 37550 14940 37556 14952
rect 37415 14912 37556 14940
rect 37415 14909 37427 14912
rect 37369 14903 37427 14909
rect 37550 14900 37556 14912
rect 37608 14900 37614 14952
rect 38286 14900 38292 14952
rect 38344 14900 38350 14952
rect 38378 14900 38384 14952
rect 38436 14940 38442 14952
rect 40788 14949 40816 14980
rect 41417 14977 41429 15011
rect 41463 14977 41475 15011
rect 41417 14971 41475 14977
rect 42613 15011 42671 15017
rect 42613 14977 42625 15011
rect 42659 14977 42671 15011
rect 42613 14971 42671 14977
rect 43257 15011 43315 15017
rect 43257 14977 43269 15011
rect 43303 15008 43315 15011
rect 43717 15011 43775 15017
rect 43717 15008 43729 15011
rect 43303 14980 43729 15008
rect 43303 14977 43315 14980
rect 43257 14971 43315 14977
rect 43717 14977 43729 14980
rect 43763 14977 43775 15011
rect 43717 14971 43775 14977
rect 40681 14943 40739 14949
rect 40681 14940 40693 14943
rect 38436 14912 40693 14940
rect 38436 14900 38442 14912
rect 40681 14909 40693 14912
rect 40727 14909 40739 14943
rect 40681 14903 40739 14909
rect 40773 14943 40831 14949
rect 40773 14909 40785 14943
rect 40819 14909 40831 14943
rect 40773 14903 40831 14909
rect 36740 14844 38148 14872
rect 37553 14807 37611 14813
rect 37553 14804 37565 14807
rect 36648 14776 37565 14804
rect 37553 14773 37565 14776
rect 37599 14804 37611 14807
rect 37826 14804 37832 14816
rect 37599 14776 37832 14804
rect 37599 14773 37611 14776
rect 37553 14767 37611 14773
rect 37826 14764 37832 14776
rect 37884 14764 37890 14816
rect 38120 14804 38148 14844
rect 39298 14832 39304 14884
rect 39356 14872 39362 14884
rect 42628 14872 42656 14971
rect 43916 14940 43944 15116
rect 44818 15104 44824 15156
rect 44876 15144 44882 15156
rect 45833 15147 45891 15153
rect 45833 15144 45845 15147
rect 44876 15116 45845 15144
rect 44876 15104 44882 15116
rect 45833 15113 45845 15116
rect 45879 15113 45891 15147
rect 45833 15107 45891 15113
rect 47670 15104 47676 15156
rect 47728 15144 47734 15156
rect 47949 15147 48007 15153
rect 47949 15144 47961 15147
rect 47728 15116 47961 15144
rect 47728 15104 47734 15116
rect 47949 15113 47961 15116
rect 47995 15113 48007 15147
rect 47949 15107 48007 15113
rect 49234 15104 49240 15156
rect 49292 15104 49298 15156
rect 44358 15036 44364 15088
rect 44416 15076 44422 15088
rect 44634 15076 44640 15088
rect 44416 15048 44640 15076
rect 44416 15036 44422 15048
rect 44634 15036 44640 15048
rect 44692 15076 44698 15088
rect 44913 15079 44971 15085
rect 44913 15076 44925 15079
rect 44692 15048 44925 15076
rect 44692 15036 44698 15048
rect 44913 15045 44925 15048
rect 44959 15045 44971 15079
rect 48682 15076 48688 15088
rect 44913 15039 44971 15045
rect 46584 15048 48688 15076
rect 43990 14968 43996 15020
rect 44048 15008 44054 15020
rect 45189 15011 45247 15017
rect 45189 15008 45201 15011
rect 44048 14980 45201 15008
rect 44048 14968 44054 14980
rect 45189 14977 45201 14980
rect 45235 14977 45247 15011
rect 45189 14971 45247 14977
rect 45646 14968 45652 15020
rect 45704 15008 45710 15020
rect 45922 15008 45928 15020
rect 45704 14980 45928 15008
rect 45704 14968 45710 14980
rect 45922 14968 45928 14980
rect 45980 14968 45986 15020
rect 46584 15017 46612 15048
rect 48682 15036 48688 15048
rect 48740 15036 48746 15088
rect 46569 15011 46627 15017
rect 46569 14977 46581 15011
rect 46615 14977 46627 15011
rect 46569 14971 46627 14977
rect 47670 14968 47676 15020
rect 47728 15008 47734 15020
rect 47765 15011 47823 15017
rect 47765 15008 47777 15011
rect 47728 14980 47777 15008
rect 47728 14968 47734 14980
rect 47765 14977 47777 14980
rect 47811 15008 47823 15011
rect 47854 15008 47860 15020
rect 47811 14980 47860 15008
rect 47811 14977 47823 14980
rect 47765 14971 47823 14977
rect 47854 14968 47860 14980
rect 47912 14968 47918 15020
rect 48590 14968 48596 15020
rect 48648 14968 48654 15020
rect 47026 14940 47032 14952
rect 43916 14912 47032 14940
rect 47026 14900 47032 14912
rect 47084 14900 47090 14952
rect 46385 14875 46443 14881
rect 46385 14872 46397 14875
rect 39356 14844 42656 14872
rect 44100 14844 46397 14872
rect 39356 14832 39362 14844
rect 39758 14804 39764 14816
rect 38120 14776 39764 14804
rect 39758 14764 39764 14776
rect 39816 14764 39822 14816
rect 39850 14764 39856 14816
rect 39908 14804 39914 14816
rect 41966 14804 41972 14816
rect 39908 14776 41972 14804
rect 39908 14764 39914 14776
rect 41966 14764 41972 14776
rect 42024 14764 42030 14816
rect 42058 14764 42064 14816
rect 42116 14764 42122 14816
rect 42426 14764 42432 14816
rect 42484 14804 42490 14816
rect 44100 14804 44128 14844
rect 46385 14841 46397 14844
rect 46431 14872 46443 14875
rect 47213 14875 47271 14881
rect 47213 14872 47225 14875
rect 46431 14844 47225 14872
rect 46431 14841 46443 14844
rect 46385 14835 46443 14841
rect 47213 14841 47225 14844
rect 47259 14872 47271 14875
rect 47305 14875 47363 14881
rect 47305 14872 47317 14875
rect 47259 14844 47317 14872
rect 47259 14841 47271 14844
rect 47213 14835 47271 14841
rect 47305 14841 47317 14844
rect 47351 14841 47363 14875
rect 47305 14835 47363 14841
rect 42484 14776 44128 14804
rect 42484 14764 42490 14776
rect 44174 14764 44180 14816
rect 44232 14804 44238 14816
rect 44361 14807 44419 14813
rect 44361 14804 44373 14807
rect 44232 14776 44373 14804
rect 44232 14764 44238 14776
rect 44361 14773 44373 14776
rect 44407 14773 44419 14807
rect 44361 14767 44419 14773
rect 44729 14807 44787 14813
rect 44729 14773 44741 14807
rect 44775 14804 44787 14807
rect 45186 14804 45192 14816
rect 44775 14776 45192 14804
rect 44775 14773 44787 14776
rect 44729 14767 44787 14773
rect 45186 14764 45192 14776
rect 45244 14804 45250 14816
rect 45462 14804 45468 14816
rect 45244 14776 45468 14804
rect 45244 14764 45250 14776
rect 45462 14764 45468 14776
rect 45520 14764 45526 14816
rect 45646 14764 45652 14816
rect 45704 14804 45710 14816
rect 46109 14807 46167 14813
rect 46109 14804 46121 14807
rect 45704 14776 46121 14804
rect 45704 14764 45710 14776
rect 46109 14773 46121 14776
rect 46155 14773 46167 14807
rect 46109 14767 46167 14773
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 50908 14680 50936 15524
rect 1104 14640 49864 14662
rect 50890 14628 50896 14680
rect 50948 14628 50954 14680
rect 3510 14560 3516 14612
rect 3568 14560 3574 14612
rect 5718 14560 5724 14612
rect 5776 14600 5782 14612
rect 7469 14603 7527 14609
rect 7469 14600 7481 14603
rect 5776 14572 7481 14600
rect 5776 14560 5782 14572
rect 7469 14569 7481 14572
rect 7515 14569 7527 14603
rect 7469 14563 7527 14569
rect 7926 14560 7932 14612
rect 7984 14600 7990 14612
rect 8573 14603 8631 14609
rect 8573 14600 8585 14603
rect 7984 14572 8585 14600
rect 7984 14560 7990 14572
rect 8573 14569 8585 14572
rect 8619 14569 8631 14603
rect 8573 14563 8631 14569
rect 8662 14560 8668 14612
rect 8720 14600 8726 14612
rect 9398 14600 9404 14612
rect 8720 14572 9404 14600
rect 8720 14560 8726 14572
rect 9398 14560 9404 14572
rect 9456 14600 9462 14612
rect 9950 14600 9956 14612
rect 9456 14572 9956 14600
rect 9456 14560 9462 14572
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 10045 14603 10103 14609
rect 10045 14569 10057 14603
rect 10091 14600 10103 14603
rect 13814 14600 13820 14612
rect 10091 14572 13820 14600
rect 10091 14569 10103 14572
rect 10045 14563 10103 14569
rect 13814 14560 13820 14572
rect 13872 14560 13878 14612
rect 13906 14560 13912 14612
rect 13964 14560 13970 14612
rect 13998 14560 14004 14612
rect 14056 14600 14062 14612
rect 14550 14600 14556 14612
rect 14056 14572 14556 14600
rect 14056 14560 14062 14572
rect 14550 14560 14556 14572
rect 14608 14560 14614 14612
rect 14642 14560 14648 14612
rect 14700 14600 14706 14612
rect 16022 14600 16028 14612
rect 14700 14572 16028 14600
rect 14700 14560 14706 14572
rect 16022 14560 16028 14572
rect 16080 14560 16086 14612
rect 16761 14603 16819 14609
rect 16761 14569 16773 14603
rect 16807 14600 16819 14603
rect 16850 14600 16856 14612
rect 16807 14572 16856 14600
rect 16807 14569 16819 14572
rect 16761 14563 16819 14569
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 17678 14560 17684 14612
rect 17736 14600 17742 14612
rect 18141 14603 18199 14609
rect 18141 14600 18153 14603
rect 17736 14572 18153 14600
rect 17736 14560 17742 14572
rect 18141 14569 18153 14572
rect 18187 14569 18199 14603
rect 19613 14603 19671 14609
rect 19613 14600 19625 14603
rect 18141 14563 18199 14569
rect 18248 14572 19625 14600
rect 1946 14492 1952 14544
rect 2004 14532 2010 14544
rect 2222 14532 2228 14544
rect 2004 14504 2228 14532
rect 2004 14492 2010 14504
rect 2222 14492 2228 14504
rect 2280 14492 2286 14544
rect 3970 14492 3976 14544
rect 4028 14492 4034 14544
rect 5258 14492 5264 14544
rect 5316 14532 5322 14544
rect 6365 14535 6423 14541
rect 6365 14532 6377 14535
rect 5316 14504 6377 14532
rect 5316 14492 5322 14504
rect 6365 14501 6377 14504
rect 6411 14501 6423 14535
rect 6365 14495 6423 14501
rect 6730 14492 6736 14544
rect 6788 14532 6794 14544
rect 11146 14532 11152 14544
rect 6788 14504 11152 14532
rect 6788 14492 6794 14504
rect 11146 14492 11152 14504
rect 11204 14492 11210 14544
rect 17862 14492 17868 14544
rect 17920 14532 17926 14544
rect 18248 14532 18276 14572
rect 19613 14569 19625 14572
rect 19659 14569 19671 14603
rect 19613 14563 19671 14569
rect 19702 14560 19708 14612
rect 19760 14600 19766 14612
rect 23293 14603 23351 14609
rect 23293 14600 23305 14603
rect 19760 14572 23305 14600
rect 19760 14560 19766 14572
rect 23293 14569 23305 14572
rect 23339 14569 23351 14603
rect 25130 14600 25136 14612
rect 23293 14563 23351 14569
rect 23400 14572 25136 14600
rect 17920 14504 18276 14532
rect 17920 14492 17926 14504
rect 18690 14492 18696 14544
rect 18748 14532 18754 14544
rect 18874 14532 18880 14544
rect 18748 14504 18880 14532
rect 18748 14492 18754 14504
rect 18874 14492 18880 14504
rect 18932 14492 18938 14544
rect 19242 14492 19248 14544
rect 19300 14532 19306 14544
rect 19300 14504 20208 14532
rect 19300 14492 19306 14504
rect 1302 14424 1308 14476
rect 1360 14464 1366 14476
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1360 14436 2053 14464
rect 1360 14424 1366 14436
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 7006 14464 7012 14476
rect 2041 14427 2099 14433
rect 4172 14436 7012 14464
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 1946 14396 1952 14408
rect 1811 14368 1952 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 1946 14356 1952 14368
rect 2004 14356 2010 14408
rect 4172 14405 4200 14436
rect 7006 14424 7012 14436
rect 7064 14424 7070 14476
rect 7558 14424 7564 14476
rect 7616 14464 7622 14476
rect 11238 14464 11244 14476
rect 7616 14436 11244 14464
rect 7616 14424 7622 14436
rect 11238 14424 11244 14436
rect 11296 14424 11302 14476
rect 12434 14424 12440 14476
rect 12492 14464 12498 14476
rect 14642 14464 14648 14476
rect 12492 14436 14648 14464
rect 12492 14424 12498 14436
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14396 3479 14399
rect 4157 14399 4215 14405
rect 4157 14396 4169 14399
rect 3467 14368 4169 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 4157 14365 4169 14368
rect 4203 14365 4215 14399
rect 4157 14359 4215 14365
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14396 4675 14399
rect 4890 14396 4896 14408
rect 4663 14368 4896 14396
rect 4663 14365 4675 14368
rect 4617 14359 4675 14365
rect 4890 14356 4896 14368
rect 4948 14356 4954 14408
rect 5721 14399 5779 14405
rect 5721 14365 5733 14399
rect 5767 14396 5779 14399
rect 5994 14396 6000 14408
rect 5767 14368 6000 14396
rect 5767 14365 5779 14368
rect 5721 14359 5779 14365
rect 5994 14356 6000 14368
rect 6052 14356 6058 14408
rect 6813 14399 6871 14405
rect 6813 14396 6825 14399
rect 6748 14368 6825 14396
rect 4798 14288 4804 14340
rect 4856 14328 4862 14340
rect 5261 14331 5319 14337
rect 5261 14328 5273 14331
rect 4856 14300 5273 14328
rect 4856 14288 4862 14300
rect 5261 14297 5273 14300
rect 5307 14297 5319 14331
rect 6748 14328 6776 14368
rect 6813 14365 6825 14368
rect 6859 14365 6871 14399
rect 6813 14359 6871 14365
rect 7929 14399 7987 14405
rect 7929 14365 7941 14399
rect 7975 14396 7987 14399
rect 8754 14396 8760 14408
rect 7975 14368 8760 14396
rect 7975 14365 7987 14368
rect 7929 14359 7987 14365
rect 8754 14356 8760 14368
rect 8812 14396 8818 14408
rect 8938 14396 8944 14408
rect 8812 14368 8944 14396
rect 8812 14356 8818 14368
rect 8938 14356 8944 14368
rect 8996 14356 9002 14408
rect 9401 14399 9459 14405
rect 9401 14365 9413 14399
rect 9447 14396 9459 14399
rect 10042 14396 10048 14408
rect 9447 14368 10048 14396
rect 9447 14365 9459 14368
rect 9401 14359 9459 14365
rect 10042 14356 10048 14368
rect 10100 14356 10106 14408
rect 10502 14356 10508 14408
rect 10560 14356 10566 14408
rect 10778 14356 10784 14408
rect 10836 14396 10842 14408
rect 11609 14399 11667 14405
rect 11609 14396 11621 14399
rect 10836 14368 11621 14396
rect 10836 14356 10842 14368
rect 11609 14365 11621 14368
rect 11655 14365 11667 14399
rect 13004 14382 13032 14436
rect 14642 14424 14648 14436
rect 14700 14424 14706 14476
rect 14826 14424 14832 14476
rect 14884 14424 14890 14476
rect 16117 14467 16175 14473
rect 16117 14433 16129 14467
rect 16163 14433 16175 14467
rect 16117 14427 16175 14433
rect 11609 14359 11667 14365
rect 13354 14356 13360 14408
rect 13412 14396 13418 14408
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 13412 14368 15853 14396
rect 13412 14356 13418 14368
rect 15841 14365 15853 14368
rect 15887 14365 15899 14399
rect 16132 14396 16160 14427
rect 16758 14424 16764 14476
rect 16816 14464 16822 14476
rect 17681 14467 17739 14473
rect 17681 14464 17693 14467
rect 16816 14436 17693 14464
rect 16816 14424 16822 14436
rect 17681 14433 17693 14436
rect 17727 14433 17739 14467
rect 17681 14427 17739 14433
rect 18782 14424 18788 14476
rect 18840 14424 18846 14476
rect 20180 14473 20208 14504
rect 20165 14467 20223 14473
rect 20165 14433 20177 14467
rect 20211 14464 20223 14467
rect 21450 14464 21456 14476
rect 20211 14436 21456 14464
rect 20211 14433 20223 14436
rect 20165 14427 20223 14433
rect 21450 14424 21456 14436
rect 21508 14424 21514 14476
rect 21818 14424 21824 14476
rect 21876 14464 21882 14476
rect 22833 14467 22891 14473
rect 22833 14464 22845 14467
rect 21876 14436 22845 14464
rect 21876 14424 21882 14436
rect 22833 14433 22845 14436
rect 22879 14464 22891 14467
rect 23400 14464 23428 14572
rect 25130 14560 25136 14572
rect 25188 14560 25194 14612
rect 25501 14603 25559 14609
rect 25501 14569 25513 14603
rect 25547 14600 25559 14603
rect 27706 14600 27712 14612
rect 25547 14572 27712 14600
rect 25547 14569 25559 14572
rect 25501 14563 25559 14569
rect 27706 14560 27712 14572
rect 27764 14560 27770 14612
rect 27890 14560 27896 14612
rect 27948 14600 27954 14612
rect 27985 14603 28043 14609
rect 27985 14600 27997 14603
rect 27948 14572 27997 14600
rect 27948 14560 27954 14572
rect 27985 14569 27997 14572
rect 28031 14569 28043 14603
rect 27985 14563 28043 14569
rect 28258 14560 28264 14612
rect 28316 14560 28322 14612
rect 28445 14603 28503 14609
rect 28445 14569 28457 14603
rect 28491 14600 28503 14603
rect 33137 14603 33195 14609
rect 28491 14572 32904 14600
rect 28491 14569 28503 14572
rect 28445 14563 28503 14569
rect 24302 14492 24308 14544
rect 24360 14532 24366 14544
rect 24489 14535 24547 14541
rect 24489 14532 24501 14535
rect 24360 14504 24501 14532
rect 24360 14492 24366 14504
rect 24489 14501 24501 14504
rect 24535 14532 24547 14535
rect 24762 14532 24768 14544
rect 24535 14504 24768 14532
rect 24535 14501 24547 14504
rect 24489 14495 24547 14501
rect 24762 14492 24768 14504
rect 24820 14492 24826 14544
rect 28074 14492 28080 14544
rect 28132 14532 28138 14544
rect 29546 14532 29552 14544
rect 28132 14504 29552 14532
rect 28132 14492 28138 14504
rect 29546 14492 29552 14504
rect 29604 14492 29610 14544
rect 31481 14535 31539 14541
rect 31481 14501 31493 14535
rect 31527 14532 31539 14535
rect 31570 14532 31576 14544
rect 31527 14504 31576 14532
rect 31527 14501 31539 14504
rect 31481 14495 31539 14501
rect 31570 14492 31576 14504
rect 31628 14532 31634 14544
rect 32214 14532 32220 14544
rect 31628 14504 32220 14532
rect 31628 14492 31634 14504
rect 32214 14492 32220 14504
rect 32272 14492 32278 14544
rect 32306 14492 32312 14544
rect 32364 14532 32370 14544
rect 32876 14532 32904 14572
rect 33137 14569 33149 14603
rect 33183 14600 33195 14603
rect 33318 14600 33324 14612
rect 33183 14572 33324 14600
rect 33183 14569 33195 14572
rect 33137 14563 33195 14569
rect 33318 14560 33324 14572
rect 33376 14560 33382 14612
rect 33962 14600 33968 14612
rect 33428 14572 33968 14600
rect 33428 14532 33456 14572
rect 33962 14560 33968 14572
rect 34020 14560 34026 14612
rect 35148 14603 35206 14609
rect 35148 14569 35160 14603
rect 35194 14600 35206 14603
rect 42058 14600 42064 14612
rect 35194 14572 42064 14600
rect 35194 14569 35206 14572
rect 35148 14563 35206 14569
rect 42058 14560 42064 14572
rect 42116 14560 42122 14612
rect 42794 14560 42800 14612
rect 42852 14600 42858 14612
rect 45833 14603 45891 14609
rect 45833 14600 45845 14603
rect 42852 14572 45845 14600
rect 42852 14560 42858 14572
rect 45833 14569 45845 14572
rect 45879 14569 45891 14603
rect 45833 14563 45891 14569
rect 46937 14603 46995 14609
rect 46937 14569 46949 14603
rect 46983 14600 46995 14603
rect 47486 14600 47492 14612
rect 46983 14572 47492 14600
rect 46983 14569 46995 14572
rect 46937 14563 46995 14569
rect 47486 14560 47492 14572
rect 47544 14560 47550 14612
rect 49326 14560 49332 14612
rect 49384 14560 49390 14612
rect 32364 14504 32444 14532
rect 32876 14504 33456 14532
rect 32364 14492 32370 14504
rect 22879 14436 23428 14464
rect 23937 14467 23995 14473
rect 22879 14433 22891 14436
rect 22833 14427 22891 14433
rect 23937 14433 23949 14467
rect 23983 14464 23995 14467
rect 24578 14464 24584 14476
rect 23983 14436 24584 14464
rect 23983 14433 23995 14436
rect 23937 14427 23995 14433
rect 24578 14424 24584 14436
rect 24636 14424 24642 14476
rect 26237 14467 26295 14473
rect 26237 14433 26249 14467
rect 26283 14464 26295 14467
rect 28718 14464 28724 14476
rect 26283 14436 28724 14464
rect 26283 14433 26295 14436
rect 26237 14427 26295 14433
rect 28718 14424 28724 14436
rect 28776 14424 28782 14476
rect 29089 14467 29147 14473
rect 29089 14433 29101 14467
rect 29135 14464 29147 14467
rect 29638 14464 29644 14476
rect 29135 14436 29644 14464
rect 29135 14433 29147 14436
rect 29089 14427 29147 14433
rect 29638 14424 29644 14436
rect 29696 14424 29702 14476
rect 29733 14467 29791 14473
rect 29733 14433 29745 14467
rect 29779 14464 29791 14467
rect 30098 14464 30104 14476
rect 29779 14436 30104 14464
rect 29779 14433 29791 14436
rect 29733 14427 29791 14433
rect 16206 14396 16212 14408
rect 16132 14368 16212 14396
rect 15841 14359 15899 14365
rect 6748 14300 11836 14328
rect 5261 14291 5319 14297
rect 1762 14220 1768 14272
rect 1820 14260 1826 14272
rect 7558 14260 7564 14272
rect 1820 14232 7564 14260
rect 1820 14220 1826 14232
rect 7558 14220 7564 14232
rect 7616 14220 7622 14272
rect 8294 14220 8300 14272
rect 8352 14260 8358 14272
rect 9033 14263 9091 14269
rect 9033 14260 9045 14263
rect 8352 14232 9045 14260
rect 8352 14220 8358 14232
rect 9033 14229 9045 14232
rect 9079 14229 9091 14263
rect 9033 14223 9091 14229
rect 11149 14263 11207 14269
rect 11149 14229 11161 14263
rect 11195 14260 11207 14263
rect 11698 14260 11704 14272
rect 11195 14232 11704 14260
rect 11195 14229 11207 14232
rect 11149 14223 11207 14229
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 11808 14260 11836 14300
rect 11882 14288 11888 14340
rect 11940 14288 11946 14340
rect 13998 14288 14004 14340
rect 14056 14328 14062 14340
rect 14737 14331 14795 14337
rect 14737 14328 14749 14331
rect 14056 14300 14749 14328
rect 14056 14288 14062 14300
rect 14737 14297 14749 14300
rect 14783 14297 14795 14331
rect 14737 14291 14795 14297
rect 15286 14288 15292 14340
rect 15344 14328 15350 14340
rect 15856 14328 15884 14359
rect 16206 14356 16212 14368
rect 16264 14396 16270 14408
rect 16850 14396 16856 14408
rect 16264 14368 16856 14396
rect 16264 14356 16270 14368
rect 16850 14356 16856 14368
rect 16908 14356 16914 14408
rect 17034 14356 17040 14408
rect 17092 14396 17098 14408
rect 20530 14396 20536 14408
rect 17092 14368 20536 14396
rect 17092 14356 17098 14368
rect 20530 14356 20536 14368
rect 20588 14356 20594 14408
rect 20806 14356 20812 14408
rect 20864 14356 20870 14408
rect 22186 14356 22192 14408
rect 22244 14356 22250 14408
rect 23753 14399 23811 14405
rect 23753 14365 23765 14399
rect 23799 14396 23811 14399
rect 24486 14396 24492 14408
rect 23799 14368 24492 14396
rect 23799 14365 23811 14368
rect 23753 14359 23811 14365
rect 24486 14356 24492 14368
rect 24544 14356 24550 14408
rect 24857 14399 24915 14405
rect 24857 14365 24869 14399
rect 24903 14396 24915 14399
rect 25590 14396 25596 14408
rect 24903 14368 25596 14396
rect 24903 14365 24915 14368
rect 24857 14359 24915 14365
rect 25590 14356 25596 14368
rect 25648 14396 25654 14408
rect 25774 14396 25780 14408
rect 25648 14368 25780 14396
rect 25648 14356 25654 14368
rect 25774 14356 25780 14368
rect 25832 14356 25838 14408
rect 25958 14356 25964 14408
rect 26016 14356 26022 14408
rect 27338 14356 27344 14408
rect 27396 14356 27402 14408
rect 29362 14356 29368 14408
rect 29420 14396 29426 14408
rect 29748 14396 29776 14427
rect 30098 14424 30104 14436
rect 30156 14424 30162 14476
rect 30650 14424 30656 14476
rect 30708 14464 30714 14476
rect 32416 14473 32444 14504
rect 38378 14492 38384 14544
rect 38436 14532 38442 14544
rect 38841 14535 38899 14541
rect 38436 14504 38654 14532
rect 38436 14492 38442 14504
rect 32401 14467 32459 14473
rect 30708 14436 32352 14464
rect 30708 14424 30714 14436
rect 32324 14405 32352 14436
rect 32401 14433 32413 14467
rect 32447 14433 32459 14467
rect 32401 14427 32459 14433
rect 32582 14424 32588 14476
rect 32640 14424 32646 14476
rect 32766 14424 32772 14476
rect 32824 14464 32830 14476
rect 33689 14467 33747 14473
rect 33689 14464 33701 14467
rect 32824 14436 33701 14464
rect 32824 14424 32830 14436
rect 33689 14433 33701 14436
rect 33735 14464 33747 14467
rect 34149 14467 34207 14473
rect 34149 14464 34161 14467
rect 33735 14436 34161 14464
rect 33735 14433 33747 14436
rect 33689 14427 33747 14433
rect 34149 14433 34161 14436
rect 34195 14433 34207 14467
rect 34149 14427 34207 14433
rect 35710 14424 35716 14476
rect 35768 14464 35774 14476
rect 36633 14467 36691 14473
rect 36633 14464 36645 14467
rect 35768 14436 36645 14464
rect 35768 14424 35774 14436
rect 36633 14433 36645 14436
rect 36679 14433 36691 14467
rect 36633 14427 36691 14433
rect 29420 14368 29776 14396
rect 32309 14399 32367 14405
rect 29420 14356 29426 14368
rect 32309 14365 32321 14399
rect 32355 14365 32367 14399
rect 32309 14359 32367 14365
rect 33597 14399 33655 14405
rect 33597 14365 33609 14399
rect 33643 14396 33655 14399
rect 33778 14396 33784 14408
rect 33643 14368 33784 14396
rect 33643 14365 33655 14368
rect 33597 14359 33655 14365
rect 33778 14356 33784 14368
rect 33836 14356 33842 14408
rect 34054 14356 34060 14408
rect 34112 14396 34118 14408
rect 34885 14399 34943 14405
rect 34885 14396 34897 14399
rect 34112 14368 34897 14396
rect 34112 14356 34118 14368
rect 34885 14365 34897 14368
rect 34931 14365 34943 14399
rect 34885 14359 34943 14365
rect 16758 14328 16764 14340
rect 15344 14300 15608 14328
rect 15856 14300 16764 14328
rect 15344 14288 15350 14300
rect 13357 14263 13415 14269
rect 13357 14260 13369 14263
rect 11808 14232 13369 14260
rect 13357 14229 13369 14232
rect 13403 14260 13415 14263
rect 13630 14260 13636 14272
rect 13403 14232 13636 14260
rect 13403 14229 13415 14232
rect 13357 14223 13415 14229
rect 13630 14220 13636 14232
rect 13688 14220 13694 14272
rect 13906 14220 13912 14272
rect 13964 14260 13970 14272
rect 14277 14263 14335 14269
rect 14277 14260 14289 14263
rect 13964 14232 14289 14260
rect 13964 14220 13970 14232
rect 14277 14229 14289 14232
rect 14323 14229 14335 14263
rect 14277 14223 14335 14229
rect 14642 14220 14648 14272
rect 14700 14220 14706 14272
rect 15470 14220 15476 14272
rect 15528 14220 15534 14272
rect 15580 14260 15608 14300
rect 16758 14288 16764 14300
rect 16816 14288 16822 14340
rect 17678 14288 17684 14340
rect 17736 14328 17742 14340
rect 18509 14331 18567 14337
rect 18509 14328 18521 14331
rect 17736 14300 18521 14328
rect 17736 14288 17742 14300
rect 18509 14297 18521 14300
rect 18555 14297 18567 14331
rect 18509 14291 18567 14297
rect 21082 14288 21088 14340
rect 21140 14288 21146 14340
rect 23661 14331 23719 14337
rect 23661 14297 23673 14331
rect 23707 14328 23719 14331
rect 25222 14328 25228 14340
rect 23707 14300 25228 14328
rect 23707 14297 23719 14300
rect 23661 14291 23719 14297
rect 25222 14288 25228 14300
rect 25280 14288 25286 14340
rect 28813 14331 28871 14337
rect 28813 14297 28825 14331
rect 28859 14328 28871 14331
rect 29546 14328 29552 14340
rect 28859 14300 29552 14328
rect 28859 14297 28871 14300
rect 28813 14291 28871 14297
rect 29546 14288 29552 14300
rect 29604 14288 29610 14340
rect 30006 14288 30012 14340
rect 30064 14288 30070 14340
rect 31478 14328 31484 14340
rect 31234 14300 31484 14328
rect 15746 14260 15752 14272
rect 15580 14232 15752 14260
rect 15746 14220 15752 14232
rect 15804 14260 15810 14272
rect 15933 14263 15991 14269
rect 15933 14260 15945 14263
rect 15804 14232 15945 14260
rect 15804 14220 15810 14232
rect 15933 14229 15945 14232
rect 15979 14229 15991 14263
rect 15933 14223 15991 14229
rect 16577 14263 16635 14269
rect 16577 14229 16589 14263
rect 16623 14260 16635 14263
rect 17586 14260 17592 14272
rect 16623 14232 17592 14260
rect 16623 14229 16635 14232
rect 16577 14223 16635 14229
rect 17586 14220 17592 14232
rect 17644 14260 17650 14272
rect 18414 14260 18420 14272
rect 17644 14232 18420 14260
rect 17644 14220 17650 14232
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 18601 14263 18659 14269
rect 18601 14229 18613 14263
rect 18647 14260 18659 14263
rect 18874 14260 18880 14272
rect 18647 14232 18880 14260
rect 18647 14229 18659 14232
rect 18601 14223 18659 14229
rect 18874 14220 18880 14232
rect 18932 14220 18938 14272
rect 19337 14263 19395 14269
rect 19337 14229 19349 14263
rect 19383 14260 19395 14263
rect 19518 14260 19524 14272
rect 19383 14232 19524 14260
rect 19383 14229 19395 14232
rect 19337 14223 19395 14229
rect 19518 14220 19524 14232
rect 19576 14220 19582 14272
rect 19978 14220 19984 14272
rect 20036 14220 20042 14272
rect 20073 14263 20131 14269
rect 20073 14229 20085 14263
rect 20119 14260 20131 14263
rect 22554 14260 22560 14272
rect 20119 14232 22560 14260
rect 20119 14229 20131 14232
rect 20073 14223 20131 14229
rect 22554 14220 22560 14232
rect 22612 14220 22618 14272
rect 25774 14220 25780 14272
rect 25832 14260 25838 14272
rect 26510 14260 26516 14272
rect 25832 14232 26516 14260
rect 25832 14220 25838 14232
rect 26510 14220 26516 14232
rect 26568 14220 26574 14272
rect 27706 14220 27712 14272
rect 27764 14220 27770 14272
rect 28258 14220 28264 14272
rect 28316 14260 28322 14272
rect 28902 14260 28908 14272
rect 28316 14232 28908 14260
rect 28316 14220 28322 14232
rect 28902 14220 28908 14232
rect 28960 14220 28966 14272
rect 30742 14220 30748 14272
rect 30800 14260 30806 14272
rect 31312 14260 31340 14300
rect 31478 14288 31484 14300
rect 31536 14328 31542 14340
rect 32674 14328 32680 14340
rect 31536 14300 32680 14328
rect 31536 14288 31542 14300
rect 32674 14288 32680 14300
rect 32732 14288 32738 14340
rect 34790 14328 34796 14340
rect 33428 14300 34796 14328
rect 30800 14232 31340 14260
rect 31941 14263 31999 14269
rect 30800 14220 30806 14232
rect 31941 14229 31953 14263
rect 31987 14260 31999 14263
rect 33428 14260 33456 14300
rect 34790 14288 34796 14300
rect 34848 14288 34854 14340
rect 35618 14288 35624 14340
rect 35676 14288 35682 14340
rect 31987 14232 33456 14260
rect 33505 14263 33563 14269
rect 31987 14229 31999 14232
rect 31941 14223 31999 14229
rect 33505 14229 33517 14263
rect 33551 14260 33563 14263
rect 34330 14260 34336 14272
rect 33551 14232 34336 14260
rect 33551 14229 33563 14232
rect 33505 14223 33563 14229
rect 34330 14220 34336 14232
rect 34388 14220 34394 14272
rect 34517 14263 34575 14269
rect 34517 14229 34529 14263
rect 34563 14260 34575 14263
rect 34606 14260 34612 14272
rect 34563 14232 34612 14260
rect 34563 14229 34575 14232
rect 34517 14223 34575 14229
rect 34606 14220 34612 14232
rect 34664 14220 34670 14272
rect 36648 14260 36676 14427
rect 36814 14424 36820 14476
rect 36872 14464 36878 14476
rect 37093 14467 37151 14473
rect 37093 14464 37105 14467
rect 36872 14436 37105 14464
rect 36872 14424 36878 14436
rect 37093 14433 37105 14436
rect 37139 14464 37151 14467
rect 37458 14464 37464 14476
rect 37139 14436 37464 14464
rect 37139 14433 37151 14436
rect 37093 14427 37151 14433
rect 37458 14424 37464 14436
rect 37516 14424 37522 14476
rect 38626 14464 38654 14504
rect 38841 14501 38853 14535
rect 38887 14532 38899 14535
rect 39206 14532 39212 14544
rect 38887 14504 39212 14532
rect 38887 14501 38899 14504
rect 38841 14495 38899 14501
rect 39206 14492 39212 14504
rect 39264 14492 39270 14544
rect 39298 14492 39304 14544
rect 39356 14492 39362 14544
rect 39390 14492 39396 14544
rect 39448 14532 39454 14544
rect 39850 14532 39856 14544
rect 39448 14504 39856 14532
rect 39448 14492 39454 14504
rect 39850 14492 39856 14504
rect 39908 14492 39914 14544
rect 40218 14492 40224 14544
rect 40276 14532 40282 14544
rect 43993 14535 44051 14541
rect 43993 14532 44005 14535
rect 40276 14504 44005 14532
rect 40276 14492 40282 14504
rect 43993 14501 44005 14504
rect 44039 14501 44051 14535
rect 43993 14495 44051 14501
rect 44082 14492 44088 14544
rect 44140 14532 44146 14544
rect 48041 14535 48099 14541
rect 48041 14532 48053 14535
rect 44140 14504 48053 14532
rect 44140 14492 44146 14504
rect 48041 14501 48053 14504
rect 48087 14501 48099 14535
rect 48041 14495 48099 14501
rect 39758 14464 39764 14476
rect 38626 14436 39764 14464
rect 39758 14424 39764 14436
rect 39816 14424 39822 14476
rect 41785 14467 41843 14473
rect 41785 14464 41797 14467
rect 40052 14436 41797 14464
rect 38838 14396 38844 14408
rect 38764 14368 38844 14396
rect 37366 14288 37372 14340
rect 37424 14288 37430 14340
rect 38764 14328 38792 14368
rect 38838 14356 38844 14368
rect 38896 14356 38902 14408
rect 38930 14356 38936 14408
rect 38988 14396 38994 14408
rect 40052 14405 40080 14436
rect 41785 14433 41797 14436
rect 41831 14433 41843 14467
rect 41785 14427 41843 14433
rect 43162 14424 43168 14476
rect 43220 14464 43226 14476
rect 44269 14467 44327 14473
rect 44269 14464 44281 14467
rect 43220 14436 44281 14464
rect 43220 14424 43226 14436
rect 44269 14433 44281 14436
rect 44315 14464 44327 14467
rect 44453 14467 44511 14473
rect 44453 14464 44465 14467
rect 44315 14436 44465 14464
rect 44315 14433 44327 14436
rect 44269 14427 44327 14433
rect 44453 14433 44465 14436
rect 44499 14433 44511 14467
rect 48317 14467 48375 14473
rect 48317 14464 48329 14467
rect 44453 14427 44511 14433
rect 46308 14436 48329 14464
rect 39485 14399 39543 14405
rect 39485 14396 39497 14399
rect 38988 14368 39497 14396
rect 38988 14356 38994 14368
rect 39485 14365 39497 14368
rect 39531 14365 39543 14399
rect 39485 14359 39543 14365
rect 40037 14399 40095 14405
rect 40037 14365 40049 14399
rect 40083 14365 40095 14399
rect 40037 14359 40095 14365
rect 41141 14399 41199 14405
rect 41141 14365 41153 14399
rect 41187 14396 41199 14399
rect 41506 14396 41512 14408
rect 41187 14368 41512 14396
rect 41187 14365 41199 14368
rect 41141 14359 41199 14365
rect 41506 14356 41512 14368
rect 41564 14356 41570 14408
rect 42245 14399 42303 14405
rect 42245 14365 42257 14399
rect 42291 14396 42303 14399
rect 43254 14396 43260 14408
rect 42291 14368 43260 14396
rect 42291 14365 42303 14368
rect 42245 14359 42303 14365
rect 43254 14356 43260 14368
rect 43312 14356 43318 14408
rect 43349 14399 43407 14405
rect 43349 14365 43361 14399
rect 43395 14365 43407 14399
rect 43349 14359 43407 14365
rect 39114 14328 39120 14340
rect 38594 14300 38792 14328
rect 38856 14300 39120 14328
rect 38856 14260 38884 14300
rect 39114 14288 39120 14300
rect 39172 14288 39178 14340
rect 39206 14288 39212 14340
rect 39264 14328 39270 14340
rect 39850 14328 39856 14340
rect 39264 14300 39856 14328
rect 39264 14288 39270 14300
rect 39850 14288 39856 14300
rect 39908 14288 39914 14340
rect 40126 14288 40132 14340
rect 40184 14328 40190 14340
rect 40681 14331 40739 14337
rect 40681 14328 40693 14331
rect 40184 14300 40693 14328
rect 40184 14288 40190 14300
rect 40681 14297 40693 14300
rect 40727 14297 40739 14331
rect 42889 14331 42947 14337
rect 42889 14328 42901 14331
rect 40681 14291 40739 14297
rect 41708 14300 42901 14328
rect 36648 14232 38884 14260
rect 38930 14220 38936 14272
rect 38988 14260 38994 14272
rect 41708 14260 41736 14300
rect 42889 14297 42901 14300
rect 42935 14297 42947 14331
rect 42889 14291 42947 14297
rect 38988 14232 41736 14260
rect 38988 14220 38994 14232
rect 41966 14220 41972 14272
rect 42024 14260 42030 14272
rect 43364 14260 43392 14359
rect 44358 14356 44364 14408
rect 44416 14396 44422 14408
rect 45189 14399 45247 14405
rect 45189 14396 45201 14399
rect 44416 14368 45201 14396
rect 44416 14356 44422 14368
rect 45189 14365 45201 14368
rect 45235 14365 45247 14399
rect 45189 14359 45247 14365
rect 45370 14356 45376 14408
rect 45428 14396 45434 14408
rect 46308 14405 46336 14436
rect 48317 14433 48329 14436
rect 48363 14433 48375 14467
rect 48317 14427 48375 14433
rect 46293 14399 46351 14405
rect 46293 14396 46305 14399
rect 45428 14368 46305 14396
rect 45428 14356 45434 14368
rect 46293 14365 46305 14368
rect 46339 14365 46351 14399
rect 46293 14359 46351 14365
rect 47302 14356 47308 14408
rect 47360 14396 47366 14408
rect 47397 14399 47455 14405
rect 47397 14396 47409 14399
rect 47360 14368 47409 14396
rect 47360 14356 47366 14368
rect 47397 14365 47409 14368
rect 47443 14365 47455 14399
rect 47397 14359 47455 14365
rect 47762 14356 47768 14408
rect 47820 14396 47826 14408
rect 48685 14399 48743 14405
rect 48685 14396 48697 14399
rect 47820 14368 48697 14396
rect 47820 14356 47826 14368
rect 48685 14365 48697 14368
rect 48731 14365 48743 14399
rect 48685 14359 48743 14365
rect 42024 14232 43392 14260
rect 42024 14220 42030 14232
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 3602 14016 3608 14068
rect 3660 14016 3666 14068
rect 4890 14016 4896 14068
rect 4948 14016 4954 14068
rect 5994 14016 6000 14068
rect 6052 14016 6058 14068
rect 6362 14016 6368 14068
rect 6420 14056 6426 14068
rect 6549 14059 6607 14065
rect 6549 14056 6561 14059
rect 6420 14028 6561 14056
rect 6420 14016 6426 14028
rect 6549 14025 6561 14028
rect 6595 14025 6607 14059
rect 6549 14019 6607 14025
rect 6822 14016 6828 14068
rect 6880 14056 6886 14068
rect 7837 14059 7895 14065
rect 7837 14056 7849 14059
rect 6880 14028 7849 14056
rect 6880 14016 6886 14028
rect 7837 14025 7849 14028
rect 7883 14025 7895 14059
rect 7837 14019 7895 14025
rect 10042 14016 10048 14068
rect 10100 14016 10106 14068
rect 10502 14016 10508 14068
rect 10560 14056 10566 14068
rect 11149 14059 11207 14065
rect 11149 14056 11161 14059
rect 10560 14028 11161 14056
rect 10560 14016 10566 14028
rect 11149 14025 11161 14028
rect 11195 14025 11207 14059
rect 11149 14019 11207 14025
rect 12345 14059 12403 14065
rect 12345 14025 12357 14059
rect 12391 14056 12403 14059
rect 13722 14056 13728 14068
rect 12391 14028 13728 14056
rect 12391 14025 12403 14028
rect 12345 14019 12403 14025
rect 13722 14016 13728 14028
rect 13780 14016 13786 14068
rect 14458 14016 14464 14068
rect 14516 14016 14522 14068
rect 14550 14016 14556 14068
rect 14608 14056 14614 14068
rect 15197 14059 15255 14065
rect 15197 14056 15209 14059
rect 14608 14028 15209 14056
rect 14608 14016 14614 14028
rect 15197 14025 15209 14028
rect 15243 14025 15255 14059
rect 15197 14019 15255 14025
rect 15470 14016 15476 14068
rect 15528 14016 15534 14068
rect 15654 14016 15660 14068
rect 15712 14016 15718 14068
rect 15930 14016 15936 14068
rect 15988 14056 15994 14068
rect 16206 14056 16212 14068
rect 15988 14028 16212 14056
rect 15988 14016 15994 14028
rect 16206 14016 16212 14028
rect 16264 14016 16270 14068
rect 16390 14016 16396 14068
rect 16448 14056 16454 14068
rect 17221 14059 17279 14065
rect 17221 14056 17233 14059
rect 16448 14028 17233 14056
rect 16448 14016 16454 14028
rect 17221 14025 17233 14028
rect 17267 14025 17279 14059
rect 17221 14019 17279 14025
rect 17589 14059 17647 14065
rect 17589 14025 17601 14059
rect 17635 14056 17647 14059
rect 19058 14056 19064 14068
rect 17635 14028 19064 14056
rect 17635 14025 17647 14028
rect 17589 14019 17647 14025
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 20806 14056 20812 14068
rect 19812 14028 20812 14056
rect 5902 13948 5908 14000
rect 5960 13988 5966 14000
rect 5960 13960 7236 13988
rect 5960 13948 5966 13960
rect 1762 13880 1768 13932
rect 1820 13880 1826 13932
rect 2774 13880 2780 13932
rect 2832 13880 2838 13932
rect 2866 13880 2872 13932
rect 2924 13920 2930 13932
rect 3602 13920 3608 13932
rect 2924 13892 3608 13920
rect 2924 13880 2930 13892
rect 3602 13880 3608 13892
rect 3660 13880 3666 13932
rect 3789 13923 3847 13929
rect 3789 13889 3801 13923
rect 3835 13920 3847 13923
rect 4062 13920 4068 13932
rect 3835 13892 4068 13920
rect 3835 13889 3847 13892
rect 3789 13883 3847 13889
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 4249 13923 4307 13929
rect 4249 13889 4261 13923
rect 4295 13889 4307 13923
rect 4249 13883 4307 13889
rect 5353 13923 5411 13929
rect 5353 13889 5365 13923
rect 5399 13920 5411 13923
rect 5399 13892 6592 13920
rect 5399 13889 5411 13892
rect 5353 13883 5411 13889
rect 934 13812 940 13864
rect 992 13852 998 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 992 13824 2053 13852
rect 992 13812 998 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2792 13852 2820 13880
rect 3329 13855 3387 13861
rect 3329 13852 3341 13855
rect 2792 13824 3341 13852
rect 2041 13815 2099 13821
rect 3329 13821 3341 13824
rect 3375 13821 3387 13855
rect 4264 13852 4292 13883
rect 5994 13852 6000 13864
rect 4264 13824 6000 13852
rect 3329 13815 3387 13821
rect 3344 13784 3372 13815
rect 5994 13812 6000 13824
rect 6052 13812 6058 13864
rect 6564 13852 6592 13892
rect 6638 13880 6644 13932
rect 6696 13920 6702 13932
rect 7208 13929 7236 13960
rect 9950 13948 9956 14000
rect 10008 13988 10014 14000
rect 12434 13988 12440 14000
rect 10008 13960 12440 13988
rect 10008 13948 10014 13960
rect 12434 13948 12440 13960
rect 12492 13948 12498 14000
rect 13173 13991 13231 13997
rect 13173 13957 13185 13991
rect 13219 13988 13231 13991
rect 15488 13988 15516 14016
rect 13219 13960 15516 13988
rect 15565 13991 15623 13997
rect 13219 13957 13231 13960
rect 13173 13951 13231 13957
rect 15565 13957 15577 13991
rect 15611 13988 15623 13991
rect 15746 13988 15752 14000
rect 15611 13960 15752 13988
rect 15611 13957 15623 13960
rect 15565 13951 15623 13957
rect 15746 13948 15752 13960
rect 15804 13948 15810 14000
rect 16298 13948 16304 14000
rect 16356 13988 16362 14000
rect 17681 13991 17739 13997
rect 17681 13988 17693 13991
rect 16356 13960 17693 13988
rect 16356 13948 16362 13960
rect 17681 13957 17693 13960
rect 17727 13957 17739 13991
rect 17681 13951 17739 13957
rect 18322 13948 18328 14000
rect 18380 13948 18386 14000
rect 19812 13988 19840 14028
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 21450 14016 21456 14068
rect 21508 14016 21514 14068
rect 22002 14016 22008 14068
rect 22060 14016 22066 14068
rect 22465 14059 22523 14065
rect 22465 14025 22477 14059
rect 22511 14056 22523 14059
rect 22830 14056 22836 14068
rect 22511 14028 22836 14056
rect 22511 14025 22523 14028
rect 22465 14019 22523 14025
rect 22830 14016 22836 14028
rect 22888 14016 22894 14068
rect 23293 14059 23351 14065
rect 23293 14025 23305 14059
rect 23339 14056 23351 14059
rect 23658 14056 23664 14068
rect 23339 14028 23664 14056
rect 23339 14025 23351 14028
rect 23293 14019 23351 14025
rect 23658 14016 23664 14028
rect 23716 14016 23722 14068
rect 23753 14059 23811 14065
rect 23753 14025 23765 14059
rect 23799 14056 23811 14059
rect 25958 14056 25964 14068
rect 23799 14028 24440 14056
rect 23799 14025 23811 14028
rect 23753 14019 23811 14025
rect 19720 13960 19840 13988
rect 6733 13923 6791 13929
rect 6733 13920 6745 13923
rect 6696 13892 6745 13920
rect 6696 13880 6702 13892
rect 6733 13889 6745 13892
rect 6779 13889 6791 13923
rect 6733 13883 6791 13889
rect 7193 13923 7251 13929
rect 7193 13889 7205 13923
rect 7239 13889 7251 13923
rect 7193 13883 7251 13889
rect 8297 13923 8355 13929
rect 8297 13889 8309 13923
rect 8343 13889 8355 13923
rect 8297 13883 8355 13889
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13920 8999 13923
rect 9401 13923 9459 13929
rect 9401 13920 9413 13923
rect 8987 13892 9413 13920
rect 8987 13889 8999 13892
rect 8941 13883 8999 13889
rect 9401 13889 9413 13892
rect 9447 13889 9459 13923
rect 9401 13883 9459 13889
rect 10505 13923 10563 13929
rect 10505 13889 10517 13923
rect 10551 13920 10563 13923
rect 11238 13920 11244 13932
rect 10551 13892 11244 13920
rect 10551 13889 10563 13892
rect 10505 13883 10563 13889
rect 7834 13852 7840 13864
rect 6564 13824 7840 13852
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 8312 13852 8340 13883
rect 11238 13880 11244 13892
rect 11296 13880 11302 13932
rect 11698 13880 11704 13932
rect 11756 13880 11762 13932
rect 13265 13923 13323 13929
rect 13265 13889 13277 13923
rect 13311 13920 13323 13923
rect 13538 13920 13544 13932
rect 13311 13892 13544 13920
rect 13311 13889 13323 13892
rect 13265 13883 13323 13889
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 14369 13923 14427 13929
rect 14369 13889 14381 13923
rect 14415 13920 14427 13923
rect 15194 13920 15200 13932
rect 14415 13892 15200 13920
rect 14415 13889 14427 13892
rect 14369 13883 14427 13889
rect 15194 13880 15200 13892
rect 15252 13880 15258 13932
rect 15654 13880 15660 13932
rect 15712 13920 15718 13932
rect 16485 13923 16543 13929
rect 16485 13920 16497 13923
rect 15712 13892 16497 13920
rect 15712 13880 15718 13892
rect 16485 13889 16497 13892
rect 16531 13920 16543 13923
rect 17126 13920 17132 13932
rect 16531 13892 17132 13920
rect 16531 13889 16543 13892
rect 16485 13883 16543 13889
rect 17126 13880 17132 13892
rect 17184 13880 17190 13932
rect 18506 13880 18512 13932
rect 18564 13920 18570 13932
rect 19720 13929 19748 13960
rect 22186 13948 22192 14000
rect 22244 13988 22250 14000
rect 22738 13988 22744 14000
rect 22244 13960 22744 13988
rect 22244 13948 22250 13960
rect 22738 13948 22744 13960
rect 22796 13988 22802 14000
rect 22796 13960 23980 13988
rect 22796 13948 22802 13960
rect 18601 13923 18659 13929
rect 18601 13920 18613 13923
rect 18564 13892 18613 13920
rect 18564 13880 18570 13892
rect 18601 13889 18613 13892
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 19705 13923 19763 13929
rect 19705 13889 19717 13923
rect 19751 13889 19763 13923
rect 22094 13920 22100 13932
rect 21114 13906 22100 13920
rect 19705 13883 19763 13889
rect 21100 13892 22100 13906
rect 12802 13852 12808 13864
rect 8312 13824 12808 13852
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 13449 13855 13507 13861
rect 13449 13821 13461 13855
rect 13495 13821 13507 13855
rect 13449 13815 13507 13821
rect 14553 13855 14611 13861
rect 14553 13821 14565 13855
rect 14599 13821 14611 13855
rect 14553 13815 14611 13821
rect 9214 13784 9220 13796
rect 3344 13756 9220 13784
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 9306 13744 9312 13796
rect 9364 13784 9370 13796
rect 13464 13784 13492 13815
rect 13538 13784 13544 13796
rect 9364 13756 13400 13784
rect 13464 13756 13544 13784
rect 9364 13744 9370 13756
rect 6546 13676 6552 13728
rect 6604 13716 6610 13728
rect 6822 13716 6828 13728
rect 6604 13688 6828 13716
rect 6604 13676 6610 13688
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 7558 13676 7564 13728
rect 7616 13716 7622 13728
rect 9858 13716 9864 13728
rect 7616 13688 9864 13716
rect 7616 13676 7622 13688
rect 9858 13676 9864 13688
rect 9916 13716 9922 13728
rect 12158 13716 12164 13728
rect 9916 13688 12164 13716
rect 9916 13676 9922 13688
rect 12158 13676 12164 13688
rect 12216 13676 12222 13728
rect 12342 13676 12348 13728
rect 12400 13716 12406 13728
rect 12710 13716 12716 13728
rect 12400 13688 12716 13716
rect 12400 13676 12406 13688
rect 12710 13676 12716 13688
rect 12768 13676 12774 13728
rect 12802 13676 12808 13728
rect 12860 13676 12866 13728
rect 13372 13716 13400 13756
rect 13538 13744 13544 13756
rect 13596 13744 13602 13796
rect 14568 13784 14596 13815
rect 15010 13812 15016 13864
rect 15068 13852 15074 13864
rect 15749 13855 15807 13861
rect 15749 13852 15761 13855
rect 15068 13824 15761 13852
rect 15068 13812 15074 13824
rect 15749 13821 15761 13824
rect 15795 13821 15807 13855
rect 15749 13815 15807 13821
rect 16945 13855 17003 13861
rect 16945 13821 16957 13855
rect 16991 13852 17003 13855
rect 17034 13852 17040 13864
rect 16991 13824 17040 13852
rect 16991 13821 17003 13824
rect 16945 13815 17003 13821
rect 17034 13812 17040 13824
rect 17092 13812 17098 13864
rect 17773 13855 17831 13861
rect 17773 13821 17785 13855
rect 17819 13821 17831 13855
rect 17773 13815 17831 13821
rect 17788 13784 17816 13815
rect 19518 13812 19524 13864
rect 19576 13852 19582 13864
rect 21100 13852 21128 13892
rect 22094 13880 22100 13892
rect 22152 13880 22158 13932
rect 22373 13923 22431 13929
rect 22373 13920 22385 13923
rect 22204 13892 22385 13920
rect 19576 13824 21128 13852
rect 19576 13812 19582 13824
rect 17862 13784 17868 13796
rect 13924 13756 14596 13784
rect 13924 13716 13952 13756
rect 13372 13688 13952 13716
rect 14001 13719 14059 13725
rect 14001 13685 14013 13719
rect 14047 13716 14059 13719
rect 14458 13716 14464 13728
rect 14047 13688 14464 13716
rect 14047 13685 14059 13688
rect 14001 13679 14059 13685
rect 14458 13676 14464 13688
rect 14516 13676 14522 13728
rect 14568 13716 14596 13756
rect 16132 13756 17868 13784
rect 16132 13716 16160 13756
rect 17862 13744 17868 13756
rect 17920 13744 17926 13796
rect 22094 13744 22100 13796
rect 22152 13784 22158 13796
rect 22204 13784 22232 13892
rect 22373 13889 22385 13892
rect 22419 13889 22431 13923
rect 22373 13883 22431 13889
rect 22646 13880 22652 13932
rect 22704 13920 22710 13932
rect 23661 13923 23719 13929
rect 23661 13920 23673 13923
rect 22704 13892 23673 13920
rect 22704 13880 22710 13892
rect 23661 13889 23673 13892
rect 23707 13889 23719 13923
rect 23661 13883 23719 13889
rect 22557 13855 22615 13861
rect 22557 13821 22569 13855
rect 22603 13821 22615 13855
rect 22557 13815 22615 13821
rect 23845 13855 23903 13861
rect 23845 13821 23857 13855
rect 23891 13821 23903 13855
rect 23952 13852 23980 13960
rect 24412 13929 24440 14028
rect 24872 14028 25964 14056
rect 24486 13948 24492 14000
rect 24544 13988 24550 14000
rect 24872 13988 24900 14028
rect 25958 14016 25964 14028
rect 26016 14016 26022 14068
rect 26510 14016 26516 14068
rect 26568 14056 26574 14068
rect 26605 14059 26663 14065
rect 26605 14056 26617 14059
rect 26568 14028 26617 14056
rect 26568 14016 26574 14028
rect 26605 14025 26617 14028
rect 26651 14025 26663 14059
rect 31754 14056 31760 14068
rect 26605 14019 26663 14025
rect 28920 14028 31760 14056
rect 27338 13988 27344 14000
rect 24544 13960 24900 13988
rect 26358 13960 27344 13988
rect 24544 13948 24550 13960
rect 24397 13923 24455 13929
rect 24397 13889 24409 13923
rect 24443 13920 24455 13923
rect 24670 13920 24676 13932
rect 24443 13892 24676 13920
rect 24443 13889 24455 13892
rect 24397 13883 24455 13889
rect 24670 13880 24676 13892
rect 24728 13880 24734 13932
rect 24872 13929 24900 13960
rect 27338 13948 27344 13960
rect 27396 13948 27402 14000
rect 28920 13997 28948 14028
rect 31754 14016 31760 14028
rect 31812 14056 31818 14068
rect 32766 14056 32772 14068
rect 31812 14028 32772 14056
rect 31812 14016 31818 14028
rect 32766 14016 32772 14028
rect 32824 14016 32830 14068
rect 33502 14016 33508 14068
rect 33560 14056 33566 14068
rect 34885 14059 34943 14065
rect 34885 14056 34897 14059
rect 33560 14028 34897 14056
rect 33560 14016 33566 14028
rect 34885 14025 34897 14028
rect 34931 14025 34943 14059
rect 34885 14019 34943 14025
rect 28905 13991 28963 13997
rect 28905 13957 28917 13991
rect 28951 13957 28963 13991
rect 28905 13951 28963 13957
rect 24857 13923 24915 13929
rect 24857 13889 24869 13923
rect 24903 13889 24915 13923
rect 24857 13883 24915 13889
rect 27154 13880 27160 13932
rect 27212 13880 27218 13932
rect 28920 13852 28948 13951
rect 31294 13948 31300 14000
rect 31352 13988 31358 14000
rect 32309 13991 32367 13997
rect 32309 13988 32321 13991
rect 31352 13960 32321 13988
rect 31352 13948 31358 13960
rect 32309 13957 32321 13960
rect 32355 13957 32367 13991
rect 32309 13951 32367 13957
rect 32674 13948 32680 14000
rect 32732 13988 32738 14000
rect 34900 13988 34928 14019
rect 35342 14016 35348 14068
rect 35400 14016 35406 14068
rect 37461 14059 37519 14065
rect 35452 14028 36952 14056
rect 35452 13988 35480 14028
rect 32732 13960 33902 13988
rect 34900 13960 35480 13988
rect 32732 13948 32738 13960
rect 35986 13948 35992 14000
rect 36044 13948 36050 14000
rect 36814 13948 36820 14000
rect 36872 13948 36878 14000
rect 36924 13988 36952 14028
rect 37461 14025 37473 14059
rect 37507 14056 37519 14059
rect 38470 14056 38476 14068
rect 37507 14028 38476 14056
rect 37507 14025 37519 14028
rect 37461 14019 37519 14025
rect 38470 14016 38476 14028
rect 38528 14016 38534 14068
rect 38657 14059 38715 14065
rect 38657 14025 38669 14059
rect 38703 14056 38715 14059
rect 38703 14028 41414 14056
rect 38703 14025 38715 14028
rect 38657 14019 38715 14025
rect 41386 13988 41414 14028
rect 41506 14016 41512 14068
rect 41564 14056 41570 14068
rect 41601 14059 41659 14065
rect 41601 14056 41613 14059
rect 41564 14028 41613 14056
rect 41564 14016 41570 14028
rect 41601 14025 41613 14028
rect 41647 14025 41659 14059
rect 41601 14019 41659 14025
rect 43254 14016 43260 14068
rect 43312 14016 43318 14068
rect 44358 14016 44364 14068
rect 44416 14016 44422 14068
rect 44542 14016 44548 14068
rect 44600 14056 44606 14068
rect 44637 14059 44695 14065
rect 44637 14056 44649 14059
rect 44600 14028 44649 14056
rect 44600 14016 44606 14028
rect 44637 14025 44649 14028
rect 44683 14056 44695 14059
rect 45554 14056 45560 14068
rect 44683 14028 45560 14056
rect 44683 14025 44695 14028
rect 44637 14019 44695 14025
rect 45554 14016 45560 14028
rect 45612 14016 45618 14068
rect 45738 14016 45744 14068
rect 45796 14056 45802 14068
rect 46937 14059 46995 14065
rect 46937 14056 46949 14059
rect 45796 14028 46949 14056
rect 45796 14016 45802 14028
rect 46937 14025 46949 14028
rect 46983 14025 46995 14059
rect 46937 14019 46995 14025
rect 47026 14016 47032 14068
rect 47084 14056 47090 14068
rect 47213 14059 47271 14065
rect 47213 14056 47225 14059
rect 47084 14028 47225 14056
rect 47084 14016 47090 14028
rect 47213 14025 47225 14028
rect 47259 14056 47271 14059
rect 47394 14056 47400 14068
rect 47259 14028 47400 14056
rect 47259 14025 47271 14028
rect 47213 14019 47271 14025
rect 47394 14016 47400 14028
rect 47452 14016 47458 14068
rect 47762 14016 47768 14068
rect 47820 14056 47826 14068
rect 47949 14059 48007 14065
rect 47949 14056 47961 14059
rect 47820 14028 47961 14056
rect 47820 14016 47826 14028
rect 47949 14025 47961 14028
rect 47995 14025 48007 14059
rect 47949 14019 48007 14025
rect 48314 14016 48320 14068
rect 48372 14056 48378 14068
rect 49329 14059 49387 14065
rect 49329 14056 49341 14059
rect 48372 14028 49341 14056
rect 48372 14016 48378 14028
rect 49329 14025 49341 14028
rect 49375 14025 49387 14059
rect 49329 14019 49387 14025
rect 43346 13988 43352 14000
rect 36924 13960 41000 13988
rect 41386 13960 43352 13988
rect 29362 13880 29368 13932
rect 29420 13880 29426 13932
rect 30742 13880 30748 13932
rect 30800 13880 30806 13932
rect 31018 13880 31024 13932
rect 31076 13920 31082 13932
rect 31076 13892 33088 13920
rect 31076 13880 31082 13892
rect 29730 13852 29736 13864
rect 23952 13824 28948 13852
rect 29012 13824 29736 13852
rect 23845 13815 23903 13821
rect 22152 13756 22232 13784
rect 22572 13784 22600 13815
rect 22646 13784 22652 13796
rect 22572 13756 22652 13784
rect 22152 13744 22158 13756
rect 22646 13744 22652 13756
rect 22704 13744 22710 13796
rect 23860 13784 23888 13815
rect 24118 13784 24124 13796
rect 23860 13756 24124 13784
rect 24118 13744 24124 13756
rect 24176 13744 24182 13796
rect 29012 13784 29040 13824
rect 29730 13812 29736 13824
rect 29788 13812 29794 13864
rect 30190 13812 30196 13864
rect 30248 13852 30254 13864
rect 31113 13855 31171 13861
rect 31113 13852 31125 13855
rect 30248 13824 31125 13852
rect 30248 13812 30254 13824
rect 31113 13821 31125 13824
rect 31159 13821 31171 13855
rect 31113 13815 31171 13821
rect 31573 13855 31631 13861
rect 31573 13821 31585 13855
rect 31619 13852 31631 13855
rect 31662 13852 31668 13864
rect 31619 13824 31668 13852
rect 31619 13821 31631 13824
rect 31573 13815 31631 13821
rect 31662 13812 31668 13824
rect 31720 13812 31726 13864
rect 33060 13852 33088 13892
rect 33134 13880 33140 13932
rect 33192 13880 33198 13932
rect 35529 13923 35587 13929
rect 35529 13889 35541 13923
rect 35575 13920 35587 13923
rect 36170 13920 36176 13932
rect 35575 13892 36176 13920
rect 35575 13889 35587 13892
rect 35529 13883 35587 13889
rect 36170 13880 36176 13892
rect 36228 13880 36234 13932
rect 37829 13923 37887 13929
rect 37829 13920 37841 13923
rect 37200 13892 37841 13920
rect 34698 13852 34704 13864
rect 33060 13824 34704 13852
rect 34698 13812 34704 13824
rect 34756 13812 34762 13864
rect 35894 13812 35900 13864
rect 35952 13852 35958 13864
rect 37090 13852 37096 13864
rect 35952 13824 37096 13852
rect 35952 13812 35958 13824
rect 37090 13812 37096 13824
rect 37148 13812 37154 13864
rect 32858 13784 32864 13796
rect 26528 13756 29040 13784
rect 30668 13756 32864 13784
rect 14568 13688 16160 13716
rect 16574 13676 16580 13728
rect 16632 13716 16638 13728
rect 16669 13719 16727 13725
rect 16669 13716 16681 13719
rect 16632 13688 16681 13716
rect 16632 13676 16638 13688
rect 16669 13685 16681 13688
rect 16715 13685 16727 13719
rect 16669 13679 16727 13685
rect 19242 13676 19248 13728
rect 19300 13676 19306 13728
rect 19968 13719 20026 13725
rect 19968 13685 19980 13719
rect 20014 13716 20026 13719
rect 21358 13716 21364 13728
rect 20014 13688 21364 13716
rect 20014 13685 20026 13688
rect 19968 13679 20026 13685
rect 21358 13676 21364 13688
rect 21416 13676 21422 13728
rect 22370 13676 22376 13728
rect 22428 13716 22434 13728
rect 22830 13716 22836 13728
rect 22428 13688 22836 13716
rect 22428 13676 22434 13688
rect 22830 13676 22836 13688
rect 22888 13676 22894 13728
rect 23474 13676 23480 13728
rect 23532 13716 23538 13728
rect 24581 13719 24639 13725
rect 24581 13716 24593 13719
rect 23532 13688 24593 13716
rect 23532 13676 23538 13688
rect 24581 13685 24593 13688
rect 24627 13716 24639 13719
rect 24946 13716 24952 13728
rect 24627 13688 24952 13716
rect 24627 13685 24639 13688
rect 24581 13679 24639 13685
rect 24946 13676 24952 13688
rect 25004 13676 25010 13728
rect 25120 13719 25178 13725
rect 25120 13685 25132 13719
rect 25166 13716 25178 13719
rect 26528 13716 26556 13756
rect 25166 13688 26556 13716
rect 29628 13719 29686 13725
rect 25166 13685 25178 13688
rect 25120 13679 25178 13685
rect 29628 13685 29640 13719
rect 29674 13716 29686 13719
rect 30668 13716 30696 13756
rect 32858 13744 32864 13756
rect 32916 13744 32922 13796
rect 35342 13744 35348 13796
rect 35400 13784 35406 13796
rect 37200 13784 37228 13892
rect 37829 13889 37841 13892
rect 37875 13889 37887 13923
rect 37829 13883 37887 13889
rect 39025 13923 39083 13929
rect 39025 13889 39037 13923
rect 39071 13920 39083 13923
rect 39758 13920 39764 13932
rect 39071 13892 39764 13920
rect 39071 13889 39083 13892
rect 39025 13883 39083 13889
rect 39758 13880 39764 13892
rect 39816 13880 39822 13932
rect 39850 13880 39856 13932
rect 39908 13880 39914 13932
rect 39942 13880 39948 13932
rect 40000 13920 40006 13932
rect 40972 13929 41000 13960
rect 43346 13948 43352 13960
rect 43404 13948 43410 14000
rect 43898 13948 43904 14000
rect 43956 13988 43962 14000
rect 44821 13991 44879 13997
rect 44821 13988 44833 13991
rect 43956 13960 44833 13988
rect 43956 13948 43962 13960
rect 44821 13957 44833 13960
rect 44867 13957 44879 13991
rect 50614 13988 50620 14000
rect 44821 13951 44879 13957
rect 45848 13960 50620 13988
rect 40957 13923 41015 13929
rect 40000 13892 40908 13920
rect 40000 13880 40006 13892
rect 37921 13855 37979 13861
rect 37921 13821 37933 13855
rect 37967 13821 37979 13855
rect 37921 13815 37979 13821
rect 38105 13855 38163 13861
rect 38105 13821 38117 13855
rect 38151 13821 38163 13855
rect 38105 13815 38163 13821
rect 35400 13756 37228 13784
rect 35400 13744 35406 13756
rect 37274 13744 37280 13796
rect 37332 13784 37338 13796
rect 37936 13784 37964 13815
rect 37332 13756 37964 13784
rect 37332 13744 37338 13756
rect 38010 13744 38016 13796
rect 38068 13784 38074 13796
rect 38120 13784 38148 13815
rect 38286 13812 38292 13864
rect 38344 13852 38350 13864
rect 39117 13855 39175 13861
rect 39117 13852 39129 13855
rect 38344 13824 39129 13852
rect 38344 13812 38350 13824
rect 39117 13821 39129 13824
rect 39163 13821 39175 13855
rect 39117 13815 39175 13821
rect 39301 13855 39359 13861
rect 39301 13821 39313 13855
rect 39347 13821 39359 13855
rect 39301 13815 39359 13821
rect 38068 13756 38148 13784
rect 38068 13744 38074 13756
rect 38194 13744 38200 13796
rect 38252 13784 38258 13796
rect 39316 13784 39344 13815
rect 40494 13812 40500 13864
rect 40552 13812 40558 13864
rect 40880 13852 40908 13892
rect 40957 13889 40969 13923
rect 41003 13889 41015 13923
rect 42613 13923 42671 13929
rect 42613 13920 42625 13923
rect 40957 13883 41015 13889
rect 41386 13892 42625 13920
rect 41386 13852 41414 13892
rect 42613 13889 42625 13892
rect 42659 13889 42671 13923
rect 42613 13883 42671 13889
rect 42702 13880 42708 13932
rect 42760 13920 42766 13932
rect 43717 13923 43775 13929
rect 43717 13920 43729 13923
rect 42760 13892 43729 13920
rect 42760 13880 42766 13892
rect 43717 13889 43729 13892
rect 43763 13889 43775 13923
rect 43717 13883 43775 13889
rect 45189 13923 45247 13929
rect 45189 13889 45201 13923
rect 45235 13920 45247 13923
rect 45278 13920 45284 13932
rect 45235 13892 45284 13920
rect 45235 13889 45247 13892
rect 45189 13883 45247 13889
rect 45278 13880 45284 13892
rect 45336 13880 45342 13932
rect 40880 13824 41414 13852
rect 41690 13812 41696 13864
rect 41748 13852 41754 13864
rect 41969 13855 42027 13861
rect 41969 13852 41981 13855
rect 41748 13824 41981 13852
rect 41748 13812 41754 13824
rect 41969 13821 41981 13824
rect 42015 13852 42027 13855
rect 42153 13855 42211 13861
rect 42153 13852 42165 13855
rect 42015 13824 42165 13852
rect 42015 13821 42027 13824
rect 41969 13815 42027 13821
rect 42153 13821 42165 13824
rect 42199 13852 42211 13855
rect 44634 13852 44640 13864
rect 42199 13824 44640 13852
rect 42199 13821 42211 13824
rect 42153 13815 42211 13821
rect 44634 13812 44640 13824
rect 44692 13812 44698 13864
rect 42610 13784 42616 13796
rect 38252 13756 42616 13784
rect 38252 13744 38258 13756
rect 42610 13744 42616 13756
rect 42668 13744 42674 13796
rect 29674 13688 30696 13716
rect 33400 13719 33458 13725
rect 29674 13685 29686 13688
rect 29628 13679 29686 13685
rect 33400 13685 33412 13719
rect 33446 13716 33458 13719
rect 34422 13716 34428 13728
rect 33446 13688 34428 13716
rect 33446 13685 33458 13688
rect 33400 13679 33458 13685
rect 34422 13676 34428 13688
rect 34480 13676 34486 13728
rect 34606 13676 34612 13728
rect 34664 13716 34670 13728
rect 38286 13716 38292 13728
rect 34664 13688 38292 13716
rect 34664 13676 34670 13688
rect 38286 13676 38292 13688
rect 38344 13676 38350 13728
rect 38562 13676 38568 13728
rect 38620 13716 38626 13728
rect 40586 13716 40592 13728
rect 38620 13688 40592 13716
rect 38620 13676 38626 13688
rect 40586 13676 40592 13688
rect 40644 13676 40650 13728
rect 42518 13676 42524 13728
rect 42576 13716 42582 13728
rect 45848 13725 45876 13960
rect 50614 13948 50620 13960
rect 50672 13948 50678 14000
rect 46290 13880 46296 13932
rect 46348 13880 46354 13932
rect 46382 13880 46388 13932
rect 46440 13920 46446 13932
rect 47765 13923 47823 13929
rect 47765 13920 47777 13923
rect 46440 13892 47777 13920
rect 46440 13880 46446 13892
rect 47765 13889 47777 13892
rect 47811 13920 47823 13923
rect 47854 13920 47860 13932
rect 47811 13892 47860 13920
rect 47811 13889 47823 13892
rect 47765 13883 47823 13889
rect 47854 13880 47860 13892
rect 47912 13880 47918 13932
rect 48590 13880 48596 13932
rect 48648 13920 48654 13932
rect 48685 13923 48743 13929
rect 48685 13920 48697 13923
rect 48648 13892 48697 13920
rect 48648 13880 48654 13892
rect 48685 13889 48697 13892
rect 48731 13920 48743 13923
rect 49142 13920 49148 13932
rect 48731 13892 49148 13920
rect 48731 13889 48743 13892
rect 48685 13883 48743 13889
rect 49142 13880 49148 13892
rect 49200 13880 49206 13932
rect 46308 13852 46336 13880
rect 48317 13855 48375 13861
rect 48317 13852 48329 13855
rect 46308 13824 48329 13852
rect 48317 13821 48329 13824
rect 48363 13821 48375 13855
rect 48317 13815 48375 13821
rect 45833 13719 45891 13725
rect 45833 13716 45845 13719
rect 42576 13688 45845 13716
rect 42576 13676 42582 13688
rect 45833 13685 45845 13688
rect 45879 13685 45891 13719
rect 45833 13679 45891 13685
rect 47486 13676 47492 13728
rect 47544 13716 47550 13728
rect 47762 13716 47768 13728
rect 47544 13688 47768 13716
rect 47544 13676 47550 13688
rect 47762 13676 47768 13688
rect 47820 13676 47826 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 3418 13472 3424 13524
rect 3476 13472 3482 13524
rect 7466 13472 7472 13524
rect 7524 13472 7530 13524
rect 8573 13515 8631 13521
rect 8573 13481 8585 13515
rect 8619 13512 8631 13515
rect 11882 13512 11888 13524
rect 8619 13484 11888 13512
rect 8619 13481 8631 13484
rect 8573 13475 8631 13481
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 12434 13472 12440 13524
rect 12492 13472 12498 13524
rect 12710 13472 12716 13524
rect 12768 13512 12774 13524
rect 16022 13512 16028 13524
rect 12768 13484 16028 13512
rect 12768 13472 12774 13484
rect 16022 13472 16028 13484
rect 16080 13472 16086 13524
rect 17862 13472 17868 13524
rect 17920 13472 17926 13524
rect 18322 13472 18328 13524
rect 18380 13512 18386 13524
rect 18782 13512 18788 13524
rect 18380 13484 18788 13512
rect 18380 13472 18386 13484
rect 18782 13472 18788 13484
rect 18840 13472 18846 13524
rect 19429 13515 19487 13521
rect 19429 13481 19441 13515
rect 19475 13512 19487 13515
rect 19518 13512 19524 13524
rect 19475 13484 19524 13512
rect 19475 13481 19487 13484
rect 19429 13475 19487 13481
rect 19518 13472 19524 13484
rect 19576 13472 19582 13524
rect 19705 13515 19763 13521
rect 19705 13481 19717 13515
rect 19751 13512 19763 13515
rect 19978 13512 19984 13524
rect 19751 13484 19984 13512
rect 19751 13481 19763 13484
rect 19705 13475 19763 13481
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 21634 13512 21640 13524
rect 20272 13484 21640 13512
rect 2130 13404 2136 13456
rect 2188 13444 2194 13456
rect 4522 13444 4528 13456
rect 2188 13416 4528 13444
rect 2188 13404 2194 13416
rect 4522 13404 4528 13416
rect 4580 13404 4586 13456
rect 8478 13444 8484 13456
rect 5736 13416 8484 13444
rect 2774 13336 2780 13388
rect 2832 13336 2838 13388
rect 3605 13379 3663 13385
rect 3605 13345 3617 13379
rect 3651 13376 3663 13379
rect 3651 13348 4660 13376
rect 3651 13345 3663 13348
rect 3605 13339 3663 13345
rect 4632 13317 4660 13348
rect 1765 13311 1823 13317
rect 1765 13277 1777 13311
rect 1811 13277 1823 13311
rect 4617 13311 4675 13317
rect 1765 13271 1823 13277
rect 2746 13280 4108 13308
rect 1780 13240 1808 13271
rect 2746 13240 2774 13280
rect 1780 13212 2774 13240
rect 3970 13200 3976 13252
rect 4028 13200 4034 13252
rect 4080 13240 4108 13280
rect 4617 13277 4629 13311
rect 4663 13308 4675 13311
rect 5074 13308 5080 13320
rect 4663 13280 5080 13308
rect 4663 13277 4675 13280
rect 4617 13271 4675 13277
rect 5074 13268 5080 13280
rect 5132 13268 5138 13320
rect 5736 13317 5764 13416
rect 8478 13404 8484 13416
rect 8536 13404 8542 13456
rect 8754 13404 8760 13456
rect 8812 13444 8818 13456
rect 9033 13447 9091 13453
rect 9033 13444 9045 13447
rect 8812 13416 9045 13444
rect 8812 13404 8818 13416
rect 9033 13413 9045 13416
rect 9079 13444 9091 13447
rect 9122 13444 9128 13456
rect 9079 13416 9128 13444
rect 9079 13413 9091 13416
rect 9033 13407 9091 13413
rect 9122 13404 9128 13416
rect 9180 13404 9186 13456
rect 9950 13404 9956 13456
rect 10008 13404 10014 13456
rect 12452 13444 12480 13472
rect 13078 13444 13084 13456
rect 12452 13416 13084 13444
rect 13078 13404 13084 13416
rect 13136 13404 13142 13456
rect 13446 13404 13452 13456
rect 13504 13444 13510 13456
rect 13909 13447 13967 13453
rect 13909 13444 13921 13447
rect 13504 13416 13921 13444
rect 13504 13404 13510 13416
rect 13909 13413 13921 13416
rect 13955 13444 13967 13447
rect 15378 13444 15384 13456
rect 13955 13416 15384 13444
rect 13955 13413 13967 13416
rect 13909 13407 13967 13413
rect 15378 13404 15384 13416
rect 15436 13404 15442 13456
rect 18509 13447 18567 13453
rect 18509 13413 18521 13447
rect 18555 13444 18567 13447
rect 20162 13444 20168 13456
rect 18555 13416 20168 13444
rect 18555 13413 18567 13416
rect 18509 13407 18567 13413
rect 20162 13404 20168 13416
rect 20220 13404 20226 13456
rect 9582 13376 9588 13388
rect 6196 13348 9588 13376
rect 5721 13311 5779 13317
rect 5721 13277 5733 13311
rect 5767 13277 5779 13311
rect 5721 13271 5779 13277
rect 6196 13240 6224 13348
rect 9582 13336 9588 13348
rect 9640 13336 9646 13388
rect 10318 13336 10324 13388
rect 10376 13376 10382 13388
rect 10413 13379 10471 13385
rect 10413 13376 10425 13379
rect 10376 13348 10425 13376
rect 10376 13336 10382 13348
rect 10413 13345 10425 13348
rect 10459 13376 10471 13379
rect 10778 13376 10784 13388
rect 10459 13348 10784 13376
rect 10459 13345 10471 13348
rect 10413 13339 10471 13345
rect 10778 13336 10784 13348
rect 10836 13336 10842 13388
rect 11146 13336 11152 13388
rect 11204 13376 11210 13388
rect 11882 13376 11888 13388
rect 11204 13348 11888 13376
rect 11204 13336 11210 13348
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 12434 13336 12440 13388
rect 12492 13376 12498 13388
rect 12986 13376 12992 13388
rect 12492 13348 12992 13376
rect 12492 13336 12498 13348
rect 12986 13336 12992 13348
rect 13044 13336 13050 13388
rect 13170 13336 13176 13388
rect 13228 13336 13234 13388
rect 13357 13379 13415 13385
rect 13357 13345 13369 13379
rect 13403 13376 13415 13379
rect 13538 13376 13544 13388
rect 13403 13348 13544 13376
rect 13403 13345 13415 13348
rect 13357 13339 13415 13345
rect 13538 13336 13544 13348
rect 13596 13336 13602 13388
rect 16393 13379 16451 13385
rect 16393 13376 16405 13379
rect 14200 13348 16405 13376
rect 6825 13311 6883 13317
rect 6825 13277 6837 13311
rect 6871 13308 6883 13311
rect 7834 13308 7840 13320
rect 6871 13280 7840 13308
rect 6871 13277 6883 13280
rect 6825 13271 6883 13277
rect 7834 13268 7840 13280
rect 7892 13268 7898 13320
rect 7929 13311 7987 13317
rect 7929 13277 7941 13311
rect 7975 13308 7987 13311
rect 8846 13308 8852 13320
rect 7975 13280 8852 13308
rect 7975 13277 7987 13280
rect 7929 13271 7987 13277
rect 8846 13268 8852 13280
rect 8904 13268 8910 13320
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13308 9367 13311
rect 9858 13308 9864 13320
rect 9355 13280 9864 13308
rect 9355 13277 9367 13280
rect 9309 13271 9367 13277
rect 9858 13268 9864 13280
rect 9916 13268 9922 13320
rect 12066 13268 12072 13320
rect 12124 13308 12130 13320
rect 13081 13311 13139 13317
rect 13081 13308 13093 13311
rect 12124 13280 13093 13308
rect 12124 13268 12130 13280
rect 13081 13277 13093 13280
rect 13127 13277 13139 13311
rect 13081 13271 13139 13277
rect 4080 13212 6224 13240
rect 6454 13200 6460 13252
rect 6512 13240 6518 13252
rect 10689 13243 10747 13249
rect 10689 13240 10701 13243
rect 6512 13212 10701 13240
rect 6512 13200 6518 13212
rect 10689 13209 10701 13212
rect 10735 13209 10747 13243
rect 10689 13203 10747 13209
rect 11698 13200 11704 13252
rect 11756 13200 11762 13252
rect 14200 13240 14228 13348
rect 16393 13345 16405 13348
rect 16439 13345 16451 13379
rect 16393 13339 16451 13345
rect 18690 13336 18696 13388
rect 18748 13336 18754 13388
rect 18874 13336 18880 13388
rect 18932 13376 18938 13388
rect 19061 13379 19119 13385
rect 19061 13376 19073 13379
rect 18932 13348 19073 13376
rect 18932 13336 18938 13348
rect 19061 13345 19073 13348
rect 19107 13376 19119 13379
rect 20070 13376 20076 13388
rect 19107 13348 20076 13376
rect 19107 13345 19119 13348
rect 19061 13339 19119 13345
rect 20070 13336 20076 13348
rect 20128 13336 20134 13388
rect 20272 13385 20300 13484
rect 21634 13472 21640 13484
rect 21692 13472 21698 13524
rect 24578 13472 24584 13524
rect 24636 13512 24642 13524
rect 26329 13515 26387 13521
rect 26329 13512 26341 13515
rect 24636 13484 26341 13512
rect 24636 13472 24642 13484
rect 26329 13481 26341 13484
rect 26375 13481 26387 13515
rect 26329 13475 26387 13481
rect 27154 13472 27160 13524
rect 27212 13512 27218 13524
rect 30098 13512 30104 13524
rect 27212 13484 30104 13512
rect 27212 13472 27218 13484
rect 30098 13472 30104 13484
rect 30156 13472 30162 13524
rect 32582 13512 32588 13524
rect 30208 13484 32588 13512
rect 23768 13416 24716 13444
rect 20257 13379 20315 13385
rect 20257 13345 20269 13379
rect 20303 13345 20315 13379
rect 20257 13339 20315 13345
rect 14274 13268 14280 13320
rect 14332 13308 14338 13320
rect 15473 13311 15531 13317
rect 15473 13308 15485 13311
rect 14332 13280 15485 13308
rect 14332 13268 14338 13280
rect 15473 13277 15485 13280
rect 15519 13308 15531 13311
rect 16117 13311 16175 13317
rect 16117 13308 16129 13311
rect 15519 13280 16129 13308
rect 15519 13277 15531 13280
rect 15473 13271 15531 13277
rect 16117 13277 16129 13280
rect 16163 13277 16175 13311
rect 16117 13271 16175 13277
rect 19610 13268 19616 13320
rect 19668 13308 19674 13320
rect 20272 13308 20300 13339
rect 20806 13336 20812 13388
rect 20864 13376 20870 13388
rect 20901 13379 20959 13385
rect 20901 13376 20913 13379
rect 20864 13348 20913 13376
rect 20864 13336 20870 13348
rect 20901 13345 20913 13348
rect 20947 13376 20959 13379
rect 21542 13376 21548 13388
rect 20947 13348 21548 13376
rect 20947 13345 20959 13348
rect 20901 13339 20959 13345
rect 21542 13336 21548 13348
rect 21600 13336 21606 13388
rect 21634 13336 21640 13388
rect 21692 13376 21698 13388
rect 22649 13379 22707 13385
rect 22649 13376 22661 13379
rect 21692 13348 22661 13376
rect 21692 13336 21698 13348
rect 22649 13345 22661 13348
rect 22695 13345 22707 13379
rect 22649 13339 22707 13345
rect 23014 13336 23020 13388
rect 23072 13336 23078 13388
rect 23768 13385 23796 13416
rect 23753 13379 23811 13385
rect 23753 13345 23765 13379
rect 23799 13345 23811 13379
rect 23753 13339 23811 13345
rect 23937 13379 23995 13385
rect 23937 13345 23949 13379
rect 23983 13376 23995 13379
rect 23983 13348 24348 13376
rect 23983 13345 23995 13348
rect 23937 13339 23995 13345
rect 23474 13308 23480 13320
rect 19668 13280 20300 13308
rect 22310 13280 23480 13308
rect 19668 13268 19674 13280
rect 23474 13268 23480 13280
rect 23532 13268 23538 13320
rect 11992 13212 14228 13240
rect 5261 13175 5319 13181
rect 5261 13141 5273 13175
rect 5307 13172 5319 13175
rect 6086 13172 6092 13184
rect 5307 13144 6092 13172
rect 5307 13141 5319 13144
rect 5261 13135 5319 13141
rect 6086 13132 6092 13144
rect 6144 13132 6150 13184
rect 6365 13175 6423 13181
rect 6365 13141 6377 13175
rect 6411 13172 6423 13175
rect 8478 13172 8484 13184
rect 6411 13144 8484 13172
rect 6411 13141 6423 13144
rect 6365 13135 6423 13141
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 10594 13132 10600 13184
rect 10652 13172 10658 13184
rect 11992 13172 12020 13212
rect 14366 13200 14372 13252
rect 14424 13200 14430 13252
rect 14737 13243 14795 13249
rect 14737 13209 14749 13243
rect 14783 13240 14795 13243
rect 14826 13240 14832 13252
rect 14783 13212 14832 13240
rect 14783 13209 14795 13212
rect 14737 13203 14795 13209
rect 14826 13200 14832 13212
rect 14884 13240 14890 13252
rect 16482 13240 16488 13252
rect 14884 13212 16488 13240
rect 14884 13200 14890 13212
rect 16482 13200 16488 13212
rect 16540 13200 16546 13252
rect 18690 13240 18696 13252
rect 17618 13212 18696 13240
rect 18690 13200 18696 13212
rect 18748 13200 18754 13252
rect 18874 13200 18880 13252
rect 18932 13240 18938 13252
rect 19794 13240 19800 13252
rect 18932 13212 19800 13240
rect 18932 13200 18938 13212
rect 19794 13200 19800 13212
rect 19852 13200 19858 13252
rect 20073 13243 20131 13249
rect 20073 13209 20085 13243
rect 20119 13240 20131 13243
rect 20898 13240 20904 13252
rect 20119 13212 20904 13240
rect 20119 13209 20131 13212
rect 20073 13203 20131 13209
rect 20898 13200 20904 13212
rect 20956 13200 20962 13252
rect 21174 13200 21180 13252
rect 21232 13200 21238 13252
rect 24320 13240 24348 13348
rect 24486 13336 24492 13388
rect 24544 13376 24550 13388
rect 24581 13379 24639 13385
rect 24581 13376 24593 13379
rect 24544 13348 24593 13376
rect 24544 13336 24550 13348
rect 24581 13345 24593 13348
rect 24627 13345 24639 13379
rect 24688 13376 24716 13416
rect 25958 13404 25964 13456
rect 26016 13444 26022 13456
rect 26016 13416 26924 13444
rect 26016 13404 26022 13416
rect 26786 13376 26792 13388
rect 24688 13348 26792 13376
rect 24581 13339 24639 13345
rect 26786 13336 26792 13348
rect 26844 13336 26850 13388
rect 26896 13385 26924 13416
rect 28902 13404 28908 13456
rect 28960 13444 28966 13456
rect 28960 13416 29500 13444
rect 28960 13404 28966 13416
rect 26881 13379 26939 13385
rect 26881 13345 26893 13379
rect 26927 13376 26939 13379
rect 29362 13376 29368 13388
rect 26927 13348 29368 13376
rect 26927 13345 26939 13348
rect 26881 13339 26939 13345
rect 29362 13336 29368 13348
rect 29420 13336 29426 13388
rect 29472 13376 29500 13416
rect 29546 13404 29552 13456
rect 29604 13404 29610 13456
rect 29638 13404 29644 13456
rect 29696 13444 29702 13456
rect 29917 13447 29975 13453
rect 29917 13444 29929 13447
rect 29696 13416 29929 13444
rect 29696 13404 29702 13416
rect 29917 13413 29929 13416
rect 29963 13413 29975 13447
rect 29917 13407 29975 13413
rect 30208 13376 30236 13484
rect 32582 13472 32588 13484
rect 32640 13472 32646 13524
rect 33318 13472 33324 13524
rect 33376 13512 33382 13524
rect 34054 13512 34060 13524
rect 33376 13484 34060 13512
rect 33376 13472 33382 13484
rect 34054 13472 34060 13484
rect 34112 13472 34118 13524
rect 34882 13472 34888 13524
rect 34940 13472 34946 13524
rect 35176 13484 37780 13512
rect 30374 13404 30380 13456
rect 30432 13404 30438 13456
rect 32493 13447 32551 13453
rect 32493 13413 32505 13447
rect 32539 13444 32551 13447
rect 32674 13444 32680 13456
rect 32539 13416 32680 13444
rect 32539 13413 32551 13416
rect 32493 13407 32551 13413
rect 32674 13404 32680 13416
rect 32732 13444 32738 13456
rect 35176 13444 35204 13484
rect 32732 13416 35204 13444
rect 35253 13447 35311 13453
rect 32732 13404 32738 13416
rect 35253 13413 35265 13447
rect 35299 13444 35311 13447
rect 36354 13444 36360 13456
rect 35299 13416 36360 13444
rect 35299 13413 35311 13416
rect 35253 13407 35311 13413
rect 36354 13404 36360 13416
rect 36412 13404 36418 13456
rect 37752 13444 37780 13484
rect 38194 13472 38200 13524
rect 38252 13472 38258 13524
rect 39666 13472 39672 13524
rect 39724 13472 39730 13524
rect 39850 13472 39856 13524
rect 39908 13512 39914 13524
rect 40681 13515 40739 13521
rect 40681 13512 40693 13515
rect 39908 13484 40693 13512
rect 39908 13472 39914 13484
rect 40681 13481 40693 13484
rect 40727 13481 40739 13515
rect 40681 13475 40739 13481
rect 42794 13472 42800 13524
rect 42852 13512 42858 13524
rect 42889 13515 42947 13521
rect 42889 13512 42901 13515
rect 42852 13484 42901 13512
rect 42852 13472 42858 13484
rect 42889 13481 42901 13484
rect 42935 13481 42947 13515
rect 42889 13475 42947 13481
rect 45002 13472 45008 13524
rect 45060 13472 45066 13524
rect 46385 13515 46443 13521
rect 46385 13481 46397 13515
rect 46431 13512 46443 13515
rect 48406 13512 48412 13524
rect 46431 13484 48412 13512
rect 46431 13481 46443 13484
rect 46385 13475 46443 13481
rect 48406 13472 48412 13484
rect 48464 13472 48470 13524
rect 37752 13416 40080 13444
rect 29472 13348 30236 13376
rect 30745 13379 30803 13385
rect 30745 13345 30757 13379
rect 30791 13376 30803 13379
rect 33502 13376 33508 13388
rect 30791 13348 33508 13376
rect 30791 13345 30803 13348
rect 30745 13339 30803 13345
rect 33502 13336 33508 13348
rect 33560 13336 33566 13388
rect 33686 13336 33692 13388
rect 33744 13376 33750 13388
rect 33744 13348 34100 13376
rect 33744 13336 33750 13348
rect 34072 13320 34100 13348
rect 34238 13336 34244 13388
rect 34296 13376 34302 13388
rect 34422 13376 34428 13388
rect 34296 13348 34428 13376
rect 34296 13336 34302 13348
rect 34422 13336 34428 13348
rect 34480 13336 34486 13388
rect 35618 13336 35624 13388
rect 35676 13376 35682 13388
rect 35805 13379 35863 13385
rect 35805 13376 35817 13379
rect 35676 13348 35817 13376
rect 35676 13336 35682 13348
rect 35805 13345 35817 13348
rect 35851 13345 35863 13379
rect 35805 13339 35863 13345
rect 36170 13336 36176 13388
rect 36228 13376 36234 13388
rect 36449 13379 36507 13385
rect 36449 13376 36461 13379
rect 36228 13348 36461 13376
rect 36228 13336 36234 13348
rect 36449 13345 36461 13348
rect 36495 13376 36507 13379
rect 36814 13376 36820 13388
rect 36495 13348 36820 13376
rect 36495 13345 36507 13348
rect 36449 13339 36507 13345
rect 36814 13336 36820 13348
rect 36872 13336 36878 13388
rect 37274 13336 37280 13388
rect 37332 13376 37338 13388
rect 38470 13376 38476 13388
rect 37332 13348 38476 13376
rect 37332 13336 37338 13348
rect 38470 13336 38476 13348
rect 38528 13336 38534 13388
rect 40052 13320 40080 13416
rect 43806 13404 43812 13456
rect 43864 13444 43870 13456
rect 43864 13416 44312 13444
rect 43864 13404 43870 13416
rect 44174 13376 44180 13388
rect 42260 13348 44180 13376
rect 28442 13268 28448 13320
rect 28500 13308 28506 13320
rect 28905 13311 28963 13317
rect 28905 13308 28917 13311
rect 28500 13280 28917 13308
rect 28500 13268 28506 13280
rect 28905 13277 28917 13280
rect 28951 13277 28963 13311
rect 28905 13271 28963 13277
rect 32306 13268 32312 13320
rect 32364 13308 32370 13320
rect 33781 13311 33839 13317
rect 33781 13308 33793 13311
rect 32364 13280 33793 13308
rect 32364 13268 32370 13280
rect 33781 13277 33793 13280
rect 33827 13277 33839 13311
rect 33781 13271 33839 13277
rect 34054 13268 34060 13320
rect 34112 13308 34118 13320
rect 34701 13311 34759 13317
rect 34701 13308 34713 13311
rect 34112 13280 34713 13308
rect 34112 13268 34118 13280
rect 34701 13277 34713 13280
rect 34747 13277 34759 13311
rect 34701 13271 34759 13277
rect 35158 13268 35164 13320
rect 35216 13308 35222 13320
rect 35713 13311 35771 13317
rect 35713 13308 35725 13311
rect 35216 13280 35725 13308
rect 35216 13268 35222 13280
rect 35713 13277 35725 13280
rect 35759 13277 35771 13311
rect 35713 13271 35771 13277
rect 38657 13311 38715 13317
rect 38657 13277 38669 13311
rect 38703 13308 38715 13311
rect 38930 13308 38936 13320
rect 38703 13280 38936 13308
rect 38703 13277 38715 13280
rect 38657 13271 38715 13277
rect 38930 13268 38936 13280
rect 38988 13268 38994 13320
rect 39666 13308 39672 13320
rect 39132 13280 39672 13308
rect 24762 13240 24768 13252
rect 22848 13212 23888 13240
rect 24320 13212 24768 13240
rect 10652 13144 12020 13172
rect 10652 13132 10658 13144
rect 12158 13132 12164 13184
rect 12216 13172 12222 13184
rect 12342 13172 12348 13184
rect 12216 13144 12348 13172
rect 12216 13132 12222 13144
rect 12342 13132 12348 13144
rect 12400 13132 12406 13184
rect 12710 13132 12716 13184
rect 12768 13132 12774 13184
rect 13170 13132 13176 13184
rect 13228 13172 13234 13184
rect 14090 13172 14096 13184
rect 13228 13144 14096 13172
rect 13228 13132 13234 13144
rect 14090 13132 14096 13144
rect 14148 13172 14154 13184
rect 14185 13175 14243 13181
rect 14185 13172 14197 13175
rect 14148 13144 14197 13172
rect 14148 13132 14154 13144
rect 14185 13141 14197 13144
rect 14231 13141 14243 13175
rect 14185 13135 14243 13141
rect 15194 13132 15200 13184
rect 15252 13172 15258 13184
rect 19426 13172 19432 13184
rect 15252 13144 19432 13172
rect 15252 13132 15258 13144
rect 19426 13132 19432 13144
rect 19484 13132 19490 13184
rect 20162 13132 20168 13184
rect 20220 13132 20226 13184
rect 20254 13132 20260 13184
rect 20312 13172 20318 13184
rect 21266 13172 21272 13184
rect 20312 13144 21272 13172
rect 20312 13132 20318 13144
rect 21266 13132 21272 13144
rect 21324 13132 21330 13184
rect 21358 13132 21364 13184
rect 21416 13172 21422 13184
rect 22848 13172 22876 13212
rect 21416 13144 22876 13172
rect 21416 13132 21422 13144
rect 23290 13132 23296 13184
rect 23348 13132 23354 13184
rect 23658 13132 23664 13184
rect 23716 13132 23722 13184
rect 23860 13172 23888 13212
rect 24762 13200 24768 13212
rect 24820 13200 24826 13252
rect 24857 13243 24915 13249
rect 24857 13209 24869 13243
rect 24903 13209 24915 13243
rect 24857 13203 24915 13209
rect 24302 13172 24308 13184
rect 23860 13144 24308 13172
rect 24302 13132 24308 13144
rect 24360 13132 24366 13184
rect 24872 13172 24900 13203
rect 24946 13200 24952 13252
rect 25004 13240 25010 13252
rect 27157 13243 27215 13249
rect 25004 13212 25346 13240
rect 25004 13200 25010 13212
rect 27157 13209 27169 13243
rect 27203 13240 27215 13243
rect 27430 13240 27436 13252
rect 27203 13212 27436 13240
rect 27203 13209 27215 13212
rect 27157 13203 27215 13209
rect 27430 13200 27436 13212
rect 27488 13200 27494 13252
rect 28534 13240 28540 13252
rect 28382 13212 28540 13240
rect 28534 13200 28540 13212
rect 28592 13200 28598 13252
rect 28994 13200 29000 13252
rect 29052 13240 29058 13252
rect 29454 13240 29460 13252
rect 29052 13212 29460 13240
rect 29052 13200 29058 13212
rect 29454 13200 29460 13212
rect 29512 13200 29518 13252
rect 31018 13200 31024 13252
rect 31076 13200 31082 13252
rect 31478 13200 31484 13252
rect 31536 13200 31542 13252
rect 32766 13200 32772 13252
rect 32824 13240 32830 13252
rect 33045 13243 33103 13249
rect 33045 13240 33057 13243
rect 32824 13212 33057 13240
rect 32824 13200 32830 13212
rect 33045 13209 33057 13212
rect 33091 13209 33103 13243
rect 33045 13203 33103 13209
rect 34425 13243 34483 13249
rect 34425 13209 34437 13243
rect 34471 13240 34483 13243
rect 34514 13240 34520 13252
rect 34471 13212 34520 13240
rect 34471 13209 34483 13212
rect 34425 13203 34483 13209
rect 34514 13200 34520 13212
rect 34572 13200 34578 13252
rect 35434 13200 35440 13252
rect 35492 13240 35498 13252
rect 35621 13243 35679 13249
rect 35621 13240 35633 13243
rect 35492 13212 35633 13240
rect 35492 13200 35498 13212
rect 35621 13209 35633 13212
rect 35667 13209 35679 13243
rect 35621 13203 35679 13209
rect 36725 13243 36783 13249
rect 36725 13209 36737 13243
rect 36771 13209 36783 13243
rect 39132 13240 39160 13280
rect 39666 13268 39672 13280
rect 39724 13268 39730 13320
rect 40034 13268 40040 13320
rect 40092 13268 40098 13320
rect 41141 13311 41199 13317
rect 41141 13277 41153 13311
rect 41187 13308 41199 13311
rect 41690 13308 41696 13320
rect 41187 13280 41696 13308
rect 41187 13277 41199 13280
rect 41141 13271 41199 13277
rect 41690 13268 41696 13280
rect 41748 13268 41754 13320
rect 42260 13317 42288 13348
rect 44174 13336 44180 13348
rect 44232 13336 44238 13388
rect 44284 13376 44312 13416
rect 44910 13404 44916 13456
rect 44968 13444 44974 13456
rect 45189 13447 45247 13453
rect 45189 13444 45201 13447
rect 44968 13416 45201 13444
rect 44968 13404 44974 13416
rect 45189 13413 45201 13416
rect 45235 13413 45247 13447
rect 46934 13444 46940 13456
rect 45189 13407 45247 13413
rect 45756 13416 46940 13444
rect 44542 13376 44548 13388
rect 44284 13348 44548 13376
rect 44542 13336 44548 13348
rect 44600 13376 44606 13388
rect 45373 13379 45431 13385
rect 45373 13376 45385 13379
rect 44600 13348 45385 13376
rect 44600 13336 44606 13348
rect 45373 13345 45385 13348
rect 45419 13345 45431 13379
rect 45373 13339 45431 13345
rect 42245 13311 42303 13317
rect 42245 13277 42257 13311
rect 42291 13277 42303 13311
rect 42245 13271 42303 13277
rect 43254 13268 43260 13320
rect 43312 13308 43318 13320
rect 43349 13311 43407 13317
rect 43349 13308 43361 13311
rect 43312 13280 43361 13308
rect 43312 13268 43318 13280
rect 43349 13277 43361 13280
rect 43395 13277 43407 13311
rect 43349 13271 43407 13277
rect 44910 13268 44916 13320
rect 44968 13308 44974 13320
rect 45756 13317 45784 13416
rect 46934 13404 46940 13416
rect 46992 13404 46998 13456
rect 47486 13404 47492 13456
rect 47544 13404 47550 13456
rect 48314 13376 48320 13388
rect 46860 13348 48320 13376
rect 46860 13317 46888 13348
rect 48314 13336 48320 13348
rect 48372 13336 48378 13388
rect 48406 13336 48412 13388
rect 48464 13376 48470 13388
rect 48682 13376 48688 13388
rect 48464 13348 48688 13376
rect 48464 13336 48470 13348
rect 48682 13336 48688 13348
rect 48740 13336 48746 13388
rect 45741 13311 45799 13317
rect 45741 13308 45753 13311
rect 44968 13280 45753 13308
rect 44968 13268 44974 13280
rect 45741 13277 45753 13280
rect 45787 13277 45799 13311
rect 45741 13271 45799 13277
rect 46845 13311 46903 13317
rect 46845 13277 46857 13311
rect 46891 13277 46903 13311
rect 46845 13271 46903 13277
rect 46934 13268 46940 13320
rect 46992 13308 46998 13320
rect 47949 13311 48007 13317
rect 47949 13308 47961 13311
rect 46992 13280 47961 13308
rect 46992 13268 46998 13280
rect 47949 13277 47961 13280
rect 47995 13277 48007 13311
rect 47949 13271 48007 13277
rect 49142 13268 49148 13320
rect 49200 13268 49206 13320
rect 40310 13240 40316 13252
rect 37950 13212 39160 13240
rect 39224 13212 40316 13240
rect 36725 13203 36783 13209
rect 25682 13172 25688 13184
rect 24872 13144 25688 13172
rect 25682 13132 25688 13144
rect 25740 13132 25746 13184
rect 28810 13132 28816 13184
rect 28868 13172 28874 13184
rect 29181 13175 29239 13181
rect 29181 13172 29193 13175
rect 28868 13144 29193 13172
rect 28868 13132 28874 13144
rect 29181 13141 29193 13144
rect 29227 13141 29239 13175
rect 29181 13135 29239 13141
rect 29822 13132 29828 13184
rect 29880 13132 29886 13184
rect 30282 13132 30288 13184
rect 30340 13172 30346 13184
rect 32674 13172 32680 13184
rect 30340 13144 32680 13172
rect 30340 13132 30346 13144
rect 32674 13132 32680 13144
rect 32732 13132 32738 13184
rect 34532 13172 34560 13200
rect 36170 13172 36176 13184
rect 34532 13144 36176 13172
rect 36170 13132 36176 13144
rect 36228 13132 36234 13184
rect 36740 13172 36768 13203
rect 39224 13172 39252 13212
rect 40310 13200 40316 13212
rect 40368 13200 40374 13252
rect 41414 13200 41420 13252
rect 41472 13240 41478 13252
rect 44453 13243 44511 13249
rect 44453 13240 44465 13243
rect 41472 13212 44465 13240
rect 41472 13200 41478 13212
rect 44453 13209 44465 13212
rect 44499 13209 44511 13243
rect 44453 13203 44511 13209
rect 36740 13144 39252 13172
rect 39298 13132 39304 13184
rect 39356 13132 39362 13184
rect 39942 13132 39948 13184
rect 40000 13172 40006 13184
rect 41785 13175 41843 13181
rect 41785 13172 41797 13175
rect 40000 13144 41797 13172
rect 40000 13132 40006 13144
rect 41785 13141 41797 13144
rect 41831 13141 41843 13175
rect 41785 13135 41843 13141
rect 43714 13132 43720 13184
rect 43772 13172 43778 13184
rect 43993 13175 44051 13181
rect 43993 13172 44005 13175
rect 43772 13144 44005 13172
rect 43772 13132 43778 13144
rect 43993 13141 44005 13144
rect 44039 13141 44051 13175
rect 43993 13135 44051 13141
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 3789 12971 3847 12977
rect 3789 12937 3801 12971
rect 3835 12968 3847 12971
rect 3878 12968 3884 12980
rect 3835 12940 3884 12968
rect 3835 12937 3847 12940
rect 3789 12931 3847 12937
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 4893 12971 4951 12977
rect 4893 12937 4905 12971
rect 4939 12968 4951 12971
rect 4982 12968 4988 12980
rect 4939 12940 4988 12968
rect 4939 12937 4951 12940
rect 4893 12931 4951 12937
rect 4982 12928 4988 12940
rect 5040 12928 5046 12980
rect 5994 12928 6000 12980
rect 6052 12928 6058 12980
rect 6362 12928 6368 12980
rect 6420 12968 6426 12980
rect 6457 12971 6515 12977
rect 6457 12968 6469 12971
rect 6420 12940 6469 12968
rect 6420 12928 6426 12940
rect 6457 12937 6469 12940
rect 6503 12937 6515 12971
rect 6457 12931 6515 12937
rect 6822 12928 6828 12980
rect 6880 12928 6886 12980
rect 8846 12928 8852 12980
rect 8904 12928 8910 12980
rect 9766 12928 9772 12980
rect 9824 12968 9830 12980
rect 10873 12971 10931 12977
rect 10873 12968 10885 12971
rect 9824 12940 10885 12968
rect 9824 12928 9830 12940
rect 10873 12937 10885 12940
rect 10919 12937 10931 12971
rect 10873 12931 10931 12937
rect 12069 12971 12127 12977
rect 12069 12937 12081 12971
rect 12115 12937 12127 12971
rect 12069 12931 12127 12937
rect 2869 12903 2927 12909
rect 2869 12869 2881 12903
rect 2915 12900 2927 12903
rect 3050 12900 3056 12912
rect 2915 12872 3056 12900
rect 2915 12869 2927 12872
rect 2869 12863 2927 12869
rect 3050 12860 3056 12872
rect 3108 12860 3114 12912
rect 4614 12860 4620 12912
rect 4672 12900 4678 12912
rect 7745 12903 7803 12909
rect 7745 12900 7757 12903
rect 4672 12872 7757 12900
rect 4672 12860 4678 12872
rect 7745 12869 7757 12872
rect 7791 12869 7803 12903
rect 7745 12863 7803 12869
rect 11146 12860 11152 12912
rect 11204 12900 11210 12912
rect 12084 12900 12112 12931
rect 13446 12928 13452 12980
rect 13504 12928 13510 12980
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 14093 12971 14151 12977
rect 14093 12968 14105 12971
rect 13872 12940 14105 12968
rect 13872 12928 13878 12940
rect 14093 12937 14105 12940
rect 14139 12968 14151 12971
rect 15102 12968 15108 12980
rect 14139 12940 15108 12968
rect 14139 12937 14151 12940
rect 14093 12931 14151 12937
rect 15102 12928 15108 12940
rect 15160 12928 15166 12980
rect 15838 12928 15844 12980
rect 15896 12968 15902 12980
rect 16301 12971 16359 12977
rect 16301 12968 16313 12971
rect 15896 12940 16313 12968
rect 15896 12928 15902 12940
rect 16301 12937 16313 12940
rect 16347 12937 16359 12971
rect 16301 12931 16359 12937
rect 16758 12928 16764 12980
rect 16816 12968 16822 12980
rect 17589 12971 17647 12977
rect 17589 12968 17601 12971
rect 16816 12940 17601 12968
rect 16816 12928 16822 12940
rect 17589 12937 17601 12940
rect 17635 12968 17647 12971
rect 18874 12968 18880 12980
rect 17635 12940 18880 12968
rect 17635 12937 17647 12940
rect 17589 12931 17647 12937
rect 18874 12928 18880 12940
rect 18932 12928 18938 12980
rect 19426 12928 19432 12980
rect 19484 12968 19490 12980
rect 20346 12968 20352 12980
rect 19484 12940 20352 12968
rect 19484 12928 19490 12940
rect 20346 12928 20352 12940
rect 20404 12928 20410 12980
rect 21836 12940 24348 12968
rect 11204 12872 11652 12900
rect 11204 12860 11210 12872
rect 11624 12856 11652 12872
rect 11900 12872 12112 12900
rect 11900 12856 11928 12872
rect 13078 12860 13084 12912
rect 13136 12900 13142 12912
rect 14829 12903 14887 12909
rect 14829 12900 14841 12903
rect 13136 12872 14841 12900
rect 13136 12860 13142 12872
rect 14829 12869 14841 12872
rect 14875 12869 14887 12903
rect 18690 12900 18696 12912
rect 14829 12863 14887 12869
rect 1302 12792 1308 12844
rect 1360 12832 1366 12844
rect 1581 12835 1639 12841
rect 1581 12832 1593 12835
rect 1360 12804 1593 12832
rect 1360 12792 1366 12804
rect 1581 12801 1593 12804
rect 1627 12801 1639 12835
rect 1581 12795 1639 12801
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12832 1915 12835
rect 2038 12832 2044 12844
rect 1903 12804 2044 12832
rect 1903 12801 1915 12804
rect 1857 12795 1915 12801
rect 1596 12764 1624 12795
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 3145 12835 3203 12841
rect 3145 12801 3157 12835
rect 3191 12801 3203 12835
rect 3145 12795 3203 12801
rect 4249 12835 4307 12841
rect 4249 12801 4261 12835
rect 4295 12832 4307 12835
rect 5353 12835 5411 12841
rect 4295 12804 5304 12832
rect 4295 12801 4307 12804
rect 4249 12795 4307 12801
rect 2774 12764 2780 12776
rect 1596 12736 2780 12764
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 3160 12764 3188 12795
rect 4798 12764 4804 12776
rect 3160 12736 4804 12764
rect 4798 12724 4804 12736
rect 4856 12724 4862 12776
rect 5276 12696 5304 12804
rect 5353 12801 5365 12835
rect 5399 12832 5411 12835
rect 5534 12832 5540 12844
rect 5399 12804 5540 12832
rect 5399 12801 5411 12804
rect 5353 12795 5411 12801
rect 5534 12792 5540 12804
rect 5592 12792 5598 12844
rect 7098 12792 7104 12844
rect 7156 12792 7162 12844
rect 8205 12835 8263 12841
rect 8205 12801 8217 12835
rect 8251 12801 8263 12835
rect 8205 12795 8263 12801
rect 6454 12724 6460 12776
rect 6512 12764 6518 12776
rect 6730 12764 6736 12776
rect 6512 12736 6736 12764
rect 6512 12724 6518 12736
rect 6730 12724 6736 12736
rect 6788 12724 6794 12776
rect 8220 12696 8248 12795
rect 9306 12792 9312 12844
rect 9364 12792 9370 12844
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12832 10839 12835
rect 10827 12804 11100 12832
rect 11624 12828 11928 12856
rect 10827 12801 10839 12804
rect 10781 12795 10839 12801
rect 9674 12724 9680 12776
rect 9732 12764 9738 12776
rect 10226 12764 10232 12776
rect 9732 12736 10232 12764
rect 9732 12724 9738 12736
rect 10226 12724 10232 12736
rect 10284 12724 10290 12776
rect 10962 12724 10968 12776
rect 11020 12724 11026 12776
rect 11072 12764 11100 12804
rect 12268 12804 12940 12832
rect 11882 12764 11888 12776
rect 11072 12736 11888 12764
rect 11882 12724 11888 12736
rect 11940 12724 11946 12776
rect 12158 12724 12164 12776
rect 12216 12724 12222 12776
rect 11606 12696 11612 12708
rect 5276 12668 8064 12696
rect 8220 12668 11612 12696
rect 5810 12588 5816 12640
rect 5868 12628 5874 12640
rect 6178 12628 6184 12640
rect 5868 12600 6184 12628
rect 5868 12588 5874 12600
rect 6178 12588 6184 12600
rect 6236 12588 6242 12640
rect 7098 12588 7104 12640
rect 7156 12628 7162 12640
rect 7742 12628 7748 12640
rect 7156 12600 7748 12628
rect 7156 12588 7162 12600
rect 7742 12588 7748 12600
rect 7800 12588 7806 12640
rect 8036 12628 8064 12668
rect 11606 12656 11612 12668
rect 11664 12656 11670 12708
rect 12066 12656 12072 12708
rect 12124 12696 12130 12708
rect 12268 12696 12296 12804
rect 12342 12724 12348 12776
rect 12400 12724 12406 12776
rect 12912 12764 12940 12804
rect 12986 12792 12992 12844
rect 13044 12832 13050 12844
rect 13357 12835 13415 12841
rect 13357 12832 13369 12835
rect 13044 12804 13369 12832
rect 13044 12792 13050 12804
rect 13357 12801 13369 12804
rect 13403 12832 13415 12835
rect 13446 12832 13452 12844
rect 13403 12804 13452 12832
rect 13403 12801 13415 12804
rect 13357 12795 13415 12801
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 14274 12792 14280 12844
rect 14332 12832 14338 12844
rect 14553 12835 14611 12841
rect 14553 12832 14565 12835
rect 14332 12804 14565 12832
rect 14332 12792 14338 12804
rect 14553 12801 14565 12804
rect 14599 12801 14611 12835
rect 14553 12795 14611 12801
rect 15856 12776 15884 12886
rect 16776 12872 18696 12900
rect 16114 12792 16120 12844
rect 16172 12832 16178 12844
rect 16669 12835 16727 12841
rect 16669 12832 16681 12835
rect 16172 12804 16681 12832
rect 16172 12792 16178 12804
rect 16669 12801 16681 12804
rect 16715 12801 16727 12835
rect 16669 12795 16727 12801
rect 13541 12767 13599 12773
rect 13541 12764 13553 12767
rect 12912 12736 13553 12764
rect 13541 12733 13553 12736
rect 13587 12764 13599 12767
rect 13722 12764 13728 12776
rect 13587 12736 13728 12764
rect 13587 12733 13599 12736
rect 13541 12727 13599 12733
rect 13722 12724 13728 12736
rect 13780 12724 13786 12776
rect 15838 12724 15844 12776
rect 15896 12764 15902 12776
rect 16776 12764 16804 12872
rect 18690 12860 18696 12872
rect 18748 12860 18754 12912
rect 19242 12860 19248 12912
rect 19300 12900 19306 12912
rect 21836 12900 21864 12940
rect 19300 12872 21864 12900
rect 19300 12860 19306 12872
rect 22186 12860 22192 12912
rect 22244 12860 22250 12912
rect 23014 12860 23020 12912
rect 23072 12900 23078 12912
rect 23293 12903 23351 12909
rect 23293 12900 23305 12903
rect 23072 12872 23305 12900
rect 23072 12860 23078 12872
rect 23293 12869 23305 12872
rect 23339 12869 23351 12903
rect 23293 12863 23351 12869
rect 23474 12860 23480 12912
rect 23532 12900 23538 12912
rect 24320 12909 24348 12940
rect 24394 12928 24400 12980
rect 24452 12968 24458 12980
rect 24670 12968 24676 12980
rect 24452 12940 24676 12968
rect 24452 12928 24458 12940
rect 24670 12928 24676 12940
rect 24728 12928 24734 12980
rect 26142 12928 26148 12980
rect 26200 12968 26206 12980
rect 27801 12971 27859 12977
rect 27801 12968 27813 12971
rect 26200 12940 27813 12968
rect 26200 12928 26206 12940
rect 27801 12937 27813 12940
rect 27847 12937 27859 12971
rect 29270 12968 29276 12980
rect 27801 12931 27859 12937
rect 29012 12940 29276 12968
rect 24305 12903 24363 12909
rect 23532 12872 24072 12900
rect 23532 12860 23538 12872
rect 17313 12835 17371 12841
rect 17313 12801 17325 12835
rect 17359 12801 17371 12835
rect 17313 12795 17371 12801
rect 15896 12736 16804 12764
rect 17328 12764 17356 12795
rect 17494 12792 17500 12844
rect 17552 12832 17558 12844
rect 17678 12832 17684 12844
rect 17552 12804 17684 12832
rect 17552 12792 17558 12804
rect 17678 12792 17684 12804
rect 17736 12832 17742 12844
rect 17957 12835 18015 12841
rect 17957 12832 17969 12835
rect 17736 12804 17969 12832
rect 17736 12792 17742 12804
rect 17957 12801 17969 12804
rect 18003 12832 18015 12835
rect 19426 12832 19432 12844
rect 18003 12804 19432 12832
rect 18003 12801 18015 12804
rect 17957 12795 18015 12801
rect 19426 12792 19432 12804
rect 19484 12792 19490 12844
rect 19518 12792 19524 12844
rect 19576 12832 19582 12844
rect 19705 12835 19763 12841
rect 19705 12832 19717 12835
rect 19576 12804 19717 12832
rect 19576 12792 19582 12804
rect 19705 12801 19717 12804
rect 19751 12801 19763 12835
rect 19705 12795 19763 12801
rect 21085 12835 21143 12841
rect 21085 12801 21097 12835
rect 21131 12832 21143 12835
rect 22002 12832 22008 12844
rect 21131 12804 22008 12832
rect 21131 12801 21143 12804
rect 21085 12795 21143 12801
rect 22002 12792 22008 12804
rect 22060 12792 22066 12844
rect 23201 12835 23259 12841
rect 23201 12801 23213 12835
rect 23247 12832 23259 12835
rect 23566 12832 23572 12844
rect 23247 12804 23572 12832
rect 23247 12801 23259 12804
rect 23201 12795 23259 12801
rect 23566 12792 23572 12804
rect 23624 12792 23630 12844
rect 24044 12841 24072 12872
rect 24305 12869 24317 12903
rect 24351 12869 24363 12903
rect 24305 12863 24363 12869
rect 28350 12860 28356 12912
rect 28408 12860 28414 12912
rect 28534 12860 28540 12912
rect 28592 12900 28598 12912
rect 29012 12900 29040 12940
rect 29270 12928 29276 12940
rect 29328 12968 29334 12980
rect 30466 12968 30472 12980
rect 29328 12940 30472 12968
rect 29328 12928 29334 12940
rect 30466 12928 30472 12940
rect 30524 12928 30530 12980
rect 31849 12971 31907 12977
rect 31849 12968 31861 12971
rect 30576 12940 31861 12968
rect 30576 12909 30604 12940
rect 31849 12937 31861 12940
rect 31895 12968 31907 12971
rect 34057 12971 34115 12977
rect 31895 12940 33916 12968
rect 31895 12937 31907 12940
rect 31849 12931 31907 12937
rect 30561 12903 30619 12909
rect 28592 12872 29118 12900
rect 28592 12860 28598 12872
rect 30561 12869 30573 12903
rect 30607 12869 30619 12903
rect 30561 12863 30619 12869
rect 31294 12860 31300 12912
rect 31352 12900 31358 12912
rect 31754 12900 31760 12912
rect 31352 12872 31760 12900
rect 31352 12860 31358 12872
rect 31754 12860 31760 12872
rect 31812 12900 31818 12912
rect 31812 12872 33074 12900
rect 31812 12860 31818 12872
rect 24029 12835 24087 12841
rect 24029 12801 24041 12835
rect 24075 12801 24087 12835
rect 24029 12795 24087 12801
rect 25406 12792 25412 12844
rect 25464 12792 25470 12844
rect 26510 12832 26516 12844
rect 26160 12804 26516 12832
rect 17328 12736 18736 12764
rect 15896 12724 15902 12736
rect 12124 12668 12296 12696
rect 12360 12696 12388 12724
rect 13630 12696 13636 12708
rect 12360 12668 13636 12696
rect 12124 12656 12130 12668
rect 13630 12656 13636 12668
rect 13688 12656 13694 12708
rect 16022 12656 16028 12708
rect 16080 12696 16086 12708
rect 17129 12699 17187 12705
rect 17129 12696 17141 12699
rect 16080 12668 17141 12696
rect 16080 12656 16086 12668
rect 17129 12665 17141 12668
rect 17175 12696 17187 12699
rect 18708 12696 18736 12736
rect 19058 12724 19064 12776
rect 19116 12764 19122 12776
rect 19797 12767 19855 12773
rect 19797 12764 19809 12767
rect 19116 12736 19809 12764
rect 19116 12724 19122 12736
rect 19797 12733 19809 12736
rect 19843 12733 19855 12767
rect 19797 12727 19855 12733
rect 19981 12767 20039 12773
rect 19981 12733 19993 12767
rect 20027 12764 20039 12767
rect 20530 12764 20536 12776
rect 20027 12736 20536 12764
rect 20027 12733 20039 12736
rect 19981 12727 20039 12733
rect 20530 12724 20536 12736
rect 20588 12724 20594 12776
rect 21177 12767 21235 12773
rect 21177 12733 21189 12767
rect 21223 12733 21235 12767
rect 21177 12727 21235 12733
rect 17175 12668 18368 12696
rect 18708 12668 19012 12696
rect 17175 12665 17187 12668
rect 17129 12659 17187 12665
rect 9582 12628 9588 12640
rect 8036 12600 9588 12628
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 9950 12588 9956 12640
rect 10008 12588 10014 12640
rect 10410 12588 10416 12640
rect 10468 12588 10474 12640
rect 11514 12588 11520 12640
rect 11572 12628 11578 12640
rect 11701 12631 11759 12637
rect 11701 12628 11713 12631
rect 11572 12600 11713 12628
rect 11572 12588 11578 12600
rect 11701 12597 11713 12600
rect 11747 12597 11759 12631
rect 11701 12591 11759 12597
rect 12989 12631 13047 12637
rect 12989 12597 13001 12631
rect 13035 12628 13047 12631
rect 13446 12628 13452 12640
rect 13035 12600 13452 12628
rect 13035 12597 13047 12600
rect 12989 12591 13047 12597
rect 13446 12588 13452 12600
rect 13504 12588 13510 12640
rect 14185 12631 14243 12637
rect 14185 12597 14197 12631
rect 14231 12628 14243 12631
rect 17678 12628 17684 12640
rect 14231 12600 17684 12628
rect 14231 12597 14243 12600
rect 14185 12591 14243 12597
rect 17678 12588 17684 12600
rect 17736 12588 17742 12640
rect 18340 12628 18368 12668
rect 18874 12628 18880 12640
rect 18340 12600 18880 12628
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 18984 12628 19012 12668
rect 19334 12656 19340 12708
rect 19392 12656 19398 12708
rect 20438 12656 20444 12708
rect 20496 12656 20502 12708
rect 21082 12696 21088 12708
rect 20640 12668 21088 12696
rect 20640 12628 20668 12668
rect 21082 12656 21088 12668
rect 21140 12656 21146 12708
rect 18984 12600 20668 12628
rect 20717 12631 20775 12637
rect 20717 12597 20729 12631
rect 20763 12628 20775 12631
rect 20806 12628 20812 12640
rect 20763 12600 20812 12628
rect 20763 12597 20775 12600
rect 20717 12591 20775 12597
rect 20806 12588 20812 12600
rect 20864 12588 20870 12640
rect 21192 12628 21220 12727
rect 21358 12724 21364 12776
rect 21416 12724 21422 12776
rect 21913 12767 21971 12773
rect 21913 12733 21925 12767
rect 21959 12764 21971 12767
rect 22738 12764 22744 12776
rect 21959 12736 22744 12764
rect 21959 12733 21971 12736
rect 21913 12727 21971 12733
rect 22738 12724 22744 12736
rect 22796 12764 22802 12776
rect 23385 12767 23443 12773
rect 23385 12764 23397 12767
rect 22796 12736 23397 12764
rect 22796 12724 22802 12736
rect 23385 12733 23397 12736
rect 23431 12764 23443 12767
rect 26160 12764 26188 12804
rect 26510 12792 26516 12804
rect 26568 12832 26574 12844
rect 26697 12835 26755 12841
rect 26697 12832 26709 12835
rect 26568 12804 26709 12832
rect 26568 12792 26574 12804
rect 26697 12801 26709 12804
rect 26743 12832 26755 12835
rect 27157 12835 27215 12841
rect 27157 12832 27169 12835
rect 26743 12804 27169 12832
rect 26743 12801 26755 12804
rect 26697 12795 26755 12801
rect 27157 12801 27169 12804
rect 27203 12832 27215 12835
rect 28368 12832 28396 12860
rect 32214 12832 32220 12844
rect 27203 12804 28396 12832
rect 30208 12804 32220 12832
rect 27203 12801 27215 12804
rect 27157 12795 27215 12801
rect 23431 12736 26188 12764
rect 23431 12733 23443 12736
rect 23385 12727 23443 12733
rect 26234 12724 26240 12776
rect 26292 12724 26298 12776
rect 26326 12724 26332 12776
rect 26384 12764 26390 12776
rect 27614 12764 27620 12776
rect 26384 12736 27620 12764
rect 26384 12724 26390 12736
rect 27614 12724 27620 12736
rect 27672 12724 27678 12776
rect 28353 12767 28411 12773
rect 28353 12733 28365 12767
rect 28399 12733 28411 12767
rect 28353 12727 28411 12733
rect 28629 12767 28687 12773
rect 28629 12733 28641 12767
rect 28675 12764 28687 12767
rect 30208 12764 30236 12804
rect 32214 12792 32220 12804
rect 32272 12792 32278 12844
rect 32306 12792 32312 12844
rect 32364 12792 32370 12844
rect 33888 12832 33916 12940
rect 34057 12937 34069 12971
rect 34103 12968 34115 12971
rect 37826 12968 37832 12980
rect 34103 12940 37832 12968
rect 34103 12937 34115 12940
rect 34057 12931 34115 12937
rect 37826 12928 37832 12940
rect 37884 12968 37890 12980
rect 37884 12940 39068 12968
rect 37884 12928 37890 12940
rect 35066 12860 35072 12912
rect 35124 12900 35130 12912
rect 35253 12903 35311 12909
rect 35253 12900 35265 12903
rect 35124 12872 35265 12900
rect 35124 12860 35130 12872
rect 35253 12869 35265 12872
rect 35299 12900 35311 12903
rect 35986 12900 35992 12912
rect 35299 12872 35992 12900
rect 35299 12869 35311 12872
rect 35253 12863 35311 12869
rect 35986 12860 35992 12872
rect 36044 12860 36050 12912
rect 36906 12900 36912 12912
rect 36648 12872 36912 12900
rect 36648 12841 36676 12872
rect 36906 12860 36912 12872
rect 36964 12860 36970 12912
rect 38746 12860 38752 12912
rect 38804 12860 38810 12912
rect 36633 12835 36691 12841
rect 36633 12832 36645 12835
rect 33888 12804 36645 12832
rect 36633 12801 36645 12804
rect 36679 12801 36691 12835
rect 36633 12795 36691 12801
rect 36814 12792 36820 12844
rect 36872 12832 36878 12844
rect 37461 12835 37519 12841
rect 37461 12832 37473 12835
rect 36872 12804 37473 12832
rect 36872 12792 36878 12804
rect 37461 12801 37473 12804
rect 37507 12801 37519 12835
rect 39040 12832 39068 12940
rect 40586 12928 40592 12980
rect 40644 12928 40650 12980
rect 41690 12928 41696 12980
rect 41748 12928 41754 12980
rect 43254 12928 43260 12980
rect 43312 12928 43318 12980
rect 44910 12928 44916 12980
rect 44968 12928 44974 12980
rect 45373 12971 45431 12977
rect 45373 12937 45385 12971
rect 45419 12968 45431 12971
rect 46934 12968 46940 12980
rect 45419 12940 46940 12968
rect 45419 12937 45431 12940
rect 45373 12931 45431 12937
rect 46934 12928 46940 12940
rect 46992 12928 46998 12980
rect 47026 12928 47032 12980
rect 47084 12968 47090 12980
rect 47581 12971 47639 12977
rect 47581 12968 47593 12971
rect 47084 12940 47593 12968
rect 47084 12928 47090 12940
rect 47581 12937 47593 12940
rect 47627 12937 47639 12971
rect 47581 12931 47639 12937
rect 40034 12860 40040 12912
rect 40092 12900 40098 12912
rect 41969 12903 42027 12909
rect 41969 12900 41981 12903
rect 40092 12872 41981 12900
rect 40092 12860 40098 12872
rect 41969 12869 41981 12872
rect 42015 12869 42027 12903
rect 41969 12863 42027 12869
rect 42245 12903 42303 12909
rect 42245 12869 42257 12903
rect 42291 12900 42303 12903
rect 44726 12900 44732 12912
rect 42291 12872 44732 12900
rect 42291 12869 42303 12872
rect 42245 12863 42303 12869
rect 39040 12804 39896 12832
rect 37461 12795 37519 12801
rect 28675 12736 30236 12764
rect 28675 12733 28687 12736
rect 28629 12727 28687 12733
rect 22370 12696 22376 12708
rect 22066 12668 22376 12696
rect 22066 12628 22094 12668
rect 22370 12656 22376 12668
rect 22428 12656 22434 12708
rect 22833 12699 22891 12705
rect 22833 12665 22845 12699
rect 22879 12696 22891 12699
rect 23750 12696 23756 12708
rect 22879 12668 23756 12696
rect 22879 12665 22891 12668
rect 22833 12659 22891 12665
rect 23750 12656 23756 12668
rect 23808 12656 23814 12708
rect 25314 12656 25320 12708
rect 25372 12696 25378 12708
rect 25777 12699 25835 12705
rect 25777 12696 25789 12699
rect 25372 12668 25789 12696
rect 25372 12656 25378 12668
rect 25777 12665 25789 12668
rect 25823 12696 25835 12699
rect 26878 12696 26884 12708
rect 25823 12668 26884 12696
rect 25823 12665 25835 12668
rect 25777 12659 25835 12665
rect 26878 12656 26884 12668
rect 26936 12656 26942 12708
rect 21192 12600 22094 12628
rect 22186 12588 22192 12640
rect 22244 12628 22250 12640
rect 25682 12628 25688 12640
rect 22244 12600 25688 12628
rect 22244 12588 22250 12600
rect 25682 12588 25688 12600
rect 25740 12588 25746 12640
rect 28368 12628 28396 12727
rect 30466 12724 30472 12776
rect 30524 12764 30530 12776
rect 31294 12764 31300 12776
rect 30524 12736 31300 12764
rect 30524 12724 30530 12736
rect 31294 12724 31300 12736
rect 31352 12724 31358 12776
rect 32585 12767 32643 12773
rect 32585 12733 32597 12767
rect 32631 12764 32643 12767
rect 32631 12736 34192 12764
rect 32631 12733 32643 12736
rect 32585 12727 32643 12733
rect 34164 12696 34192 12736
rect 34238 12724 34244 12776
rect 34296 12764 34302 12776
rect 34517 12767 34575 12773
rect 34517 12764 34529 12767
rect 34296 12736 34529 12764
rect 34296 12724 34302 12736
rect 34517 12733 34529 12736
rect 34563 12733 34575 12767
rect 34517 12727 34575 12733
rect 34606 12724 34612 12776
rect 34664 12764 34670 12776
rect 35250 12764 35256 12776
rect 34664 12736 35256 12764
rect 34664 12724 34670 12736
rect 35250 12724 35256 12736
rect 35308 12724 35314 12776
rect 35710 12724 35716 12776
rect 35768 12764 35774 12776
rect 35989 12767 36047 12773
rect 35989 12764 36001 12767
rect 35768 12736 36001 12764
rect 35768 12724 35774 12736
rect 35989 12733 36001 12736
rect 36035 12733 36047 12767
rect 35989 12727 36047 12733
rect 36722 12724 36728 12776
rect 36780 12764 36786 12776
rect 37737 12767 37795 12773
rect 36780 12736 37596 12764
rect 36780 12724 36786 12736
rect 37366 12696 37372 12708
rect 34164 12668 37372 12696
rect 37366 12656 37372 12668
rect 37424 12656 37430 12708
rect 29914 12628 29920 12640
rect 28368 12600 29920 12628
rect 29914 12588 29920 12600
rect 29972 12588 29978 12640
rect 30101 12631 30159 12637
rect 30101 12597 30113 12631
rect 30147 12628 30159 12631
rect 30834 12628 30840 12640
rect 30147 12600 30840 12628
rect 30147 12597 30159 12600
rect 30101 12591 30159 12597
rect 30834 12588 30840 12600
rect 30892 12588 30898 12640
rect 33318 12588 33324 12640
rect 33376 12628 33382 12640
rect 35342 12628 35348 12640
rect 33376 12600 35348 12628
rect 33376 12588 33382 12600
rect 35342 12588 35348 12600
rect 35400 12588 35406 12640
rect 36538 12588 36544 12640
rect 36596 12628 36602 12640
rect 36817 12631 36875 12637
rect 36817 12628 36829 12631
rect 36596 12600 36829 12628
rect 36596 12588 36602 12600
rect 36817 12597 36829 12600
rect 36863 12597 36875 12631
rect 37568 12628 37596 12736
rect 37737 12733 37749 12767
rect 37783 12764 37795 12767
rect 39485 12767 39543 12773
rect 37783 12736 39436 12764
rect 37783 12733 37795 12736
rect 37737 12727 37795 12733
rect 39408 12696 39436 12736
rect 39485 12733 39497 12767
rect 39531 12764 39543 12767
rect 39574 12764 39580 12776
rect 39531 12736 39580 12764
rect 39531 12733 39543 12736
rect 39485 12727 39543 12733
rect 39574 12724 39580 12736
rect 39632 12724 39638 12776
rect 39868 12764 39896 12804
rect 39942 12792 39948 12844
rect 40000 12792 40006 12844
rect 41049 12835 41107 12841
rect 41049 12801 41061 12835
rect 41095 12801 41107 12835
rect 41049 12795 41107 12801
rect 41064 12764 41092 12795
rect 41138 12792 41144 12844
rect 41196 12832 41202 12844
rect 42260 12832 42288 12863
rect 44726 12860 44732 12872
rect 44784 12860 44790 12912
rect 45554 12860 45560 12912
rect 45612 12900 45618 12912
rect 45612 12872 46612 12900
rect 45612 12860 45618 12872
rect 46584 12844 46612 12872
rect 46750 12860 46756 12912
rect 46808 12900 46814 12912
rect 47213 12903 47271 12909
rect 47213 12900 47225 12903
rect 46808 12872 47225 12900
rect 46808 12860 46814 12872
rect 47213 12869 47225 12872
rect 47259 12869 47271 12903
rect 47213 12863 47271 12869
rect 47320 12872 47992 12900
rect 41196 12804 42288 12832
rect 41196 12792 41202 12804
rect 42610 12792 42616 12844
rect 42668 12792 42674 12844
rect 43714 12792 43720 12844
rect 43772 12792 43778 12844
rect 45281 12835 45339 12841
rect 45281 12801 45293 12835
rect 45327 12801 45339 12835
rect 45281 12795 45339 12801
rect 39868 12736 41092 12764
rect 41874 12724 41880 12776
rect 41932 12764 41938 12776
rect 45296 12764 45324 12795
rect 45370 12792 45376 12844
rect 45428 12832 45434 12844
rect 46109 12835 46167 12841
rect 46109 12832 46121 12835
rect 45428 12804 46121 12832
rect 45428 12792 45434 12804
rect 46109 12801 46121 12804
rect 46155 12801 46167 12835
rect 46109 12795 46167 12801
rect 46566 12792 46572 12844
rect 46624 12792 46630 12844
rect 41932 12736 45324 12764
rect 41932 12724 41938 12736
rect 44361 12699 44419 12705
rect 44361 12696 44373 12699
rect 39408 12668 44373 12696
rect 44361 12665 44373 12668
rect 44407 12665 44419 12699
rect 44361 12659 44419 12665
rect 44726 12656 44732 12708
rect 44784 12696 44790 12708
rect 45186 12696 45192 12708
rect 44784 12668 45192 12696
rect 44784 12656 44790 12668
rect 45186 12656 45192 12668
rect 45244 12656 45250 12708
rect 45925 12699 45983 12705
rect 45925 12665 45937 12699
rect 45971 12696 45983 12699
rect 47320 12696 47348 12872
rect 47670 12792 47676 12844
rect 47728 12792 47734 12844
rect 47964 12841 47992 12872
rect 47949 12835 48007 12841
rect 47949 12801 47961 12835
rect 47995 12801 48007 12835
rect 47949 12795 48007 12801
rect 49142 12792 49148 12844
rect 49200 12792 49206 12844
rect 45971 12668 47348 12696
rect 45971 12665 45983 12668
rect 45925 12659 45983 12665
rect 47688 12640 47716 12792
rect 37826 12628 37832 12640
rect 37568 12600 37832 12628
rect 36817 12591 36875 12597
rect 37826 12588 37832 12600
rect 37884 12588 37890 12640
rect 39574 12588 39580 12640
rect 39632 12628 39638 12640
rect 41138 12628 41144 12640
rect 39632 12600 41144 12628
rect 39632 12588 39638 12600
rect 41138 12588 41144 12600
rect 41196 12588 41202 12640
rect 44634 12588 44640 12640
rect 44692 12588 44698 12640
rect 47670 12588 47676 12640
rect 47728 12588 47734 12640
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 2314 12384 2320 12436
rect 2372 12384 2378 12436
rect 2774 12384 2780 12436
rect 2832 12384 2838 12436
rect 6362 12384 6368 12436
rect 6420 12384 6426 12436
rect 7469 12427 7527 12433
rect 7469 12393 7481 12427
rect 7515 12424 7527 12427
rect 7650 12424 7656 12436
rect 7515 12396 7656 12424
rect 7515 12393 7527 12396
rect 7469 12387 7527 12393
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 9858 12384 9864 12436
rect 9916 12384 9922 12436
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10962 12424 10968 12436
rect 10100 12396 10968 12424
rect 10100 12384 10106 12396
rect 10962 12384 10968 12396
rect 11020 12424 11026 12436
rect 11882 12424 11888 12436
rect 11020 12396 11888 12424
rect 11020 12384 11026 12396
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 12989 12427 13047 12433
rect 12989 12424 13001 12427
rect 12032 12396 13001 12424
rect 12032 12384 12038 12396
rect 12989 12393 13001 12396
rect 13035 12393 13047 12427
rect 14642 12424 14648 12436
rect 12989 12387 13047 12393
rect 13188 12396 14648 12424
rect 3973 12359 4031 12365
rect 3973 12325 3985 12359
rect 4019 12356 4031 12359
rect 9674 12356 9680 12368
rect 4019 12328 9680 12356
rect 4019 12325 4031 12328
rect 3973 12319 4031 12325
rect 6380 12300 6408 12328
rect 9674 12316 9680 12328
rect 9732 12316 9738 12368
rect 11606 12316 11612 12368
rect 11664 12356 11670 12368
rect 12066 12356 12072 12368
rect 11664 12328 12072 12356
rect 11664 12316 11670 12328
rect 12066 12316 12072 12328
rect 12124 12316 12130 12368
rect 12713 12359 12771 12365
rect 12713 12325 12725 12359
rect 12759 12356 12771 12359
rect 13078 12356 13084 12368
rect 12759 12328 13084 12356
rect 12759 12325 12771 12328
rect 12713 12319 12771 12325
rect 13078 12316 13084 12328
rect 13136 12356 13142 12368
rect 13188 12356 13216 12396
rect 14642 12384 14648 12396
rect 14700 12384 14706 12436
rect 14734 12384 14740 12436
rect 14792 12424 14798 12436
rect 18598 12424 18604 12436
rect 14792 12396 18604 12424
rect 14792 12384 14798 12396
rect 18598 12384 18604 12396
rect 18656 12384 18662 12436
rect 19613 12427 19671 12433
rect 19613 12393 19625 12427
rect 19659 12424 19671 12427
rect 20162 12424 20168 12436
rect 19659 12396 20168 12424
rect 19659 12393 19671 12396
rect 19613 12387 19671 12393
rect 20162 12384 20168 12396
rect 20220 12384 20226 12436
rect 20438 12384 20444 12436
rect 20496 12424 20502 12436
rect 23934 12424 23940 12436
rect 20496 12396 23940 12424
rect 20496 12384 20502 12396
rect 23934 12384 23940 12396
rect 23992 12384 23998 12436
rect 27062 12424 27068 12436
rect 24688 12396 27068 12424
rect 13998 12356 14004 12368
rect 13136 12328 13216 12356
rect 13464 12328 14004 12356
rect 13136 12316 13142 12328
rect 3418 12248 3424 12300
rect 3476 12248 3482 12300
rect 6362 12248 6368 12300
rect 6420 12248 6426 12300
rect 7190 12248 7196 12300
rect 7248 12288 7254 12300
rect 7466 12288 7472 12300
rect 7248 12260 7472 12288
rect 7248 12248 7254 12260
rect 7466 12248 7472 12260
rect 7524 12248 7530 12300
rect 7558 12248 7564 12300
rect 7616 12288 7622 12300
rect 7616 12260 7972 12288
rect 7616 12248 7622 12260
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12189 1731 12223
rect 1673 12183 1731 12189
rect 3237 12223 3295 12229
rect 3237 12189 3249 12223
rect 3283 12220 3295 12223
rect 3694 12220 3700 12232
rect 3283 12192 3700 12220
rect 3283 12189 3295 12192
rect 3237 12183 3295 12189
rect 1688 12084 1716 12183
rect 3694 12180 3700 12192
rect 3752 12180 3758 12232
rect 3878 12180 3884 12232
rect 3936 12220 3942 12232
rect 4062 12220 4068 12232
rect 3936 12192 4068 12220
rect 3936 12180 3942 12192
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12189 4215 12223
rect 4157 12183 4215 12189
rect 4172 12152 4200 12183
rect 4614 12180 4620 12232
rect 4672 12180 4678 12232
rect 5721 12223 5779 12229
rect 5721 12189 5733 12223
rect 5767 12189 5779 12223
rect 5721 12183 5779 12189
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12220 6883 12223
rect 7834 12220 7840 12232
rect 6871 12192 7840 12220
rect 6871 12189 6883 12192
rect 6825 12183 6883 12189
rect 5736 12152 5764 12183
rect 7834 12180 7840 12192
rect 7892 12180 7898 12232
rect 7944 12229 7972 12260
rect 10318 12248 10324 12300
rect 10376 12288 10382 12300
rect 12986 12288 12992 12300
rect 10376 12260 12992 12288
rect 10376 12248 10382 12260
rect 12986 12248 12992 12260
rect 13044 12248 13050 12300
rect 13464 12288 13492 12328
rect 13998 12316 14004 12328
rect 14056 12316 14062 12368
rect 16025 12359 16083 12365
rect 16025 12325 16037 12359
rect 16071 12356 16083 12359
rect 16114 12356 16120 12368
rect 16071 12328 16120 12356
rect 16071 12325 16083 12328
rect 16025 12319 16083 12325
rect 16114 12316 16120 12328
rect 16172 12356 16178 12368
rect 17034 12356 17040 12368
rect 16172 12328 17040 12356
rect 16172 12316 16178 12328
rect 17034 12316 17040 12328
rect 17092 12316 17098 12368
rect 18690 12316 18696 12368
rect 18748 12356 18754 12368
rect 23661 12359 23719 12365
rect 18748 12328 23612 12356
rect 18748 12316 18754 12328
rect 13188 12260 13492 12288
rect 7929 12223 7987 12229
rect 7929 12189 7941 12223
rect 7975 12189 7987 12223
rect 7929 12183 7987 12189
rect 9217 12223 9275 12229
rect 9217 12189 9229 12223
rect 9263 12189 9275 12223
rect 9217 12183 9275 12189
rect 12529 12223 12587 12229
rect 12529 12189 12541 12223
rect 12575 12220 12587 12223
rect 13188 12220 13216 12260
rect 13538 12248 13544 12300
rect 13596 12248 13602 12300
rect 14016 12288 14044 12316
rect 14550 12288 14556 12300
rect 14016 12260 14556 12288
rect 14550 12248 14556 12260
rect 14608 12248 14614 12300
rect 15286 12248 15292 12300
rect 15344 12288 15350 12300
rect 15344 12260 15700 12288
rect 15344 12248 15350 12260
rect 14274 12220 14280 12232
rect 12575 12192 13216 12220
rect 13280 12192 14280 12220
rect 12575 12189 12587 12192
rect 12529 12183 12587 12189
rect 8846 12152 8852 12164
rect 4172 12124 4660 12152
rect 5736 12124 8852 12152
rect 4632 12096 4660 12124
rect 8846 12112 8852 12124
rect 8904 12112 8910 12164
rect 4062 12084 4068 12096
rect 1688 12056 4068 12084
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 4614 12044 4620 12096
rect 4672 12044 4678 12096
rect 5261 12087 5319 12093
rect 5261 12053 5273 12087
rect 5307 12084 5319 12087
rect 7558 12084 7564 12096
rect 5307 12056 7564 12084
rect 5307 12053 5319 12056
rect 5261 12047 5319 12053
rect 7558 12044 7564 12056
rect 7616 12044 7622 12096
rect 8570 12044 8576 12096
rect 8628 12044 8634 12096
rect 9232 12084 9260 12183
rect 10594 12112 10600 12164
rect 10652 12112 10658 12164
rect 12342 12152 12348 12164
rect 11822 12124 12348 12152
rect 12342 12112 12348 12124
rect 12400 12112 12406 12164
rect 12986 12112 12992 12164
rect 13044 12152 13050 12164
rect 13280 12152 13308 12192
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 15672 12220 15700 12260
rect 16850 12248 16856 12300
rect 16908 12288 16914 12300
rect 18414 12288 18420 12300
rect 16908 12260 18420 12288
rect 16908 12248 16914 12260
rect 18414 12248 18420 12260
rect 18472 12288 18478 12300
rect 18509 12291 18567 12297
rect 18509 12288 18521 12291
rect 18472 12260 18521 12288
rect 18472 12248 18478 12260
rect 18509 12257 18521 12260
rect 18555 12257 18567 12291
rect 18509 12251 18567 12257
rect 18782 12248 18788 12300
rect 18840 12288 18846 12300
rect 20165 12291 20223 12297
rect 20165 12288 20177 12291
rect 18840 12260 20177 12288
rect 18840 12248 18846 12260
rect 20165 12257 20177 12260
rect 20211 12257 20223 12291
rect 20165 12251 20223 12257
rect 20254 12248 20260 12300
rect 20312 12288 20318 12300
rect 23474 12288 23480 12300
rect 20312 12260 23480 12288
rect 20312 12248 20318 12260
rect 23474 12248 23480 12260
rect 23532 12248 23538 12300
rect 23584 12288 23612 12328
rect 23661 12325 23673 12359
rect 23707 12356 23719 12359
rect 24688 12356 24716 12396
rect 27062 12384 27068 12396
rect 27120 12384 27126 12436
rect 28994 12424 29000 12436
rect 27448 12396 29000 12424
rect 23707 12328 24716 12356
rect 23707 12325 23719 12328
rect 23661 12319 23719 12325
rect 24121 12291 24179 12297
rect 24121 12288 24133 12291
rect 23584 12260 24133 12288
rect 24121 12257 24133 12260
rect 24167 12288 24179 12291
rect 24394 12288 24400 12300
rect 24167 12260 24400 12288
rect 24167 12257 24179 12260
rect 24121 12251 24179 12257
rect 24394 12248 24400 12260
rect 24452 12248 24458 12300
rect 27448 12297 27476 12396
rect 28994 12384 29000 12396
rect 29052 12424 29058 12436
rect 30193 12427 30251 12433
rect 30193 12424 30205 12427
rect 29052 12396 30205 12424
rect 29052 12384 29058 12396
rect 30193 12393 30205 12396
rect 30239 12424 30251 12427
rect 30282 12424 30288 12436
rect 30239 12396 30288 12424
rect 30239 12393 30251 12396
rect 30193 12387 30251 12393
rect 30282 12384 30288 12396
rect 30340 12384 30346 12436
rect 30916 12427 30974 12433
rect 30916 12393 30928 12427
rect 30962 12424 30974 12427
rect 40681 12427 40739 12433
rect 40681 12424 40693 12427
rect 30962 12396 36216 12424
rect 30962 12393 30974 12396
rect 30916 12387 30974 12393
rect 27798 12316 27804 12368
rect 27856 12356 27862 12368
rect 30558 12356 30564 12368
rect 27856 12328 30564 12356
rect 27856 12316 27862 12328
rect 30558 12316 30564 12328
rect 30616 12316 30622 12368
rect 36188 12356 36216 12396
rect 37108 12396 40693 12424
rect 37108 12356 37136 12396
rect 40681 12393 40693 12396
rect 40727 12393 40739 12427
rect 40681 12387 40739 12393
rect 42150 12384 42156 12436
rect 42208 12424 42214 12436
rect 42426 12424 42432 12436
rect 42208 12396 42432 12424
rect 42208 12384 42214 12396
rect 42426 12384 42432 12396
rect 42484 12384 42490 12436
rect 44453 12427 44511 12433
rect 44453 12393 44465 12427
rect 44499 12424 44511 12427
rect 45370 12424 45376 12436
rect 44499 12396 45376 12424
rect 44499 12393 44511 12396
rect 44453 12387 44511 12393
rect 45370 12384 45376 12396
rect 45428 12384 45434 12436
rect 36188 12328 37136 12356
rect 37182 12316 37188 12368
rect 37240 12356 37246 12368
rect 41414 12356 41420 12368
rect 37240 12328 38792 12356
rect 37240 12316 37246 12328
rect 24857 12291 24915 12297
rect 24857 12257 24869 12291
rect 24903 12288 24915 12291
rect 27433 12291 27491 12297
rect 24903 12260 27384 12288
rect 24903 12257 24915 12260
rect 24857 12251 24915 12257
rect 15838 12220 15844 12232
rect 15672 12206 15844 12220
rect 15686 12192 15844 12206
rect 15838 12180 15844 12192
rect 15896 12180 15902 12232
rect 16482 12180 16488 12232
rect 16540 12220 16546 12232
rect 16577 12223 16635 12229
rect 16577 12220 16589 12223
rect 16540 12192 16589 12220
rect 16540 12180 16546 12192
rect 16577 12189 16589 12192
rect 16623 12220 16635 12223
rect 19337 12223 19395 12229
rect 19337 12220 19349 12223
rect 16623 12192 19349 12220
rect 16623 12189 16635 12192
rect 16577 12183 16635 12189
rect 19337 12189 19349 12192
rect 19383 12220 19395 12223
rect 20070 12220 20076 12232
rect 19383 12192 20076 12220
rect 19383 12189 19395 12192
rect 19337 12183 19395 12189
rect 20070 12180 20076 12192
rect 20128 12220 20134 12232
rect 20901 12223 20959 12229
rect 20901 12220 20913 12223
rect 20128 12192 20913 12220
rect 20128 12180 20134 12192
rect 20901 12189 20913 12192
rect 20947 12220 20959 12223
rect 22278 12220 22284 12232
rect 20947 12192 22284 12220
rect 20947 12189 20959 12192
rect 20901 12183 20959 12189
rect 22278 12180 22284 12192
rect 22336 12180 22342 12232
rect 23845 12223 23903 12229
rect 23845 12189 23857 12223
rect 23891 12220 23903 12223
rect 23934 12220 23940 12232
rect 23891 12192 23940 12220
rect 23891 12189 23903 12192
rect 23845 12183 23903 12189
rect 23934 12180 23940 12192
rect 23992 12180 23998 12232
rect 24578 12180 24584 12232
rect 24636 12180 24642 12232
rect 27356 12220 27384 12260
rect 27433 12257 27445 12291
rect 27479 12257 27491 12291
rect 27433 12251 27491 12257
rect 27614 12248 27620 12300
rect 27672 12288 27678 12300
rect 27985 12291 28043 12297
rect 27985 12288 27997 12291
rect 27672 12260 27997 12288
rect 27672 12248 27678 12260
rect 27985 12257 27997 12260
rect 28031 12257 28043 12291
rect 27985 12251 28043 12257
rect 28074 12248 28080 12300
rect 28132 12288 28138 12300
rect 28810 12288 28816 12300
rect 28132 12260 28816 12288
rect 28132 12248 28138 12260
rect 28810 12248 28816 12260
rect 28868 12248 28874 12300
rect 29089 12291 29147 12297
rect 29089 12257 29101 12291
rect 29135 12288 29147 12291
rect 29454 12288 29460 12300
rect 29135 12260 29460 12288
rect 29135 12257 29147 12260
rect 29089 12251 29147 12257
rect 29454 12248 29460 12260
rect 29512 12288 29518 12300
rect 30190 12288 30196 12300
rect 29512 12260 30196 12288
rect 29512 12248 29518 12260
rect 30190 12248 30196 12260
rect 30248 12248 30254 12300
rect 32306 12288 32312 12300
rect 30668 12260 32312 12288
rect 29546 12220 29552 12232
rect 27356 12192 29552 12220
rect 29546 12180 29552 12192
rect 29604 12180 29610 12232
rect 29638 12180 29644 12232
rect 29696 12220 29702 12232
rect 29696 12192 30236 12220
rect 29696 12180 29702 12192
rect 30208 12164 30236 12192
rect 30374 12180 30380 12232
rect 30432 12220 30438 12232
rect 30668 12229 30696 12260
rect 32306 12248 32312 12260
rect 32364 12248 32370 12300
rect 33413 12291 33471 12297
rect 33413 12257 33425 12291
rect 33459 12288 33471 12291
rect 34606 12288 34612 12300
rect 33459 12260 34612 12288
rect 33459 12257 33471 12260
rect 33413 12251 33471 12257
rect 34606 12248 34612 12260
rect 34664 12248 34670 12300
rect 35710 12288 35716 12300
rect 34900 12260 35716 12288
rect 30653 12223 30711 12229
rect 30653 12220 30665 12223
rect 30432 12192 30665 12220
rect 30432 12180 30438 12192
rect 30653 12189 30665 12192
rect 30699 12189 30711 12223
rect 30653 12183 30711 12189
rect 33502 12180 33508 12232
rect 33560 12220 33566 12232
rect 34900 12229 34928 12260
rect 35710 12248 35716 12260
rect 35768 12248 35774 12300
rect 35802 12248 35808 12300
rect 35860 12288 35866 12300
rect 36633 12291 36691 12297
rect 36633 12288 36645 12291
rect 35860 12260 36645 12288
rect 35860 12248 35866 12260
rect 36633 12257 36645 12260
rect 36679 12288 36691 12291
rect 37550 12288 37556 12300
rect 36679 12260 37556 12288
rect 36679 12257 36691 12260
rect 36633 12251 36691 12257
rect 37550 12248 37556 12260
rect 37608 12248 37614 12300
rect 37737 12291 37795 12297
rect 37737 12257 37749 12291
rect 37783 12288 37795 12291
rect 38562 12288 38568 12300
rect 37783 12260 38568 12288
rect 37783 12257 37795 12260
rect 37737 12251 37795 12257
rect 38562 12248 38568 12260
rect 38620 12248 38626 12300
rect 38764 12297 38792 12328
rect 38856 12328 41420 12356
rect 38749 12291 38807 12297
rect 38749 12257 38761 12291
rect 38795 12257 38807 12291
rect 38749 12251 38807 12257
rect 34885 12223 34943 12229
rect 34885 12220 34897 12223
rect 33560 12192 34897 12220
rect 33560 12180 33566 12192
rect 34885 12189 34897 12192
rect 34931 12189 34943 12223
rect 34885 12183 34943 12189
rect 36446 12180 36452 12232
rect 36504 12220 36510 12232
rect 37461 12223 37519 12229
rect 36504 12192 37136 12220
rect 36504 12180 36510 12192
rect 13044 12124 13308 12152
rect 13357 12155 13415 12161
rect 13044 12112 13050 12124
rect 13357 12121 13369 12155
rect 13403 12152 13415 12155
rect 13906 12152 13912 12164
rect 13403 12124 13912 12152
rect 13403 12121 13415 12124
rect 13357 12115 13415 12121
rect 13906 12112 13912 12124
rect 13964 12112 13970 12164
rect 13998 12112 14004 12164
rect 14056 12152 14062 12164
rect 14553 12155 14611 12161
rect 14553 12152 14565 12155
rect 14056 12124 14565 12152
rect 14056 12112 14062 12124
rect 14553 12121 14565 12124
rect 14599 12121 14611 12155
rect 14553 12115 14611 12121
rect 15856 12124 16160 12152
rect 10962 12084 10968 12096
rect 9232 12056 10968 12084
rect 10962 12044 10968 12056
rect 11020 12044 11026 12096
rect 11882 12044 11888 12096
rect 11940 12084 11946 12096
rect 12069 12087 12127 12093
rect 12069 12084 12081 12087
rect 11940 12056 12081 12084
rect 11940 12044 11946 12056
rect 12069 12053 12081 12056
rect 12115 12053 12127 12087
rect 12069 12047 12127 12053
rect 13449 12087 13507 12093
rect 13449 12053 13461 12087
rect 13495 12084 13507 12087
rect 15856 12084 15884 12124
rect 13495 12056 15884 12084
rect 16132 12084 16160 12124
rect 16298 12112 16304 12164
rect 16356 12152 16362 12164
rect 17313 12155 17371 12161
rect 17313 12152 17325 12155
rect 16356 12124 17325 12152
rect 16356 12112 16362 12124
rect 17313 12121 17325 12124
rect 17359 12121 17371 12155
rect 17313 12115 17371 12121
rect 18322 12112 18328 12164
rect 18380 12112 18386 12164
rect 18506 12112 18512 12164
rect 18564 12152 18570 12164
rect 19058 12152 19064 12164
rect 18564 12124 19064 12152
rect 18564 12112 18570 12124
rect 19058 12112 19064 12124
rect 19116 12112 19122 12164
rect 19978 12112 19984 12164
rect 20036 12112 20042 12164
rect 20714 12112 20720 12164
rect 20772 12152 20778 12164
rect 20990 12152 20996 12164
rect 20772 12124 20996 12152
rect 20772 12112 20778 12124
rect 20990 12112 20996 12124
rect 21048 12112 21054 12164
rect 21634 12112 21640 12164
rect 21692 12112 21698 12164
rect 23109 12155 23167 12161
rect 23109 12121 23121 12155
rect 23155 12152 23167 12155
rect 24210 12152 24216 12164
rect 23155 12124 24216 12152
rect 23155 12121 23167 12124
rect 23109 12115 23167 12121
rect 24210 12112 24216 12124
rect 24268 12112 24274 12164
rect 25314 12112 25320 12164
rect 25372 12112 25378 12164
rect 28905 12155 28963 12161
rect 28905 12152 28917 12155
rect 26804 12124 28917 12152
rect 17402 12084 17408 12096
rect 16132 12056 17408 12084
rect 13495 12053 13507 12056
rect 13449 12047 13507 12053
rect 17402 12044 17408 12056
rect 17460 12044 17466 12096
rect 17494 12044 17500 12096
rect 17552 12084 17558 12096
rect 17957 12087 18015 12093
rect 17957 12084 17969 12087
rect 17552 12056 17969 12084
rect 17552 12044 17558 12056
rect 17957 12053 17969 12056
rect 18003 12053 18015 12087
rect 17957 12047 18015 12053
rect 18417 12087 18475 12093
rect 18417 12053 18429 12087
rect 18463 12084 18475 12087
rect 18690 12084 18696 12096
rect 18463 12056 18696 12084
rect 18463 12053 18475 12056
rect 18417 12047 18475 12053
rect 18690 12044 18696 12056
rect 18748 12044 18754 12096
rect 18782 12044 18788 12096
rect 18840 12084 18846 12096
rect 18969 12087 19027 12093
rect 18969 12084 18981 12087
rect 18840 12056 18981 12084
rect 18840 12044 18846 12056
rect 18969 12053 18981 12056
rect 19015 12084 19027 12087
rect 19242 12084 19248 12096
rect 19015 12056 19248 12084
rect 19015 12053 19027 12056
rect 18969 12047 19027 12053
rect 19242 12044 19248 12056
rect 19300 12044 19306 12096
rect 20073 12087 20131 12093
rect 20073 12053 20085 12087
rect 20119 12084 20131 12087
rect 20254 12084 20260 12096
rect 20119 12056 20260 12084
rect 20119 12053 20131 12056
rect 20073 12047 20131 12053
rect 20254 12044 20260 12056
rect 20312 12044 20318 12096
rect 22554 12044 22560 12096
rect 22612 12084 22618 12096
rect 23290 12084 23296 12096
rect 22612 12056 23296 12084
rect 22612 12044 22618 12056
rect 23290 12044 23296 12056
rect 23348 12044 23354 12096
rect 24854 12044 24860 12096
rect 24912 12084 24918 12096
rect 26804 12093 26832 12124
rect 28905 12121 28917 12124
rect 28951 12121 28963 12155
rect 28905 12115 28963 12121
rect 29086 12112 29092 12164
rect 29144 12152 29150 12164
rect 29270 12152 29276 12164
rect 29144 12124 29276 12152
rect 29144 12112 29150 12124
rect 29270 12112 29276 12124
rect 29328 12112 29334 12164
rect 29362 12112 29368 12164
rect 29420 12152 29426 12164
rect 29733 12155 29791 12161
rect 29733 12152 29745 12155
rect 29420 12124 29745 12152
rect 29420 12112 29426 12124
rect 29733 12121 29745 12124
rect 29779 12121 29791 12155
rect 29733 12115 29791 12121
rect 30190 12112 30196 12164
rect 30248 12112 30254 12164
rect 31478 12112 31484 12164
rect 31536 12112 31542 12164
rect 33321 12155 33379 12161
rect 33321 12121 33333 12155
rect 33367 12152 33379 12155
rect 33778 12152 33784 12164
rect 33367 12124 33784 12152
rect 33367 12121 33379 12124
rect 33321 12115 33379 12121
rect 33778 12112 33784 12124
rect 33836 12112 33842 12164
rect 35161 12155 35219 12161
rect 35161 12121 35173 12155
rect 35207 12152 35219 12155
rect 35434 12152 35440 12164
rect 35207 12124 35440 12152
rect 35207 12121 35219 12124
rect 35161 12115 35219 12121
rect 35434 12112 35440 12124
rect 35492 12112 35498 12164
rect 36538 12152 36544 12164
rect 36386 12124 36544 12152
rect 26329 12087 26387 12093
rect 26329 12084 26341 12087
rect 24912 12056 26341 12084
rect 24912 12044 24918 12056
rect 26329 12053 26341 12056
rect 26375 12053 26387 12087
rect 26329 12047 26387 12053
rect 26789 12087 26847 12093
rect 26789 12053 26801 12087
rect 26835 12053 26847 12087
rect 26789 12047 26847 12053
rect 27062 12044 27068 12096
rect 27120 12084 27126 12096
rect 27157 12087 27215 12093
rect 27157 12084 27169 12087
rect 27120 12056 27169 12084
rect 27120 12044 27126 12056
rect 27157 12053 27169 12056
rect 27203 12053 27215 12087
rect 27157 12047 27215 12053
rect 27246 12044 27252 12096
rect 27304 12044 27310 12096
rect 27706 12044 27712 12096
rect 27764 12084 27770 12096
rect 27893 12087 27951 12093
rect 27893 12084 27905 12087
rect 27764 12056 27905 12084
rect 27764 12044 27770 12056
rect 27893 12053 27905 12056
rect 27939 12084 27951 12087
rect 28074 12084 28080 12096
rect 27939 12056 28080 12084
rect 27939 12053 27951 12056
rect 27893 12047 27951 12053
rect 28074 12044 28080 12056
rect 28132 12044 28138 12096
rect 28442 12044 28448 12096
rect 28500 12044 28506 12096
rect 28813 12087 28871 12093
rect 28813 12053 28825 12087
rect 28859 12084 28871 12087
rect 29638 12084 29644 12096
rect 28859 12056 29644 12084
rect 28859 12053 28871 12056
rect 28813 12047 28871 12053
rect 29638 12044 29644 12056
rect 29696 12044 29702 12096
rect 32398 12044 32404 12096
rect 32456 12044 32462 12096
rect 32858 12044 32864 12096
rect 32916 12044 32922 12096
rect 33229 12087 33287 12093
rect 33229 12053 33241 12087
rect 33275 12084 33287 12087
rect 33962 12084 33968 12096
rect 33275 12056 33968 12084
rect 33275 12053 33287 12056
rect 33229 12047 33287 12053
rect 33962 12044 33968 12056
rect 34020 12044 34026 12096
rect 34054 12044 34060 12096
rect 34112 12084 34118 12096
rect 34149 12087 34207 12093
rect 34149 12084 34161 12087
rect 34112 12056 34161 12084
rect 34112 12044 34118 12056
rect 34149 12053 34161 12056
rect 34195 12053 34207 12087
rect 34149 12047 34207 12053
rect 34330 12044 34336 12096
rect 34388 12084 34394 12096
rect 34425 12087 34483 12093
rect 34425 12084 34437 12087
rect 34388 12056 34437 12084
rect 34388 12044 34394 12056
rect 34425 12053 34437 12056
rect 34471 12084 34483 12087
rect 34974 12084 34980 12096
rect 34471 12056 34980 12084
rect 34471 12053 34483 12056
rect 34425 12047 34483 12053
rect 34974 12044 34980 12056
rect 35032 12044 35038 12096
rect 35342 12044 35348 12096
rect 35400 12084 35406 12096
rect 35802 12084 35808 12096
rect 35400 12056 35808 12084
rect 35400 12044 35406 12056
rect 35802 12044 35808 12056
rect 35860 12044 35866 12096
rect 35986 12044 35992 12096
rect 36044 12084 36050 12096
rect 36464 12084 36492 12124
rect 36538 12112 36544 12124
rect 36596 12112 36602 12164
rect 37108 12093 37136 12192
rect 37461 12189 37473 12223
rect 37507 12220 37519 12223
rect 38856 12220 38884 12328
rect 41414 12316 41420 12328
rect 41472 12316 41478 12368
rect 43070 12316 43076 12368
rect 43128 12356 43134 12368
rect 43128 12328 45508 12356
rect 43128 12316 43134 12328
rect 38933 12291 38991 12297
rect 38933 12257 38945 12291
rect 38979 12288 38991 12291
rect 39206 12288 39212 12300
rect 38979 12260 39212 12288
rect 38979 12257 38991 12260
rect 38933 12251 38991 12257
rect 39206 12248 39212 12260
rect 39264 12288 39270 12300
rect 45480 12297 45508 12328
rect 45646 12316 45652 12368
rect 45704 12356 45710 12368
rect 47302 12356 47308 12368
rect 45704 12328 47308 12356
rect 45704 12316 45710 12328
rect 47302 12316 47308 12328
rect 47360 12316 47366 12368
rect 45465 12291 45523 12297
rect 39264 12260 43392 12288
rect 39264 12248 39270 12260
rect 37507 12192 38884 12220
rect 39393 12223 39451 12229
rect 37507 12189 37519 12192
rect 37461 12183 37519 12189
rect 39393 12189 39405 12223
rect 39439 12220 39451 12223
rect 39666 12220 39672 12232
rect 39439 12192 39672 12220
rect 39439 12189 39451 12192
rect 39393 12183 39451 12189
rect 39666 12180 39672 12192
rect 39724 12220 39730 12232
rect 39850 12220 39856 12232
rect 39724 12192 39856 12220
rect 39724 12180 39730 12192
rect 39850 12180 39856 12192
rect 39908 12180 39914 12232
rect 40037 12223 40095 12229
rect 40037 12189 40049 12223
rect 40083 12220 40095 12223
rect 40126 12220 40132 12232
rect 40083 12192 40132 12220
rect 40083 12189 40095 12192
rect 40037 12183 40095 12189
rect 40126 12180 40132 12192
rect 40184 12180 40190 12232
rect 41138 12180 41144 12232
rect 41196 12180 41202 12232
rect 41414 12180 41420 12232
rect 41472 12220 41478 12232
rect 43364 12229 43392 12260
rect 45465 12257 45477 12291
rect 45511 12257 45523 12291
rect 45465 12251 45523 12257
rect 46750 12248 46756 12300
rect 46808 12248 46814 12300
rect 49142 12248 49148 12300
rect 49200 12248 49206 12300
rect 42245 12223 42303 12229
rect 42245 12220 42257 12223
rect 41472 12192 42257 12220
rect 41472 12180 41478 12192
rect 42245 12189 42257 12192
rect 42291 12189 42303 12223
rect 42245 12183 42303 12189
rect 43349 12223 43407 12229
rect 43349 12189 43361 12223
rect 43395 12189 43407 12223
rect 44637 12223 44695 12229
rect 44637 12220 44649 12223
rect 43349 12183 43407 12189
rect 43456 12192 44649 12220
rect 37734 12112 37740 12164
rect 37792 12152 37798 12164
rect 42889 12155 42947 12161
rect 42889 12152 42901 12155
rect 37792 12124 42901 12152
rect 37792 12112 37798 12124
rect 42889 12121 42901 12124
rect 42935 12121 42947 12155
rect 42889 12115 42947 12121
rect 36044 12056 36492 12084
rect 37093 12087 37151 12093
rect 36044 12044 36050 12056
rect 37093 12053 37105 12087
rect 37139 12053 37151 12087
rect 37093 12047 37151 12053
rect 37458 12044 37464 12096
rect 37516 12084 37522 12096
rect 37553 12087 37611 12093
rect 37553 12084 37565 12087
rect 37516 12056 37565 12084
rect 37516 12044 37522 12056
rect 37553 12053 37565 12056
rect 37599 12053 37611 12087
rect 37553 12047 37611 12053
rect 38289 12087 38347 12093
rect 38289 12053 38301 12087
rect 38335 12084 38347 12087
rect 38470 12084 38476 12096
rect 38335 12056 38476 12084
rect 38335 12053 38347 12056
rect 38289 12047 38347 12053
rect 38470 12044 38476 12056
rect 38528 12044 38534 12096
rect 38654 12044 38660 12096
rect 38712 12044 38718 12096
rect 39482 12044 39488 12096
rect 39540 12044 39546 12096
rect 39666 12044 39672 12096
rect 39724 12084 39730 12096
rect 41785 12087 41843 12093
rect 41785 12084 41797 12087
rect 39724 12056 41797 12084
rect 39724 12044 39730 12056
rect 41785 12053 41797 12056
rect 41831 12053 41843 12087
rect 41785 12047 41843 12053
rect 42978 12044 42984 12096
rect 43036 12084 43042 12096
rect 43456 12084 43484 12192
rect 44637 12189 44649 12192
rect 44683 12189 44695 12223
rect 44637 12183 44695 12189
rect 45189 12223 45247 12229
rect 45189 12189 45201 12223
rect 45235 12220 45247 12223
rect 45278 12220 45284 12232
rect 45235 12192 45284 12220
rect 45235 12189 45247 12192
rect 45189 12183 45247 12189
rect 45278 12180 45284 12192
rect 45336 12180 45342 12232
rect 46382 12180 46388 12232
rect 46440 12220 46446 12232
rect 46477 12223 46535 12229
rect 46477 12220 46489 12223
rect 46440 12192 46489 12220
rect 46440 12180 46446 12192
rect 46477 12189 46489 12192
rect 46523 12189 46535 12223
rect 46477 12183 46535 12189
rect 46842 12180 46848 12232
rect 46900 12220 46906 12232
rect 47949 12223 48007 12229
rect 47949 12220 47961 12223
rect 46900 12192 47961 12220
rect 46900 12180 46906 12192
rect 47949 12189 47961 12192
rect 47995 12189 48007 12223
rect 47949 12183 48007 12189
rect 44174 12112 44180 12164
rect 44232 12152 44238 12164
rect 45002 12152 45008 12164
rect 44232 12124 45008 12152
rect 44232 12112 44238 12124
rect 45002 12112 45008 12124
rect 45060 12152 45066 12164
rect 50706 12152 50712 12164
rect 45060 12124 50712 12152
rect 45060 12112 45066 12124
rect 50706 12112 50712 12124
rect 50764 12112 50770 12164
rect 43036 12056 43484 12084
rect 43036 12044 43042 12056
rect 43990 12044 43996 12096
rect 44048 12044 44054 12096
rect 45462 12044 45468 12096
rect 45520 12084 45526 12096
rect 47581 12087 47639 12093
rect 47581 12084 47593 12087
rect 45520 12056 47593 12084
rect 45520 12044 45526 12056
rect 47581 12053 47593 12056
rect 47627 12053 47639 12087
rect 47581 12047 47639 12053
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 1762 11840 1768 11892
rect 1820 11840 1826 11892
rect 2590 11840 2596 11892
rect 2648 11840 2654 11892
rect 3602 11880 3608 11892
rect 2746 11852 3608 11880
rect 2501 11815 2559 11821
rect 2501 11781 2513 11815
rect 2547 11812 2559 11815
rect 2746 11812 2774 11852
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 4338 11880 4344 11892
rect 3988 11852 4344 11880
rect 2547 11784 2774 11812
rect 2547 11781 2559 11784
rect 2501 11775 2559 11781
rect 2866 11772 2872 11824
rect 2924 11812 2930 11824
rect 3237 11815 3295 11821
rect 3237 11812 3249 11815
rect 2924 11784 3249 11812
rect 2924 11772 2930 11784
rect 3237 11781 3249 11784
rect 3283 11781 3295 11815
rect 3237 11775 3295 11781
rect 3421 11815 3479 11821
rect 3421 11781 3433 11815
rect 3467 11812 3479 11815
rect 3988 11812 4016 11852
rect 4338 11840 4344 11852
rect 4396 11840 4402 11892
rect 4798 11840 4804 11892
rect 4856 11880 4862 11892
rect 4893 11883 4951 11889
rect 4893 11880 4905 11883
rect 4856 11852 4905 11880
rect 4856 11840 4862 11852
rect 4893 11849 4905 11852
rect 4939 11849 4951 11883
rect 4893 11843 4951 11849
rect 5442 11840 5448 11892
rect 5500 11840 5506 11892
rect 10226 11880 10232 11892
rect 5552 11852 10232 11880
rect 3467 11784 4016 11812
rect 3467 11781 3479 11784
rect 3421 11775 3479 11781
rect 1302 11704 1308 11756
rect 1360 11744 1366 11756
rect 1581 11747 1639 11753
rect 1581 11744 1593 11747
rect 1360 11716 1593 11744
rect 1360 11704 1366 11716
rect 1581 11713 1593 11716
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 1596 11676 1624 11707
rect 1854 11704 1860 11756
rect 1912 11744 1918 11756
rect 3252 11744 3280 11775
rect 4062 11772 4068 11824
rect 4120 11812 4126 11824
rect 5552 11812 5580 11852
rect 10226 11840 10232 11852
rect 10284 11840 10290 11892
rect 13906 11880 13912 11892
rect 10520 11852 13912 11880
rect 4120 11784 5580 11812
rect 4120 11772 4126 11784
rect 6086 11772 6092 11824
rect 6144 11812 6150 11824
rect 6144 11784 7328 11812
rect 6144 11772 6150 11784
rect 3694 11744 3700 11756
rect 1912 11716 3188 11744
rect 3252 11716 3700 11744
rect 1912 11704 1918 11716
rect 2866 11676 2872 11688
rect 1596 11648 2872 11676
rect 2866 11636 2872 11648
rect 2924 11636 2930 11688
rect 3160 11676 3188 11716
rect 3694 11704 3700 11716
rect 3752 11704 3758 11756
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11744 4307 11747
rect 5258 11744 5264 11756
rect 4295 11716 5264 11744
rect 4295 11713 4307 11716
rect 4249 11707 4307 11713
rect 5258 11704 5264 11716
rect 5316 11704 5322 11756
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11744 5871 11747
rect 6457 11747 6515 11753
rect 5859 11716 6132 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 6104 11688 6132 11716
rect 6457 11713 6469 11747
rect 6503 11744 6515 11747
rect 6730 11744 6736 11756
rect 6503 11716 6736 11744
rect 6503 11713 6515 11716
rect 6457 11707 6515 11713
rect 6730 11704 6736 11716
rect 6788 11704 6794 11756
rect 7190 11704 7196 11756
rect 7248 11704 7254 11756
rect 7300 11744 7328 11784
rect 7742 11772 7748 11824
rect 7800 11812 7806 11824
rect 8941 11815 8999 11821
rect 8941 11812 8953 11815
rect 7800 11784 8953 11812
rect 7800 11772 7806 11784
rect 8941 11781 8953 11784
rect 8987 11781 8999 11815
rect 8941 11775 8999 11781
rect 9048 11784 9536 11812
rect 8297 11747 8355 11753
rect 8297 11744 8309 11747
rect 7300 11716 8309 11744
rect 8297 11713 8309 11716
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 5997 11679 6055 11685
rect 5997 11676 6009 11679
rect 3160 11648 6009 11676
rect 5997 11645 6009 11648
rect 6043 11645 6055 11679
rect 5997 11639 6055 11645
rect 6086 11636 6092 11688
rect 6144 11636 6150 11688
rect 7834 11636 7840 11688
rect 7892 11636 7898 11688
rect 3789 11611 3847 11617
rect 3789 11577 3801 11611
rect 3835 11608 3847 11611
rect 4614 11608 4620 11620
rect 3835 11580 4620 11608
rect 3835 11577 3847 11580
rect 3789 11571 3847 11577
rect 4614 11568 4620 11580
rect 4672 11568 4678 11620
rect 5258 11568 5264 11620
rect 5316 11568 5322 11620
rect 5534 11568 5540 11620
rect 5592 11608 5598 11620
rect 9048 11608 9076 11784
rect 9401 11747 9459 11753
rect 9401 11713 9413 11747
rect 9447 11713 9459 11747
rect 9508 11744 9536 11784
rect 9858 11744 9864 11756
rect 9508 11716 9864 11744
rect 9401 11707 9459 11713
rect 5592 11580 9076 11608
rect 9416 11608 9444 11707
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 10520 11753 10548 11852
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 14093 11883 14151 11889
rect 14093 11849 14105 11883
rect 14139 11880 14151 11883
rect 14458 11880 14464 11892
rect 14139 11852 14464 11880
rect 14139 11849 14151 11852
rect 14093 11843 14151 11849
rect 14458 11840 14464 11852
rect 14516 11840 14522 11892
rect 15933 11883 15991 11889
rect 15933 11849 15945 11883
rect 15979 11880 15991 11883
rect 16022 11880 16028 11892
rect 15979 11852 16028 11880
rect 15979 11849 15991 11852
rect 15933 11843 15991 11849
rect 16022 11840 16028 11852
rect 16080 11840 16086 11892
rect 19429 11883 19487 11889
rect 19429 11880 19441 11883
rect 16132 11852 19441 11880
rect 10962 11772 10968 11824
rect 11020 11812 11026 11824
rect 11149 11815 11207 11821
rect 11149 11812 11161 11815
rect 11020 11784 11161 11812
rect 11020 11772 11026 11784
rect 11149 11781 11161 11784
rect 11195 11781 11207 11815
rect 11149 11775 11207 11781
rect 11974 11772 11980 11824
rect 12032 11772 12038 11824
rect 12066 11772 12072 11824
rect 12124 11812 12130 11824
rect 12250 11812 12256 11824
rect 12124 11784 12256 11812
rect 12124 11772 12130 11784
rect 12250 11772 12256 11784
rect 12308 11772 12314 11824
rect 13722 11772 13728 11824
rect 13780 11772 13786 11824
rect 15286 11812 15292 11824
rect 14200 11784 15292 11812
rect 10505 11747 10563 11753
rect 10505 11713 10517 11747
rect 10551 11713 10563 11747
rect 14200 11744 14228 11784
rect 15286 11772 15292 11784
rect 15344 11772 15350 11824
rect 13110 11716 14228 11744
rect 10505 11707 10563 11713
rect 14274 11704 14280 11756
rect 14332 11744 14338 11756
rect 14737 11747 14795 11753
rect 14737 11744 14749 11747
rect 14332 11716 14749 11744
rect 14332 11704 14338 11716
rect 14737 11713 14749 11716
rect 14783 11713 14795 11747
rect 14737 11707 14795 11713
rect 14829 11747 14887 11753
rect 14829 11713 14841 11747
rect 14875 11744 14887 11747
rect 14918 11744 14924 11756
rect 14875 11716 14924 11744
rect 14875 11713 14887 11716
rect 14829 11707 14887 11713
rect 14918 11704 14924 11716
rect 14976 11704 14982 11756
rect 16132 11744 16160 11852
rect 19429 11849 19441 11852
rect 19475 11849 19487 11883
rect 19429 11843 19487 11849
rect 19797 11883 19855 11889
rect 19797 11849 19809 11883
rect 19843 11880 19855 11883
rect 21082 11880 21088 11892
rect 19843 11852 21088 11880
rect 19843 11849 19855 11852
rect 19797 11843 19855 11849
rect 21082 11840 21088 11852
rect 21140 11840 21146 11892
rect 24581 11883 24639 11889
rect 24581 11880 24593 11883
rect 22066 11852 24593 11880
rect 17037 11815 17095 11821
rect 17037 11781 17049 11815
rect 17083 11812 17095 11815
rect 18230 11812 18236 11824
rect 17083 11784 18236 11812
rect 17083 11781 17095 11784
rect 17037 11775 17095 11781
rect 18230 11772 18236 11784
rect 18288 11772 18294 11824
rect 20073 11815 20131 11821
rect 20073 11781 20085 11815
rect 20119 11812 20131 11815
rect 22066 11812 22094 11852
rect 24581 11849 24593 11852
rect 24627 11849 24639 11883
rect 24581 11843 24639 11849
rect 25222 11840 25228 11892
rect 25280 11880 25286 11892
rect 25409 11883 25467 11889
rect 25409 11880 25421 11883
rect 25280 11852 25421 11880
rect 25280 11840 25286 11852
rect 25409 11849 25421 11852
rect 25455 11849 25467 11883
rect 25409 11843 25467 11849
rect 25774 11840 25780 11892
rect 25832 11840 25838 11892
rect 25866 11840 25872 11892
rect 25924 11880 25930 11892
rect 29362 11880 29368 11892
rect 25924 11852 29368 11880
rect 25924 11840 25930 11852
rect 29362 11840 29368 11852
rect 29420 11840 29426 11892
rect 30101 11883 30159 11889
rect 30101 11849 30113 11883
rect 30147 11880 30159 11883
rect 30190 11880 30196 11892
rect 30147 11852 30196 11880
rect 30147 11849 30159 11852
rect 30101 11843 30159 11849
rect 30190 11840 30196 11852
rect 30248 11880 30254 11892
rect 30742 11880 30748 11892
rect 30248 11852 30748 11880
rect 30248 11840 30254 11852
rect 30742 11840 30748 11852
rect 30800 11840 30806 11892
rect 31941 11883 31999 11889
rect 31941 11880 31953 11883
rect 31726 11852 31953 11880
rect 20119 11784 22094 11812
rect 20119 11781 20131 11784
rect 20073 11775 20131 11781
rect 22278 11772 22284 11824
rect 22336 11812 22342 11824
rect 22336 11784 22770 11812
rect 22336 11772 22342 11784
rect 23750 11772 23756 11824
rect 23808 11812 23814 11824
rect 23934 11812 23940 11824
rect 23808 11784 23940 11812
rect 23808 11772 23814 11784
rect 23934 11772 23940 11784
rect 23992 11812 23998 11824
rect 24673 11815 24731 11821
rect 24673 11812 24685 11815
rect 23992 11784 24685 11812
rect 23992 11772 23998 11784
rect 24673 11781 24685 11784
rect 24719 11812 24731 11815
rect 26050 11812 26056 11824
rect 24719 11784 26056 11812
rect 24719 11781 24731 11784
rect 24673 11775 24731 11781
rect 26050 11772 26056 11784
rect 26108 11772 26114 11824
rect 26697 11815 26755 11821
rect 26697 11781 26709 11815
rect 26743 11812 26755 11815
rect 27246 11812 27252 11824
rect 26743 11784 27252 11812
rect 26743 11781 26755 11784
rect 26697 11775 26755 11781
rect 27246 11772 27252 11784
rect 27304 11772 27310 11824
rect 28350 11772 28356 11824
rect 28408 11812 28414 11824
rect 28629 11815 28687 11821
rect 28629 11812 28641 11815
rect 28408 11784 28641 11812
rect 28408 11772 28414 11784
rect 28629 11781 28641 11784
rect 28675 11781 28687 11815
rect 28629 11775 28687 11781
rect 29086 11772 29092 11824
rect 29144 11772 29150 11824
rect 30653 11815 30711 11821
rect 30653 11781 30665 11815
rect 30699 11812 30711 11815
rect 31726 11812 31754 11852
rect 31941 11849 31953 11852
rect 31987 11880 31999 11883
rect 32766 11880 32772 11892
rect 31987 11852 32772 11880
rect 31987 11849 31999 11852
rect 31941 11843 31999 11849
rect 32766 11840 32772 11852
rect 32824 11840 32830 11892
rect 32858 11840 32864 11892
rect 32916 11880 32922 11892
rect 36265 11883 36323 11889
rect 36265 11880 36277 11883
rect 32916 11852 36277 11880
rect 32916 11840 32922 11852
rect 36265 11849 36277 11852
rect 36311 11849 36323 11883
rect 36265 11843 36323 11849
rect 36906 11840 36912 11892
rect 36964 11880 36970 11892
rect 37001 11883 37059 11889
rect 37001 11880 37013 11883
rect 36964 11852 37013 11880
rect 36964 11840 36970 11852
rect 37001 11849 37013 11852
rect 37047 11849 37059 11883
rect 37001 11843 37059 11849
rect 37246 11852 39160 11880
rect 35986 11812 35992 11824
rect 30699 11784 31754 11812
rect 35006 11784 35992 11812
rect 30699 11781 30711 11784
rect 30653 11775 30711 11781
rect 35986 11772 35992 11784
rect 36044 11772 36050 11824
rect 36817 11815 36875 11821
rect 36817 11781 36829 11815
rect 36863 11812 36875 11815
rect 37246 11812 37274 11852
rect 36863 11784 37274 11812
rect 36863 11781 36875 11784
rect 36817 11775 36875 11781
rect 37734 11772 37740 11824
rect 37792 11772 37798 11824
rect 39132 11812 39160 11852
rect 39206 11840 39212 11892
rect 39264 11840 39270 11892
rect 40310 11840 40316 11892
rect 40368 11840 40374 11892
rect 41414 11840 41420 11892
rect 41472 11840 41478 11892
rect 41874 11840 41880 11892
rect 41932 11840 41938 11892
rect 42426 11840 42432 11892
rect 42484 11880 42490 11892
rect 44266 11880 44272 11892
rect 42484 11852 44272 11880
rect 42484 11840 42490 11852
rect 44266 11840 44272 11852
rect 44324 11840 44330 11892
rect 44358 11840 44364 11892
rect 44416 11840 44422 11892
rect 44726 11840 44732 11892
rect 44784 11880 44790 11892
rect 45097 11883 45155 11889
rect 45097 11880 45109 11883
rect 44784 11852 45109 11880
rect 44784 11840 44790 11852
rect 45097 11849 45109 11852
rect 45143 11849 45155 11883
rect 45097 11843 45155 11849
rect 47118 11840 47124 11892
rect 47176 11840 47182 11892
rect 39850 11812 39856 11824
rect 39132 11784 39856 11812
rect 39850 11772 39856 11784
rect 39908 11772 39914 11824
rect 43364 11784 46060 11812
rect 17494 11744 17500 11756
rect 15028 11716 16160 11744
rect 16316 11716 17500 11744
rect 15028 11688 15056 11716
rect 10318 11636 10324 11688
rect 10376 11676 10382 11688
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 10376 11648 11713 11676
rect 10376 11636 10382 11648
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 13354 11676 13360 11688
rect 11701 11639 11759 11645
rect 11808 11648 13360 11676
rect 10778 11608 10784 11620
rect 9416 11580 10784 11608
rect 5592 11568 5598 11580
rect 10778 11568 10784 11580
rect 10836 11568 10842 11620
rect 10962 11568 10968 11620
rect 11020 11608 11026 11620
rect 11808 11608 11836 11648
rect 13354 11636 13360 11648
rect 13412 11636 13418 11688
rect 15010 11636 15016 11688
rect 15068 11636 15074 11688
rect 15562 11636 15568 11688
rect 15620 11676 15626 11688
rect 16025 11679 16083 11685
rect 16025 11676 16037 11679
rect 15620 11648 16037 11676
rect 15620 11636 15626 11648
rect 16025 11645 16037 11648
rect 16071 11645 16083 11679
rect 16025 11639 16083 11645
rect 16206 11636 16212 11688
rect 16264 11636 16270 11688
rect 11020 11580 11836 11608
rect 11020 11568 11026 11580
rect 14182 11568 14188 11620
rect 14240 11608 14246 11620
rect 14369 11611 14427 11617
rect 14369 11608 14381 11611
rect 14240 11580 14381 11608
rect 14240 11568 14246 11580
rect 14369 11577 14381 11580
rect 14415 11577 14427 11611
rect 16316 11608 16344 11716
rect 17494 11704 17500 11716
rect 17552 11704 17558 11756
rect 20714 11744 20720 11756
rect 19090 11716 20720 11744
rect 20714 11704 20720 11716
rect 20772 11704 20778 11756
rect 21082 11704 21088 11756
rect 21140 11704 21146 11756
rect 21818 11744 21824 11756
rect 21376 11716 21824 11744
rect 21376 11688 21404 11716
rect 21818 11704 21824 11716
rect 21876 11704 21882 11756
rect 24394 11704 24400 11756
rect 24452 11744 24458 11756
rect 24452 11716 25544 11744
rect 24452 11704 24458 11716
rect 17681 11679 17739 11685
rect 17681 11645 17693 11679
rect 17727 11645 17739 11679
rect 17681 11639 17739 11645
rect 17957 11679 18015 11685
rect 17957 11645 17969 11679
rect 18003 11676 18015 11679
rect 18003 11648 19104 11676
rect 18003 11645 18015 11648
rect 17957 11639 18015 11645
rect 17696 11608 17724 11639
rect 19076 11620 19104 11648
rect 19242 11636 19248 11688
rect 19300 11676 19306 11688
rect 21177 11679 21235 11685
rect 21177 11676 21189 11679
rect 19300 11648 21189 11676
rect 19300 11636 19306 11648
rect 21177 11645 21189 11648
rect 21223 11676 21235 11679
rect 21266 11676 21272 11688
rect 21223 11648 21272 11676
rect 21223 11645 21235 11648
rect 21177 11639 21235 11645
rect 21266 11636 21272 11648
rect 21324 11636 21330 11688
rect 21358 11636 21364 11688
rect 21416 11636 21422 11688
rect 21634 11636 21640 11688
rect 21692 11676 21698 11688
rect 22005 11679 22063 11685
rect 22005 11676 22017 11679
rect 21692 11648 22017 11676
rect 21692 11636 21698 11648
rect 22005 11645 22017 11648
rect 22051 11645 22063 11679
rect 22005 11639 22063 11645
rect 22281 11679 22339 11685
rect 22281 11645 22293 11679
rect 22327 11676 22339 11679
rect 23934 11676 23940 11688
rect 22327 11648 23940 11676
rect 22327 11645 22339 11648
rect 22281 11639 22339 11645
rect 23934 11636 23940 11648
rect 23992 11636 23998 11688
rect 24765 11679 24823 11685
rect 24765 11645 24777 11679
rect 24811 11676 24823 11679
rect 25038 11676 25044 11688
rect 24811 11648 25044 11676
rect 24811 11645 24823 11648
rect 24765 11639 24823 11645
rect 25038 11636 25044 11648
rect 25096 11676 25102 11688
rect 25406 11676 25412 11688
rect 25096 11648 25412 11676
rect 25096 11636 25102 11648
rect 25406 11636 25412 11648
rect 25464 11636 25470 11688
rect 25516 11676 25544 11716
rect 25590 11704 25596 11756
rect 25648 11744 25654 11756
rect 27525 11747 27583 11753
rect 25648 11716 26004 11744
rect 25648 11704 25654 11716
rect 25976 11685 26004 11716
rect 27525 11713 27537 11747
rect 27571 11713 27583 11747
rect 27525 11707 27583 11713
rect 25869 11679 25927 11685
rect 25869 11676 25881 11679
rect 25516 11648 25881 11676
rect 25869 11645 25881 11648
rect 25915 11645 25927 11679
rect 25869 11639 25927 11645
rect 25961 11679 26019 11685
rect 25961 11645 25973 11679
rect 26007 11645 26019 11679
rect 25961 11639 26019 11645
rect 14369 11571 14427 11577
rect 14936 11580 16344 11608
rect 16776 11580 17724 11608
rect 3878 11500 3884 11552
rect 3936 11500 3942 11552
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 6549 11543 6607 11549
rect 6549 11540 6561 11543
rect 4396 11512 6561 11540
rect 4396 11500 4402 11512
rect 6549 11509 6561 11512
rect 6595 11540 6607 11543
rect 7374 11540 7380 11552
rect 6595 11512 7380 11540
rect 6595 11509 6607 11512
rect 6549 11503 6607 11509
rect 7374 11500 7380 11512
rect 7432 11500 7438 11552
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 10045 11543 10103 11549
rect 10045 11540 10057 11543
rect 9456 11512 10057 11540
rect 9456 11500 9462 11512
rect 10045 11509 10057 11512
rect 10091 11509 10103 11543
rect 10045 11503 10103 11509
rect 11054 11500 11060 11552
rect 11112 11540 11118 11552
rect 11330 11540 11336 11552
rect 11112 11512 11336 11540
rect 11112 11500 11118 11512
rect 11330 11500 11336 11512
rect 11388 11500 11394 11552
rect 12434 11500 12440 11552
rect 12492 11540 12498 11552
rect 13078 11540 13084 11552
rect 12492 11512 13084 11540
rect 12492 11500 12498 11512
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 13354 11500 13360 11552
rect 13412 11540 13418 11552
rect 14936 11540 14964 11580
rect 16776 11552 16804 11580
rect 19058 11568 19064 11620
rect 19116 11568 19122 11620
rect 20438 11608 20444 11620
rect 19168 11580 20444 11608
rect 13412 11512 14964 11540
rect 15565 11543 15623 11549
rect 13412 11500 13418 11512
rect 15565 11509 15577 11543
rect 15611 11540 15623 11543
rect 16666 11540 16672 11552
rect 15611 11512 16672 11540
rect 15611 11509 15623 11512
rect 15565 11503 15623 11509
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 16758 11500 16764 11552
rect 16816 11500 16822 11552
rect 17218 11500 17224 11552
rect 17276 11540 17282 11552
rect 17770 11540 17776 11552
rect 17276 11512 17776 11540
rect 17276 11500 17282 11512
rect 17770 11500 17776 11512
rect 17828 11500 17834 11552
rect 17954 11500 17960 11552
rect 18012 11540 18018 11552
rect 19168 11540 19196 11580
rect 20438 11568 20444 11580
rect 20496 11568 20502 11620
rect 20717 11611 20775 11617
rect 20717 11577 20729 11611
rect 20763 11608 20775 11611
rect 20990 11608 20996 11620
rect 20763 11580 20996 11608
rect 20763 11577 20775 11580
rect 20717 11571 20775 11577
rect 20990 11568 20996 11580
rect 21048 11568 21054 11620
rect 23658 11568 23664 11620
rect 23716 11608 23722 11620
rect 24213 11611 24271 11617
rect 24213 11608 24225 11611
rect 23716 11580 24225 11608
rect 23716 11568 23722 11580
rect 24213 11577 24225 11580
rect 24259 11577 24271 11611
rect 25884 11608 25912 11639
rect 26418 11608 26424 11620
rect 25884 11580 26424 11608
rect 24213 11571 24271 11577
rect 26418 11568 26424 11580
rect 26476 11568 26482 11620
rect 27338 11568 27344 11620
rect 27396 11608 27402 11620
rect 27540 11608 27568 11707
rect 29914 11704 29920 11756
rect 29972 11744 29978 11756
rect 31389 11747 31447 11753
rect 31389 11744 31401 11747
rect 29972 11716 31401 11744
rect 29972 11704 29978 11716
rect 31389 11713 31401 11716
rect 31435 11713 31447 11747
rect 31389 11707 31447 11713
rect 32674 11704 32680 11756
rect 32732 11704 32738 11756
rect 35802 11704 35808 11756
rect 35860 11744 35866 11756
rect 36173 11747 36231 11753
rect 36173 11744 36185 11747
rect 35860 11716 36185 11744
rect 35860 11704 35866 11716
rect 36173 11713 36185 11716
rect 36219 11713 36231 11747
rect 36173 11707 36231 11713
rect 38838 11704 38844 11756
rect 38896 11704 38902 11756
rect 39669 11747 39727 11753
rect 39669 11713 39681 11747
rect 39715 11744 39727 11747
rect 40218 11744 40224 11756
rect 39715 11716 40224 11744
rect 39715 11713 39727 11716
rect 39669 11707 39727 11713
rect 40218 11704 40224 11716
rect 40276 11704 40282 11756
rect 40586 11704 40592 11756
rect 40644 11744 40650 11756
rect 40773 11747 40831 11753
rect 40773 11744 40785 11747
rect 40644 11716 40785 11744
rect 40644 11704 40650 11716
rect 40773 11713 40785 11716
rect 40819 11713 40831 11747
rect 40773 11707 40831 11713
rect 41506 11704 41512 11756
rect 41564 11744 41570 11756
rect 42061 11747 42119 11753
rect 42061 11744 42073 11747
rect 41564 11716 42073 11744
rect 41564 11704 41570 11716
rect 42061 11713 42073 11716
rect 42107 11713 42119 11747
rect 42061 11707 42119 11713
rect 42150 11704 42156 11756
rect 42208 11744 42214 11756
rect 42705 11747 42763 11753
rect 42705 11744 42717 11747
rect 42208 11716 42717 11744
rect 42208 11704 42214 11716
rect 42705 11713 42717 11716
rect 42751 11713 42763 11747
rect 42705 11707 42763 11713
rect 42889 11747 42947 11753
rect 42889 11713 42901 11747
rect 42935 11744 42947 11747
rect 43364 11744 43392 11784
rect 42935 11716 43392 11744
rect 43441 11747 43499 11753
rect 42935 11713 42947 11716
rect 42889 11707 42947 11713
rect 43441 11713 43453 11747
rect 43487 11744 43499 11747
rect 43487 11716 43852 11744
rect 43487 11713 43499 11716
rect 43441 11707 43499 11713
rect 27614 11636 27620 11688
rect 27672 11636 27678 11688
rect 27798 11636 27804 11688
rect 27856 11636 27862 11688
rect 28353 11679 28411 11685
rect 28353 11645 28365 11679
rect 28399 11645 28411 11679
rect 28353 11639 28411 11645
rect 27706 11608 27712 11620
rect 27396 11580 27712 11608
rect 27396 11568 27402 11580
rect 27706 11568 27712 11580
rect 27764 11568 27770 11620
rect 18012 11512 19196 11540
rect 18012 11500 18018 11512
rect 19334 11500 19340 11552
rect 19392 11540 19398 11552
rect 19610 11540 19616 11552
rect 19392 11512 19616 11540
rect 19392 11500 19398 11512
rect 19610 11500 19616 11512
rect 19668 11500 19674 11552
rect 19886 11500 19892 11552
rect 19944 11540 19950 11552
rect 22278 11540 22284 11552
rect 19944 11512 22284 11540
rect 19944 11500 19950 11512
rect 22278 11500 22284 11512
rect 22336 11500 22342 11552
rect 22462 11500 22468 11552
rect 22520 11540 22526 11552
rect 23753 11543 23811 11549
rect 23753 11540 23765 11543
rect 22520 11512 23765 11540
rect 22520 11500 22526 11512
rect 23753 11509 23765 11512
rect 23799 11509 23811 11543
rect 23753 11503 23811 11509
rect 24946 11500 24952 11552
rect 25004 11540 25010 11552
rect 26513 11543 26571 11549
rect 26513 11540 26525 11543
rect 25004 11512 26525 11540
rect 25004 11500 25010 11512
rect 26513 11509 26525 11512
rect 26559 11540 26571 11543
rect 27062 11540 27068 11552
rect 26559 11512 27068 11540
rect 26559 11509 26571 11512
rect 26513 11503 26571 11509
rect 27062 11500 27068 11512
rect 27120 11500 27126 11552
rect 27154 11500 27160 11552
rect 27212 11500 27218 11552
rect 27246 11500 27252 11552
rect 27304 11540 27310 11552
rect 28368 11540 28396 11639
rect 28626 11636 28632 11688
rect 28684 11676 28690 11688
rect 30190 11676 30196 11688
rect 28684 11648 30196 11676
rect 28684 11636 28690 11648
rect 30190 11636 30196 11648
rect 30248 11636 30254 11688
rect 31846 11636 31852 11688
rect 31904 11676 31910 11688
rect 32769 11679 32827 11685
rect 32769 11676 32781 11679
rect 31904 11648 32781 11676
rect 31904 11636 31910 11648
rect 32769 11645 32781 11648
rect 32815 11645 32827 11679
rect 32769 11639 32827 11645
rect 32861 11679 32919 11685
rect 32861 11645 32873 11679
rect 32907 11645 32919 11679
rect 32861 11639 32919 11645
rect 29914 11568 29920 11620
rect 29972 11608 29978 11620
rect 32876 11608 32904 11639
rect 33502 11636 33508 11688
rect 33560 11636 33566 11688
rect 33778 11636 33784 11688
rect 33836 11636 33842 11688
rect 34514 11636 34520 11688
rect 34572 11676 34578 11688
rect 35253 11679 35311 11685
rect 35253 11676 35265 11679
rect 34572 11648 35265 11676
rect 34572 11636 34578 11648
rect 35253 11645 35265 11648
rect 35299 11645 35311 11679
rect 35253 11639 35311 11645
rect 35894 11636 35900 11688
rect 35952 11676 35958 11688
rect 36449 11679 36507 11685
rect 36449 11676 36461 11679
rect 35952 11648 36461 11676
rect 35952 11636 35958 11648
rect 36449 11645 36461 11648
rect 36495 11645 36507 11679
rect 36449 11639 36507 11645
rect 36538 11636 36544 11688
rect 36596 11676 36602 11688
rect 37182 11676 37188 11688
rect 36596 11648 37188 11676
rect 36596 11636 36602 11648
rect 37182 11636 37188 11648
rect 37240 11636 37246 11688
rect 37461 11679 37519 11685
rect 37461 11645 37473 11679
rect 37507 11645 37519 11679
rect 37461 11639 37519 11645
rect 29972 11580 32904 11608
rect 29972 11568 29978 11580
rect 35710 11568 35716 11620
rect 35768 11608 35774 11620
rect 37476 11608 37504 11639
rect 37734 11636 37740 11688
rect 37792 11676 37798 11688
rect 42978 11676 42984 11688
rect 37792 11648 42984 11676
rect 37792 11636 37798 11648
rect 42978 11636 42984 11648
rect 43036 11636 43042 11688
rect 43824 11676 43852 11716
rect 44174 11704 44180 11756
rect 44232 11704 44238 11756
rect 44910 11704 44916 11756
rect 44968 11704 44974 11756
rect 45370 11704 45376 11756
rect 45428 11744 45434 11756
rect 45925 11747 45983 11753
rect 45925 11744 45937 11747
rect 45428 11716 45937 11744
rect 45428 11704 45434 11716
rect 45925 11713 45937 11716
rect 45971 11713 45983 11747
rect 46032 11744 46060 11784
rect 46106 11772 46112 11824
rect 46164 11812 46170 11824
rect 47581 11815 47639 11821
rect 47581 11812 47593 11815
rect 46164 11784 47593 11812
rect 46164 11772 46170 11784
rect 47581 11781 47593 11784
rect 47627 11781 47639 11815
rect 47581 11775 47639 11781
rect 49142 11772 49148 11824
rect 49200 11772 49206 11824
rect 46842 11744 46848 11756
rect 46032 11716 46848 11744
rect 45925 11707 45983 11713
rect 46842 11704 46848 11716
rect 46900 11704 46906 11756
rect 46934 11704 46940 11756
rect 46992 11704 46998 11756
rect 47026 11704 47032 11756
rect 47084 11744 47090 11756
rect 47949 11747 48007 11753
rect 47949 11744 47961 11747
rect 47084 11716 47961 11744
rect 47084 11704 47090 11716
rect 47949 11713 47961 11716
rect 47995 11713 48007 11747
rect 47949 11707 48007 11713
rect 45186 11676 45192 11688
rect 43824 11648 45192 11676
rect 45186 11636 45192 11648
rect 45244 11636 45250 11688
rect 45649 11679 45707 11685
rect 45649 11645 45661 11679
rect 45695 11645 45707 11679
rect 46952 11676 46980 11704
rect 50798 11676 50804 11688
rect 46952 11648 50804 11676
rect 45649 11639 45707 11645
rect 35768 11580 37504 11608
rect 35768 11568 35774 11580
rect 41690 11568 41696 11620
rect 41748 11608 41754 11620
rect 43070 11608 43076 11620
rect 41748 11580 43076 11608
rect 41748 11568 41754 11580
rect 43070 11568 43076 11580
rect 43128 11568 43134 11620
rect 45462 11608 45468 11620
rect 43732 11580 45468 11608
rect 29730 11540 29736 11552
rect 27304 11512 29736 11540
rect 27304 11500 27310 11512
rect 29730 11500 29736 11512
rect 29788 11500 29794 11552
rect 30926 11500 30932 11552
rect 30984 11540 30990 11552
rect 31110 11540 31116 11552
rect 30984 11512 31116 11540
rect 30984 11500 30990 11512
rect 31110 11500 31116 11512
rect 31168 11500 31174 11552
rect 32309 11543 32367 11549
rect 32309 11509 32321 11543
rect 32355 11540 32367 11543
rect 35618 11540 35624 11552
rect 32355 11512 35624 11540
rect 32355 11509 32367 11512
rect 32309 11503 32367 11509
rect 35618 11500 35624 11512
rect 35676 11500 35682 11552
rect 35805 11543 35863 11549
rect 35805 11509 35817 11543
rect 35851 11540 35863 11543
rect 39758 11540 39764 11552
rect 35851 11512 39764 11540
rect 35851 11509 35863 11512
rect 35805 11503 35863 11509
rect 39758 11500 39764 11512
rect 39816 11500 39822 11552
rect 42426 11500 42432 11552
rect 42484 11540 42490 11552
rect 43625 11543 43683 11549
rect 43625 11540 43637 11543
rect 42484 11512 43637 11540
rect 42484 11500 42490 11512
rect 43625 11509 43637 11512
rect 43671 11540 43683 11543
rect 43732 11540 43760 11580
rect 45462 11568 45468 11580
rect 45520 11568 45526 11620
rect 43671 11512 43760 11540
rect 43671 11509 43683 11512
rect 43625 11503 43683 11509
rect 44266 11500 44272 11552
rect 44324 11540 44330 11552
rect 45664 11540 45692 11639
rect 50798 11636 50804 11648
rect 50856 11636 50862 11688
rect 47118 11540 47124 11552
rect 44324 11512 47124 11540
rect 44324 11500 44330 11512
rect 47118 11500 47124 11512
rect 47176 11500 47182 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 1765 11339 1823 11345
rect 1765 11305 1777 11339
rect 1811 11336 1823 11339
rect 1811 11308 3280 11336
rect 1811 11305 1823 11308
rect 1765 11299 1823 11305
rect 2682 11228 2688 11280
rect 2740 11228 2746 11280
rect 3252 11268 3280 11308
rect 3326 11296 3332 11348
rect 3384 11296 3390 11348
rect 3694 11296 3700 11348
rect 3752 11336 3758 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 3752 11308 3801 11336
rect 3752 11296 3758 11308
rect 3789 11305 3801 11308
rect 3835 11305 3847 11339
rect 3789 11299 3847 11305
rect 4430 11296 4436 11348
rect 4488 11296 4494 11348
rect 5166 11296 5172 11348
rect 5224 11296 5230 11348
rect 5718 11296 5724 11348
rect 5776 11296 5782 11348
rect 6270 11296 6276 11348
rect 6328 11296 6334 11348
rect 8938 11296 8944 11348
rect 8996 11296 9002 11348
rect 9306 11296 9312 11348
rect 9364 11296 9370 11348
rect 10321 11339 10379 11345
rect 10321 11305 10333 11339
rect 10367 11336 10379 11339
rect 13998 11336 14004 11348
rect 10367 11308 14004 11336
rect 10367 11305 10379 11308
rect 10321 11299 10379 11305
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 14277 11339 14335 11345
rect 14277 11305 14289 11339
rect 14323 11336 14335 11339
rect 14458 11336 14464 11348
rect 14323 11308 14464 11336
rect 14323 11305 14335 11308
rect 14277 11299 14335 11305
rect 14458 11296 14464 11308
rect 14516 11336 14522 11348
rect 14826 11336 14832 11348
rect 14516 11308 14832 11336
rect 14516 11296 14522 11308
rect 14826 11296 14832 11308
rect 14884 11296 14890 11348
rect 18141 11339 18199 11345
rect 18141 11305 18153 11339
rect 18187 11336 18199 11339
rect 18506 11336 18512 11348
rect 18187 11308 18512 11336
rect 18187 11305 18199 11308
rect 18141 11299 18199 11305
rect 18506 11296 18512 11308
rect 18564 11296 18570 11348
rect 18598 11296 18604 11348
rect 18656 11296 18662 11348
rect 18782 11336 18788 11348
rect 18708 11308 18788 11336
rect 5534 11268 5540 11280
rect 3252 11240 5540 11268
rect 5534 11228 5540 11240
rect 5592 11228 5598 11280
rect 5629 11271 5687 11277
rect 5629 11237 5641 11271
rect 5675 11268 5687 11271
rect 9858 11268 9864 11280
rect 5675 11240 9864 11268
rect 5675 11237 5687 11240
rect 5629 11231 5687 11237
rect 2516 11172 5028 11200
rect 1578 11092 1584 11144
rect 1636 11092 1642 11144
rect 2516 11141 2544 11172
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11101 2559 11135
rect 2501 11095 2559 11101
rect 4338 11092 4344 11144
rect 4396 11092 4402 11144
rect 2774 11024 2780 11076
rect 2832 11064 2838 11076
rect 3237 11067 3295 11073
rect 3237 11064 3249 11067
rect 2832 11036 3249 11064
rect 2832 11024 2838 11036
rect 3237 11033 3249 11036
rect 3283 11033 3295 11067
rect 5000 11064 5028 11172
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11132 5135 11135
rect 5644 11132 5672 11231
rect 9858 11228 9864 11240
rect 9916 11228 9922 11280
rect 12989 11271 13047 11277
rect 12989 11237 13001 11271
rect 13035 11268 13047 11271
rect 14918 11268 14924 11280
rect 13035 11240 14924 11268
rect 13035 11237 13047 11240
rect 12989 11231 13047 11237
rect 14918 11228 14924 11240
rect 14976 11228 14982 11280
rect 15194 11228 15200 11280
rect 15252 11268 15258 11280
rect 15252 11240 16344 11268
rect 15252 11228 15258 11240
rect 8573 11203 8631 11209
rect 8573 11200 8585 11203
rect 6840 11172 8585 11200
rect 5123 11104 5672 11132
rect 6181 11135 6239 11141
rect 5123 11101 5135 11104
rect 5077 11095 5135 11101
rect 6181 11101 6193 11135
rect 6227 11132 6239 11135
rect 6454 11132 6460 11144
rect 6227 11104 6460 11132
rect 6227 11101 6239 11104
rect 6181 11095 6239 11101
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 6840 11141 6868 11172
rect 8573 11169 8585 11172
rect 8619 11169 8631 11203
rect 8573 11163 8631 11169
rect 8938 11160 8944 11212
rect 8996 11200 9002 11212
rect 9122 11200 9128 11212
rect 8996 11172 9128 11200
rect 8996 11160 9002 11172
rect 9122 11160 9128 11172
rect 9180 11160 9186 11212
rect 10042 11200 10048 11212
rect 9600 11172 10048 11200
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11101 6883 11135
rect 6825 11095 6883 11101
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11132 7987 11135
rect 9600 11132 9628 11172
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 12250 11160 12256 11212
rect 12308 11200 12314 11212
rect 12529 11203 12587 11209
rect 12529 11200 12541 11203
rect 12308 11172 12541 11200
rect 12308 11160 12314 11172
rect 12529 11169 12541 11172
rect 12575 11169 12587 11203
rect 12529 11163 12587 11169
rect 12710 11160 12716 11212
rect 12768 11200 12774 11212
rect 13449 11203 13507 11209
rect 13449 11200 13461 11203
rect 12768 11172 13461 11200
rect 12768 11160 12774 11172
rect 13449 11169 13461 11172
rect 13495 11169 13507 11203
rect 13449 11163 13507 11169
rect 13633 11203 13691 11209
rect 13633 11169 13645 11203
rect 13679 11200 13691 11203
rect 13722 11200 13728 11212
rect 13679 11172 13728 11200
rect 13679 11169 13691 11172
rect 13633 11163 13691 11169
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 14642 11160 14648 11212
rect 14700 11200 14706 11212
rect 15013 11203 15071 11209
rect 15013 11200 15025 11203
rect 14700 11172 15025 11200
rect 14700 11160 14706 11172
rect 15013 11169 15025 11172
rect 15059 11169 15071 11203
rect 15013 11163 15071 11169
rect 15105 11203 15163 11209
rect 15105 11169 15117 11203
rect 15151 11200 15163 11203
rect 15470 11200 15476 11212
rect 15151 11172 15476 11200
rect 15151 11169 15163 11172
rect 15105 11163 15163 11169
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 16316 11209 16344 11240
rect 16850 11228 16856 11280
rect 16908 11268 16914 11280
rect 16945 11271 17003 11277
rect 16945 11268 16957 11271
rect 16908 11240 16957 11268
rect 16908 11228 16914 11240
rect 16945 11237 16957 11240
rect 16991 11237 17003 11271
rect 16945 11231 17003 11237
rect 18414 11228 18420 11280
rect 18472 11268 18478 11280
rect 18616 11268 18644 11296
rect 18472 11240 18644 11268
rect 18472 11228 18478 11240
rect 16301 11203 16359 11209
rect 16301 11169 16313 11203
rect 16347 11169 16359 11203
rect 16301 11163 16359 11169
rect 17589 11203 17647 11209
rect 17589 11169 17601 11203
rect 17635 11200 17647 11203
rect 18506 11200 18512 11212
rect 17635 11172 18512 11200
rect 17635 11169 17647 11172
rect 17589 11163 17647 11169
rect 18506 11160 18512 11172
rect 18564 11160 18570 11212
rect 18598 11160 18604 11212
rect 18656 11160 18662 11212
rect 18708 11209 18736 11308
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 19426 11296 19432 11348
rect 19484 11336 19490 11348
rect 19886 11336 19892 11348
rect 19484 11308 19892 11336
rect 19484 11296 19490 11308
rect 19886 11296 19892 11308
rect 19944 11296 19950 11348
rect 20070 11296 20076 11348
rect 20128 11296 20134 11348
rect 20441 11339 20499 11345
rect 20441 11305 20453 11339
rect 20487 11336 20499 11339
rect 20622 11336 20628 11348
rect 20487 11308 20628 11336
rect 20487 11305 20499 11308
rect 20441 11299 20499 11305
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 24946 11336 24952 11348
rect 21744 11308 24952 11336
rect 21744 11268 21772 11308
rect 24946 11296 24952 11308
rect 25004 11296 25010 11348
rect 25222 11296 25228 11348
rect 25280 11336 25286 11348
rect 26326 11336 26332 11348
rect 25280 11308 26332 11336
rect 25280 11296 25286 11308
rect 26326 11296 26332 11308
rect 26384 11296 26390 11348
rect 27144 11339 27202 11345
rect 27144 11305 27156 11339
rect 27190 11336 27202 11339
rect 27706 11336 27712 11348
rect 27190 11308 27712 11336
rect 27190 11305 27202 11308
rect 27144 11299 27202 11305
rect 27706 11296 27712 11308
rect 27764 11296 27770 11348
rect 29546 11296 29552 11348
rect 29604 11336 29610 11348
rect 30377 11339 30435 11345
rect 30377 11336 30389 11339
rect 29604 11308 30389 11336
rect 29604 11296 29610 11308
rect 30377 11305 30389 11308
rect 30423 11305 30435 11339
rect 32766 11336 32772 11348
rect 30377 11299 30435 11305
rect 30484 11308 32772 11336
rect 19306 11240 21772 11268
rect 18693 11203 18751 11209
rect 18693 11169 18705 11203
rect 18739 11169 18751 11203
rect 19306 11200 19334 11240
rect 23382 11228 23388 11280
rect 23440 11228 23446 11280
rect 28629 11271 28687 11277
rect 28629 11237 28641 11271
rect 28675 11268 28687 11271
rect 29914 11268 29920 11280
rect 28675 11240 29920 11268
rect 28675 11237 28687 11240
rect 28629 11231 28687 11237
rect 29914 11228 29920 11240
rect 29972 11228 29978 11280
rect 18693 11163 18751 11169
rect 18800 11172 19334 11200
rect 21085 11203 21143 11209
rect 7975 11104 9628 11132
rect 9677 11135 9735 11141
rect 7975 11101 7987 11104
rect 7929 11095 7987 11101
rect 9677 11101 9689 11135
rect 9723 11132 9735 11135
rect 10226 11132 10232 11144
rect 9723 11104 10232 11132
rect 9723 11101 9735 11104
rect 9677 11095 9735 11101
rect 10226 11092 10232 11104
rect 10284 11092 10290 11144
rect 10778 11092 10784 11144
rect 10836 11092 10842 11144
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 13357 11135 13415 11141
rect 13357 11132 13369 11135
rect 12860 11104 13369 11132
rect 12860 11092 12866 11104
rect 13357 11101 13369 11104
rect 13403 11101 13415 11135
rect 13357 11095 13415 11101
rect 14921 11135 14979 11141
rect 14921 11101 14933 11135
rect 14967 11132 14979 11135
rect 16390 11132 16396 11144
rect 14967 11104 16396 11132
rect 14967 11101 14979 11104
rect 14921 11095 14979 11101
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 17954 11132 17960 11144
rect 17236 11104 17960 11132
rect 7374 11064 7380 11076
rect 5000 11036 7380 11064
rect 3237 11027 3295 11033
rect 7374 11024 7380 11036
rect 7432 11024 7438 11076
rect 7469 11067 7527 11073
rect 7469 11033 7481 11067
rect 7515 11064 7527 11067
rect 11057 11067 11115 11073
rect 11057 11064 11069 11067
rect 7515 11036 11069 11064
rect 7515 11033 7527 11036
rect 7469 11027 7527 11033
rect 11057 11033 11069 11036
rect 11103 11033 11115 11067
rect 12342 11064 12348 11076
rect 12282 11036 12348 11064
rect 11057 11027 11115 11033
rect 12342 11024 12348 11036
rect 12400 11064 12406 11076
rect 13906 11064 13912 11076
rect 12400 11036 13912 11064
rect 12400 11024 12406 11036
rect 13906 11024 13912 11036
rect 13964 11024 13970 11076
rect 14182 11024 14188 11076
rect 14240 11064 14246 11076
rect 14240 11036 16068 11064
rect 14240 11024 14246 11036
rect 1946 10956 1952 11008
rect 2004 10996 2010 11008
rect 5258 10996 5264 11008
rect 2004 10968 5264 10996
rect 2004 10956 2010 10968
rect 5258 10956 5264 10968
rect 5316 10956 5322 11008
rect 6914 10956 6920 11008
rect 6972 10996 6978 11008
rect 12434 10996 12440 11008
rect 6972 10968 12440 10996
rect 6972 10956 6978 10968
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 14553 10999 14611 11005
rect 14553 10965 14565 10999
rect 14599 10996 14611 10999
rect 14642 10996 14648 11008
rect 14599 10968 14648 10996
rect 14599 10965 14611 10968
rect 14553 10959 14611 10965
rect 14642 10956 14648 10968
rect 14700 10956 14706 11008
rect 15746 10956 15752 11008
rect 15804 10956 15810 11008
rect 16040 10996 16068 11036
rect 16114 11024 16120 11076
rect 16172 11024 16178 11076
rect 17236 11064 17264 11104
rect 17954 11092 17960 11104
rect 18012 11092 18018 11144
rect 18800 11132 18828 11172
rect 21085 11169 21097 11203
rect 21131 11200 21143 11203
rect 21358 11200 21364 11212
rect 21131 11172 21364 11200
rect 21131 11169 21143 11172
rect 21085 11163 21143 11169
rect 21358 11160 21364 11172
rect 21416 11160 21422 11212
rect 22646 11160 22652 11212
rect 22704 11200 22710 11212
rect 23400 11200 23428 11228
rect 22704 11172 23428 11200
rect 22704 11160 22710 11172
rect 24578 11160 24584 11212
rect 24636 11200 24642 11212
rect 26786 11200 26792 11212
rect 24636 11172 26792 11200
rect 24636 11160 24642 11172
rect 26786 11160 26792 11172
rect 26844 11200 26850 11212
rect 26881 11203 26939 11209
rect 26881 11200 26893 11203
rect 26844 11172 26893 11200
rect 26844 11160 26850 11172
rect 26881 11169 26893 11172
rect 26927 11200 26939 11203
rect 27246 11200 27252 11212
rect 26927 11172 27252 11200
rect 26927 11169 26939 11172
rect 26881 11163 26939 11169
rect 27246 11160 27252 11172
rect 27304 11160 27310 11212
rect 29086 11200 29092 11212
rect 28644 11172 29092 11200
rect 28644 11144 28672 11172
rect 29086 11160 29092 11172
rect 29144 11160 29150 11212
rect 29270 11160 29276 11212
rect 29328 11200 29334 11212
rect 30484 11200 30512 11308
rect 32766 11296 32772 11308
rect 32824 11296 32830 11348
rect 34882 11336 34888 11348
rect 32968 11308 34888 11336
rect 32214 11228 32220 11280
rect 32272 11268 32278 11280
rect 32968 11268 32996 11308
rect 34882 11296 34888 11308
rect 34940 11296 34946 11348
rect 35066 11296 35072 11348
rect 35124 11296 35130 11348
rect 35158 11296 35164 11348
rect 35216 11336 35222 11348
rect 35253 11339 35311 11345
rect 35253 11336 35265 11339
rect 35216 11308 35265 11336
rect 35216 11296 35222 11308
rect 35253 11305 35265 11308
rect 35299 11305 35311 11339
rect 35253 11299 35311 11305
rect 35529 11339 35587 11345
rect 35529 11305 35541 11339
rect 35575 11336 35587 11339
rect 35986 11336 35992 11348
rect 35575 11308 35992 11336
rect 35575 11305 35587 11308
rect 35529 11299 35587 11305
rect 35986 11296 35992 11308
rect 36044 11296 36050 11348
rect 38562 11336 38568 11348
rect 36096 11308 38568 11336
rect 32272 11240 32996 11268
rect 33045 11271 33103 11277
rect 32272 11228 32278 11240
rect 33045 11237 33057 11271
rect 33091 11268 33103 11271
rect 34054 11268 34060 11280
rect 33091 11240 34060 11268
rect 33091 11237 33103 11240
rect 33045 11231 33103 11237
rect 34054 11228 34060 11240
rect 34112 11228 34118 11280
rect 29328 11172 30512 11200
rect 29328 11160 29334 11172
rect 32122 11160 32128 11212
rect 32180 11200 32186 11212
rect 33505 11203 33563 11209
rect 33505 11200 33517 11203
rect 32180 11172 33517 11200
rect 32180 11160 32186 11172
rect 33505 11169 33517 11172
rect 33551 11169 33563 11203
rect 33505 11163 33563 11169
rect 33597 11203 33655 11209
rect 33597 11169 33609 11203
rect 33643 11169 33655 11203
rect 34900 11200 34928 11296
rect 34974 11228 34980 11280
rect 35032 11268 35038 11280
rect 36096 11268 36124 11308
rect 38562 11296 38568 11308
rect 38620 11296 38626 11348
rect 39114 11296 39120 11348
rect 39172 11296 39178 11348
rect 39485 11339 39543 11345
rect 39485 11305 39497 11339
rect 39531 11336 39543 11339
rect 39850 11336 39856 11348
rect 39531 11308 39856 11336
rect 39531 11305 39543 11308
rect 39485 11299 39543 11305
rect 39850 11296 39856 11308
rect 39908 11296 39914 11348
rect 40586 11336 40592 11348
rect 40052 11308 40592 11336
rect 35032 11240 36124 11268
rect 35032 11228 35038 11240
rect 37550 11228 37556 11280
rect 37608 11268 37614 11280
rect 40052 11268 40080 11308
rect 40586 11296 40592 11308
rect 40644 11296 40650 11348
rect 41782 11296 41788 11348
rect 41840 11336 41846 11348
rect 42702 11336 42708 11348
rect 41840 11308 42708 11336
rect 41840 11296 41846 11308
rect 42702 11296 42708 11308
rect 42760 11296 42766 11348
rect 42981 11339 43039 11345
rect 42981 11305 42993 11339
rect 43027 11336 43039 11339
rect 43438 11336 43444 11348
rect 43027 11308 43444 11336
rect 43027 11305 43039 11308
rect 42981 11299 43039 11305
rect 43438 11296 43444 11308
rect 43496 11296 43502 11348
rect 44542 11336 44548 11348
rect 44008 11308 44548 11336
rect 37608 11240 40080 11268
rect 37608 11228 37614 11240
rect 41874 11228 41880 11280
rect 41932 11268 41938 11280
rect 44008 11268 44036 11308
rect 44542 11296 44548 11308
rect 44600 11336 44606 11348
rect 44821 11339 44879 11345
rect 44821 11336 44833 11339
rect 44600 11308 44833 11336
rect 44600 11296 44606 11308
rect 44821 11305 44833 11308
rect 44867 11305 44879 11339
rect 45278 11336 45284 11348
rect 44821 11299 44879 11305
rect 45020 11308 45284 11336
rect 41932 11240 44036 11268
rect 41932 11228 41938 11240
rect 44726 11228 44732 11280
rect 44784 11268 44790 11280
rect 45020 11277 45048 11308
rect 45278 11296 45284 11308
rect 45336 11296 45342 11348
rect 46566 11296 46572 11348
rect 46624 11336 46630 11348
rect 46753 11339 46811 11345
rect 46753 11336 46765 11339
rect 46624 11308 46765 11336
rect 46624 11296 46630 11308
rect 46753 11305 46765 11308
rect 46799 11305 46811 11339
rect 46753 11299 46811 11305
rect 47394 11296 47400 11348
rect 47452 11296 47458 11348
rect 45005 11271 45063 11277
rect 45005 11268 45017 11271
rect 44784 11240 45017 11268
rect 44784 11228 44790 11240
rect 45005 11237 45017 11240
rect 45051 11237 45063 11271
rect 45005 11231 45063 11237
rect 45186 11228 45192 11280
rect 45244 11268 45250 11280
rect 48498 11268 48504 11280
rect 45244 11240 48504 11268
rect 45244 11228 45250 11240
rect 48498 11228 48504 11240
rect 48556 11228 48562 11280
rect 35250 11200 35256 11212
rect 34900 11172 35256 11200
rect 33597 11163 33655 11169
rect 18156 11104 18828 11132
rect 16224 11036 17264 11064
rect 16224 11005 16252 11036
rect 17310 11024 17316 11076
rect 17368 11024 17374 11076
rect 16209 10999 16267 11005
rect 16209 10996 16221 10999
rect 16040 10968 16221 10996
rect 16209 10965 16221 10968
rect 16255 10965 16267 10999
rect 16209 10959 16267 10965
rect 16942 10956 16948 11008
rect 17000 10996 17006 11008
rect 17405 10999 17463 11005
rect 17405 10996 17417 10999
rect 17000 10968 17417 10996
rect 17000 10956 17006 10968
rect 17405 10965 17417 10968
rect 17451 10965 17463 10999
rect 17405 10959 17463 10965
rect 17678 10956 17684 11008
rect 17736 10996 17742 11008
rect 18156 10996 18184 11104
rect 18966 11092 18972 11144
rect 19024 11132 19030 11144
rect 19426 11132 19432 11144
rect 19024 11104 19432 11132
rect 19024 11092 19030 11104
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 19613 11135 19671 11141
rect 19613 11101 19625 11135
rect 19659 11132 19671 11135
rect 19702 11132 19708 11144
rect 19659 11104 19708 11132
rect 19659 11101 19671 11104
rect 19613 11095 19671 11101
rect 19702 11092 19708 11104
rect 19760 11092 19766 11144
rect 21634 11092 21640 11144
rect 21692 11092 21698 11144
rect 28626 11132 28632 11144
rect 28290 11104 28632 11132
rect 28626 11092 28632 11104
rect 28684 11092 28690 11144
rect 29733 11135 29791 11141
rect 29733 11101 29745 11135
rect 29779 11101 29791 11135
rect 29733 11095 29791 11101
rect 18230 11024 18236 11076
rect 18288 11064 18294 11076
rect 20809 11067 20867 11073
rect 20809 11064 20821 11067
rect 18288 11036 20821 11064
rect 18288 11024 18294 11036
rect 20809 11033 20821 11036
rect 20855 11033 20867 11067
rect 20809 11027 20867 11033
rect 20901 11067 20959 11073
rect 20901 11033 20913 11067
rect 20947 11064 20959 11067
rect 21818 11064 21824 11076
rect 20947 11036 21824 11064
rect 20947 11033 20959 11036
rect 20901 11027 20959 11033
rect 21818 11024 21824 11036
rect 21876 11024 21882 11076
rect 21910 11024 21916 11076
rect 21968 11024 21974 11076
rect 22370 11064 22376 11076
rect 22066 11036 22376 11064
rect 18509 10999 18567 11005
rect 18509 10996 18521 10999
rect 17736 10968 18521 10996
rect 17736 10956 17742 10968
rect 18509 10965 18521 10968
rect 18555 10965 18567 10999
rect 18509 10959 18567 10965
rect 19242 10956 19248 11008
rect 19300 10996 19306 11008
rect 19429 10999 19487 11005
rect 19429 10996 19441 10999
rect 19300 10968 19441 10996
rect 19300 10956 19306 10968
rect 19429 10965 19441 10968
rect 19475 10965 19487 10999
rect 19429 10959 19487 10965
rect 20714 10956 20720 11008
rect 20772 10996 20778 11008
rect 22066 10996 22094 11036
rect 22370 11024 22376 11036
rect 22428 11024 22434 11076
rect 23845 11067 23903 11073
rect 23845 11033 23857 11067
rect 23891 11064 23903 11067
rect 24857 11067 24915 11073
rect 23891 11036 24808 11064
rect 23891 11033 23903 11036
rect 23845 11027 23903 11033
rect 20772 10968 22094 10996
rect 24780 10996 24808 11036
rect 24857 11033 24869 11067
rect 24903 11064 24915 11067
rect 25130 11064 25136 11076
rect 24903 11036 25136 11064
rect 24903 11033 24915 11036
rect 24857 11027 24915 11033
rect 25130 11024 25136 11036
rect 25188 11024 25194 11076
rect 25406 11024 25412 11076
rect 25464 11024 25470 11076
rect 29748 11064 29776 11095
rect 29822 11092 29828 11144
rect 29880 11132 29886 11144
rect 30282 11132 30288 11144
rect 29880 11104 30288 11132
rect 29880 11092 29886 11104
rect 30282 11092 30288 11104
rect 30340 11132 30346 11144
rect 30837 11135 30895 11141
rect 30837 11132 30849 11135
rect 30340 11104 30849 11132
rect 30340 11092 30346 11104
rect 30837 11101 30849 11104
rect 30883 11101 30895 11135
rect 30837 11095 30895 11101
rect 33410 11092 33416 11144
rect 33468 11092 33474 11144
rect 29012 11036 29776 11064
rect 29012 11008 29040 11036
rect 30742 11024 30748 11076
rect 30800 11064 30806 11076
rect 31113 11067 31171 11073
rect 31113 11064 31125 11067
rect 30800 11036 31125 11064
rect 30800 11024 30806 11036
rect 31113 11033 31125 11036
rect 31159 11033 31171 11067
rect 31113 11027 31171 11033
rect 31754 11024 31760 11076
rect 31812 11024 31818 11076
rect 33612 11064 33640 11163
rect 35250 11160 35256 11172
rect 35308 11200 35314 11212
rect 35621 11203 35679 11209
rect 35621 11200 35633 11203
rect 35308 11172 35633 11200
rect 35308 11160 35314 11172
rect 35621 11169 35633 11172
rect 35667 11169 35679 11203
rect 35621 11163 35679 11169
rect 35710 11160 35716 11212
rect 35768 11200 35774 11212
rect 35989 11203 36047 11209
rect 35989 11200 36001 11203
rect 35768 11172 36001 11200
rect 35768 11160 35774 11172
rect 35989 11169 36001 11172
rect 36035 11169 36047 11203
rect 35989 11163 36047 11169
rect 36265 11203 36323 11209
rect 36265 11169 36277 11203
rect 36311 11200 36323 11203
rect 41785 11203 41843 11209
rect 41785 11200 41797 11203
rect 36311 11172 41797 11200
rect 36311 11169 36323 11172
rect 36265 11163 36323 11169
rect 41785 11169 41797 11172
rect 41831 11169 41843 11203
rect 41785 11163 41843 11169
rect 41966 11160 41972 11212
rect 42024 11200 42030 11212
rect 43901 11203 43959 11209
rect 43901 11200 43913 11203
rect 42024 11172 43913 11200
rect 42024 11160 42030 11172
rect 43901 11169 43913 11172
rect 43947 11169 43959 11203
rect 43901 11163 43959 11169
rect 44174 11160 44180 11212
rect 44232 11200 44238 11212
rect 45925 11203 45983 11209
rect 45925 11200 45937 11203
rect 44232 11172 45937 11200
rect 44232 11160 44238 11172
rect 45925 11169 45937 11172
rect 45971 11169 45983 11203
rect 45925 11163 45983 11169
rect 46842 11160 46848 11212
rect 46900 11200 46906 11212
rect 46900 11172 47992 11200
rect 46900 11160 46906 11172
rect 34146 11092 34152 11144
rect 34204 11092 34210 11144
rect 35158 11092 35164 11144
rect 35216 11132 35222 11144
rect 35802 11132 35808 11144
rect 35216 11104 35808 11132
rect 35216 11092 35222 11104
rect 35802 11092 35808 11104
rect 35860 11092 35866 11144
rect 37274 11092 37280 11144
rect 37332 11132 37338 11144
rect 37332 11104 38148 11132
rect 37332 11092 37338 11104
rect 32784 11036 33640 11064
rect 24946 10996 24952 11008
rect 24780 10968 24952 10996
rect 20772 10956 20778 10968
rect 24946 10956 24952 10968
rect 25004 10956 25010 11008
rect 28994 10956 29000 11008
rect 29052 10956 29058 11008
rect 32582 10956 32588 11008
rect 32640 10996 32646 11008
rect 32784 10996 32812 11036
rect 37642 11024 37648 11076
rect 37700 11064 37706 11076
rect 38013 11067 38071 11073
rect 38013 11064 38025 11067
rect 37700 11036 38025 11064
rect 37700 11024 37706 11036
rect 38013 11033 38025 11036
rect 38059 11033 38071 11067
rect 38120 11064 38148 11104
rect 38286 11092 38292 11144
rect 38344 11132 38350 11144
rect 38473 11135 38531 11141
rect 38473 11132 38485 11135
rect 38344 11104 38485 11132
rect 38344 11092 38350 11104
rect 38473 11101 38485 11104
rect 38519 11101 38531 11135
rect 38473 11095 38531 11101
rect 38562 11092 38568 11144
rect 38620 11132 38626 11144
rect 39666 11132 39672 11144
rect 38620 11104 39672 11132
rect 38620 11092 38626 11104
rect 39666 11092 39672 11104
rect 39724 11092 39730 11144
rect 40037 11135 40095 11141
rect 40037 11101 40049 11135
rect 40083 11101 40095 11135
rect 40037 11095 40095 11101
rect 38838 11064 38844 11076
rect 38120 11036 38844 11064
rect 38013 11027 38071 11033
rect 32640 10968 32812 10996
rect 32640 10956 32646 10968
rect 36170 10956 36176 11008
rect 36228 10996 36234 11008
rect 36538 10996 36544 11008
rect 36228 10968 36544 10996
rect 36228 10956 36234 10968
rect 36538 10956 36544 10968
rect 36596 10956 36602 11008
rect 38028 10996 38056 11027
rect 38838 11024 38844 11036
rect 38896 11024 38902 11076
rect 40052 11064 40080 11095
rect 40126 11092 40132 11144
rect 40184 11132 40190 11144
rect 40681 11135 40739 11141
rect 40681 11132 40693 11135
rect 40184 11104 40693 11132
rect 40184 11092 40190 11104
rect 40681 11101 40693 11104
rect 40727 11101 40739 11135
rect 40681 11095 40739 11101
rect 41138 11092 41144 11144
rect 41196 11092 41202 11144
rect 42058 11092 42064 11144
rect 42116 11132 42122 11144
rect 42337 11135 42395 11141
rect 42337 11132 42349 11135
rect 42116 11104 42349 11132
rect 42116 11092 42122 11104
rect 42337 11101 42349 11104
rect 42383 11101 42395 11135
rect 42337 11095 42395 11101
rect 43165 11135 43223 11141
rect 43165 11101 43177 11135
rect 43211 11132 43223 11135
rect 43346 11132 43352 11144
rect 43211 11104 43352 11132
rect 43211 11101 43223 11104
rect 43165 11095 43223 11101
rect 43346 11092 43352 11104
rect 43404 11092 43410 11144
rect 43438 11092 43444 11144
rect 43496 11132 43502 11144
rect 43625 11135 43683 11141
rect 43625 11132 43637 11135
rect 43496 11104 43637 11132
rect 43496 11092 43502 11104
rect 43625 11101 43637 11104
rect 43671 11101 43683 11135
rect 43625 11095 43683 11101
rect 44542 11092 44548 11144
rect 44600 11132 44606 11144
rect 45462 11132 45468 11144
rect 44600 11104 45468 11132
rect 44600 11092 44606 11104
rect 45462 11092 45468 11104
rect 45520 11092 45526 11144
rect 45557 11135 45615 11141
rect 45557 11101 45569 11135
rect 45603 11132 45615 11135
rect 45649 11135 45707 11141
rect 45649 11132 45661 11135
rect 45603 11104 45661 11132
rect 45603 11101 45615 11104
rect 45557 11095 45615 11101
rect 45649 11101 45661 11104
rect 45695 11132 45707 11135
rect 46106 11132 46112 11144
rect 45695 11104 46112 11132
rect 45695 11101 45707 11104
rect 45649 11095 45707 11101
rect 46106 11092 46112 11104
rect 46164 11092 46170 11144
rect 47213 11135 47271 11141
rect 47213 11101 47225 11135
rect 47259 11132 47271 11135
rect 47394 11132 47400 11144
rect 47259 11104 47400 11132
rect 47259 11101 47271 11104
rect 47213 11095 47271 11101
rect 47394 11092 47400 11104
rect 47452 11092 47458 11144
rect 47964 11141 47992 11172
rect 49142 11160 49148 11212
rect 49200 11160 49206 11212
rect 47949 11135 48007 11141
rect 47949 11101 47961 11135
rect 47995 11101 48007 11135
rect 47949 11095 48007 11101
rect 41598 11064 41604 11076
rect 38948 11036 41604 11064
rect 38948 10996 38976 11036
rect 41598 11024 41604 11036
rect 41656 11024 41662 11076
rect 42521 11067 42579 11073
rect 42521 11033 42533 11067
rect 42567 11064 42579 11067
rect 42702 11064 42708 11076
rect 42567 11036 42708 11064
rect 42567 11033 42579 11036
rect 42521 11027 42579 11033
rect 42702 11024 42708 11036
rect 42760 11024 42766 11076
rect 43254 11024 43260 11076
rect 43312 11064 43318 11076
rect 45189 11067 45247 11073
rect 45189 11064 45201 11067
rect 43312 11036 45201 11064
rect 43312 11024 43318 11036
rect 45189 11033 45201 11036
rect 45235 11064 45247 11067
rect 45278 11064 45284 11076
rect 45235 11036 45284 11064
rect 45235 11033 45247 11036
rect 45189 11027 45247 11033
rect 45278 11024 45284 11036
rect 45336 11024 45342 11076
rect 47412 11064 47440 11092
rect 49418 11064 49424 11076
rect 47412 11036 49424 11064
rect 49418 11024 49424 11036
rect 49476 11024 49482 11076
rect 38028 10968 38976 10996
rect 39022 10956 39028 11008
rect 39080 10996 39086 11008
rect 44542 10996 44548 11008
rect 39080 10968 44548 10996
rect 39080 10956 39086 10968
rect 44542 10956 44548 10968
rect 44600 10956 44606 11008
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 2866 10752 2872 10804
rect 2924 10752 2930 10804
rect 3145 10795 3203 10801
rect 3145 10761 3157 10795
rect 3191 10792 3203 10795
rect 4062 10792 4068 10804
rect 3191 10764 4068 10792
rect 3191 10761 3203 10764
rect 3145 10755 3203 10761
rect 4062 10752 4068 10764
rect 4120 10752 4126 10804
rect 4522 10752 4528 10804
rect 4580 10792 4586 10804
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 4580 10764 5641 10792
rect 4580 10752 4586 10764
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 7745 10795 7803 10801
rect 7745 10792 7757 10795
rect 5629 10755 5687 10761
rect 5736 10764 7757 10792
rect 3326 10724 3332 10736
rect 1596 10696 3332 10724
rect 1210 10616 1216 10668
rect 1268 10656 1274 10668
rect 1596 10665 1624 10696
rect 3326 10684 3332 10696
rect 3384 10684 3390 10736
rect 5258 10684 5264 10736
rect 5316 10724 5322 10736
rect 5736 10724 5764 10764
rect 7745 10761 7757 10764
rect 7791 10761 7803 10795
rect 7745 10755 7803 10761
rect 8846 10752 8852 10804
rect 8904 10792 8910 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8904 10764 8953 10792
rect 8904 10752 8910 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 8941 10755 8999 10761
rect 9306 10752 9312 10804
rect 9364 10792 9370 10804
rect 11606 10792 11612 10804
rect 9364 10764 11612 10792
rect 9364 10752 9370 10764
rect 11606 10752 11612 10764
rect 11664 10752 11670 10804
rect 11698 10752 11704 10804
rect 11756 10792 11762 10804
rect 12345 10795 12403 10801
rect 12345 10792 12357 10795
rect 11756 10764 12357 10792
rect 11756 10752 11762 10764
rect 12345 10761 12357 10764
rect 12391 10761 12403 10795
rect 12345 10755 12403 10761
rect 12710 10752 12716 10804
rect 12768 10792 12774 10804
rect 15562 10792 15568 10804
rect 12768 10764 15568 10792
rect 12768 10752 12774 10764
rect 15562 10752 15568 10764
rect 15620 10752 15626 10804
rect 17310 10792 17316 10804
rect 15660 10764 17316 10792
rect 5316 10696 5764 10724
rect 6089 10727 6147 10733
rect 5316 10684 5322 10696
rect 6089 10693 6101 10727
rect 6135 10724 6147 10727
rect 6135 10696 6960 10724
rect 6135 10693 6147 10696
rect 6089 10687 6147 10693
rect 6932 10668 6960 10696
rect 7098 10684 7104 10736
rect 7156 10684 7162 10736
rect 10778 10684 10784 10736
rect 10836 10724 10842 10736
rect 13354 10724 13360 10736
rect 10836 10696 13360 10724
rect 10836 10684 10842 10696
rect 1581 10659 1639 10665
rect 1581 10656 1593 10659
rect 1268 10628 1593 10656
rect 1268 10616 1274 10628
rect 1581 10625 1593 10628
rect 1627 10625 1639 10659
rect 1581 10619 1639 10625
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10625 2375 10659
rect 2317 10619 2375 10625
rect 1302 10548 1308 10600
rect 1360 10588 1366 10600
rect 2332 10588 2360 10619
rect 3694 10616 3700 10668
rect 3752 10616 3758 10668
rect 3786 10616 3792 10668
rect 3844 10656 3850 10668
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 3844 10628 4445 10656
rect 3844 10616 3850 10628
rect 4433 10625 4445 10628
rect 4479 10625 4491 10659
rect 4433 10619 4491 10625
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10656 5595 10659
rect 6178 10656 6184 10668
rect 5583 10628 6184 10656
rect 5583 10625 5595 10628
rect 5537 10619 5595 10625
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 6914 10616 6920 10668
rect 6972 10616 6978 10668
rect 7653 10659 7711 10665
rect 7653 10625 7665 10659
rect 7699 10625 7711 10659
rect 7653 10619 7711 10625
rect 2406 10588 2412 10600
rect 1360 10560 2412 10588
rect 1360 10548 1366 10560
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 4157 10591 4215 10597
rect 4157 10557 4169 10591
rect 4203 10588 4215 10591
rect 4338 10588 4344 10600
rect 4203 10560 4344 10588
rect 4203 10557 4215 10560
rect 4157 10551 4215 10557
rect 4338 10548 4344 10560
rect 4396 10588 4402 10600
rect 5994 10588 6000 10600
rect 4396 10560 6000 10588
rect 4396 10548 4402 10560
rect 5994 10548 6000 10560
rect 6052 10548 6058 10600
rect 6549 10591 6607 10597
rect 6549 10557 6561 10591
rect 6595 10588 6607 10591
rect 7668 10588 7696 10619
rect 8294 10616 8300 10668
rect 8352 10656 8358 10668
rect 9030 10656 9036 10668
rect 8352 10628 9036 10656
rect 8352 10616 8358 10628
rect 9030 10616 9036 10628
rect 9088 10616 9094 10668
rect 9398 10616 9404 10668
rect 9456 10616 9462 10668
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 10505 10659 10563 10665
rect 10505 10656 10517 10659
rect 10008 10628 10517 10656
rect 10008 10616 10014 10628
rect 10505 10625 10517 10628
rect 10551 10625 10563 10659
rect 10505 10619 10563 10625
rect 11422 10616 11428 10668
rect 11480 10656 11486 10668
rect 12158 10656 12164 10668
rect 11480 10628 12164 10656
rect 11480 10616 11486 10628
rect 12158 10616 12164 10628
rect 12216 10616 12222 10668
rect 12250 10616 12256 10668
rect 12308 10656 12314 10668
rect 13188 10665 13216 10696
rect 13354 10684 13360 10696
rect 13412 10684 13418 10736
rect 15286 10724 15292 10736
rect 14674 10696 15292 10724
rect 15286 10684 15292 10696
rect 15344 10684 15350 10736
rect 15660 10724 15688 10764
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 17770 10752 17776 10804
rect 17828 10792 17834 10804
rect 18141 10795 18199 10801
rect 18141 10792 18153 10795
rect 17828 10764 18153 10792
rect 17828 10752 17834 10764
rect 18141 10761 18153 10764
rect 18187 10761 18199 10795
rect 18141 10755 18199 10761
rect 18506 10752 18512 10804
rect 18564 10792 18570 10804
rect 19334 10792 19340 10804
rect 18564 10764 19340 10792
rect 18564 10752 18570 10764
rect 19334 10752 19340 10764
rect 19392 10752 19398 10804
rect 19426 10752 19432 10804
rect 19484 10752 19490 10804
rect 21634 10792 21640 10804
rect 19720 10764 21640 10792
rect 15396 10696 15688 10724
rect 16301 10727 16359 10733
rect 12437 10659 12495 10665
rect 12437 10656 12449 10659
rect 12308 10628 12449 10656
rect 12308 10616 12314 10628
rect 12437 10625 12449 10628
rect 12483 10625 12495 10659
rect 12437 10619 12495 10625
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10625 13231 10659
rect 13173 10619 13231 10625
rect 15102 10616 15108 10668
rect 15160 10656 15166 10668
rect 15396 10656 15424 10696
rect 16301 10693 16313 10727
rect 16347 10724 16359 10727
rect 19610 10724 19616 10736
rect 16347 10696 18276 10724
rect 16347 10693 16359 10696
rect 16301 10687 16359 10693
rect 15160 10628 15424 10656
rect 15657 10659 15715 10665
rect 15160 10616 15166 10628
rect 15657 10625 15669 10659
rect 15703 10625 15715 10659
rect 15657 10619 15715 10625
rect 10962 10588 10968 10600
rect 6595 10560 10968 10588
rect 6595 10557 6607 10560
rect 6549 10551 6607 10557
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 12526 10548 12532 10600
rect 12584 10548 12590 10600
rect 12802 10548 12808 10600
rect 12860 10588 12866 10600
rect 13449 10591 13507 10597
rect 13449 10588 13461 10591
rect 12860 10560 13461 10588
rect 12860 10548 12866 10560
rect 13449 10557 13461 10560
rect 13495 10557 13507 10591
rect 13449 10551 13507 10557
rect 14458 10548 14464 10600
rect 14516 10588 14522 10600
rect 15194 10588 15200 10600
rect 14516 10560 15200 10588
rect 14516 10548 14522 10560
rect 15194 10548 15200 10560
rect 15252 10548 15258 10600
rect 1762 10480 1768 10532
rect 1820 10480 1826 10532
rect 2501 10523 2559 10529
rect 2501 10489 2513 10523
rect 2547 10520 2559 10523
rect 8018 10520 8024 10532
rect 2547 10492 8024 10520
rect 2547 10489 2559 10492
rect 2501 10483 2559 10489
rect 8018 10480 8024 10492
rect 8076 10480 8082 10532
rect 10686 10520 10692 10532
rect 9646 10492 10692 10520
rect 3513 10455 3571 10461
rect 3513 10421 3525 10455
rect 3559 10452 3571 10455
rect 5718 10452 5724 10464
rect 3559 10424 5724 10452
rect 3559 10421 3571 10424
rect 3513 10415 3571 10421
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 9646 10452 9674 10492
rect 10686 10480 10692 10492
rect 10744 10480 10750 10532
rect 11149 10523 11207 10529
rect 11149 10489 11161 10523
rect 11195 10520 11207 10523
rect 15672 10520 15700 10619
rect 17310 10616 17316 10668
rect 17368 10616 17374 10668
rect 17405 10659 17463 10665
rect 17405 10625 17417 10659
rect 17451 10656 17463 10659
rect 17770 10656 17776 10668
rect 17451 10628 17776 10656
rect 17451 10625 17463 10628
rect 17405 10619 17463 10625
rect 16574 10548 16580 10600
rect 16632 10588 16638 10600
rect 17420 10588 17448 10619
rect 17770 10616 17776 10628
rect 17828 10616 17834 10668
rect 18248 10656 18276 10696
rect 18432 10696 19616 10724
rect 18432 10656 18460 10696
rect 19610 10684 19616 10696
rect 19668 10684 19674 10736
rect 18248 10628 18460 10656
rect 18509 10659 18567 10665
rect 18509 10625 18521 10659
rect 18555 10656 18567 10659
rect 18966 10656 18972 10668
rect 18555 10628 18972 10656
rect 18555 10625 18567 10628
rect 18509 10619 18567 10625
rect 18966 10616 18972 10628
rect 19024 10616 19030 10668
rect 19720 10600 19748 10764
rect 21634 10752 21640 10764
rect 21692 10752 21698 10804
rect 22097 10795 22155 10801
rect 22097 10761 22109 10795
rect 22143 10792 22155 10795
rect 24026 10792 24032 10804
rect 22143 10764 24032 10792
rect 22143 10761 22155 10764
rect 22097 10755 22155 10761
rect 24026 10752 24032 10764
rect 24084 10752 24090 10804
rect 26234 10792 26240 10804
rect 24320 10764 26240 10792
rect 20714 10684 20720 10736
rect 20772 10684 20778 10736
rect 21818 10684 21824 10736
rect 21876 10724 21882 10736
rect 22465 10727 22523 10733
rect 21876 10696 22094 10724
rect 21876 10684 21882 10696
rect 16632 10560 17448 10588
rect 17589 10591 17647 10597
rect 16632 10548 16638 10560
rect 17589 10557 17601 10591
rect 17635 10588 17647 10591
rect 17862 10588 17868 10600
rect 17635 10560 17868 10588
rect 17635 10557 17647 10560
rect 17589 10551 17647 10557
rect 17862 10548 17868 10560
rect 17920 10548 17926 10600
rect 18601 10591 18659 10597
rect 18601 10557 18613 10591
rect 18647 10557 18659 10591
rect 18601 10551 18659 10557
rect 18506 10520 18512 10532
rect 11195 10492 13308 10520
rect 15672 10492 18512 10520
rect 11195 10489 11207 10492
rect 11149 10483 11207 10489
rect 6052 10424 9674 10452
rect 10045 10455 10103 10461
rect 6052 10412 6058 10424
rect 10045 10421 10057 10455
rect 10091 10452 10103 10455
rect 11238 10452 11244 10464
rect 10091 10424 11244 10452
rect 10091 10421 10103 10424
rect 10045 10415 10103 10421
rect 11238 10412 11244 10424
rect 11296 10412 11302 10464
rect 11977 10455 12035 10461
rect 11977 10421 11989 10455
rect 12023 10452 12035 10455
rect 12158 10452 12164 10464
rect 12023 10424 12164 10452
rect 12023 10421 12035 10424
rect 11977 10415 12035 10421
rect 12158 10412 12164 10424
rect 12216 10412 12222 10464
rect 13280 10452 13308 10492
rect 18506 10480 18512 10492
rect 18564 10480 18570 10532
rect 18616 10520 18644 10551
rect 18690 10548 18696 10600
rect 18748 10548 18754 10600
rect 19702 10548 19708 10600
rect 19760 10548 19766 10600
rect 19978 10548 19984 10600
rect 20036 10548 20042 10600
rect 20622 10548 20628 10600
rect 20680 10588 20686 10600
rect 21453 10591 21511 10597
rect 21453 10588 21465 10591
rect 20680 10560 21465 10588
rect 20680 10548 20686 10560
rect 21453 10557 21465 10560
rect 21499 10557 21511 10591
rect 22066 10588 22094 10696
rect 22465 10693 22477 10727
rect 22511 10724 22523 10727
rect 24320 10724 24348 10764
rect 26234 10752 26240 10764
rect 26292 10752 26298 10804
rect 26510 10752 26516 10804
rect 26568 10752 26574 10804
rect 27798 10752 27804 10804
rect 27856 10792 27862 10804
rect 28261 10795 28319 10801
rect 28261 10792 28273 10795
rect 27856 10764 28273 10792
rect 27856 10752 27862 10764
rect 28261 10761 28273 10764
rect 28307 10761 28319 10795
rect 28261 10755 28319 10761
rect 28718 10752 28724 10804
rect 28776 10792 28782 10804
rect 29273 10795 29331 10801
rect 29273 10792 29285 10795
rect 28776 10764 29285 10792
rect 28776 10752 28782 10764
rect 29273 10761 29285 10764
rect 29319 10761 29331 10795
rect 29273 10755 29331 10761
rect 30392 10764 31524 10792
rect 22511 10696 24348 10724
rect 22511 10693 22523 10696
rect 22465 10687 22523 10693
rect 24394 10684 24400 10736
rect 24452 10724 24458 10736
rect 24452 10696 24978 10724
rect 24452 10684 24458 10696
rect 27154 10684 27160 10736
rect 27212 10724 27218 10736
rect 30392 10724 30420 10764
rect 27212 10696 30420 10724
rect 31496 10724 31524 10764
rect 31662 10752 31668 10804
rect 31720 10792 31726 10804
rect 32953 10795 33011 10801
rect 32953 10792 32965 10795
rect 31720 10764 32965 10792
rect 31720 10752 31726 10764
rect 32953 10761 32965 10764
rect 32999 10761 33011 10795
rect 35066 10792 35072 10804
rect 32953 10755 33011 10761
rect 33796 10764 35072 10792
rect 33045 10727 33103 10733
rect 33045 10724 33057 10727
rect 31496 10696 33057 10724
rect 27212 10684 27218 10696
rect 33045 10693 33057 10696
rect 33091 10693 33103 10727
rect 33045 10687 33103 10693
rect 23474 10616 23480 10668
rect 23532 10656 23538 10668
rect 24210 10656 24216 10668
rect 23532 10628 24216 10656
rect 23532 10616 23538 10628
rect 24210 10616 24216 10628
rect 24268 10616 24274 10668
rect 27617 10659 27675 10665
rect 27617 10625 27629 10659
rect 27663 10656 27675 10659
rect 28074 10656 28080 10668
rect 27663 10628 28080 10656
rect 27663 10625 27675 10628
rect 27617 10619 27675 10625
rect 28074 10616 28080 10628
rect 28132 10616 28138 10668
rect 28629 10659 28687 10665
rect 28629 10625 28641 10659
rect 28675 10656 28687 10659
rect 29178 10656 29184 10668
rect 28675 10628 29184 10656
rect 28675 10625 28687 10628
rect 28629 10619 28687 10625
rect 29178 10616 29184 10628
rect 29236 10616 29242 10668
rect 31478 10656 31484 10668
rect 31326 10628 31484 10656
rect 31478 10616 31484 10628
rect 31536 10616 31542 10668
rect 32398 10616 32404 10668
rect 32456 10656 32462 10668
rect 32456 10628 32812 10656
rect 32456 10616 32462 10628
rect 32784 10600 32812 10628
rect 32858 10616 32864 10668
rect 32916 10656 32922 10668
rect 33796 10656 33824 10764
rect 35066 10752 35072 10764
rect 35124 10752 35130 10804
rect 35526 10752 35532 10804
rect 35584 10752 35590 10804
rect 36449 10795 36507 10801
rect 36449 10761 36461 10795
rect 36495 10792 36507 10795
rect 36630 10792 36636 10804
rect 36495 10764 36636 10792
rect 36495 10761 36507 10764
rect 36449 10755 36507 10761
rect 36630 10752 36636 10764
rect 36688 10792 36694 10804
rect 36998 10792 37004 10804
rect 36688 10764 37004 10792
rect 36688 10752 36694 10764
rect 36998 10752 37004 10764
rect 37056 10752 37062 10804
rect 37090 10752 37096 10804
rect 37148 10752 37154 10804
rect 37550 10752 37556 10804
rect 37608 10792 37614 10804
rect 38010 10792 38016 10804
rect 37608 10764 38016 10792
rect 37608 10752 37614 10764
rect 38010 10752 38016 10764
rect 38068 10752 38074 10804
rect 42058 10752 42064 10804
rect 42116 10752 42122 10804
rect 43438 10752 43444 10804
rect 43496 10792 43502 10804
rect 46937 10795 46995 10801
rect 46937 10792 46949 10795
rect 43496 10764 46949 10792
rect 43496 10752 43502 10764
rect 46937 10761 46949 10764
rect 46983 10761 46995 10795
rect 46937 10755 46995 10761
rect 47670 10752 47676 10804
rect 47728 10752 47734 10804
rect 35434 10684 35440 10736
rect 35492 10724 35498 10736
rect 35492 10696 36860 10724
rect 35492 10684 35498 10696
rect 36170 10656 36176 10668
rect 32916 10628 33824 10656
rect 35190 10628 36176 10656
rect 32916 10616 32922 10628
rect 36170 10616 36176 10628
rect 36228 10616 36234 10668
rect 36357 10659 36415 10665
rect 36357 10625 36369 10659
rect 36403 10625 36415 10659
rect 36357 10619 36415 10625
rect 22557 10591 22615 10597
rect 22557 10588 22569 10591
rect 22066 10560 22569 10588
rect 21453 10551 21511 10557
rect 22557 10557 22569 10560
rect 22603 10557 22615 10591
rect 22557 10551 22615 10557
rect 22572 10520 22600 10551
rect 22738 10548 22744 10600
rect 22796 10548 22802 10600
rect 23290 10548 23296 10600
rect 23348 10548 23354 10600
rect 24489 10591 24547 10597
rect 24489 10557 24501 10591
rect 24535 10588 24547 10591
rect 25866 10588 25872 10600
rect 24535 10560 25872 10588
rect 24535 10557 24547 10560
rect 24489 10551 24547 10557
rect 25866 10548 25872 10560
rect 25924 10548 25930 10600
rect 26050 10548 26056 10600
rect 26108 10588 26114 10600
rect 26237 10591 26295 10597
rect 26237 10588 26249 10591
rect 26108 10560 26249 10588
rect 26108 10548 26114 10560
rect 26237 10557 26249 10560
rect 26283 10557 26295 10591
rect 26237 10551 26295 10557
rect 26789 10591 26847 10597
rect 26789 10557 26801 10591
rect 26835 10588 26847 10591
rect 26970 10588 26976 10600
rect 26835 10560 26976 10588
rect 26835 10557 26847 10560
rect 26789 10551 26847 10557
rect 26970 10548 26976 10560
rect 27028 10588 27034 10600
rect 27709 10591 27767 10597
rect 27709 10588 27721 10591
rect 27028 10560 27721 10588
rect 27028 10548 27034 10560
rect 27709 10557 27721 10560
rect 27755 10588 27767 10591
rect 27798 10588 27804 10600
rect 27755 10560 27804 10588
rect 27755 10557 27767 10560
rect 27709 10551 27767 10557
rect 27798 10548 27804 10560
rect 27856 10548 27862 10600
rect 27893 10591 27951 10597
rect 27893 10557 27905 10591
rect 27939 10588 27951 10591
rect 28534 10588 28540 10600
rect 27939 10560 28540 10588
rect 27939 10557 27951 10560
rect 27893 10551 27951 10557
rect 28534 10548 28540 10560
rect 28592 10548 28598 10600
rect 29730 10548 29736 10600
rect 29788 10588 29794 10600
rect 29917 10591 29975 10597
rect 29917 10588 29929 10591
rect 29788 10560 29929 10588
rect 29788 10548 29794 10560
rect 29917 10557 29929 10560
rect 29963 10557 29975 10591
rect 29917 10551 29975 10557
rect 30193 10591 30251 10597
rect 30193 10557 30205 10591
rect 30239 10588 30251 10591
rect 30650 10588 30656 10600
rect 30239 10560 30656 10588
rect 30239 10557 30251 10560
rect 30193 10551 30251 10557
rect 30650 10548 30656 10560
rect 30708 10548 30714 10600
rect 32674 10588 32680 10600
rect 31220 10560 32680 10588
rect 23566 10520 23572 10532
rect 18616 10492 19840 10520
rect 22572 10492 23572 10520
rect 15194 10452 15200 10464
rect 13280 10424 15200 10452
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 16945 10455 17003 10461
rect 16945 10421 16957 10455
rect 16991 10452 17003 10455
rect 17126 10452 17132 10464
rect 16991 10424 17132 10452
rect 16991 10421 17003 10424
rect 16945 10415 17003 10421
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 17954 10412 17960 10464
rect 18012 10452 18018 10464
rect 19150 10452 19156 10464
rect 18012 10424 19156 10452
rect 18012 10412 18018 10424
rect 19150 10412 19156 10424
rect 19208 10412 19214 10464
rect 19812 10452 19840 10492
rect 23566 10480 23572 10492
rect 23624 10480 23630 10532
rect 27249 10523 27307 10529
rect 27249 10489 27261 10523
rect 27295 10520 27307 10523
rect 27295 10492 29868 10520
rect 27295 10489 27307 10492
rect 27249 10483 27307 10489
rect 21358 10452 21364 10464
rect 19812 10424 21364 10452
rect 21358 10412 21364 10424
rect 21416 10412 21422 10464
rect 23658 10412 23664 10464
rect 23716 10452 23722 10464
rect 23937 10455 23995 10461
rect 23937 10452 23949 10455
rect 23716 10424 23949 10452
rect 23716 10412 23722 10424
rect 23937 10421 23949 10424
rect 23983 10452 23995 10455
rect 24026 10452 24032 10464
rect 23983 10424 24032 10452
rect 23983 10421 23995 10424
rect 23937 10415 23995 10421
rect 24026 10412 24032 10424
rect 24084 10412 24090 10464
rect 24302 10412 24308 10464
rect 24360 10452 24366 10464
rect 24670 10452 24676 10464
rect 24360 10424 24676 10452
rect 24360 10412 24366 10424
rect 24670 10412 24676 10424
rect 24728 10452 24734 10464
rect 25961 10455 26019 10461
rect 25961 10452 25973 10455
rect 24728 10424 25973 10452
rect 24728 10412 24734 10424
rect 25961 10421 25973 10424
rect 26007 10421 26019 10455
rect 25961 10415 26019 10421
rect 29546 10412 29552 10464
rect 29604 10412 29610 10464
rect 29840 10452 29868 10492
rect 31220 10452 31248 10560
rect 32674 10548 32680 10560
rect 32732 10548 32738 10600
rect 32766 10548 32772 10600
rect 32824 10588 32830 10600
rect 33137 10591 33195 10597
rect 33137 10588 33149 10591
rect 32824 10560 33149 10588
rect 32824 10548 32830 10560
rect 33137 10557 33149 10560
rect 33183 10557 33195 10591
rect 33137 10551 33195 10557
rect 33781 10591 33839 10597
rect 33781 10557 33793 10591
rect 33827 10557 33839 10591
rect 33781 10551 33839 10557
rect 34057 10591 34115 10597
rect 34057 10557 34069 10591
rect 34103 10588 34115 10591
rect 36262 10588 36268 10600
rect 34103 10560 36268 10588
rect 34103 10557 34115 10560
rect 34057 10551 34115 10557
rect 31386 10480 31392 10532
rect 31444 10520 31450 10532
rect 31665 10523 31723 10529
rect 31665 10520 31677 10523
rect 31444 10492 31677 10520
rect 31444 10480 31450 10492
rect 31665 10489 31677 10492
rect 31711 10489 31723 10523
rect 31665 10483 31723 10489
rect 29840 10424 31248 10452
rect 31680 10452 31708 10483
rect 31938 10480 31944 10532
rect 31996 10520 32002 10532
rect 33502 10520 33508 10532
rect 31996 10492 33508 10520
rect 31996 10480 32002 10492
rect 33502 10480 33508 10492
rect 33560 10520 33566 10532
rect 33796 10520 33824 10551
rect 36262 10548 36268 10560
rect 36320 10548 36326 10600
rect 36372 10588 36400 10619
rect 36538 10588 36544 10600
rect 36372 10560 36544 10588
rect 36538 10548 36544 10560
rect 36596 10548 36602 10600
rect 36630 10548 36636 10600
rect 36688 10548 36694 10600
rect 36832 10588 36860 10696
rect 37458 10684 37464 10736
rect 37516 10724 37522 10736
rect 37516 10696 40908 10724
rect 37516 10684 37522 10696
rect 36906 10616 36912 10668
rect 36964 10656 36970 10668
rect 37642 10656 37648 10668
rect 36964 10628 37648 10656
rect 36964 10616 36970 10628
rect 37642 10616 37648 10628
rect 37700 10616 37706 10668
rect 37826 10616 37832 10668
rect 37884 10616 37890 10668
rect 37921 10659 37979 10665
rect 37921 10625 37933 10659
rect 37967 10656 37979 10659
rect 38562 10656 38568 10668
rect 37967 10628 38568 10656
rect 37967 10625 37979 10628
rect 37921 10619 37979 10625
rect 38562 10616 38568 10628
rect 38620 10616 38626 10668
rect 38657 10660 38715 10665
rect 38657 10659 38884 10660
rect 38657 10625 38669 10659
rect 38703 10656 38884 10659
rect 39574 10656 39580 10668
rect 38703 10632 39580 10656
rect 38703 10625 38715 10632
rect 38856 10628 39580 10632
rect 38657 10619 38715 10625
rect 39574 10616 39580 10628
rect 39632 10616 39638 10668
rect 40880 10665 40908 10696
rect 43622 10684 43628 10736
rect 43680 10724 43686 10736
rect 45554 10724 45560 10736
rect 43680 10696 45560 10724
rect 43680 10684 43686 10696
rect 45554 10684 45560 10696
rect 45612 10684 45618 10736
rect 46198 10724 46204 10736
rect 45848 10696 46204 10724
rect 39761 10659 39819 10665
rect 39761 10625 39773 10659
rect 39807 10625 39819 10659
rect 39761 10619 39819 10625
rect 40865 10659 40923 10665
rect 40865 10625 40877 10659
rect 40911 10625 40923 10659
rect 40865 10619 40923 10625
rect 37660 10588 37688 10616
rect 38013 10591 38071 10597
rect 38013 10588 38025 10591
rect 36832 10560 37596 10588
rect 37660 10560 38025 10588
rect 33560 10492 33824 10520
rect 33560 10480 33566 10492
rect 35342 10480 35348 10532
rect 35400 10520 35406 10532
rect 37461 10523 37519 10529
rect 37461 10520 37473 10523
rect 35400 10492 37473 10520
rect 35400 10480 35406 10492
rect 37461 10489 37473 10492
rect 37507 10489 37519 10523
rect 37461 10483 37519 10489
rect 32030 10452 32036 10464
rect 31680 10424 32036 10452
rect 32030 10412 32036 10424
rect 32088 10412 32094 10464
rect 32585 10455 32643 10461
rect 32585 10421 32597 10455
rect 32631 10452 32643 10455
rect 33318 10452 33324 10464
rect 32631 10424 33324 10452
rect 32631 10421 32643 10424
rect 32585 10415 32643 10421
rect 33318 10412 33324 10424
rect 33376 10412 33382 10464
rect 35989 10455 36047 10461
rect 35989 10421 36001 10455
rect 36035 10452 36047 10455
rect 36906 10452 36912 10464
rect 36035 10424 36912 10452
rect 36035 10421 36047 10424
rect 35989 10415 36047 10421
rect 36906 10412 36912 10424
rect 36964 10412 36970 10464
rect 37568 10452 37596 10560
rect 38013 10557 38025 10560
rect 38059 10588 38071 10591
rect 38102 10588 38108 10600
rect 38059 10560 38108 10588
rect 38059 10557 38071 10560
rect 38013 10551 38071 10557
rect 38102 10548 38108 10560
rect 38160 10548 38166 10600
rect 38286 10548 38292 10600
rect 38344 10588 38350 10600
rect 39776 10588 39804 10619
rect 40954 10616 40960 10668
rect 41012 10656 41018 10668
rect 42797 10659 42855 10665
rect 42797 10656 42809 10659
rect 41012 10628 42809 10656
rect 41012 10616 41018 10628
rect 42797 10625 42809 10628
rect 42843 10625 42855 10659
rect 42797 10619 42855 10625
rect 43533 10659 43591 10665
rect 43533 10625 43545 10659
rect 43579 10656 43591 10659
rect 44082 10656 44088 10668
rect 43579 10628 44088 10656
rect 43579 10625 43591 10628
rect 43533 10619 43591 10625
rect 44082 10616 44088 10628
rect 44140 10616 44146 10668
rect 44542 10616 44548 10668
rect 44600 10616 44606 10668
rect 45848 10665 45876 10696
rect 46198 10684 46204 10696
rect 46256 10684 46262 10736
rect 47397 10727 47455 10733
rect 47397 10693 47409 10727
rect 47443 10724 47455 10727
rect 48590 10724 48596 10736
rect 47443 10696 48596 10724
rect 47443 10693 47455 10696
rect 47397 10687 47455 10693
rect 48590 10684 48596 10696
rect 48648 10684 48654 10736
rect 49145 10727 49203 10733
rect 49145 10693 49157 10727
rect 49191 10724 49203 10727
rect 49326 10724 49332 10736
rect 49191 10696 49332 10724
rect 49191 10693 49203 10696
rect 49145 10687 49203 10693
rect 49326 10684 49332 10696
rect 49384 10684 49390 10736
rect 45833 10659 45891 10665
rect 45833 10625 45845 10659
rect 45879 10625 45891 10659
rect 45833 10619 45891 10625
rect 46106 10616 46112 10668
rect 46164 10616 46170 10668
rect 47949 10659 48007 10665
rect 47949 10656 47961 10659
rect 46216 10628 47961 10656
rect 38344 10560 39804 10588
rect 38344 10548 38350 10560
rect 39850 10548 39856 10600
rect 39908 10588 39914 10600
rect 41785 10591 41843 10597
rect 41785 10588 41797 10591
rect 39908 10560 41797 10588
rect 39908 10548 39914 10560
rect 41785 10557 41797 10560
rect 41831 10557 41843 10591
rect 41785 10551 41843 10557
rect 41874 10548 41880 10600
rect 41932 10588 41938 10600
rect 42150 10588 42156 10600
rect 41932 10560 42156 10588
rect 41932 10548 41938 10560
rect 42150 10548 42156 10560
rect 42208 10548 42214 10600
rect 42610 10548 42616 10600
rect 42668 10588 42674 10600
rect 43257 10591 43315 10597
rect 43257 10588 43269 10591
rect 42668 10560 43269 10588
rect 42668 10548 42674 10560
rect 43257 10557 43269 10560
rect 43303 10588 43315 10591
rect 43714 10588 43720 10600
rect 43303 10560 43720 10588
rect 43303 10557 43315 10560
rect 43257 10551 43315 10557
rect 43714 10548 43720 10560
rect 43772 10548 43778 10600
rect 44726 10548 44732 10600
rect 44784 10588 44790 10600
rect 44821 10591 44879 10597
rect 44821 10588 44833 10591
rect 44784 10560 44833 10588
rect 44784 10548 44790 10560
rect 44821 10557 44833 10560
rect 44867 10557 44879 10591
rect 44821 10551 44879 10557
rect 38562 10480 38568 10532
rect 38620 10520 38626 10532
rect 41509 10523 41567 10529
rect 41509 10520 41521 10523
rect 38620 10492 41521 10520
rect 38620 10480 38626 10492
rect 41509 10489 41521 10492
rect 41555 10489 41567 10523
rect 43990 10520 43996 10532
rect 41509 10483 41567 10489
rect 42076 10492 43996 10520
rect 39301 10455 39359 10461
rect 39301 10452 39313 10455
rect 37568 10424 39313 10452
rect 39301 10421 39313 10424
rect 39347 10421 39359 10455
rect 39301 10415 39359 10421
rect 40402 10412 40408 10464
rect 40460 10412 40466 10464
rect 40678 10412 40684 10464
rect 40736 10452 40742 10464
rect 42076 10452 42104 10492
rect 43990 10480 43996 10492
rect 44048 10480 44054 10532
rect 45370 10480 45376 10532
rect 45428 10520 45434 10532
rect 46216 10520 46244 10628
rect 47949 10625 47961 10628
rect 47995 10625 48007 10659
rect 47949 10619 48007 10625
rect 47213 10591 47271 10597
rect 47213 10557 47225 10591
rect 47259 10588 47271 10591
rect 48866 10588 48872 10600
rect 47259 10560 48872 10588
rect 47259 10557 47271 10560
rect 47213 10551 47271 10557
rect 48866 10548 48872 10560
rect 48924 10548 48930 10600
rect 45428 10492 46244 10520
rect 45428 10480 45434 10492
rect 40736 10424 42104 10452
rect 42613 10455 42671 10461
rect 40736 10412 40742 10424
rect 42613 10421 42625 10455
rect 42659 10452 42671 10455
rect 44082 10452 44088 10464
rect 42659 10424 44088 10452
rect 42659 10421 42671 10424
rect 42613 10415 42671 10421
rect 44082 10412 44088 10424
rect 44140 10412 44146 10464
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 1578 10208 1584 10260
rect 1636 10248 1642 10260
rect 3329 10251 3387 10257
rect 3329 10248 3341 10251
rect 1636 10220 3341 10248
rect 1636 10208 1642 10220
rect 3329 10217 3341 10220
rect 3375 10217 3387 10251
rect 3329 10211 3387 10217
rect 3605 10251 3663 10257
rect 3605 10217 3617 10251
rect 3651 10248 3663 10251
rect 3694 10248 3700 10260
rect 3651 10220 3700 10248
rect 3651 10217 3663 10220
rect 3605 10211 3663 10217
rect 3694 10208 3700 10220
rect 3752 10208 3758 10260
rect 5166 10208 5172 10260
rect 5224 10208 5230 10260
rect 5902 10208 5908 10260
rect 5960 10208 5966 10260
rect 7374 10208 7380 10260
rect 7432 10208 7438 10260
rect 8662 10248 8668 10260
rect 7760 10220 8668 10248
rect 1872 10152 5764 10180
rect 1872 10121 1900 10152
rect 1857 10115 1915 10121
rect 1857 10081 1869 10115
rect 1903 10081 1915 10115
rect 1857 10075 1915 10081
rect 4246 10072 4252 10124
rect 4304 10072 4310 10124
rect 5736 10112 5764 10152
rect 5810 10140 5816 10192
rect 5868 10180 5874 10192
rect 6733 10183 6791 10189
rect 6733 10180 6745 10183
rect 5868 10152 6745 10180
rect 5868 10140 5874 10152
rect 6733 10149 6745 10152
rect 6779 10149 6791 10183
rect 6733 10143 6791 10149
rect 7760 10112 7788 10220
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 9122 10208 9128 10260
rect 9180 10208 9186 10260
rect 9582 10208 9588 10260
rect 9640 10248 9646 10260
rect 10229 10251 10287 10257
rect 10229 10248 10241 10251
rect 9640 10220 10241 10248
rect 9640 10208 9646 10220
rect 10229 10217 10241 10220
rect 10275 10217 10287 10251
rect 10229 10211 10287 10217
rect 11333 10251 11391 10257
rect 11333 10217 11345 10251
rect 11379 10248 11391 10251
rect 12802 10248 12808 10260
rect 11379 10220 12808 10248
rect 11379 10217 11391 10220
rect 11333 10211 11391 10217
rect 12802 10208 12808 10220
rect 12860 10208 12866 10260
rect 13906 10208 13912 10260
rect 13964 10248 13970 10260
rect 15286 10248 15292 10260
rect 13964 10220 15292 10248
rect 13964 10208 13970 10220
rect 15286 10208 15292 10220
rect 15344 10248 15350 10260
rect 16206 10248 16212 10260
rect 15344 10220 16212 10248
rect 15344 10208 15350 10220
rect 16206 10208 16212 10220
rect 16264 10208 16270 10260
rect 16485 10251 16543 10257
rect 16485 10217 16497 10251
rect 16531 10248 16543 10251
rect 16574 10248 16580 10260
rect 16531 10220 16580 10248
rect 16531 10217 16543 10220
rect 16485 10211 16543 10217
rect 16574 10208 16580 10220
rect 16632 10208 16638 10260
rect 16942 10208 16948 10260
rect 17000 10208 17006 10260
rect 17402 10248 17408 10260
rect 17328 10220 17408 10248
rect 8386 10140 8392 10192
rect 8444 10180 8450 10192
rect 9217 10183 9275 10189
rect 9217 10180 9229 10183
rect 8444 10152 9229 10180
rect 8444 10140 8450 10152
rect 9217 10149 9229 10152
rect 9263 10149 9275 10183
rect 10870 10180 10876 10192
rect 9217 10143 9275 10149
rect 9646 10152 10876 10180
rect 9646 10112 9674 10152
rect 10870 10140 10876 10152
rect 10928 10140 10934 10192
rect 12066 10140 12072 10192
rect 12124 10180 12130 10192
rect 12989 10183 13047 10189
rect 12989 10180 13001 10183
rect 12124 10152 13001 10180
rect 12124 10140 12130 10152
rect 12989 10149 13001 10152
rect 13035 10149 13047 10183
rect 12989 10143 13047 10149
rect 15562 10140 15568 10192
rect 15620 10180 15626 10192
rect 16025 10183 16083 10189
rect 16025 10180 16037 10183
rect 15620 10152 16037 10180
rect 15620 10140 15626 10152
rect 16025 10149 16037 10152
rect 16071 10149 16083 10183
rect 16025 10143 16083 10149
rect 5736 10084 7788 10112
rect 7852 10084 9674 10112
rect 1578 10004 1584 10056
rect 1636 10004 1642 10056
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10013 4031 10047
rect 3973 10007 4031 10013
rect 2685 9979 2743 9985
rect 2685 9945 2697 9979
rect 2731 9976 2743 9979
rect 3988 9976 4016 10007
rect 5534 10004 5540 10056
rect 5592 10044 5598 10056
rect 7285 10047 7343 10053
rect 7285 10044 7297 10047
rect 5592 10016 7297 10044
rect 5592 10004 5598 10016
rect 7285 10013 7297 10016
rect 7331 10013 7343 10047
rect 7285 10007 7343 10013
rect 5626 9976 5632 9988
rect 2731 9948 2912 9976
rect 3988 9948 5632 9976
rect 2731 9945 2743 9948
rect 2685 9939 2743 9945
rect 2884 9917 2912 9948
rect 5626 9936 5632 9948
rect 5684 9936 5690 9988
rect 5813 9979 5871 9985
rect 5813 9945 5825 9979
rect 5859 9976 5871 9979
rect 6362 9976 6368 9988
rect 5859 9948 6368 9976
rect 5859 9945 5871 9948
rect 5813 9939 5871 9945
rect 6362 9936 6368 9948
rect 6420 9936 6426 9988
rect 6549 9979 6607 9985
rect 6549 9945 6561 9979
rect 6595 9976 6607 9979
rect 7852 9976 7880 10084
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 12253 10115 12311 10121
rect 12253 10112 12265 10115
rect 10468 10084 12265 10112
rect 10468 10072 10474 10084
rect 12253 10081 12265 10084
rect 12299 10081 12311 10115
rect 12253 10075 12311 10081
rect 12342 10072 12348 10124
rect 12400 10072 12406 10124
rect 13446 10072 13452 10124
rect 13504 10072 13510 10124
rect 13630 10072 13636 10124
rect 13688 10072 13694 10124
rect 14277 10115 14335 10121
rect 14277 10081 14289 10115
rect 14323 10112 14335 10115
rect 16298 10112 16304 10124
rect 14323 10084 16304 10112
rect 14323 10081 14335 10084
rect 14277 10075 14335 10081
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 6595 9948 7880 9976
rect 6595 9945 6607 9948
rect 6549 9939 6607 9945
rect 2869 9911 2927 9917
rect 2869 9877 2881 9911
rect 2915 9908 2927 9911
rect 5994 9908 6000 9920
rect 2915 9880 6000 9908
rect 2915 9877 2927 9880
rect 2869 9871 2927 9877
rect 5994 9868 6000 9880
rect 6052 9868 6058 9920
rect 7944 9908 7972 10007
rect 8018 10004 8024 10056
rect 8076 10044 8082 10056
rect 8386 10044 8392 10056
rect 8076 10016 8392 10044
rect 8076 10004 8082 10016
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 8478 10004 8484 10056
rect 8536 10044 8542 10056
rect 9585 10047 9643 10053
rect 9585 10044 9597 10047
rect 8536 10016 9597 10044
rect 8536 10004 8542 10016
rect 9585 10013 9597 10016
rect 9631 10013 9643 10047
rect 9585 10007 9643 10013
rect 10686 10004 10692 10056
rect 10744 10004 10750 10056
rect 12158 10004 12164 10056
rect 12216 10004 12222 10056
rect 12360 10044 12388 10072
rect 12268 10016 12388 10044
rect 8573 9979 8631 9985
rect 8573 9945 8585 9979
rect 8619 9976 8631 9979
rect 9674 9976 9680 9988
rect 8619 9948 9680 9976
rect 8619 9945 8631 9948
rect 8573 9939 8631 9945
rect 9674 9936 9680 9948
rect 9732 9936 9738 9988
rect 12268 9976 12296 10016
rect 13262 10004 13268 10056
rect 13320 10044 13326 10056
rect 14292 10044 14320 10075
rect 16298 10072 16304 10084
rect 16356 10072 16362 10124
rect 13320 10016 14320 10044
rect 13320 10004 13326 10016
rect 16114 10004 16120 10056
rect 16172 10044 16178 10056
rect 17328 10053 17356 10220
rect 17402 10208 17408 10220
rect 17460 10208 17466 10260
rect 18046 10208 18052 10260
rect 18104 10248 18110 10260
rect 18598 10248 18604 10260
rect 18104 10220 18604 10248
rect 18104 10208 18110 10220
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 22925 10251 22983 10257
rect 22925 10248 22937 10251
rect 18708 10220 22937 10248
rect 18708 10180 18736 10220
rect 22925 10217 22937 10220
rect 22971 10217 22983 10251
rect 22925 10211 22983 10217
rect 23750 10208 23756 10260
rect 23808 10248 23814 10260
rect 24029 10251 24087 10257
rect 24029 10248 24041 10251
rect 23808 10220 24041 10248
rect 23808 10208 23814 10220
rect 24029 10217 24041 10220
rect 24075 10217 24087 10251
rect 24029 10211 24087 10217
rect 24210 10208 24216 10260
rect 24268 10248 24274 10260
rect 25593 10251 25651 10257
rect 25593 10248 25605 10251
rect 24268 10220 25605 10248
rect 24268 10208 24274 10220
rect 25593 10217 25605 10220
rect 25639 10217 25651 10251
rect 25593 10211 25651 10217
rect 25958 10208 25964 10260
rect 26016 10208 26022 10260
rect 26053 10251 26111 10257
rect 26053 10217 26065 10251
rect 26099 10248 26111 10251
rect 28537 10251 28595 10257
rect 26099 10220 26924 10248
rect 26099 10217 26111 10220
rect 26053 10211 26111 10217
rect 18616 10152 18736 10180
rect 21729 10183 21787 10189
rect 17405 10115 17463 10121
rect 17405 10081 17417 10115
rect 17451 10112 17463 10115
rect 17494 10112 17500 10124
rect 17451 10084 17500 10112
rect 17451 10081 17463 10084
rect 17405 10075 17463 10081
rect 17494 10072 17500 10084
rect 17552 10072 17558 10124
rect 17589 10115 17647 10121
rect 17589 10081 17601 10115
rect 17635 10112 17647 10115
rect 18506 10112 18512 10124
rect 17635 10084 18512 10112
rect 17635 10081 17647 10084
rect 17589 10075 17647 10081
rect 18506 10072 18512 10084
rect 18564 10072 18570 10124
rect 18616 10121 18644 10152
rect 21729 10149 21741 10183
rect 21775 10180 21787 10183
rect 22094 10180 22100 10192
rect 21775 10152 22100 10180
rect 21775 10149 21787 10152
rect 21729 10143 21787 10149
rect 22094 10140 22100 10152
rect 22152 10140 22158 10192
rect 24581 10183 24639 10189
rect 24581 10180 24593 10183
rect 22296 10152 24593 10180
rect 18601 10115 18659 10121
rect 18601 10081 18613 10115
rect 18647 10081 18659 10115
rect 18601 10075 18659 10081
rect 18785 10115 18843 10121
rect 18785 10081 18797 10115
rect 18831 10112 18843 10115
rect 19429 10115 19487 10121
rect 18831 10084 19288 10112
rect 18831 10081 18843 10084
rect 18785 10075 18843 10081
rect 17313 10047 17371 10053
rect 16172 10016 17264 10044
rect 16172 10004 16178 10016
rect 11716 9948 12296 9976
rect 11716 9908 11744 9948
rect 13170 9936 13176 9988
rect 13228 9976 13234 9988
rect 14458 9976 14464 9988
rect 13228 9948 14464 9976
rect 13228 9936 13234 9948
rect 14458 9936 14464 9948
rect 14516 9936 14522 9988
rect 14553 9979 14611 9985
rect 14553 9945 14565 9979
rect 14599 9976 14611 9979
rect 14826 9976 14832 9988
rect 14599 9948 14832 9976
rect 14599 9945 14611 9948
rect 14553 9939 14611 9945
rect 14826 9936 14832 9948
rect 14884 9936 14890 9988
rect 15286 9936 15292 9988
rect 15344 9936 15350 9988
rect 17236 9976 17264 10016
rect 17313 10013 17325 10047
rect 17359 10013 17371 10047
rect 17512 10044 17540 10072
rect 17770 10044 17776 10056
rect 17512 10016 17776 10044
rect 17313 10007 17371 10013
rect 17770 10004 17776 10016
rect 17828 10004 17834 10056
rect 17954 9976 17960 9988
rect 17236 9948 17960 9976
rect 17954 9936 17960 9948
rect 18012 9936 18018 9988
rect 7944 9880 11744 9908
rect 11790 9868 11796 9920
rect 11848 9868 11854 9920
rect 13354 9868 13360 9920
rect 13412 9868 13418 9920
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 16577 9911 16635 9917
rect 16577 9908 16589 9911
rect 13872 9880 16589 9908
rect 13872 9868 13878 9880
rect 16577 9877 16589 9880
rect 16623 9908 16635 9911
rect 18046 9908 18052 9920
rect 16623 9880 18052 9908
rect 16623 9877 16635 9880
rect 16577 9871 16635 9877
rect 18046 9868 18052 9880
rect 18104 9868 18110 9920
rect 18138 9868 18144 9920
rect 18196 9868 18202 9920
rect 18509 9911 18567 9917
rect 18509 9877 18521 9911
rect 18555 9908 18567 9911
rect 19150 9908 19156 9920
rect 18555 9880 19156 9908
rect 18555 9877 18567 9880
rect 18509 9871 18567 9877
rect 19150 9868 19156 9880
rect 19208 9868 19214 9920
rect 19260 9908 19288 10084
rect 19429 10081 19441 10115
rect 19475 10112 19487 10115
rect 19702 10112 19708 10124
rect 19475 10084 19708 10112
rect 19475 10081 19487 10084
rect 19429 10075 19487 10081
rect 19702 10072 19708 10084
rect 19760 10072 19766 10124
rect 20346 10072 20352 10124
rect 20404 10112 20410 10124
rect 21177 10115 21235 10121
rect 21177 10112 21189 10115
rect 20404 10084 21189 10112
rect 20404 10072 20410 10084
rect 21177 10081 21189 10084
rect 21223 10081 21235 10115
rect 21177 10075 21235 10081
rect 22002 10072 22008 10124
rect 22060 10112 22066 10124
rect 22296 10112 22324 10152
rect 24581 10149 24593 10152
rect 24627 10149 24639 10183
rect 24762 10180 24768 10192
rect 24581 10143 24639 10149
rect 24688 10152 24768 10180
rect 22060 10084 22324 10112
rect 22373 10115 22431 10121
rect 22060 10072 22066 10084
rect 22373 10081 22385 10115
rect 22419 10112 22431 10115
rect 22646 10112 22652 10124
rect 22419 10084 22652 10112
rect 22419 10081 22431 10084
rect 22373 10075 22431 10081
rect 22646 10072 22652 10084
rect 22704 10072 22710 10124
rect 23382 10072 23388 10124
rect 23440 10072 23446 10124
rect 23477 10115 23535 10121
rect 23477 10081 23489 10115
rect 23523 10081 23535 10115
rect 23477 10075 23535 10081
rect 22097 10047 22155 10053
rect 22097 10013 22109 10047
rect 22143 10044 22155 10047
rect 23290 10044 23296 10056
rect 22143 10016 23296 10044
rect 22143 10013 22155 10016
rect 22097 10007 22155 10013
rect 23290 10004 23296 10016
rect 23348 10004 23354 10056
rect 19334 9936 19340 9988
rect 19392 9976 19398 9988
rect 19705 9979 19763 9985
rect 19705 9976 19717 9979
rect 19392 9948 19717 9976
rect 19392 9936 19398 9948
rect 19705 9945 19717 9948
rect 19751 9945 19763 9979
rect 19705 9939 19763 9945
rect 20714 9936 20720 9988
rect 20772 9936 20778 9988
rect 21266 9936 21272 9988
rect 21324 9976 21330 9988
rect 22002 9976 22008 9988
rect 21324 9948 22008 9976
rect 21324 9936 21330 9948
rect 22002 9936 22008 9948
rect 22060 9936 22066 9988
rect 22646 9936 22652 9988
rect 22704 9976 22710 9988
rect 23492 9976 23520 10075
rect 23566 10072 23572 10124
rect 23624 10112 23630 10124
rect 24688 10112 24716 10152
rect 24762 10140 24768 10152
rect 24820 10180 24826 10192
rect 25976 10180 26004 10208
rect 24820 10152 26004 10180
rect 24820 10140 24826 10152
rect 23624 10084 24716 10112
rect 23624 10072 23630 10084
rect 25222 10072 25228 10124
rect 25280 10072 25286 10124
rect 25869 10115 25927 10121
rect 25869 10081 25881 10115
rect 25915 10112 25927 10115
rect 25958 10112 25964 10124
rect 25915 10084 25964 10112
rect 25915 10081 25927 10084
rect 25869 10075 25927 10081
rect 24946 10004 24952 10056
rect 25004 10004 25010 10056
rect 25041 10047 25099 10053
rect 25041 10013 25053 10047
rect 25087 10044 25099 10047
rect 25314 10044 25320 10056
rect 25087 10016 25320 10044
rect 25087 10013 25099 10016
rect 25041 10007 25099 10013
rect 25314 10004 25320 10016
rect 25372 10044 25378 10056
rect 25884 10044 25912 10075
rect 25958 10072 25964 10084
rect 26016 10072 26022 10124
rect 25372 10016 25912 10044
rect 25372 10004 25378 10016
rect 22704 9948 23520 9976
rect 22704 9936 22710 9948
rect 24394 9936 24400 9988
rect 24452 9976 24458 9988
rect 25406 9976 25412 9988
rect 24452 9948 25412 9976
rect 24452 9936 24458 9948
rect 25406 9936 25412 9948
rect 25464 9936 25470 9988
rect 20070 9908 20076 9920
rect 19260 9880 20076 9908
rect 20070 9868 20076 9880
rect 20128 9868 20134 9920
rect 22186 9868 22192 9920
rect 22244 9868 22250 9920
rect 22922 9868 22928 9920
rect 22980 9908 22986 9920
rect 23293 9911 23351 9917
rect 23293 9908 23305 9911
rect 22980 9880 23305 9908
rect 22980 9868 22986 9880
rect 23293 9877 23305 9880
rect 23339 9908 23351 9911
rect 26068 9908 26096 10211
rect 26786 10072 26792 10124
rect 26844 10072 26850 10124
rect 26896 10112 26924 10220
rect 28537 10217 28549 10251
rect 28583 10248 28595 10251
rect 28902 10248 28908 10260
rect 28583 10220 28908 10248
rect 28583 10217 28595 10220
rect 28537 10211 28595 10217
rect 28902 10208 28908 10220
rect 28960 10208 28966 10260
rect 30926 10208 30932 10260
rect 30984 10248 30990 10260
rect 30984 10220 32444 10248
rect 30984 10208 30990 10220
rect 28442 10140 28448 10192
rect 28500 10180 28506 10192
rect 28500 10152 32352 10180
rect 28500 10140 28506 10152
rect 29178 10112 29184 10124
rect 26896 10084 29184 10112
rect 29178 10072 29184 10084
rect 29236 10072 29242 10124
rect 29546 10072 29552 10124
rect 29604 10112 29610 10124
rect 30193 10115 30251 10121
rect 30193 10112 30205 10115
rect 29604 10084 30205 10112
rect 29604 10072 29610 10084
rect 30193 10081 30205 10084
rect 30239 10081 30251 10115
rect 30193 10075 30251 10081
rect 30374 10072 30380 10124
rect 30432 10072 30438 10124
rect 31386 10072 31392 10124
rect 31444 10112 31450 10124
rect 31757 10115 31815 10121
rect 31757 10112 31769 10115
rect 31444 10084 31769 10112
rect 31444 10072 31450 10084
rect 31757 10081 31769 10084
rect 31803 10081 31815 10115
rect 31757 10075 31815 10081
rect 30101 10047 30159 10053
rect 30101 10013 30113 10047
rect 30147 10044 30159 10047
rect 32324 10044 32352 10152
rect 32416 10112 32444 10220
rect 33778 10208 33784 10260
rect 33836 10248 33842 10260
rect 36446 10248 36452 10260
rect 33836 10220 36452 10248
rect 33836 10208 33842 10220
rect 36446 10208 36452 10220
rect 36504 10208 36510 10260
rect 36630 10208 36636 10260
rect 36688 10248 36694 10260
rect 36909 10251 36967 10257
rect 36909 10248 36921 10251
rect 36688 10220 36921 10248
rect 36688 10208 36694 10220
rect 36909 10217 36921 10220
rect 36955 10217 36967 10251
rect 36909 10211 36967 10217
rect 37461 10251 37519 10257
rect 37461 10217 37473 10251
rect 37507 10248 37519 10251
rect 38654 10248 38660 10260
rect 37507 10220 38660 10248
rect 37507 10217 37519 10220
rect 37461 10211 37519 10217
rect 38654 10208 38660 10220
rect 38712 10208 38718 10260
rect 40681 10251 40739 10257
rect 40681 10217 40693 10251
rect 40727 10248 40739 10251
rect 41138 10248 41144 10260
rect 40727 10220 41144 10248
rect 40727 10217 40739 10220
rect 40681 10211 40739 10217
rect 41138 10208 41144 10220
rect 41196 10208 41202 10260
rect 43714 10208 43720 10260
rect 43772 10208 43778 10260
rect 45097 10251 45155 10257
rect 45097 10217 45109 10251
rect 45143 10248 45155 10251
rect 45186 10248 45192 10260
rect 45143 10220 45192 10248
rect 45143 10217 45155 10220
rect 45097 10211 45155 10217
rect 45186 10208 45192 10220
rect 45244 10208 45250 10260
rect 45557 10251 45615 10257
rect 45557 10217 45569 10251
rect 45603 10248 45615 10251
rect 48406 10248 48412 10260
rect 45603 10220 48412 10248
rect 45603 10217 45615 10220
rect 45557 10211 45615 10217
rect 48406 10208 48412 10220
rect 48464 10208 48470 10260
rect 32585 10183 32643 10189
rect 32585 10149 32597 10183
rect 32631 10180 32643 10183
rect 34514 10180 34520 10192
rect 32631 10152 34520 10180
rect 32631 10149 32643 10152
rect 32585 10143 32643 10149
rect 34514 10140 34520 10152
rect 34572 10140 34578 10192
rect 40402 10180 40408 10192
rect 36832 10152 40408 10180
rect 33137 10115 33195 10121
rect 33137 10112 33149 10115
rect 32416 10084 33149 10112
rect 33137 10081 33149 10084
rect 33183 10081 33195 10115
rect 33137 10075 33195 10081
rect 33502 10072 33508 10124
rect 33560 10112 33566 10124
rect 34885 10115 34943 10121
rect 34885 10112 34897 10115
rect 33560 10084 34897 10112
rect 33560 10072 33566 10084
rect 34885 10081 34897 10084
rect 34931 10081 34943 10115
rect 34885 10075 34943 10081
rect 35161 10115 35219 10121
rect 35161 10081 35173 10115
rect 35207 10112 35219 10115
rect 36832 10112 36860 10152
rect 40402 10140 40408 10152
rect 40460 10140 40466 10192
rect 41417 10183 41475 10189
rect 41417 10149 41429 10183
rect 41463 10180 41475 10183
rect 41463 10152 46152 10180
rect 41463 10149 41475 10152
rect 41417 10143 41475 10149
rect 35207 10084 36860 10112
rect 35207 10081 35219 10084
rect 35161 10075 35219 10081
rect 36906 10072 36912 10124
rect 36964 10112 36970 10124
rect 37921 10115 37979 10121
rect 37921 10112 37933 10115
rect 36964 10084 37933 10112
rect 36964 10072 36970 10084
rect 37921 10081 37933 10084
rect 37967 10081 37979 10115
rect 37921 10075 37979 10081
rect 38010 10072 38016 10124
rect 38068 10072 38074 10124
rect 39301 10115 39359 10121
rect 39301 10112 39313 10115
rect 38120 10084 39313 10112
rect 32953 10047 33011 10053
rect 32953 10044 32965 10047
rect 30147 10016 31754 10044
rect 32324 10016 32965 10044
rect 30147 10013 30159 10016
rect 30101 10007 30159 10013
rect 27065 9979 27123 9985
rect 27065 9945 27077 9979
rect 27111 9945 27123 9979
rect 28626 9976 28632 9988
rect 28290 9948 28632 9976
rect 27065 9939 27123 9945
rect 23339 9880 26096 9908
rect 27080 9908 27108 9939
rect 28626 9936 28632 9948
rect 28684 9976 28690 9988
rect 29270 9976 29276 9988
rect 28684 9948 29276 9976
rect 28684 9936 28690 9948
rect 29270 9936 29276 9948
rect 29328 9936 29334 9988
rect 31573 9979 31631 9985
rect 31573 9976 31585 9979
rect 29748 9948 31585 9976
rect 27798 9908 27804 9920
rect 27080 9880 27804 9908
rect 23339 9877 23351 9880
rect 23293 9871 23351 9877
rect 27798 9868 27804 9880
rect 27856 9868 27862 9920
rect 28074 9868 28080 9920
rect 28132 9908 28138 9920
rect 29748 9917 29776 9948
rect 31573 9945 31585 9948
rect 31619 9945 31631 9979
rect 31726 9976 31754 10016
rect 32953 10013 32965 10016
rect 32999 10013 33011 10047
rect 32953 10007 33011 10013
rect 36446 10004 36452 10056
rect 36504 10044 36510 10056
rect 38120 10044 38148 10084
rect 39301 10081 39313 10084
rect 39347 10081 39359 10115
rect 39301 10075 39359 10081
rect 39390 10072 39396 10124
rect 39448 10112 39454 10124
rect 39448 10084 42012 10112
rect 39448 10072 39454 10084
rect 36504 10016 38148 10044
rect 36504 10004 36510 10016
rect 38654 10004 38660 10056
rect 38712 10004 38718 10056
rect 40037 10047 40095 10053
rect 40037 10013 40049 10047
rect 40083 10044 40095 10047
rect 40678 10044 40684 10056
rect 40083 10016 40684 10044
rect 40083 10013 40095 10016
rect 40037 10007 40095 10013
rect 40678 10004 40684 10016
rect 40736 10004 40742 10056
rect 41984 10053 42012 10084
rect 42058 10072 42064 10124
rect 42116 10112 42122 10124
rect 42889 10115 42947 10121
rect 42889 10112 42901 10115
rect 42116 10084 42901 10112
rect 42116 10072 42122 10084
rect 42889 10081 42901 10084
rect 42935 10081 42947 10115
rect 42889 10075 42947 10081
rect 41969 10047 42027 10053
rect 41969 10013 41981 10047
rect 42015 10013 42027 10047
rect 41969 10007 42027 10013
rect 31726 9948 32352 9976
rect 31573 9939 31631 9945
rect 28997 9911 29055 9917
rect 28997 9908 29009 9911
rect 28132 9880 29009 9908
rect 28132 9868 28138 9880
rect 28997 9877 29009 9880
rect 29043 9877 29055 9911
rect 28997 9871 29055 9877
rect 29733 9911 29791 9917
rect 29733 9877 29745 9911
rect 29779 9877 29791 9911
rect 29733 9871 29791 9877
rect 30650 9868 30656 9920
rect 30708 9908 30714 9920
rect 30834 9908 30840 9920
rect 30708 9880 30840 9908
rect 30708 9868 30714 9880
rect 30834 9868 30840 9880
rect 30892 9868 30898 9920
rect 31110 9868 31116 9920
rect 31168 9908 31174 9920
rect 31205 9911 31263 9917
rect 31205 9908 31217 9911
rect 31168 9880 31217 9908
rect 31168 9868 31174 9880
rect 31205 9877 31217 9880
rect 31251 9877 31263 9911
rect 31205 9871 31263 9877
rect 31294 9868 31300 9920
rect 31352 9908 31358 9920
rect 31665 9911 31723 9917
rect 31665 9908 31677 9911
rect 31352 9880 31677 9908
rect 31352 9868 31358 9880
rect 31665 9877 31677 9880
rect 31711 9877 31723 9911
rect 32324 9908 32352 9948
rect 32398 9936 32404 9988
rect 32456 9976 32462 9988
rect 33045 9979 33103 9985
rect 33045 9976 33057 9979
rect 32456 9948 33057 9976
rect 32456 9936 32462 9948
rect 33045 9945 33057 9948
rect 33091 9945 33103 9979
rect 33045 9939 33103 9945
rect 36170 9936 36176 9988
rect 36228 9936 36234 9988
rect 37829 9979 37887 9985
rect 37829 9976 37841 9979
rect 36464 9948 37841 9976
rect 34146 9908 34152 9920
rect 32324 9880 34152 9908
rect 31665 9871 31723 9877
rect 34146 9868 34152 9880
rect 34204 9868 34210 9920
rect 34974 9868 34980 9920
rect 35032 9908 35038 9920
rect 36464 9908 36492 9948
rect 37829 9945 37841 9948
rect 37875 9945 37887 9979
rect 37829 9939 37887 9945
rect 37936 9948 39804 9976
rect 35032 9880 36492 9908
rect 35032 9868 35038 9880
rect 36630 9868 36636 9920
rect 36688 9868 36694 9920
rect 37090 9868 37096 9920
rect 37148 9868 37154 9920
rect 37182 9868 37188 9920
rect 37240 9908 37246 9920
rect 37936 9908 37964 9948
rect 37240 9880 37964 9908
rect 37240 9868 37246 9880
rect 38102 9868 38108 9920
rect 38160 9908 38166 9920
rect 39577 9911 39635 9917
rect 39577 9908 39589 9911
rect 38160 9880 39589 9908
rect 38160 9868 38166 9880
rect 39577 9877 39589 9880
rect 39623 9877 39635 9911
rect 39776 9908 39804 9948
rect 39850 9936 39856 9988
rect 39908 9976 39914 9988
rect 41233 9979 41291 9985
rect 41233 9976 41245 9979
rect 39908 9948 41245 9976
rect 39908 9936 39914 9948
rect 41233 9945 41245 9948
rect 41279 9945 41291 9979
rect 41984 9976 42012 10007
rect 42610 10004 42616 10056
rect 42668 10044 42674 10056
rect 43806 10044 43812 10056
rect 42668 10016 43812 10044
rect 42668 10004 42674 10016
rect 43806 10004 43812 10016
rect 43864 10004 43870 10056
rect 44450 10004 44456 10056
rect 44508 10004 44514 10056
rect 45373 10047 45431 10053
rect 45373 10013 45385 10047
rect 45419 10044 45431 10047
rect 45554 10044 45560 10056
rect 45419 10016 45560 10044
rect 45419 10013 45431 10016
rect 45373 10007 45431 10013
rect 45554 10004 45560 10016
rect 45612 10004 45618 10056
rect 46124 10053 46152 10152
rect 46198 10140 46204 10192
rect 46256 10180 46262 10192
rect 47670 10180 47676 10192
rect 46256 10152 47676 10180
rect 46256 10140 46262 10152
rect 47670 10140 47676 10152
rect 47728 10140 47734 10192
rect 46842 10072 46848 10124
rect 46900 10072 46906 10124
rect 49142 10072 49148 10124
rect 49200 10072 49206 10124
rect 46109 10047 46167 10053
rect 46109 10013 46121 10047
rect 46155 10013 46167 10047
rect 46109 10007 46167 10013
rect 47949 10047 48007 10053
rect 47949 10013 47961 10047
rect 47995 10013 48007 10047
rect 47949 10007 48007 10013
rect 43901 9979 43959 9985
rect 43901 9976 43913 9979
rect 41984 9948 43913 9976
rect 41233 9939 41291 9945
rect 43901 9945 43913 9948
rect 43947 9945 43959 9979
rect 43901 9939 43959 9945
rect 44637 9979 44695 9985
rect 44637 9945 44649 9979
rect 44683 9976 44695 9979
rect 47964 9976 47992 10007
rect 44683 9948 47992 9976
rect 44683 9945 44695 9948
rect 44637 9939 44695 9945
rect 41966 9908 41972 9920
rect 39776 9880 41972 9908
rect 39577 9871 39635 9877
rect 41966 9868 41972 9880
rect 42024 9868 42030 9920
rect 42058 9868 42064 9920
rect 42116 9868 42122 9920
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 2406 9664 2412 9716
rect 2464 9664 2470 9716
rect 3421 9707 3479 9713
rect 3421 9673 3433 9707
rect 3467 9704 3479 9707
rect 3602 9704 3608 9716
rect 3467 9676 3608 9704
rect 3467 9673 3479 9676
rect 3421 9667 3479 9673
rect 3602 9664 3608 9676
rect 3660 9664 3666 9716
rect 4065 9707 4123 9713
rect 4065 9673 4077 9707
rect 4111 9673 4123 9707
rect 4065 9667 4123 9673
rect 1210 9528 1216 9580
rect 1268 9568 1274 9580
rect 1581 9571 1639 9577
rect 1581 9568 1593 9571
rect 1268 9540 1593 9568
rect 1268 9528 1274 9540
rect 1581 9537 1593 9540
rect 1627 9568 1639 9571
rect 2130 9568 2136 9580
rect 1627 9540 2136 9568
rect 1627 9537 1639 9540
rect 1581 9531 1639 9537
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9568 2375 9571
rect 2961 9571 3019 9577
rect 2961 9568 2973 9571
rect 2363 9540 2973 9568
rect 2363 9537 2375 9540
rect 2317 9531 2375 9537
rect 2961 9537 2973 9540
rect 3007 9568 3019 9571
rect 3510 9568 3516 9580
rect 3007 9540 3516 9568
rect 3007 9537 3019 9540
rect 2961 9531 3019 9537
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 3602 9528 3608 9580
rect 3660 9568 3666 9580
rect 3970 9568 3976 9580
rect 3660 9540 3976 9568
rect 3660 9528 3666 9540
rect 3970 9528 3976 9540
rect 4028 9528 4034 9580
rect 4080 9500 4108 9667
rect 8294 9664 8300 9716
rect 8352 9704 8358 9716
rect 13170 9704 13176 9716
rect 8352 9676 13176 9704
rect 8352 9664 8358 9676
rect 13170 9664 13176 9676
rect 13228 9664 13234 9716
rect 13446 9664 13452 9716
rect 13504 9704 13510 9716
rect 15746 9704 15752 9716
rect 13504 9676 15752 9704
rect 13504 9664 13510 9676
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 16206 9664 16212 9716
rect 16264 9704 16270 9716
rect 16942 9704 16948 9716
rect 16264 9676 16948 9704
rect 16264 9664 16270 9676
rect 16942 9664 16948 9676
rect 17000 9664 17006 9716
rect 17126 9664 17132 9716
rect 17184 9704 17190 9716
rect 17494 9704 17500 9716
rect 17184 9676 17500 9704
rect 17184 9664 17190 9676
rect 17494 9664 17500 9676
rect 17552 9664 17558 9716
rect 17770 9664 17776 9716
rect 17828 9704 17834 9716
rect 18138 9704 18144 9716
rect 17828 9676 18144 9704
rect 17828 9664 17834 9676
rect 18138 9664 18144 9676
rect 18196 9664 18202 9716
rect 18414 9664 18420 9716
rect 18472 9664 18478 9716
rect 18506 9664 18512 9716
rect 18564 9704 18570 9716
rect 20438 9704 20444 9716
rect 18564 9676 20444 9704
rect 18564 9664 18570 9676
rect 20438 9664 20444 9676
rect 20496 9664 20502 9716
rect 21358 9664 21364 9716
rect 21416 9704 21422 9716
rect 22005 9707 22063 9713
rect 22005 9704 22017 9707
rect 21416 9676 22017 9704
rect 21416 9664 21422 9676
rect 22005 9673 22017 9676
rect 22051 9673 22063 9707
rect 22005 9667 22063 9673
rect 23201 9707 23259 9713
rect 23201 9673 23213 9707
rect 23247 9704 23259 9707
rect 23382 9704 23388 9716
rect 23247 9676 23388 9704
rect 23247 9673 23259 9676
rect 23201 9667 23259 9673
rect 23382 9664 23388 9676
rect 23440 9664 23446 9716
rect 27816 9676 29500 9704
rect 4706 9596 4712 9648
rect 4764 9596 4770 9648
rect 5718 9596 5724 9648
rect 5776 9636 5782 9648
rect 7929 9639 7987 9645
rect 7929 9636 7941 9639
rect 5776 9608 7941 9636
rect 5776 9596 5782 9608
rect 7929 9605 7941 9608
rect 7975 9605 7987 9639
rect 7929 9599 7987 9605
rect 8665 9639 8723 9645
rect 8665 9605 8677 9639
rect 8711 9636 8723 9639
rect 8757 9639 8815 9645
rect 8757 9636 8769 9639
rect 8711 9608 8769 9636
rect 8711 9605 8723 9608
rect 8665 9599 8723 9605
rect 8757 9605 8769 9608
rect 8803 9636 8815 9639
rect 11054 9636 11060 9648
rect 8803 9608 11060 9636
rect 8803 9605 8815 9608
rect 8757 9599 8815 9605
rect 11054 9596 11060 9608
rect 11112 9596 11118 9648
rect 11238 9596 11244 9648
rect 11296 9636 11302 9648
rect 13541 9639 13599 9645
rect 13541 9636 13553 9639
rect 11296 9608 13553 9636
rect 11296 9596 11302 9608
rect 13541 9605 13553 9608
rect 13587 9605 13599 9639
rect 13541 9599 13599 9605
rect 13998 9596 14004 9648
rect 14056 9596 14062 9648
rect 16960 9636 16988 9664
rect 16960 9608 17618 9636
rect 4154 9528 4160 9580
rect 4212 9568 4218 9580
rect 4249 9571 4307 9577
rect 4249 9568 4261 9571
rect 4212 9540 4261 9568
rect 4212 9528 4218 9540
rect 4249 9537 4261 9540
rect 4295 9568 4307 9571
rect 4525 9571 4583 9577
rect 4525 9568 4537 9571
rect 4295 9540 4537 9568
rect 4295 9537 4307 9540
rect 4249 9531 4307 9537
rect 4525 9537 4537 9540
rect 4571 9537 4583 9571
rect 4525 9531 4583 9537
rect 5350 9528 5356 9580
rect 5408 9528 5414 9580
rect 5994 9528 6000 9580
rect 6052 9528 6058 9580
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9568 6607 9571
rect 9214 9568 9220 9580
rect 6595 9540 9220 9568
rect 6595 9537 6607 9540
rect 6549 9531 6607 9537
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 9401 9571 9459 9577
rect 9401 9537 9413 9571
rect 9447 9568 9459 9571
rect 10318 9568 10324 9580
rect 9447 9540 10324 9568
rect 9447 9537 9459 9540
rect 9401 9531 9459 9537
rect 10318 9528 10324 9540
rect 10376 9528 10382 9580
rect 10502 9528 10508 9580
rect 10560 9528 10566 9580
rect 12158 9528 12164 9580
rect 12216 9528 12222 9580
rect 13262 9528 13268 9580
rect 13320 9528 13326 9580
rect 15010 9528 15016 9580
rect 15068 9568 15074 9580
rect 15470 9568 15476 9580
rect 15068 9540 15476 9568
rect 15068 9528 15074 9540
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 15841 9571 15899 9577
rect 15841 9537 15853 9571
rect 15887 9568 15899 9571
rect 16390 9568 16396 9580
rect 15887 9540 16396 9568
rect 15887 9537 15899 9540
rect 15841 9531 15899 9537
rect 16390 9528 16396 9540
rect 16448 9528 16454 9580
rect 16758 9528 16764 9580
rect 16816 9568 16822 9580
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16816 9540 16865 9568
rect 16816 9528 16822 9540
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 6178 9500 6184 9512
rect 4080 9472 6184 9500
rect 6178 9460 6184 9472
rect 6236 9460 6242 9512
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9469 6883 9503
rect 6825 9463 6883 9469
rect 1762 9392 1768 9444
rect 1820 9392 1826 9444
rect 2774 9392 2780 9444
rect 2832 9392 2838 9444
rect 6840 9432 6868 9463
rect 6914 9460 6920 9512
rect 6972 9500 6978 9512
rect 9950 9500 9956 9512
rect 6972 9472 9956 9500
rect 6972 9460 6978 9472
rect 9950 9460 9956 9472
rect 10008 9460 10014 9512
rect 10045 9503 10103 9509
rect 10045 9469 10057 9503
rect 10091 9500 10103 9503
rect 11974 9500 11980 9512
rect 10091 9472 11980 9500
rect 10091 9469 10103 9472
rect 10045 9463 10103 9469
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 13538 9460 13544 9512
rect 13596 9500 13602 9512
rect 15933 9503 15991 9509
rect 15933 9500 15945 9503
rect 13596 9472 15945 9500
rect 13596 9460 13602 9472
rect 15933 9469 15945 9472
rect 15979 9469 15991 9503
rect 15933 9463 15991 9469
rect 16025 9503 16083 9509
rect 16025 9469 16037 9503
rect 16071 9469 16083 9503
rect 16025 9463 16083 9469
rect 3344 9404 6868 9432
rect 2498 9324 2504 9376
rect 2556 9364 2562 9376
rect 3344 9364 3372 9404
rect 7190 9392 7196 9444
rect 7248 9432 7254 9444
rect 11149 9435 11207 9441
rect 11149 9432 11161 9435
rect 7248 9404 9674 9432
rect 7248 9392 7254 9404
rect 2556 9336 3372 9364
rect 5169 9367 5227 9373
rect 2556 9324 2562 9336
rect 5169 9333 5181 9367
rect 5215 9364 5227 9367
rect 5534 9364 5540 9376
rect 5215 9336 5540 9364
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 5813 9367 5871 9373
rect 5813 9333 5825 9367
rect 5859 9364 5871 9367
rect 7742 9364 7748 9376
rect 5859 9336 7748 9364
rect 5859 9333 5871 9336
rect 5813 9327 5871 9333
rect 7742 9324 7748 9336
rect 7800 9324 7806 9376
rect 8018 9324 8024 9376
rect 8076 9324 8082 9376
rect 9646 9364 9674 9404
rect 9876 9404 11161 9432
rect 9876 9364 9904 9404
rect 11149 9401 11161 9404
rect 11195 9401 11207 9435
rect 11885 9435 11943 9441
rect 11885 9432 11897 9435
rect 11149 9395 11207 9401
rect 11256 9404 11897 9432
rect 9646 9336 9904 9364
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 11256 9364 11284 9404
rect 11885 9401 11897 9404
rect 11931 9432 11943 9435
rect 13262 9432 13268 9444
rect 11931 9404 13268 9432
rect 11931 9401 11943 9404
rect 11885 9395 11943 9401
rect 13262 9392 13268 9404
rect 13320 9392 13326 9444
rect 16040 9432 16068 9463
rect 16206 9460 16212 9512
rect 16264 9500 16270 9512
rect 16776 9500 16804 9528
rect 18432 9512 18460 9664
rect 18782 9596 18788 9648
rect 18840 9636 18846 9648
rect 19702 9636 19708 9648
rect 18840 9608 19708 9636
rect 18840 9596 18846 9608
rect 19702 9596 19708 9608
rect 19760 9596 19766 9648
rect 21542 9596 21548 9648
rect 21600 9596 21606 9648
rect 22094 9596 22100 9648
rect 22152 9636 22158 9648
rect 22152 9608 22508 9636
rect 22152 9596 22158 9608
rect 20714 9528 20720 9580
rect 20772 9528 20778 9580
rect 22186 9528 22192 9580
rect 22244 9568 22250 9580
rect 22480 9577 22508 9608
rect 24394 9596 24400 9648
rect 24452 9596 24458 9648
rect 27816 9636 27844 9676
rect 28442 9636 28448 9648
rect 26344 9608 27844 9636
rect 27908 9608 28448 9636
rect 22373 9571 22431 9577
rect 22373 9568 22385 9571
rect 22244 9540 22385 9568
rect 22244 9528 22250 9540
rect 22373 9537 22385 9540
rect 22419 9537 22431 9571
rect 22373 9531 22431 9537
rect 22465 9571 22523 9577
rect 22465 9537 22477 9571
rect 22511 9568 22523 9571
rect 23290 9568 23296 9580
rect 22511 9540 23296 9568
rect 22511 9537 22523 9540
rect 22465 9531 22523 9537
rect 23290 9528 23296 9540
rect 23348 9528 23354 9580
rect 23474 9528 23480 9580
rect 23532 9528 23538 9580
rect 25958 9528 25964 9580
rect 26016 9568 26022 9580
rect 26237 9571 26295 9577
rect 26237 9568 26249 9571
rect 26016 9540 26249 9568
rect 26016 9528 26022 9540
rect 26237 9537 26249 9540
rect 26283 9537 26295 9571
rect 26237 9531 26295 9537
rect 16264 9472 16804 9500
rect 16264 9460 16270 9472
rect 17126 9460 17132 9512
rect 17184 9460 17190 9512
rect 18414 9460 18420 9512
rect 18472 9460 18478 9512
rect 18506 9460 18512 9512
rect 18564 9500 18570 9512
rect 18877 9503 18935 9509
rect 18877 9500 18889 9503
rect 18564 9472 18889 9500
rect 18564 9460 18570 9472
rect 18877 9469 18889 9472
rect 18923 9469 18935 9503
rect 18877 9463 18935 9469
rect 19242 9460 19248 9512
rect 19300 9500 19306 9512
rect 19337 9503 19395 9509
rect 19337 9500 19349 9503
rect 19300 9472 19349 9500
rect 19300 9460 19306 9472
rect 19337 9469 19349 9472
rect 19383 9469 19395 9503
rect 19613 9503 19671 9509
rect 19613 9500 19625 9503
rect 19337 9463 19395 9469
rect 19444 9472 19625 9500
rect 15304 9404 16068 9432
rect 15304 9376 15332 9404
rect 18322 9392 18328 9444
rect 18380 9432 18386 9444
rect 19444 9432 19472 9472
rect 19613 9469 19625 9472
rect 19659 9469 19671 9503
rect 19613 9463 19671 9469
rect 20070 9460 20076 9512
rect 20128 9500 20134 9512
rect 22278 9500 22284 9512
rect 20128 9472 22284 9500
rect 20128 9460 20134 9472
rect 22278 9460 22284 9472
rect 22336 9460 22342 9512
rect 22557 9503 22615 9509
rect 22557 9469 22569 9503
rect 22603 9469 22615 9503
rect 22557 9463 22615 9469
rect 18380 9404 19472 9432
rect 21453 9435 21511 9441
rect 18380 9392 18386 9404
rect 21453 9401 21465 9435
rect 21499 9432 21511 9435
rect 21818 9432 21824 9444
rect 21499 9404 21824 9432
rect 21499 9401 21511 9404
rect 21453 9395 21511 9401
rect 21818 9392 21824 9404
rect 21876 9392 21882 9444
rect 22002 9392 22008 9444
rect 22060 9432 22066 9444
rect 22572 9432 22600 9463
rect 23750 9460 23756 9512
rect 23808 9460 23814 9512
rect 24302 9460 24308 9512
rect 24360 9500 24366 9512
rect 26344 9509 26372 9608
rect 27908 9577 27936 9608
rect 28442 9596 28448 9608
rect 28500 9596 28506 9648
rect 27893 9571 27951 9577
rect 27893 9537 27905 9571
rect 27939 9537 27951 9571
rect 27893 9531 27951 9537
rect 29270 9528 29276 9580
rect 29328 9528 29334 9580
rect 29472 9568 29500 9676
rect 30006 9664 30012 9716
rect 30064 9704 30070 9716
rect 32398 9704 32404 9716
rect 30064 9676 32404 9704
rect 30064 9664 30070 9676
rect 32398 9664 32404 9676
rect 32456 9664 32462 9716
rect 32858 9664 32864 9716
rect 32916 9704 32922 9716
rect 34238 9704 34244 9716
rect 32916 9676 34244 9704
rect 32916 9664 32922 9676
rect 34238 9664 34244 9676
rect 34296 9664 34302 9716
rect 36372 9676 36860 9704
rect 29638 9596 29644 9648
rect 29696 9636 29702 9648
rect 30101 9639 30159 9645
rect 30101 9636 30113 9639
rect 29696 9608 30113 9636
rect 29696 9596 29702 9608
rect 30101 9605 30113 9608
rect 30147 9605 30159 9639
rect 30101 9599 30159 9605
rect 30208 9608 32260 9636
rect 30208 9568 30236 9608
rect 29472 9540 30236 9568
rect 30466 9528 30472 9580
rect 30524 9568 30530 9580
rect 30653 9571 30711 9577
rect 30653 9568 30665 9571
rect 30524 9540 30665 9568
rect 30524 9528 30530 9540
rect 30653 9537 30665 9540
rect 30699 9537 30711 9571
rect 30653 9531 30711 9537
rect 25501 9503 25559 9509
rect 25501 9500 25513 9503
rect 24360 9472 25513 9500
rect 24360 9460 24366 9472
rect 25501 9469 25513 9472
rect 25547 9500 25559 9503
rect 26329 9503 26387 9509
rect 26329 9500 26341 9503
rect 25547 9472 26341 9500
rect 25547 9469 25559 9472
rect 25501 9463 25559 9469
rect 26329 9469 26341 9472
rect 26375 9469 26387 9503
rect 26329 9463 26387 9469
rect 26513 9503 26571 9509
rect 26513 9469 26525 9503
rect 26559 9500 26571 9503
rect 26602 9500 26608 9512
rect 26559 9472 26608 9500
rect 26559 9469 26571 9472
rect 26513 9463 26571 9469
rect 26602 9460 26608 9472
rect 26660 9460 26666 9512
rect 27246 9460 27252 9512
rect 27304 9460 27310 9512
rect 28169 9503 28227 9509
rect 28169 9469 28181 9503
rect 28215 9500 28227 9503
rect 30558 9500 30564 9512
rect 28215 9472 30564 9500
rect 28215 9469 28227 9472
rect 28169 9463 28227 9469
rect 30558 9460 30564 9472
rect 30616 9460 30622 9512
rect 30668 9500 30696 9531
rect 31386 9528 31392 9580
rect 31444 9528 31450 9580
rect 31481 9503 31539 9509
rect 31481 9500 31493 9503
rect 30668 9472 31493 9500
rect 31481 9469 31493 9472
rect 31527 9469 31539 9503
rect 31481 9463 31539 9469
rect 31665 9503 31723 9509
rect 31665 9469 31677 9503
rect 31711 9500 31723 9503
rect 31754 9500 31760 9512
rect 31711 9472 31760 9500
rect 31711 9469 31723 9472
rect 31665 9463 31723 9469
rect 31754 9460 31760 9472
rect 31812 9460 31818 9512
rect 32232 9500 32260 9608
rect 32582 9596 32588 9648
rect 32640 9596 32646 9648
rect 33318 9596 33324 9648
rect 33376 9596 33382 9648
rect 34790 9596 34796 9648
rect 34848 9636 34854 9648
rect 34977 9639 35035 9645
rect 34977 9636 34989 9639
rect 34848 9608 34989 9636
rect 34848 9596 34854 9608
rect 34977 9605 34989 9608
rect 35023 9605 35035 9639
rect 34977 9599 35035 9605
rect 35066 9596 35072 9648
rect 35124 9636 35130 9648
rect 36372 9636 36400 9676
rect 36832 9674 36860 9676
rect 35124 9608 36400 9636
rect 35124 9596 35130 9608
rect 36446 9596 36452 9648
rect 36504 9596 36510 9648
rect 36832 9646 36952 9674
rect 36998 9664 37004 9716
rect 37056 9704 37062 9716
rect 37826 9704 37832 9716
rect 37056 9676 37832 9704
rect 37056 9664 37062 9676
rect 37826 9664 37832 9676
rect 37884 9664 37890 9716
rect 38654 9664 38660 9716
rect 38712 9704 38718 9716
rect 39209 9707 39267 9713
rect 39209 9704 39221 9707
rect 38712 9676 39221 9704
rect 38712 9664 38718 9676
rect 39209 9673 39221 9676
rect 39255 9673 39267 9707
rect 40126 9704 40132 9716
rect 39209 9667 39267 9673
rect 39316 9676 40132 9704
rect 32306 9528 32312 9580
rect 32364 9528 32370 9580
rect 33870 9528 33876 9580
rect 33928 9568 33934 9580
rect 33928 9540 34376 9568
rect 33928 9528 33934 9540
rect 33778 9500 33784 9512
rect 32232 9472 33784 9500
rect 33778 9460 33784 9472
rect 33836 9460 33842 9512
rect 22060 9404 22600 9432
rect 22060 9392 22066 9404
rect 29270 9392 29276 9444
rect 29328 9432 29334 9444
rect 29822 9432 29828 9444
rect 29328 9404 29828 9432
rect 29328 9392 29334 9404
rect 29822 9392 29828 9404
rect 29880 9392 29886 9444
rect 10008 9336 11284 9364
rect 10008 9324 10014 9336
rect 11698 9324 11704 9376
rect 11756 9324 11762 9376
rect 12805 9367 12863 9373
rect 12805 9333 12817 9367
rect 12851 9364 12863 9367
rect 14550 9364 14556 9376
rect 12851 9336 14556 9364
rect 12851 9333 12863 9336
rect 12805 9327 12863 9333
rect 14550 9324 14556 9336
rect 14608 9324 14614 9376
rect 15013 9367 15071 9373
rect 15013 9333 15025 9367
rect 15059 9364 15071 9367
rect 15286 9364 15292 9376
rect 15059 9336 15292 9364
rect 15059 9333 15071 9336
rect 15013 9327 15071 9333
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 15378 9324 15384 9376
rect 15436 9364 15442 9376
rect 15473 9367 15531 9373
rect 15473 9364 15485 9367
rect 15436 9336 15485 9364
rect 15436 9324 15442 9336
rect 15473 9333 15485 9336
rect 15519 9333 15531 9367
rect 15473 9327 15531 9333
rect 17770 9324 17776 9376
rect 17828 9364 17834 9376
rect 18230 9364 18236 9376
rect 17828 9336 18236 9364
rect 17828 9324 17834 9336
rect 18230 9324 18236 9336
rect 18288 9324 18294 9376
rect 19702 9324 19708 9376
rect 19760 9364 19766 9376
rect 21085 9367 21143 9373
rect 21085 9364 21097 9367
rect 19760 9336 21097 9364
rect 19760 9324 19766 9336
rect 21085 9333 21097 9336
rect 21131 9333 21143 9367
rect 21085 9327 21143 9333
rect 22094 9324 22100 9376
rect 22152 9364 22158 9376
rect 22370 9364 22376 9376
rect 22152 9336 22376 9364
rect 22152 9324 22158 9336
rect 22370 9324 22376 9336
rect 22428 9324 22434 9376
rect 22646 9324 22652 9376
rect 22704 9364 22710 9376
rect 25225 9367 25283 9373
rect 25225 9364 25237 9367
rect 22704 9336 25237 9364
rect 22704 9324 22710 9336
rect 25225 9333 25237 9336
rect 25271 9333 25283 9367
rect 25225 9327 25283 9333
rect 25869 9367 25927 9373
rect 25869 9333 25881 9367
rect 25915 9364 25927 9367
rect 28718 9364 28724 9376
rect 25915 9336 28724 9364
rect 25915 9333 25927 9336
rect 25869 9327 25927 9333
rect 28718 9324 28724 9336
rect 28776 9324 28782 9376
rect 28810 9324 28816 9376
rect 28868 9364 28874 9376
rect 29641 9367 29699 9373
rect 29641 9364 29653 9367
rect 28868 9336 29653 9364
rect 28868 9324 28874 9336
rect 29641 9333 29653 9336
rect 29687 9333 29699 9367
rect 29641 9327 29699 9333
rect 31021 9367 31079 9373
rect 31021 9333 31033 9367
rect 31067 9364 31079 9367
rect 33962 9364 33968 9376
rect 31067 9336 33968 9364
rect 31067 9333 31079 9336
rect 31021 9327 31079 9333
rect 33962 9324 33968 9336
rect 34020 9324 34026 9376
rect 34057 9367 34115 9373
rect 34057 9333 34069 9367
rect 34103 9364 34115 9367
rect 34238 9364 34244 9376
rect 34103 9336 34244 9364
rect 34103 9333 34115 9336
rect 34057 9327 34115 9333
rect 34238 9324 34244 9336
rect 34296 9324 34302 9376
rect 34348 9364 34376 9540
rect 34882 9528 34888 9580
rect 34940 9528 34946 9580
rect 35894 9568 35900 9580
rect 34992 9540 35900 9568
rect 34422 9460 34428 9512
rect 34480 9500 34486 9512
rect 34992 9500 35020 9540
rect 35894 9528 35900 9540
rect 35952 9528 35958 9580
rect 36354 9528 36360 9580
rect 36412 9528 36418 9580
rect 36630 9568 36636 9580
rect 36556 9540 36636 9568
rect 34480 9472 35020 9500
rect 34480 9460 34486 9472
rect 35066 9460 35072 9512
rect 35124 9460 35130 9512
rect 35526 9460 35532 9512
rect 35584 9460 35590 9512
rect 36556 9509 36584 9540
rect 36630 9528 36636 9540
rect 36688 9528 36694 9580
rect 36541 9503 36599 9509
rect 36541 9469 36553 9503
rect 36587 9469 36599 9503
rect 36924 9500 36952 9646
rect 37182 9596 37188 9648
rect 37240 9636 37246 9648
rect 39114 9636 39120 9648
rect 37240 9608 39120 9636
rect 37240 9596 37246 9608
rect 39114 9596 39120 9608
rect 39172 9596 39178 9648
rect 37274 9528 37280 9580
rect 37332 9568 37338 9580
rect 37461 9571 37519 9577
rect 37461 9568 37473 9571
rect 37332 9540 37473 9568
rect 37332 9528 37338 9540
rect 37461 9537 37473 9540
rect 37507 9537 37519 9571
rect 37461 9531 37519 9537
rect 37826 9528 37832 9580
rect 37884 9568 37890 9580
rect 37884 9540 38516 9568
rect 37884 9528 37890 9540
rect 38488 9500 38516 9540
rect 38562 9528 38568 9580
rect 38620 9528 38626 9580
rect 38930 9528 38936 9580
rect 38988 9568 38994 9580
rect 39316 9568 39344 9676
rect 40126 9664 40132 9676
rect 40184 9664 40190 9716
rect 39850 9596 39856 9648
rect 39908 9636 39914 9648
rect 39908 9608 44220 9636
rect 39908 9596 39914 9608
rect 38988 9540 39344 9568
rect 38988 9528 38994 9540
rect 39758 9528 39764 9580
rect 39816 9528 39822 9580
rect 40586 9568 40592 9580
rect 39868 9540 40592 9568
rect 36924 9472 38240 9500
rect 38488 9472 39620 9500
rect 36541 9463 36599 9469
rect 34517 9435 34575 9441
rect 34517 9401 34529 9435
rect 34563 9432 34575 9435
rect 35710 9432 35716 9444
rect 34563 9404 35716 9432
rect 34563 9401 34575 9404
rect 34517 9395 34575 9401
rect 35710 9392 35716 9404
rect 35768 9392 35774 9444
rect 37550 9432 37556 9444
rect 35820 9404 37556 9432
rect 35820 9364 35848 9404
rect 37550 9392 37556 9404
rect 37608 9392 37614 9444
rect 34348 9336 35848 9364
rect 35986 9324 35992 9376
rect 36044 9324 36050 9376
rect 36998 9324 37004 9376
rect 37056 9324 37062 9376
rect 37274 9324 37280 9376
rect 37332 9364 37338 9376
rect 38105 9367 38163 9373
rect 38105 9364 38117 9367
rect 37332 9336 38117 9364
rect 37332 9324 37338 9336
rect 38105 9333 38117 9336
rect 38151 9333 38163 9367
rect 38212 9364 38240 9472
rect 38470 9392 38476 9444
rect 38528 9432 38534 9444
rect 38654 9432 38660 9444
rect 38528 9404 38660 9432
rect 38528 9392 38534 9404
rect 38654 9392 38660 9404
rect 38712 9392 38718 9444
rect 39592 9432 39620 9472
rect 39868 9432 39896 9540
rect 40586 9528 40592 9540
rect 40644 9528 40650 9580
rect 40696 9540 41368 9568
rect 39942 9460 39948 9512
rect 40000 9500 40006 9512
rect 40696 9500 40724 9540
rect 40000 9472 40724 9500
rect 40000 9460 40006 9472
rect 41230 9460 41236 9512
rect 41288 9460 41294 9512
rect 41340 9500 41368 9540
rect 41414 9528 41420 9580
rect 41472 9568 41478 9580
rect 41509 9571 41567 9577
rect 41509 9568 41521 9571
rect 41472 9540 41521 9568
rect 41472 9528 41478 9540
rect 41509 9537 41521 9540
rect 41555 9537 41567 9571
rect 41509 9531 41567 9537
rect 42886 9528 42892 9580
rect 42944 9528 42950 9580
rect 43254 9528 43260 9580
rect 43312 9568 43318 9580
rect 43714 9568 43720 9580
rect 43312 9540 43720 9568
rect 43312 9528 43318 9540
rect 43714 9528 43720 9540
rect 43772 9528 43778 9580
rect 44192 9577 44220 9608
rect 44542 9596 44548 9648
rect 44600 9636 44606 9648
rect 46293 9639 46351 9645
rect 46293 9636 46305 9639
rect 44600 9608 46305 9636
rect 44600 9596 44606 9608
rect 46293 9605 46305 9608
rect 46339 9605 46351 9639
rect 46293 9599 46351 9605
rect 47210 9596 47216 9648
rect 47268 9636 47274 9648
rect 47305 9639 47363 9645
rect 47305 9636 47317 9639
rect 47268 9608 47317 9636
rect 47268 9596 47274 9608
rect 47305 9605 47317 9608
rect 47351 9605 47363 9639
rect 47305 9599 47363 9605
rect 47673 9639 47731 9645
rect 47673 9605 47685 9639
rect 47719 9636 47731 9639
rect 47854 9636 47860 9648
rect 47719 9608 47860 9636
rect 47719 9605 47731 9608
rect 47673 9599 47731 9605
rect 47854 9596 47860 9608
rect 47912 9596 47918 9648
rect 49145 9639 49203 9645
rect 49145 9605 49157 9639
rect 49191 9636 49203 9639
rect 49418 9636 49424 9648
rect 49191 9608 49424 9636
rect 49191 9605 49203 9608
rect 49145 9599 49203 9605
rect 49418 9596 49424 9608
rect 49476 9596 49482 9648
rect 44177 9571 44235 9577
rect 44177 9537 44189 9571
rect 44223 9537 44235 9571
rect 44177 9531 44235 9537
rect 45094 9528 45100 9580
rect 45152 9568 45158 9580
rect 45465 9571 45523 9577
rect 45465 9568 45477 9571
rect 45152 9540 45477 9568
rect 45152 9528 45158 9540
rect 45465 9537 45477 9540
rect 45511 9537 45523 9571
rect 45465 9531 45523 9537
rect 45738 9528 45744 9580
rect 45796 9568 45802 9580
rect 46474 9568 46480 9580
rect 45796 9540 46480 9568
rect 45796 9528 45802 9540
rect 46474 9528 46480 9540
rect 46532 9568 46538 9580
rect 46753 9571 46811 9577
rect 46753 9568 46765 9571
rect 46532 9540 46765 9568
rect 46532 9528 46538 9540
rect 46753 9537 46765 9540
rect 46799 9537 46811 9571
rect 47949 9571 48007 9577
rect 47949 9568 47961 9571
rect 46753 9531 46811 9537
rect 46860 9540 47961 9568
rect 42518 9500 42524 9512
rect 41340 9472 42524 9500
rect 42518 9460 42524 9472
rect 42576 9460 42582 9512
rect 42610 9460 42616 9512
rect 42668 9460 42674 9512
rect 42702 9460 42708 9512
rect 42760 9500 42766 9512
rect 42760 9472 43852 9500
rect 42760 9460 42766 9472
rect 39592 9404 39896 9432
rect 43824 9432 43852 9472
rect 43898 9460 43904 9512
rect 43956 9460 43962 9512
rect 45186 9460 45192 9512
rect 45244 9460 45250 9512
rect 46860 9432 46888 9540
rect 47949 9537 47961 9540
rect 47995 9537 48007 9571
rect 47949 9531 48007 9537
rect 43824 9404 46888 9432
rect 46937 9435 46995 9441
rect 46937 9401 46949 9435
rect 46983 9432 46995 9435
rect 47486 9432 47492 9444
rect 46983 9404 47492 9432
rect 46983 9401 46995 9404
rect 46937 9395 46995 9401
rect 47486 9392 47492 9404
rect 47544 9392 47550 9444
rect 38930 9364 38936 9376
rect 38212 9336 38936 9364
rect 38105 9327 38163 9333
rect 38930 9324 38936 9336
rect 38988 9324 38994 9376
rect 39850 9324 39856 9376
rect 39908 9324 39914 9376
rect 40681 9367 40739 9373
rect 40681 9333 40693 9367
rect 40727 9364 40739 9367
rect 47118 9364 47124 9376
rect 40727 9336 47124 9364
rect 40727 9333 40739 9336
rect 40681 9327 40739 9333
rect 47118 9324 47124 9336
rect 47176 9324 47182 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 3602 9120 3608 9172
rect 3660 9120 3666 9172
rect 8478 9160 8484 9172
rect 5276 9132 8484 9160
rect 2501 9095 2559 9101
rect 2501 9061 2513 9095
rect 2547 9092 2559 9095
rect 5276 9092 5304 9132
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 10318 9120 10324 9172
rect 10376 9120 10382 9172
rect 10594 9120 10600 9172
rect 10652 9160 10658 9172
rect 11425 9163 11483 9169
rect 11425 9160 11437 9163
rect 10652 9132 11437 9160
rect 10652 9120 10658 9132
rect 11425 9129 11437 9132
rect 11471 9129 11483 9163
rect 11425 9123 11483 9129
rect 12250 9120 12256 9172
rect 12308 9160 12314 9172
rect 12989 9163 13047 9169
rect 12989 9160 13001 9163
rect 12308 9132 13001 9160
rect 12308 9120 12314 9132
rect 12989 9129 13001 9132
rect 13035 9129 13047 9163
rect 12989 9123 13047 9129
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 15286 9160 15292 9172
rect 13780 9132 15292 9160
rect 13780 9120 13786 9132
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 15470 9120 15476 9172
rect 15528 9160 15534 9172
rect 15528 9132 16344 9160
rect 15528 9120 15534 9132
rect 8018 9092 8024 9104
rect 2547 9064 5304 9092
rect 5368 9064 8024 9092
rect 2547 9061 2559 9064
rect 2501 9055 2559 9061
rect 2222 8984 2228 9036
rect 2280 9024 2286 9036
rect 5368 9024 5396 9064
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 16022 9092 16028 9104
rect 8496 9064 16028 9092
rect 2280 8996 5396 9024
rect 6181 9027 6239 9033
rect 2280 8984 2286 8996
rect 6181 8993 6193 9027
rect 6227 9024 6239 9027
rect 7282 9024 7288 9036
rect 6227 8996 7288 9024
rect 6227 8993 6239 8996
rect 6181 8987 6239 8993
rect 7282 8984 7288 8996
rect 7340 8984 7346 9036
rect 7742 8984 7748 9036
rect 7800 8984 7806 9036
rect 1302 8916 1308 8968
rect 1360 8956 1366 8968
rect 1581 8959 1639 8965
rect 1581 8956 1593 8959
rect 1360 8928 1593 8956
rect 1360 8916 1366 8928
rect 1581 8925 1593 8928
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8925 2375 8959
rect 2317 8919 2375 8925
rect 3237 8959 3295 8965
rect 3237 8925 3249 8959
rect 3283 8956 3295 8959
rect 3418 8956 3424 8968
rect 3283 8928 3424 8956
rect 3283 8925 3295 8928
rect 3237 8919 3295 8925
rect 1210 8848 1216 8900
rect 1268 8888 1274 8900
rect 2332 8888 2360 8919
rect 3418 8916 3424 8928
rect 3476 8956 3482 8968
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 3476 8928 3801 8956
rect 3476 8916 3482 8928
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 1268 8860 2360 8888
rect 5920 8888 5948 8919
rect 7650 8916 7656 8968
rect 7708 8956 7714 8968
rect 8021 8959 8079 8965
rect 8021 8956 8033 8959
rect 7708 8928 8033 8956
rect 7708 8916 7714 8928
rect 8021 8925 8033 8928
rect 8067 8925 8079 8959
rect 8021 8919 8079 8925
rect 8386 8888 8392 8900
rect 5920 8860 8392 8888
rect 1268 8848 1274 8860
rect 8386 8848 8392 8860
rect 8444 8848 8450 8900
rect 1762 8780 1768 8832
rect 1820 8780 1826 8832
rect 3053 8823 3111 8829
rect 3053 8789 3065 8823
rect 3099 8820 3111 8823
rect 4338 8820 4344 8832
rect 3099 8792 4344 8820
rect 3099 8789 3111 8792
rect 3053 8783 3111 8789
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 5350 8780 5356 8832
rect 5408 8820 5414 8832
rect 5537 8823 5595 8829
rect 5537 8820 5549 8823
rect 5408 8792 5549 8820
rect 5408 8780 5414 8792
rect 5537 8789 5549 8792
rect 5583 8820 5595 8823
rect 8496 8820 8524 9064
rect 16022 9052 16028 9064
rect 16080 9052 16086 9104
rect 8570 8984 8576 9036
rect 8628 9024 8634 9036
rect 8628 8996 10824 9024
rect 8628 8984 8634 8996
rect 9674 8916 9680 8968
rect 9732 8916 9738 8968
rect 10796 8965 10824 8996
rect 13446 8984 13452 9036
rect 13504 8984 13510 9036
rect 13630 8984 13636 9036
rect 13688 8984 13694 9036
rect 14918 8984 14924 9036
rect 14976 9024 14982 9036
rect 15473 9027 15531 9033
rect 15473 9024 15485 9027
rect 14976 8996 15485 9024
rect 14976 8984 14982 8996
rect 15473 8993 15485 8996
rect 15519 8993 15531 9027
rect 15473 8987 15531 8993
rect 15562 8984 15568 9036
rect 15620 8984 15626 9036
rect 16206 8984 16212 9036
rect 16264 8984 16270 9036
rect 16316 9024 16344 9132
rect 17678 9120 17684 9172
rect 17736 9160 17742 9172
rect 18233 9163 18291 9169
rect 18233 9160 18245 9163
rect 17736 9132 18245 9160
rect 17736 9120 17742 9132
rect 18233 9129 18245 9132
rect 18279 9129 18291 9163
rect 18233 9123 18291 9129
rect 19337 9163 19395 9169
rect 19337 9129 19349 9163
rect 19383 9160 19395 9163
rect 19426 9160 19432 9172
rect 19383 9132 19432 9160
rect 19383 9129 19395 9132
rect 19337 9123 19395 9129
rect 19426 9120 19432 9132
rect 19484 9120 19490 9172
rect 20806 9160 20812 9172
rect 20088 9132 20812 9160
rect 18690 9052 18696 9104
rect 18748 9052 18754 9104
rect 20088 9092 20116 9132
rect 20806 9120 20812 9132
rect 20864 9120 20870 9172
rect 22278 9120 22284 9172
rect 22336 9160 22342 9172
rect 23937 9163 23995 9169
rect 23937 9160 23949 9163
rect 22336 9132 23949 9160
rect 22336 9120 22342 9132
rect 23937 9129 23949 9132
rect 23983 9129 23995 9163
rect 23937 9123 23995 9129
rect 25130 9120 25136 9172
rect 25188 9160 25194 9172
rect 27709 9163 27767 9169
rect 27709 9160 27721 9163
rect 25188 9132 27721 9160
rect 25188 9120 25194 9132
rect 27709 9129 27721 9132
rect 27755 9129 27767 9163
rect 27709 9123 27767 9129
rect 28261 9163 28319 9169
rect 28261 9129 28273 9163
rect 28307 9160 28319 9163
rect 34882 9160 34888 9172
rect 28307 9132 34888 9160
rect 28307 9129 28319 9132
rect 28261 9123 28319 9129
rect 34882 9120 34888 9132
rect 34940 9120 34946 9172
rect 36538 9160 36544 9172
rect 35452 9132 36544 9160
rect 18892 9064 20116 9092
rect 16316 8996 18000 9024
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8925 10839 8959
rect 10781 8919 10839 8925
rect 11885 8959 11943 8965
rect 11885 8925 11897 8959
rect 11931 8956 11943 8959
rect 13262 8956 13268 8968
rect 11931 8928 13268 8956
rect 11931 8925 11943 8928
rect 11885 8919 11943 8925
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 14369 8959 14427 8965
rect 14369 8925 14381 8959
rect 14415 8956 14427 8959
rect 15102 8956 15108 8968
rect 14415 8928 15108 8956
rect 14415 8925 14427 8928
rect 14369 8919 14427 8925
rect 15102 8916 15108 8928
rect 15160 8916 15166 8968
rect 15378 8916 15384 8968
rect 15436 8916 15442 8968
rect 8846 8848 8852 8900
rect 8904 8888 8910 8900
rect 11698 8888 11704 8900
rect 8904 8860 11704 8888
rect 8904 8848 8910 8860
rect 11698 8848 11704 8860
rect 11756 8888 11762 8900
rect 12529 8891 12587 8897
rect 11756 8860 12434 8888
rect 11756 8848 11762 8860
rect 5583 8792 8524 8820
rect 5583 8789 5595 8792
rect 5537 8783 5595 8789
rect 8570 8780 8576 8832
rect 8628 8820 8634 8832
rect 11606 8820 11612 8832
rect 8628 8792 11612 8820
rect 8628 8780 8634 8792
rect 11606 8780 11612 8792
rect 11664 8780 11670 8832
rect 12406 8820 12434 8860
rect 12529 8857 12541 8891
rect 12575 8888 12587 8891
rect 13630 8888 13636 8900
rect 12575 8860 13636 8888
rect 12575 8857 12587 8860
rect 12529 8851 12587 8857
rect 13630 8848 13636 8860
rect 13688 8848 13694 8900
rect 15194 8848 15200 8900
rect 15252 8888 15258 8900
rect 16485 8891 16543 8897
rect 16485 8888 16497 8891
rect 15252 8860 16497 8888
rect 15252 8848 15258 8860
rect 16485 8857 16497 8860
rect 16531 8857 16543 8891
rect 16485 8851 16543 8857
rect 16942 8848 16948 8900
rect 17000 8848 17006 8900
rect 13170 8820 13176 8832
rect 12406 8792 13176 8820
rect 13170 8780 13176 8792
rect 13228 8820 13234 8832
rect 13357 8823 13415 8829
rect 13357 8820 13369 8823
rect 13228 8792 13369 8820
rect 13228 8780 13234 8792
rect 13357 8789 13369 8792
rect 13403 8789 13415 8823
rect 13357 8783 13415 8789
rect 13446 8780 13452 8832
rect 13504 8820 13510 8832
rect 14918 8820 14924 8832
rect 13504 8792 14924 8820
rect 13504 8780 13510 8792
rect 14918 8780 14924 8792
rect 14976 8780 14982 8832
rect 15010 8780 15016 8832
rect 15068 8780 15074 8832
rect 17972 8829 18000 8996
rect 18506 8916 18512 8968
rect 18564 8956 18570 8968
rect 18690 8956 18696 8968
rect 18564 8928 18696 8956
rect 18564 8916 18570 8928
rect 18690 8916 18696 8928
rect 18748 8916 18754 8968
rect 18892 8965 18920 9064
rect 25958 9052 25964 9104
rect 26016 9052 26022 9104
rect 28534 9052 28540 9104
rect 28592 9092 28598 9104
rect 28810 9092 28816 9104
rect 28592 9064 28816 9092
rect 28592 9052 28598 9064
rect 28810 9052 28816 9064
rect 28868 9052 28874 9104
rect 31294 9052 31300 9104
rect 31352 9092 31358 9104
rect 31481 9095 31539 9101
rect 31481 9092 31493 9095
rect 31352 9064 31493 9092
rect 31352 9052 31358 9064
rect 31481 9061 31493 9064
rect 31527 9061 31539 9095
rect 31481 9055 31539 9061
rect 31726 9064 32076 9092
rect 19242 8984 19248 9036
rect 19300 9024 19306 9036
rect 19521 9027 19579 9033
rect 19521 9024 19533 9027
rect 19300 8996 19533 9024
rect 19300 8984 19306 8996
rect 19521 8993 19533 8996
rect 19567 9024 19579 9027
rect 19981 9027 20039 9033
rect 19981 9024 19993 9027
rect 19567 8996 19993 9024
rect 19567 8993 19579 8996
rect 19521 8987 19579 8993
rect 19981 8993 19993 8996
rect 20027 9024 20039 9027
rect 21818 9024 21824 9036
rect 20027 8996 21824 9024
rect 20027 8993 20039 8996
rect 19981 8987 20039 8993
rect 21818 8984 21824 8996
rect 21876 9024 21882 9036
rect 22189 9027 22247 9033
rect 22189 9024 22201 9027
rect 21876 8996 22201 9024
rect 21876 8984 21882 8996
rect 22189 8993 22201 8996
rect 22235 9024 22247 9027
rect 23474 9024 23480 9036
rect 22235 8996 23480 9024
rect 22235 8993 22247 8996
rect 22189 8987 22247 8993
rect 23474 8984 23480 8996
rect 23532 8984 23538 9036
rect 25593 9027 25651 9033
rect 25593 8993 25605 9027
rect 25639 9024 25651 9027
rect 25976 9024 26004 9052
rect 27614 9024 27620 9036
rect 25639 8996 27620 9024
rect 25639 8993 25651 8996
rect 25593 8987 25651 8993
rect 27614 8984 27620 8996
rect 27672 8984 27678 9036
rect 28718 8984 28724 9036
rect 28776 8984 28782 9036
rect 28902 8984 28908 9036
rect 28960 8984 28966 9036
rect 30009 9027 30067 9033
rect 30009 8993 30021 9027
rect 30055 9024 30067 9027
rect 30742 9024 30748 9036
rect 30055 8996 30748 9024
rect 30055 8993 30067 8996
rect 30009 8987 30067 8993
rect 30742 8984 30748 8996
rect 30800 8984 30806 9036
rect 18877 8959 18935 8965
rect 18877 8925 18889 8959
rect 18923 8925 18935 8959
rect 18877 8919 18935 8925
rect 19702 8916 19708 8968
rect 19760 8916 19766 8968
rect 24486 8916 24492 8968
rect 24544 8956 24550 8968
rect 24581 8959 24639 8965
rect 24581 8956 24593 8959
rect 24544 8928 24593 8956
rect 24544 8916 24550 8928
rect 24581 8925 24593 8928
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 25038 8916 25044 8968
rect 25096 8956 25102 8968
rect 25961 8959 26019 8965
rect 25961 8956 25973 8959
rect 25096 8928 25973 8956
rect 25096 8916 25102 8928
rect 25961 8925 25973 8928
rect 26007 8925 26019 8959
rect 25961 8919 26019 8925
rect 27062 8916 27068 8968
rect 27120 8916 27126 8968
rect 28442 8916 28448 8968
rect 28500 8956 28506 8968
rect 29730 8956 29736 8968
rect 28500 8928 29736 8956
rect 28500 8916 28506 8928
rect 29730 8916 29736 8928
rect 29788 8916 29794 8968
rect 31478 8956 31484 8968
rect 31142 8928 31484 8956
rect 31478 8916 31484 8928
rect 31536 8956 31542 8968
rect 31726 8956 31754 9064
rect 31938 8984 31944 9036
rect 31996 8984 32002 9036
rect 32048 9024 32076 9064
rect 33686 9052 33692 9104
rect 33744 9052 33750 9104
rect 34698 9052 34704 9104
rect 34756 9092 34762 9104
rect 35250 9092 35256 9104
rect 34756 9064 35256 9092
rect 34756 9052 34762 9064
rect 35250 9052 35256 9064
rect 35308 9052 35314 9104
rect 32048 8996 33364 9024
rect 33336 8968 33364 8996
rect 34146 8984 34152 9036
rect 34204 8984 34210 9036
rect 35158 8984 35164 9036
rect 35216 9024 35222 9036
rect 35452 9033 35480 9132
rect 36538 9120 36544 9132
rect 36596 9160 36602 9172
rect 37001 9163 37059 9169
rect 37001 9160 37013 9163
rect 36596 9132 37013 9160
rect 36596 9120 36602 9132
rect 37001 9129 37013 9132
rect 37047 9129 37059 9163
rect 37001 9123 37059 9129
rect 37182 9120 37188 9172
rect 37240 9160 37246 9172
rect 38562 9160 38568 9172
rect 37240 9132 38568 9160
rect 37240 9120 37246 9132
rect 38562 9120 38568 9132
rect 38620 9120 38626 9172
rect 38749 9163 38807 9169
rect 38749 9129 38761 9163
rect 38795 9160 38807 9163
rect 38838 9160 38844 9172
rect 38795 9132 38844 9160
rect 38795 9129 38807 9132
rect 38749 9123 38807 9129
rect 38838 9120 38844 9132
rect 38896 9160 38902 9172
rect 39758 9160 39764 9172
rect 38896 9132 39764 9160
rect 38896 9120 38902 9132
rect 39758 9120 39764 9132
rect 39816 9120 39822 9172
rect 43806 9120 43812 9172
rect 43864 9120 43870 9172
rect 45002 9120 45008 9172
rect 45060 9160 45066 9172
rect 45189 9163 45247 9169
rect 45189 9160 45201 9163
rect 45060 9132 45201 9160
rect 45060 9120 45066 9132
rect 45189 9129 45201 9132
rect 45235 9129 45247 9163
rect 45189 9123 45247 9129
rect 45922 9120 45928 9172
rect 45980 9160 45986 9172
rect 46661 9163 46719 9169
rect 46661 9160 46673 9163
rect 45980 9132 46673 9160
rect 45980 9120 45986 9132
rect 46661 9129 46673 9132
rect 46707 9129 46719 9163
rect 46661 9123 46719 9129
rect 47397 9163 47455 9169
rect 47397 9129 47409 9163
rect 47443 9160 47455 9163
rect 47578 9160 47584 9172
rect 47443 9132 47584 9160
rect 47443 9129 47455 9132
rect 47397 9123 47455 9129
rect 47578 9120 47584 9132
rect 47636 9120 47642 9172
rect 35618 9052 35624 9104
rect 35676 9092 35682 9104
rect 36630 9092 36636 9104
rect 35676 9064 36636 9092
rect 35676 9052 35682 9064
rect 36630 9052 36636 9064
rect 36688 9052 36694 9104
rect 37366 9052 37372 9104
rect 37424 9092 37430 9104
rect 38378 9092 38384 9104
rect 37424 9064 38384 9092
rect 37424 9052 37430 9064
rect 38378 9052 38384 9064
rect 38436 9052 38442 9104
rect 38930 9052 38936 9104
rect 38988 9092 38994 9104
rect 39577 9095 39635 9101
rect 39577 9092 39589 9095
rect 38988 9064 39589 9092
rect 38988 9052 38994 9064
rect 39577 9061 39589 9064
rect 39623 9061 39635 9095
rect 39577 9055 39635 9061
rect 39850 9052 39856 9104
rect 39908 9092 39914 9104
rect 39908 9064 47992 9092
rect 39908 9052 39914 9064
rect 35345 9027 35403 9033
rect 35345 9024 35357 9027
rect 35216 8996 35357 9024
rect 35216 8984 35222 8996
rect 35345 8993 35357 8996
rect 35391 8993 35403 9027
rect 35345 8987 35403 8993
rect 35437 9027 35495 9033
rect 35437 8993 35449 9027
rect 35483 8993 35495 9027
rect 35437 8987 35495 8993
rect 35526 8984 35532 9036
rect 35584 9024 35590 9036
rect 38105 9027 38163 9033
rect 38105 9024 38117 9027
rect 35584 8996 38117 9024
rect 35584 8984 35590 8996
rect 38105 8993 38117 8996
rect 38151 8993 38163 9027
rect 38105 8987 38163 8993
rect 39114 8984 39120 9036
rect 39172 9024 39178 9036
rect 40773 9027 40831 9033
rect 40773 9024 40785 9027
rect 39172 8996 40785 9024
rect 39172 8984 39178 8996
rect 40773 8993 40785 8996
rect 40819 8993 40831 9027
rect 40773 8987 40831 8993
rect 40862 8984 40868 9036
rect 40920 9024 40926 9036
rect 42337 9027 42395 9033
rect 42337 9024 42349 9027
rect 40920 8996 42349 9024
rect 40920 8984 40926 8996
rect 42337 8993 42349 8996
rect 42383 8993 42395 9027
rect 42337 8987 42395 8993
rect 42426 8984 42432 9036
rect 42484 9024 42490 9036
rect 42484 8996 44496 9024
rect 42484 8984 42490 8996
rect 31536 8928 31754 8956
rect 31536 8916 31542 8928
rect 33318 8916 33324 8968
rect 33376 8916 33382 8968
rect 33502 8916 33508 8968
rect 33560 8956 33566 8968
rect 35253 8959 35311 8965
rect 35253 8956 35265 8959
rect 33560 8928 35265 8956
rect 33560 8916 33566 8928
rect 35253 8925 35265 8928
rect 35299 8925 35311 8959
rect 35253 8919 35311 8925
rect 35618 8916 35624 8968
rect 35676 8956 35682 8968
rect 35802 8956 35808 8968
rect 35676 8928 35808 8956
rect 35676 8916 35682 8928
rect 35802 8916 35808 8928
rect 35860 8916 35866 8968
rect 36078 8916 36084 8968
rect 36136 8916 36142 8968
rect 36446 8916 36452 8968
rect 36504 8956 36510 8968
rect 36725 8959 36783 8965
rect 36725 8956 36737 8959
rect 36504 8928 36737 8956
rect 36504 8916 36510 8928
rect 36725 8925 36737 8928
rect 36771 8925 36783 8959
rect 36725 8919 36783 8925
rect 37461 8959 37519 8965
rect 37461 8925 37473 8959
rect 37507 8925 37519 8959
rect 37461 8919 37519 8925
rect 18598 8848 18604 8900
rect 18656 8888 18662 8900
rect 20257 8891 20315 8897
rect 18656 8860 19748 8888
rect 18656 8848 18662 8860
rect 17957 8823 18015 8829
rect 17957 8789 17969 8823
rect 18003 8820 18015 8823
rect 18506 8820 18512 8832
rect 18003 8792 18512 8820
rect 18003 8789 18015 8792
rect 17957 8783 18015 8789
rect 18506 8780 18512 8792
rect 18564 8780 18570 8832
rect 19720 8820 19748 8860
rect 20257 8857 20269 8891
rect 20303 8888 20315 8891
rect 20530 8888 20536 8900
rect 20303 8860 20536 8888
rect 20303 8857 20315 8860
rect 20257 8851 20315 8857
rect 20530 8848 20536 8860
rect 20588 8848 20594 8900
rect 20714 8848 20720 8900
rect 20772 8848 20778 8900
rect 22465 8891 22523 8897
rect 22465 8857 22477 8891
rect 22511 8888 22523 8891
rect 22511 8860 22876 8888
rect 22511 8857 22523 8860
rect 22465 8851 22523 8857
rect 21729 8823 21787 8829
rect 21729 8820 21741 8823
rect 19720 8792 21741 8820
rect 21729 8789 21741 8792
rect 21775 8789 21787 8823
rect 22848 8820 22876 8860
rect 22922 8848 22928 8900
rect 22980 8848 22986 8900
rect 27246 8848 27252 8900
rect 27304 8888 27310 8900
rect 28629 8891 28687 8897
rect 28629 8888 28641 8891
rect 27304 8860 28641 8888
rect 27304 8848 27310 8860
rect 28629 8857 28641 8860
rect 28675 8857 28687 8891
rect 28629 8851 28687 8857
rect 32214 8848 32220 8900
rect 32272 8848 32278 8900
rect 34238 8848 34244 8900
rect 34296 8888 34302 8900
rect 37476 8888 37504 8919
rect 37550 8916 37556 8968
rect 37608 8956 37614 8968
rect 41049 8959 41107 8965
rect 41049 8956 41061 8959
rect 37608 8928 41061 8956
rect 37608 8916 37614 8928
rect 41049 8925 41061 8928
rect 41095 8925 41107 8959
rect 41049 8919 41107 8925
rect 41966 8916 41972 8968
rect 42024 8956 42030 8968
rect 42061 8959 42119 8965
rect 42061 8956 42073 8959
rect 42024 8928 42073 8956
rect 42024 8916 42030 8928
rect 42061 8925 42073 8928
rect 42107 8925 42119 8959
rect 42061 8919 42119 8925
rect 43530 8916 43536 8968
rect 43588 8916 43594 8968
rect 44082 8916 44088 8968
rect 44140 8956 44146 8968
rect 44361 8959 44419 8965
rect 44361 8956 44373 8959
rect 44140 8928 44373 8956
rect 44140 8916 44146 8928
rect 44361 8925 44373 8928
rect 44407 8925 44419 8959
rect 44468 8956 44496 8996
rect 44542 8984 44548 9036
rect 44600 9024 44606 9036
rect 45557 9027 45615 9033
rect 45557 9024 45569 9027
rect 44600 8996 45569 9024
rect 44600 8984 44606 8996
rect 45557 8993 45569 8996
rect 45603 8993 45615 9027
rect 45557 8987 45615 8993
rect 45833 8959 45891 8965
rect 45833 8956 45845 8959
rect 44468 8928 45845 8956
rect 44361 8919 44419 8925
rect 45833 8925 45845 8928
rect 45879 8925 45891 8959
rect 45833 8919 45891 8925
rect 46750 8916 46756 8968
rect 46808 8956 46814 8968
rect 47964 8965 47992 9064
rect 49145 9027 49203 9033
rect 49145 8993 49157 9027
rect 49191 9024 49203 9027
rect 49234 9024 49240 9036
rect 49191 8996 49240 9024
rect 49191 8993 49203 8996
rect 49145 8987 49203 8993
rect 49234 8984 49240 8996
rect 49292 8984 49298 9036
rect 47213 8959 47271 8965
rect 47213 8956 47225 8959
rect 46808 8928 47225 8956
rect 46808 8916 46814 8928
rect 47213 8925 47225 8928
rect 47259 8925 47271 8959
rect 47213 8919 47271 8925
rect 47949 8959 48007 8965
rect 47949 8925 47961 8959
rect 47995 8925 48007 8959
rect 47949 8919 48007 8925
rect 34296 8860 37504 8888
rect 37568 8860 38608 8888
rect 34296 8848 34302 8860
rect 24210 8820 24216 8832
rect 22848 8792 24216 8820
rect 21729 8783 21787 8789
rect 24210 8780 24216 8792
rect 24268 8780 24274 8832
rect 24486 8780 24492 8832
rect 24544 8820 24550 8832
rect 25225 8823 25283 8829
rect 25225 8820 25237 8823
rect 24544 8792 25237 8820
rect 24544 8780 24550 8792
rect 25225 8789 25237 8792
rect 25271 8789 25283 8823
rect 25225 8783 25283 8789
rect 25958 8780 25964 8832
rect 26016 8820 26022 8832
rect 26605 8823 26663 8829
rect 26605 8820 26617 8823
rect 26016 8792 26617 8820
rect 26016 8780 26022 8792
rect 26605 8789 26617 8792
rect 26651 8789 26663 8823
rect 26605 8783 26663 8789
rect 34885 8823 34943 8829
rect 34885 8789 34897 8823
rect 34931 8820 34943 8823
rect 34974 8820 34980 8832
rect 34931 8792 34980 8820
rect 34931 8789 34943 8792
rect 34885 8783 34943 8789
rect 34974 8780 34980 8792
rect 35032 8780 35038 8832
rect 35250 8780 35256 8832
rect 35308 8820 35314 8832
rect 37568 8820 37596 8860
rect 35308 8792 37596 8820
rect 35308 8780 35314 8792
rect 37642 8780 37648 8832
rect 37700 8820 37706 8832
rect 38470 8820 38476 8832
rect 37700 8792 38476 8820
rect 37700 8780 37706 8792
rect 38470 8780 38476 8792
rect 38528 8780 38534 8832
rect 38580 8820 38608 8860
rect 38930 8848 38936 8900
rect 38988 8888 38994 8900
rect 39117 8891 39175 8897
rect 39117 8888 39129 8891
rect 38988 8860 39129 8888
rect 38988 8848 38994 8860
rect 39117 8857 39129 8860
rect 39163 8857 39175 8891
rect 39117 8851 39175 8857
rect 39298 8848 39304 8900
rect 39356 8848 39362 8900
rect 39574 8848 39580 8900
rect 39632 8888 39638 8900
rect 40129 8891 40187 8897
rect 40129 8888 40141 8891
rect 39632 8860 40141 8888
rect 39632 8848 39638 8860
rect 40129 8857 40141 8860
rect 40175 8857 40187 8891
rect 40129 8851 40187 8857
rect 40310 8848 40316 8900
rect 40368 8848 40374 8900
rect 44545 8891 44603 8897
rect 44545 8857 44557 8891
rect 44591 8888 44603 8891
rect 47854 8888 47860 8900
rect 44591 8860 47860 8888
rect 44591 8857 44603 8860
rect 44545 8851 44603 8857
rect 47854 8848 47860 8860
rect 47912 8848 47918 8900
rect 41966 8820 41972 8832
rect 38580 8792 41972 8820
rect 41966 8780 41972 8792
rect 42024 8780 42030 8832
rect 43349 8823 43407 8829
rect 43349 8789 43361 8823
rect 43395 8820 43407 8823
rect 43714 8820 43720 8832
rect 43395 8792 43720 8820
rect 43395 8789 43407 8792
rect 43349 8783 43407 8789
rect 43714 8780 43720 8792
rect 43772 8780 43778 8832
rect 43898 8780 43904 8832
rect 43956 8820 43962 8832
rect 45005 8823 45063 8829
rect 45005 8820 45017 8823
rect 43956 8792 45017 8820
rect 43956 8780 43962 8792
rect 45005 8789 45017 8792
rect 45051 8789 45063 8823
rect 45005 8783 45063 8789
rect 46937 8823 46995 8829
rect 46937 8789 46949 8823
rect 46983 8820 46995 8823
rect 48314 8820 48320 8832
rect 46983 8792 48320 8820
rect 46983 8789 46995 8792
rect 46937 8783 46995 8789
rect 48314 8780 48320 8792
rect 48372 8780 48378 8832
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 1302 8576 1308 8628
rect 1360 8616 1366 8628
rect 3237 8619 3295 8625
rect 3237 8616 3249 8619
rect 1360 8588 3249 8616
rect 1360 8576 1366 8588
rect 3237 8585 3249 8588
rect 3283 8585 3295 8619
rect 3237 8579 3295 8585
rect 5626 8576 5632 8628
rect 5684 8616 5690 8628
rect 7469 8619 7527 8625
rect 7469 8616 7481 8619
rect 5684 8588 7481 8616
rect 5684 8576 5690 8588
rect 7469 8585 7481 8588
rect 7515 8585 7527 8619
rect 7469 8579 7527 8585
rect 7558 8576 7564 8628
rect 7616 8616 7622 8628
rect 12989 8619 13047 8625
rect 7616 8588 10548 8616
rect 7616 8576 7622 8588
rect 1210 8508 1216 8560
rect 1268 8548 1274 8560
rect 3421 8551 3479 8557
rect 3421 8548 3433 8551
rect 1268 8520 3433 8548
rect 1268 8508 1274 8520
rect 3421 8517 3433 8520
rect 3467 8517 3479 8551
rect 3421 8511 3479 8517
rect 5994 8508 6000 8560
rect 6052 8548 6058 8560
rect 6089 8551 6147 8557
rect 6089 8548 6101 8551
rect 6052 8520 6101 8548
rect 6052 8508 6058 8520
rect 6089 8517 6101 8520
rect 6135 8517 6147 8551
rect 10134 8548 10140 8560
rect 6089 8511 6147 8517
rect 7668 8520 10140 8548
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 1903 8452 3004 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 1578 8372 1584 8424
rect 1636 8412 1642 8424
rect 2866 8412 2872 8424
rect 1636 8384 2872 8412
rect 1636 8372 1642 8384
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 2976 8412 3004 8452
rect 3142 8440 3148 8492
rect 3200 8440 3206 8492
rect 7668 8489 7696 8520
rect 10134 8508 10140 8520
rect 10192 8508 10198 8560
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8480 8355 8483
rect 8343 8452 9352 8480
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 8570 8412 8576 8424
rect 2976 8384 8576 8412
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 9125 8415 9183 8421
rect 9125 8381 9137 8415
rect 9171 8381 9183 8415
rect 9324 8412 9352 8452
rect 9398 8440 9404 8492
rect 9456 8440 9462 8492
rect 10520 8489 10548 8588
rect 12989 8585 13001 8619
rect 13035 8616 13047 8619
rect 13538 8616 13544 8628
rect 13035 8588 13544 8616
rect 13035 8585 13047 8588
rect 12989 8579 13047 8585
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14093 8619 14151 8625
rect 14093 8616 14105 8619
rect 14056 8588 14105 8616
rect 14056 8576 14062 8588
rect 14093 8585 14105 8588
rect 14139 8616 14151 8619
rect 14182 8616 14188 8628
rect 14139 8588 14188 8616
rect 14139 8585 14151 8588
rect 14093 8579 14151 8585
rect 14182 8576 14188 8588
rect 14240 8576 14246 8628
rect 14277 8619 14335 8625
rect 14277 8585 14289 8619
rect 14323 8616 14335 8619
rect 14366 8616 14372 8628
rect 14323 8588 14372 8616
rect 14323 8585 14335 8588
rect 14277 8579 14335 8585
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 15562 8616 15568 8628
rect 15120 8588 15568 8616
rect 15120 8548 15148 8588
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 16390 8576 16396 8628
rect 16448 8616 16454 8628
rect 16945 8619 17003 8625
rect 16945 8616 16957 8619
rect 16448 8588 16957 8616
rect 16448 8576 16454 8588
rect 16945 8585 16957 8588
rect 16991 8585 17003 8619
rect 16945 8579 17003 8585
rect 18049 8619 18107 8625
rect 18049 8585 18061 8619
rect 18095 8616 18107 8619
rect 18138 8616 18144 8628
rect 18095 8588 18144 8616
rect 18095 8585 18107 8588
rect 18049 8579 18107 8585
rect 18138 8576 18144 8588
rect 18196 8576 18202 8628
rect 18230 8576 18236 8628
rect 18288 8616 18294 8628
rect 18782 8616 18788 8628
rect 18288 8588 18788 8616
rect 18288 8576 18294 8588
rect 18782 8576 18788 8588
rect 18840 8576 18846 8628
rect 19886 8616 19892 8628
rect 18892 8588 19892 8616
rect 11900 8520 15148 8548
rect 15197 8551 15255 8557
rect 11900 8489 11928 8520
rect 15197 8517 15209 8551
rect 15243 8548 15255 8551
rect 18322 8548 18328 8560
rect 15243 8520 18328 8548
rect 15243 8517 15255 8520
rect 15197 8511 15255 8517
rect 18322 8508 18328 8520
rect 18380 8508 18386 8560
rect 18892 8548 18920 8588
rect 19886 8576 19892 8588
rect 19944 8576 19950 8628
rect 20898 8576 20904 8628
rect 20956 8616 20962 8628
rect 21177 8619 21235 8625
rect 21177 8616 21189 8619
rect 20956 8588 21189 8616
rect 20956 8576 20962 8588
rect 21177 8585 21189 8588
rect 21223 8585 21235 8619
rect 22922 8616 22928 8628
rect 21177 8579 21235 8585
rect 22664 8588 22928 8616
rect 20714 8548 20720 8560
rect 18616 8520 18920 8548
rect 20470 8520 20720 8548
rect 10505 8483 10563 8489
rect 10505 8449 10517 8483
rect 10551 8449 10563 8483
rect 10505 8443 10563 8449
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8449 11943 8483
rect 13357 8483 13415 8489
rect 13357 8480 13369 8483
rect 11885 8443 11943 8449
rect 12406 8452 13369 8480
rect 11514 8412 11520 8424
rect 9324 8384 11520 8412
rect 9125 8375 9183 8381
rect 2774 8304 2780 8356
rect 2832 8304 2838 8356
rect 3326 8344 3332 8356
rect 3068 8316 3332 8344
rect 2869 8279 2927 8285
rect 2869 8245 2881 8279
rect 2915 8276 2927 8279
rect 3068 8276 3096 8316
rect 3326 8304 3332 8316
rect 3384 8304 3390 8356
rect 8113 8347 8171 8353
rect 8113 8313 8125 8347
rect 8159 8344 8171 8347
rect 9140 8344 9168 8375
rect 11514 8372 11520 8384
rect 11572 8372 11578 8424
rect 11606 8372 11612 8424
rect 11664 8412 11670 8424
rect 12406 8412 12434 8452
rect 13357 8449 13369 8452
rect 13403 8480 13415 8483
rect 13403 8452 13860 8480
rect 13403 8449 13415 8452
rect 13357 8443 13415 8449
rect 11664 8384 12434 8412
rect 11664 8372 11670 8384
rect 12710 8372 12716 8424
rect 12768 8412 12774 8424
rect 13449 8415 13507 8421
rect 13449 8412 13461 8415
rect 12768 8384 13461 8412
rect 12768 8372 12774 8384
rect 13449 8381 13461 8384
rect 13495 8381 13507 8415
rect 13449 8375 13507 8381
rect 13633 8415 13691 8421
rect 13633 8381 13645 8415
rect 13679 8412 13691 8415
rect 13722 8412 13728 8424
rect 13679 8384 13728 8412
rect 13679 8381 13691 8384
rect 13633 8375 13691 8381
rect 13722 8372 13728 8384
rect 13780 8372 13786 8424
rect 13832 8412 13860 8452
rect 14550 8440 14556 8492
rect 14608 8440 14614 8492
rect 15657 8483 15715 8489
rect 15657 8449 15669 8483
rect 15703 8449 15715 8483
rect 15657 8443 15715 8449
rect 15562 8412 15568 8424
rect 13832 8384 15568 8412
rect 15562 8372 15568 8384
rect 15620 8372 15626 8424
rect 15672 8412 15700 8443
rect 15838 8440 15844 8492
rect 15896 8480 15902 8492
rect 17313 8483 17371 8489
rect 17313 8480 17325 8483
rect 15896 8452 17325 8480
rect 15896 8440 15902 8452
rect 17313 8449 17325 8452
rect 17359 8449 17371 8483
rect 17313 8443 17371 8449
rect 17405 8483 17463 8489
rect 17405 8449 17417 8483
rect 17451 8480 17463 8483
rect 18046 8480 18052 8492
rect 17451 8452 18052 8480
rect 17451 8449 17463 8452
rect 17405 8443 17463 8449
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 18233 8483 18291 8489
rect 18233 8449 18245 8483
rect 18279 8480 18291 8483
rect 18616 8480 18644 8520
rect 20714 8508 20720 8520
rect 20772 8548 20778 8560
rect 22664 8548 22692 8588
rect 22922 8576 22928 8588
rect 22980 8616 22986 8628
rect 24394 8616 24400 8628
rect 22980 8588 24400 8616
rect 22980 8576 22986 8588
rect 24394 8576 24400 8588
rect 24452 8576 24458 8628
rect 24762 8576 24768 8628
rect 24820 8616 24826 8628
rect 25133 8619 25191 8625
rect 25133 8616 25145 8619
rect 24820 8588 25145 8616
rect 24820 8576 24826 8588
rect 25133 8585 25145 8588
rect 25179 8585 25191 8619
rect 25133 8579 25191 8585
rect 26605 8619 26663 8625
rect 26605 8585 26617 8619
rect 26651 8616 26663 8619
rect 28994 8616 29000 8628
rect 26651 8588 29000 8616
rect 26651 8585 26663 8588
rect 26605 8579 26663 8585
rect 28994 8576 29000 8588
rect 29052 8576 29058 8628
rect 30653 8619 30711 8625
rect 30653 8616 30665 8619
rect 29104 8588 30665 8616
rect 20772 8520 22770 8548
rect 20772 8508 20778 8520
rect 23842 8508 23848 8560
rect 23900 8548 23906 8560
rect 29104 8548 29132 8588
rect 30653 8585 30665 8588
rect 30699 8585 30711 8619
rect 30653 8579 30711 8585
rect 31021 8619 31079 8625
rect 31021 8585 31033 8619
rect 31067 8616 31079 8619
rect 32401 8619 32459 8625
rect 31067 8588 31754 8616
rect 31067 8585 31079 8588
rect 31021 8579 31079 8585
rect 23900 8520 29132 8548
rect 30668 8548 30696 8579
rect 31481 8551 31539 8557
rect 31481 8548 31493 8551
rect 30668 8520 31493 8548
rect 23900 8508 23906 8520
rect 31481 8517 31493 8520
rect 31527 8517 31539 8551
rect 31726 8548 31754 8588
rect 32401 8585 32413 8619
rect 32447 8616 32459 8619
rect 32490 8616 32496 8628
rect 32447 8588 32496 8616
rect 32447 8585 32459 8588
rect 32401 8579 32459 8585
rect 32490 8576 32496 8588
rect 32548 8576 32554 8628
rect 32769 8619 32827 8625
rect 32769 8585 32781 8619
rect 32815 8616 32827 8619
rect 32858 8616 32864 8628
rect 32815 8588 32864 8616
rect 32815 8585 32827 8588
rect 32769 8579 32827 8585
rect 32858 8576 32864 8588
rect 32916 8576 32922 8628
rect 33962 8576 33968 8628
rect 34020 8576 34026 8628
rect 34054 8576 34060 8628
rect 34112 8576 34118 8628
rect 34885 8619 34943 8625
rect 34885 8585 34897 8619
rect 34931 8616 34943 8619
rect 36354 8616 36360 8628
rect 34931 8588 36360 8616
rect 34931 8585 34943 8588
rect 34885 8579 34943 8585
rect 36354 8576 36360 8588
rect 36412 8576 36418 8628
rect 38105 8619 38163 8625
rect 38105 8585 38117 8619
rect 38151 8616 38163 8619
rect 38286 8616 38292 8628
rect 38151 8588 38292 8616
rect 38151 8585 38163 8588
rect 38105 8579 38163 8585
rect 38286 8576 38292 8588
rect 38344 8576 38350 8628
rect 38378 8576 38384 8628
rect 38436 8616 38442 8628
rect 38565 8619 38623 8625
rect 38565 8616 38577 8619
rect 38436 8588 38577 8616
rect 38436 8576 38442 8588
rect 38565 8585 38577 8588
rect 38611 8585 38623 8619
rect 38565 8579 38623 8585
rect 39022 8576 39028 8628
rect 39080 8576 39086 8628
rect 39574 8576 39580 8628
rect 39632 8616 39638 8628
rect 41509 8619 41567 8625
rect 41509 8616 41521 8619
rect 39632 8588 41521 8616
rect 39632 8576 39638 8588
rect 41509 8585 41521 8588
rect 41555 8585 41567 8619
rect 41509 8579 41567 8585
rect 41785 8619 41843 8625
rect 41785 8585 41797 8619
rect 41831 8616 41843 8619
rect 41831 8588 42288 8616
rect 41831 8585 41843 8588
rect 41785 8579 41843 8585
rect 35253 8551 35311 8557
rect 35253 8548 35265 8551
rect 31726 8520 35265 8548
rect 31481 8511 31539 8517
rect 35253 8517 35265 8520
rect 35299 8517 35311 8551
rect 35253 8511 35311 8517
rect 18279 8452 18644 8480
rect 18279 8449 18291 8452
rect 18233 8443 18291 8449
rect 23566 8440 23572 8492
rect 23624 8480 23630 8492
rect 24029 8483 24087 8489
rect 24029 8480 24041 8483
rect 23624 8452 24041 8480
rect 23624 8440 23630 8452
rect 24029 8449 24041 8452
rect 24075 8480 24087 8483
rect 24394 8480 24400 8492
rect 24075 8452 24400 8480
rect 24075 8449 24087 8452
rect 24029 8443 24087 8449
rect 24394 8440 24400 8452
rect 24452 8440 24458 8492
rect 24486 8440 24492 8492
rect 24544 8440 24550 8492
rect 25958 8440 25964 8492
rect 26016 8440 26022 8492
rect 26602 8440 26608 8492
rect 26660 8480 26666 8492
rect 27341 8483 27399 8489
rect 27341 8480 27353 8483
rect 26660 8452 27353 8480
rect 26660 8440 26666 8452
rect 27341 8449 27353 8452
rect 27387 8449 27399 8483
rect 27341 8443 27399 8449
rect 29822 8440 29828 8492
rect 29880 8440 29886 8492
rect 31386 8440 31392 8492
rect 31444 8440 31450 8492
rect 31496 8480 31524 8511
rect 35342 8508 35348 8560
rect 35400 8508 35406 8560
rect 36630 8508 36636 8560
rect 36688 8548 36694 8560
rect 38010 8548 38016 8560
rect 36688 8520 38016 8548
rect 36688 8508 36694 8520
rect 38010 8508 38016 8520
rect 38068 8508 38074 8560
rect 38930 8508 38936 8560
rect 38988 8548 38994 8560
rect 38988 8520 39988 8548
rect 38988 8508 38994 8520
rect 32674 8480 32680 8492
rect 31496 8452 32680 8480
rect 32674 8440 32680 8452
rect 32732 8440 32738 8492
rect 36081 8483 36139 8489
rect 36081 8449 36093 8483
rect 36127 8449 36139 8483
rect 36081 8443 36139 8449
rect 15672 8384 17540 8412
rect 8159 8316 9168 8344
rect 11149 8347 11207 8353
rect 8159 8313 8171 8316
rect 8113 8307 8171 8313
rect 11149 8313 11161 8347
rect 11195 8344 11207 8347
rect 11974 8344 11980 8356
rect 11195 8316 11980 8344
rect 11195 8313 11207 8316
rect 11149 8307 11207 8313
rect 11974 8304 11980 8316
rect 12032 8304 12038 8356
rect 13170 8304 13176 8356
rect 13228 8344 13234 8356
rect 16301 8347 16359 8353
rect 13228 8316 16252 8344
rect 13228 8304 13234 8316
rect 2915 8248 3096 8276
rect 12529 8279 12587 8285
rect 2915 8245 2927 8248
rect 2869 8239 2927 8245
rect 12529 8245 12541 8279
rect 12575 8276 12587 8279
rect 12802 8276 12808 8288
rect 12575 8248 12808 8276
rect 12575 8245 12587 8248
rect 12529 8239 12587 8245
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 16224 8276 16252 8316
rect 16301 8313 16313 8347
rect 16347 8344 16359 8347
rect 16482 8344 16488 8356
rect 16347 8316 16488 8344
rect 16347 8313 16359 8316
rect 16301 8307 16359 8313
rect 16482 8304 16488 8316
rect 16540 8304 16546 8356
rect 17512 8344 17540 8384
rect 17586 8372 17592 8424
rect 17644 8372 17650 8424
rect 17954 8372 17960 8424
rect 18012 8412 18018 8424
rect 18969 8415 19027 8421
rect 18012 8384 18736 8412
rect 18012 8372 18018 8384
rect 18230 8344 18236 8356
rect 17512 8316 18236 8344
rect 18230 8304 18236 8316
rect 18288 8304 18294 8356
rect 17402 8276 17408 8288
rect 16224 8248 17408 8276
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 17770 8236 17776 8288
rect 17828 8276 17834 8288
rect 18325 8279 18383 8285
rect 18325 8276 18337 8279
rect 17828 8248 18337 8276
rect 17828 8236 17834 8248
rect 18325 8245 18337 8248
rect 18371 8245 18383 8279
rect 18325 8239 18383 8245
rect 18414 8236 18420 8288
rect 18472 8276 18478 8288
rect 18601 8279 18659 8285
rect 18601 8276 18613 8279
rect 18472 8248 18613 8276
rect 18472 8236 18478 8248
rect 18601 8245 18613 8248
rect 18647 8245 18659 8279
rect 18708 8276 18736 8384
rect 18969 8381 18981 8415
rect 19015 8412 19027 8415
rect 19242 8412 19248 8424
rect 19015 8384 19248 8412
rect 19015 8381 19027 8384
rect 18969 8375 19027 8381
rect 19242 8372 19248 8384
rect 19300 8372 19306 8424
rect 20438 8372 20444 8424
rect 20496 8412 20502 8424
rect 20717 8415 20775 8421
rect 20717 8412 20729 8415
rect 20496 8384 20729 8412
rect 20496 8372 20502 8384
rect 20717 8381 20729 8384
rect 20763 8381 20775 8415
rect 20717 8375 20775 8381
rect 21818 8372 21824 8424
rect 21876 8412 21882 8424
rect 22005 8415 22063 8421
rect 22005 8412 22017 8415
rect 21876 8384 22017 8412
rect 21876 8372 21882 8384
rect 22005 8381 22017 8384
rect 22051 8381 22063 8415
rect 23753 8415 23811 8421
rect 23753 8412 23765 8415
rect 22005 8375 22063 8381
rect 22112 8384 23765 8412
rect 20806 8304 20812 8356
rect 20864 8344 20870 8356
rect 22112 8344 22140 8384
rect 23753 8381 23765 8384
rect 23799 8381 23811 8415
rect 23753 8375 23811 8381
rect 28442 8372 28448 8424
rect 28500 8372 28506 8424
rect 28721 8415 28779 8421
rect 28721 8381 28733 8415
rect 28767 8412 28779 8415
rect 30282 8412 30288 8424
rect 28767 8384 30288 8412
rect 28767 8381 28779 8384
rect 28721 8375 28779 8381
rect 30282 8372 30288 8384
rect 30340 8372 30346 8424
rect 31665 8415 31723 8421
rect 31665 8381 31677 8415
rect 31711 8412 31723 8415
rect 31754 8412 31760 8424
rect 31711 8384 31760 8412
rect 31711 8381 31723 8384
rect 31665 8375 31723 8381
rect 31754 8372 31760 8384
rect 31812 8412 31818 8424
rect 32122 8412 32128 8424
rect 31812 8384 32128 8412
rect 31812 8372 31818 8384
rect 32122 8372 32128 8384
rect 32180 8372 32186 8424
rect 32858 8372 32864 8424
rect 32916 8372 32922 8424
rect 33042 8372 33048 8424
rect 33100 8372 33106 8424
rect 34238 8372 34244 8424
rect 34296 8372 34302 8424
rect 35434 8372 35440 8424
rect 35492 8412 35498 8424
rect 35529 8415 35587 8421
rect 35529 8412 35541 8415
rect 35492 8384 35541 8412
rect 35492 8372 35498 8384
rect 35529 8381 35541 8384
rect 35575 8412 35587 8415
rect 36096 8412 36124 8443
rect 36262 8440 36268 8492
rect 36320 8480 36326 8492
rect 36725 8483 36783 8489
rect 36725 8480 36737 8483
rect 36320 8452 36737 8480
rect 36320 8440 36326 8452
rect 36725 8449 36737 8452
rect 36771 8449 36783 8483
rect 36725 8443 36783 8449
rect 37458 8440 37464 8492
rect 37516 8440 37522 8492
rect 39960 8489 39988 8520
rect 40034 8508 40040 8560
rect 40092 8548 40098 8560
rect 41230 8548 41236 8560
rect 40092 8520 41236 8548
rect 40092 8508 40098 8520
rect 41230 8508 41236 8520
rect 41288 8548 41294 8560
rect 42061 8551 42119 8557
rect 42061 8548 42073 8551
rect 41288 8520 42073 8548
rect 41288 8508 41294 8520
rect 42061 8517 42073 8520
rect 42107 8517 42119 8551
rect 42260 8548 42288 8588
rect 42334 8576 42340 8628
rect 42392 8616 42398 8628
rect 42613 8619 42671 8625
rect 42613 8616 42625 8619
rect 42392 8588 42625 8616
rect 42392 8576 42398 8588
rect 42613 8585 42625 8588
rect 42659 8585 42671 8619
rect 42613 8579 42671 8585
rect 44174 8576 44180 8628
rect 44232 8616 44238 8628
rect 44637 8619 44695 8625
rect 44637 8616 44649 8619
rect 44232 8588 44649 8616
rect 44232 8576 44238 8588
rect 44637 8585 44649 8588
rect 44683 8585 44695 8619
rect 44637 8579 44695 8585
rect 43806 8548 43812 8560
rect 42260 8520 43812 8548
rect 42061 8511 42119 8517
rect 43806 8508 43812 8520
rect 43864 8508 43870 8560
rect 43990 8508 43996 8560
rect 44048 8548 44054 8560
rect 45189 8551 45247 8557
rect 45189 8548 45201 8551
rect 44048 8520 45201 8548
rect 44048 8508 44054 8520
rect 45189 8517 45201 8520
rect 45235 8517 45247 8551
rect 45189 8511 45247 8517
rect 45370 8508 45376 8560
rect 45428 8508 45434 8560
rect 47762 8548 47768 8560
rect 45756 8520 47768 8548
rect 38749 8483 38807 8489
rect 38749 8449 38761 8483
rect 38795 8449 38807 8483
rect 39669 8483 39727 8489
rect 39669 8480 39681 8483
rect 38749 8443 38807 8449
rect 38948 8452 39681 8480
rect 37826 8412 37832 8424
rect 35575 8384 36032 8412
rect 36096 8384 37832 8412
rect 35575 8381 35587 8384
rect 35529 8375 35587 8381
rect 20864 8316 22140 8344
rect 30193 8347 30251 8353
rect 20864 8304 20870 8316
rect 22020 8288 22048 8316
rect 30193 8313 30205 8347
rect 30239 8344 30251 8347
rect 33597 8347 33655 8353
rect 30239 8316 33548 8344
rect 30239 8313 30251 8316
rect 30193 8307 30251 8313
rect 19226 8279 19284 8285
rect 19226 8276 19238 8279
rect 18708 8248 19238 8276
rect 18601 8239 18659 8245
rect 19226 8245 19238 8248
rect 19272 8245 19284 8279
rect 19226 8239 19284 8245
rect 22002 8236 22008 8288
rect 22060 8236 22066 8288
rect 22268 8279 22326 8285
rect 22268 8245 22280 8279
rect 22314 8276 22326 8279
rect 23474 8276 23480 8288
rect 22314 8248 23480 8276
rect 22314 8245 22326 8248
rect 22268 8239 22326 8245
rect 23474 8236 23480 8248
rect 23532 8236 23538 8288
rect 27982 8236 27988 8288
rect 28040 8236 28046 8288
rect 33520 8276 33548 8316
rect 33597 8313 33609 8347
rect 33643 8344 33655 8347
rect 35802 8344 35808 8356
rect 33643 8316 35808 8344
rect 33643 8313 33655 8316
rect 33597 8307 33655 8313
rect 35802 8304 35808 8316
rect 35860 8304 35866 8356
rect 36004 8344 36032 8384
rect 37826 8372 37832 8384
rect 37884 8372 37890 8424
rect 38764 8412 38792 8443
rect 38580 8384 38792 8412
rect 37458 8344 37464 8356
rect 36004 8316 37464 8344
rect 37458 8304 37464 8316
rect 37516 8304 37522 8356
rect 38010 8304 38016 8356
rect 38068 8344 38074 8356
rect 38580 8344 38608 8384
rect 38948 8356 38976 8452
rect 39669 8449 39681 8452
rect 39715 8449 39727 8483
rect 39669 8443 39727 8449
rect 39945 8483 40003 8489
rect 39945 8449 39957 8483
rect 39991 8449 40003 8483
rect 39945 8443 40003 8449
rect 41049 8483 41107 8489
rect 41049 8449 41061 8483
rect 41095 8449 41107 8483
rect 41049 8443 41107 8449
rect 39114 8372 39120 8424
rect 39172 8412 39178 8424
rect 39301 8415 39359 8421
rect 39301 8412 39313 8415
rect 39172 8384 39313 8412
rect 39172 8372 39178 8384
rect 39301 8381 39313 8384
rect 39347 8381 39359 8415
rect 39301 8375 39359 8381
rect 39482 8372 39488 8424
rect 39540 8412 39546 8424
rect 40862 8412 40868 8424
rect 39540 8384 40868 8412
rect 39540 8372 39546 8384
rect 40862 8372 40868 8384
rect 40920 8412 40926 8424
rect 41064 8412 41092 8443
rect 42150 8440 42156 8492
rect 42208 8480 42214 8492
rect 42797 8483 42855 8489
rect 42797 8480 42809 8483
rect 42208 8452 42809 8480
rect 42208 8440 42214 8452
rect 42797 8449 42809 8452
rect 42843 8449 42855 8483
rect 42797 8443 42855 8449
rect 44174 8440 44180 8492
rect 44232 8440 44238 8492
rect 44361 8483 44419 8489
rect 44361 8449 44373 8483
rect 44407 8480 44419 8483
rect 45756 8480 45784 8520
rect 47762 8508 47768 8520
rect 47820 8508 47826 8560
rect 49142 8508 49148 8560
rect 49200 8508 49206 8560
rect 44407 8452 45784 8480
rect 45833 8483 45891 8489
rect 44407 8449 44419 8452
rect 44361 8443 44419 8449
rect 45833 8449 45845 8483
rect 45879 8449 45891 8483
rect 45833 8443 45891 8449
rect 40920 8384 41092 8412
rect 41233 8415 41291 8421
rect 40920 8372 40926 8384
rect 41233 8381 41245 8415
rect 41279 8412 41291 8415
rect 42518 8412 42524 8424
rect 41279 8384 42524 8412
rect 41279 8381 41291 8384
rect 41233 8375 41291 8381
rect 42518 8372 42524 8384
rect 42576 8372 42582 8424
rect 42702 8372 42708 8424
rect 42760 8412 42766 8424
rect 43073 8415 43131 8421
rect 43073 8412 43085 8415
rect 42760 8384 43085 8412
rect 42760 8372 42766 8384
rect 43073 8381 43085 8384
rect 43119 8381 43131 8415
rect 43073 8375 43131 8381
rect 43438 8372 43444 8424
rect 43496 8372 43502 8424
rect 38068 8316 38608 8344
rect 38068 8304 38074 8316
rect 38930 8304 38936 8356
rect 38988 8304 38994 8356
rect 41322 8304 41328 8356
rect 41380 8344 41386 8356
rect 41877 8347 41935 8353
rect 41877 8344 41889 8347
rect 41380 8316 41889 8344
rect 41380 8304 41386 8316
rect 41877 8313 41889 8316
rect 41923 8313 41935 8347
rect 41877 8307 41935 8313
rect 42058 8304 42064 8356
rect 42116 8344 42122 8356
rect 45848 8344 45876 8443
rect 47854 8440 47860 8492
rect 47912 8480 47918 8492
rect 47949 8483 48007 8489
rect 47949 8480 47961 8483
rect 47912 8452 47961 8480
rect 47912 8440 47918 8452
rect 47949 8449 47961 8452
rect 47995 8449 48007 8483
rect 47949 8443 48007 8449
rect 46842 8372 46848 8424
rect 46900 8372 46906 8424
rect 46382 8344 46388 8356
rect 42116 8316 45876 8344
rect 45940 8316 46388 8344
rect 42116 8304 42122 8316
rect 34882 8276 34888 8288
rect 33520 8248 34888 8276
rect 34882 8236 34888 8248
rect 34940 8236 34946 8288
rect 35894 8236 35900 8288
rect 35952 8276 35958 8288
rect 39942 8276 39948 8288
rect 35952 8248 39948 8276
rect 35952 8236 35958 8248
rect 39942 8236 39948 8248
rect 40000 8236 40006 8288
rect 41414 8236 41420 8288
rect 41472 8276 41478 8288
rect 45940 8276 45968 8316
rect 46382 8304 46388 8316
rect 46440 8344 46446 8356
rect 47581 8347 47639 8353
rect 47581 8344 47593 8347
rect 46440 8316 47593 8344
rect 46440 8304 46446 8316
rect 47581 8313 47593 8316
rect 47627 8313 47639 8347
rect 47581 8307 47639 8313
rect 41472 8248 45968 8276
rect 41472 8236 41478 8248
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 2130 8032 2136 8084
rect 2188 8032 2194 8084
rect 8386 8032 8392 8084
rect 8444 8032 8450 8084
rect 9766 8072 9772 8084
rect 8496 8044 9772 8072
rect 1765 8007 1823 8013
rect 1765 7973 1777 8007
rect 1811 8004 1823 8007
rect 8496 8004 8524 8044
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 11333 8075 11391 8081
rect 11333 8041 11345 8075
rect 11379 8072 11391 8075
rect 11422 8072 11428 8084
rect 11379 8044 11428 8072
rect 11379 8041 11391 8044
rect 11333 8035 11391 8041
rect 11422 8032 11428 8044
rect 11480 8032 11486 8084
rect 13725 8075 13783 8081
rect 13725 8072 13737 8075
rect 11532 8044 13737 8072
rect 1811 7976 8524 8004
rect 1811 7973 1823 7976
rect 1765 7967 1823 7973
rect 10042 7896 10048 7948
rect 10100 7896 10106 7948
rect 10689 7939 10747 7945
rect 10689 7905 10701 7939
rect 10735 7936 10747 7939
rect 11146 7936 11152 7948
rect 10735 7908 11152 7936
rect 10735 7905 10747 7908
rect 10689 7899 10747 7905
rect 11146 7896 11152 7908
rect 11204 7896 11210 7948
rect 11532 7936 11560 8044
rect 13725 8041 13737 8044
rect 13771 8041 13783 8075
rect 13725 8035 13783 8041
rect 14553 8075 14611 8081
rect 14553 8041 14565 8075
rect 14599 8072 14611 8075
rect 14734 8072 14740 8084
rect 14599 8044 14740 8072
rect 14599 8041 14611 8044
rect 14553 8035 14611 8041
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 15841 8075 15899 8081
rect 15841 8041 15853 8075
rect 15887 8072 15899 8075
rect 17954 8072 17960 8084
rect 15887 8044 17960 8072
rect 15887 8041 15899 8044
rect 15841 8035 15899 8041
rect 17954 8032 17960 8044
rect 18012 8032 18018 8084
rect 18414 8032 18420 8084
rect 18472 8072 18478 8084
rect 18969 8075 19027 8081
rect 18969 8072 18981 8075
rect 18472 8044 18981 8072
rect 18472 8032 18478 8044
rect 18969 8041 18981 8044
rect 19015 8072 19027 8075
rect 19242 8072 19248 8084
rect 19015 8044 19248 8072
rect 19015 8041 19027 8044
rect 18969 8035 19027 8041
rect 19242 8032 19248 8044
rect 19300 8032 19306 8084
rect 21269 8075 21327 8081
rect 21269 8041 21281 8075
rect 21315 8072 21327 8075
rect 21450 8072 21456 8084
rect 21315 8044 21456 8072
rect 21315 8041 21327 8044
rect 21269 8035 21327 8041
rect 21450 8032 21456 8044
rect 21508 8032 21514 8084
rect 22186 8032 22192 8084
rect 22244 8072 22250 8084
rect 22244 8044 22784 8072
rect 22244 8032 22250 8044
rect 15194 8004 15200 8016
rect 11256 7908 11560 7936
rect 11624 7976 15200 8004
rect 1302 7828 1308 7880
rect 1360 7868 1366 7880
rect 1581 7871 1639 7877
rect 1581 7868 1593 7871
rect 1360 7840 1593 7868
rect 1360 7828 1366 7840
rect 1581 7837 1593 7840
rect 1627 7868 1639 7871
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 1627 7840 2329 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 2317 7837 2329 7840
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 8570 7828 8576 7880
rect 8628 7828 8634 7880
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7868 9367 7871
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 9355 7840 9597 7868
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 9585 7837 9597 7840
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 9600 7800 9628 7831
rect 10226 7828 10232 7880
rect 10284 7868 10290 7880
rect 11256 7868 11284 7908
rect 10284 7840 11284 7868
rect 10284 7828 10290 7840
rect 11330 7828 11336 7880
rect 11388 7868 11394 7880
rect 11517 7871 11575 7877
rect 11517 7868 11529 7871
rect 11388 7840 11529 7868
rect 11388 7828 11394 7840
rect 11517 7837 11529 7840
rect 11563 7837 11575 7871
rect 11517 7831 11575 7837
rect 11624 7800 11652 7976
rect 15194 7964 15200 7976
rect 15252 7964 15258 8016
rect 17770 7964 17776 8016
rect 17828 8004 17834 8016
rect 18049 8007 18107 8013
rect 18049 8004 18061 8007
rect 17828 7976 18061 8004
rect 17828 7964 17834 7976
rect 18049 7973 18061 7976
rect 18095 7973 18107 8007
rect 18049 7967 18107 7973
rect 21174 7964 21180 8016
rect 21232 8004 21238 8016
rect 22756 8013 22784 8044
rect 23750 8032 23756 8084
rect 23808 8072 23814 8084
rect 24029 8075 24087 8081
rect 24029 8072 24041 8075
rect 23808 8044 24041 8072
rect 23808 8032 23814 8044
rect 24029 8041 24041 8044
rect 24075 8041 24087 8075
rect 24029 8035 24087 8041
rect 24394 8032 24400 8084
rect 24452 8032 24458 8084
rect 26789 8075 26847 8081
rect 26789 8041 26801 8075
rect 26835 8072 26847 8075
rect 27062 8072 27068 8084
rect 26835 8044 27068 8072
rect 26835 8041 26847 8044
rect 26789 8035 26847 8041
rect 27062 8032 27068 8044
rect 27120 8032 27126 8084
rect 27798 8032 27804 8084
rect 27856 8072 27862 8084
rect 28077 8075 28135 8081
rect 28077 8072 28089 8075
rect 27856 8044 28089 8072
rect 27856 8032 27862 8044
rect 28077 8041 28089 8044
rect 28123 8041 28135 8075
rect 28077 8035 28135 8041
rect 28350 8032 28356 8084
rect 28408 8072 28414 8084
rect 32953 8075 33011 8081
rect 32953 8072 32965 8075
rect 28408 8044 32965 8072
rect 28408 8032 28414 8044
rect 32953 8041 32965 8044
rect 32999 8041 33011 8075
rect 32953 8035 33011 8041
rect 34241 8075 34299 8081
rect 34241 8041 34253 8075
rect 34287 8072 34299 8075
rect 35894 8072 35900 8084
rect 34287 8044 35900 8072
rect 34287 8041 34299 8044
rect 34241 8035 34299 8041
rect 35894 8032 35900 8044
rect 35952 8032 35958 8084
rect 35986 8032 35992 8084
rect 36044 8072 36050 8084
rect 36044 8044 44128 8072
rect 36044 8032 36050 8044
rect 22373 8007 22431 8013
rect 22373 8004 22385 8007
rect 21232 7976 22385 8004
rect 21232 7964 21238 7976
rect 22373 7973 22385 7976
rect 22419 7973 22431 8007
rect 22373 7967 22431 7973
rect 22741 8007 22799 8013
rect 22741 7973 22753 8007
rect 22787 8004 22799 8007
rect 23842 8004 23848 8016
rect 22787 7976 23848 8004
rect 22787 7973 22799 7976
rect 22741 7967 22799 7973
rect 23842 7964 23848 7976
rect 23900 7964 23906 8016
rect 27430 7964 27436 8016
rect 27488 8004 27494 8016
rect 29181 8007 29239 8013
rect 29181 8004 29193 8007
rect 27488 7976 29193 8004
rect 27488 7964 27494 7976
rect 29181 7973 29193 7976
rect 29227 7973 29239 8007
rect 29181 7967 29239 7973
rect 31110 7964 31116 8016
rect 31168 8004 31174 8016
rect 31168 7976 35112 8004
rect 31168 7964 31174 7976
rect 12066 7896 12072 7948
rect 12124 7936 12130 7948
rect 12621 7939 12679 7945
rect 12621 7936 12633 7939
rect 12124 7908 12633 7936
rect 12124 7896 12130 7908
rect 12621 7905 12633 7908
rect 12667 7905 12679 7939
rect 22554 7936 22560 7948
rect 12621 7899 12679 7905
rect 14752 7908 22560 7936
rect 11974 7828 11980 7880
rect 12032 7828 12038 7880
rect 14752 7877 14780 7908
rect 22554 7896 22560 7908
rect 22612 7896 22618 7948
rect 31754 7896 31760 7948
rect 31812 7936 31818 7948
rect 31849 7939 31907 7945
rect 31849 7936 31861 7939
rect 31812 7908 31861 7936
rect 31812 7896 31818 7908
rect 31849 7905 31861 7908
rect 31895 7905 31907 7939
rect 31849 7899 31907 7905
rect 13081 7871 13139 7877
rect 13081 7837 13093 7871
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 14737 7871 14795 7877
rect 14737 7837 14749 7871
rect 14783 7837 14795 7871
rect 14737 7831 14795 7837
rect 9600 7772 11652 7800
rect 13096 7800 13124 7831
rect 15194 7828 15200 7880
rect 15252 7828 15258 7880
rect 16298 7828 16304 7880
rect 16356 7828 16362 7880
rect 19521 7871 19579 7877
rect 19521 7837 19533 7871
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 13096 7772 16528 7800
rect 7466 7692 7472 7744
rect 7524 7732 7530 7744
rect 9401 7735 9459 7741
rect 9401 7732 9413 7735
rect 7524 7704 9413 7732
rect 7524 7692 7530 7704
rect 9401 7701 9413 7704
rect 9447 7701 9459 7735
rect 9401 7695 9459 7701
rect 14182 7692 14188 7744
rect 14240 7692 14246 7744
rect 16500 7732 16528 7772
rect 16574 7760 16580 7812
rect 16632 7760 16638 7812
rect 17034 7760 17040 7812
rect 17092 7760 17098 7812
rect 18690 7800 18696 7812
rect 18432 7772 18696 7800
rect 18432 7732 18460 7772
rect 18690 7760 18696 7772
rect 18748 7760 18754 7812
rect 19536 7800 19564 7831
rect 19610 7828 19616 7880
rect 19668 7868 19674 7880
rect 20625 7871 20683 7877
rect 20625 7868 20637 7871
rect 19668 7840 20637 7868
rect 19668 7828 19674 7840
rect 20625 7837 20637 7840
rect 20671 7837 20683 7871
rect 20625 7831 20683 7837
rect 21726 7828 21732 7880
rect 21784 7828 21790 7880
rect 23385 7871 23443 7877
rect 23385 7837 23397 7871
rect 23431 7868 23443 7871
rect 24946 7868 24952 7880
rect 23431 7840 24952 7868
rect 23431 7837 23443 7840
rect 23385 7831 23443 7837
rect 24946 7828 24952 7840
rect 25004 7828 25010 7880
rect 25038 7828 25044 7880
rect 25096 7828 25102 7880
rect 25685 7871 25743 7877
rect 25685 7837 25697 7871
rect 25731 7868 25743 7871
rect 26145 7871 26203 7877
rect 26145 7868 26157 7871
rect 25731 7840 26157 7868
rect 25731 7837 25743 7840
rect 25685 7831 25743 7837
rect 26145 7837 26157 7840
rect 26191 7837 26203 7871
rect 26145 7831 26203 7837
rect 27433 7871 27491 7877
rect 27433 7837 27445 7871
rect 27479 7868 27491 7871
rect 27982 7868 27988 7880
rect 27479 7840 27988 7868
rect 27479 7837 27491 7840
rect 27433 7831 27491 7837
rect 27982 7828 27988 7840
rect 28040 7828 28046 7880
rect 28537 7871 28595 7877
rect 28537 7837 28549 7871
rect 28583 7868 28595 7871
rect 29362 7868 29368 7880
rect 28583 7840 29368 7868
rect 28583 7837 28595 7840
rect 28537 7831 28595 7837
rect 29362 7828 29368 7840
rect 29420 7828 29426 7880
rect 29454 7828 29460 7880
rect 29512 7868 29518 7880
rect 29733 7871 29791 7877
rect 29733 7868 29745 7871
rect 29512 7840 29745 7868
rect 29512 7828 29518 7840
rect 29733 7837 29745 7840
rect 29779 7837 29791 7871
rect 29733 7831 29791 7837
rect 30837 7871 30895 7877
rect 30837 7837 30849 7871
rect 30883 7868 30895 7871
rect 30926 7868 30932 7880
rect 30883 7840 30932 7868
rect 30883 7837 30895 7840
rect 30837 7831 30895 7837
rect 30926 7828 30932 7840
rect 30984 7828 30990 7880
rect 31570 7828 31576 7880
rect 31628 7868 31634 7880
rect 32309 7871 32367 7877
rect 32309 7868 32321 7871
rect 31628 7840 32321 7868
rect 31628 7828 31634 7840
rect 32309 7837 32321 7840
rect 32355 7837 32367 7871
rect 32309 7831 32367 7837
rect 32950 7828 32956 7880
rect 33008 7868 33014 7880
rect 33318 7868 33324 7880
rect 33008 7840 33324 7868
rect 33008 7828 33014 7840
rect 33318 7828 33324 7840
rect 33376 7828 33382 7880
rect 33597 7871 33655 7877
rect 33597 7837 33609 7871
rect 33643 7868 33655 7871
rect 34514 7868 34520 7880
rect 33643 7840 34520 7868
rect 33643 7837 33655 7840
rect 33597 7831 33655 7837
rect 34514 7828 34520 7840
rect 34572 7828 34578 7880
rect 34882 7828 34888 7880
rect 34940 7828 34946 7880
rect 35084 7868 35112 7976
rect 37476 7976 39436 8004
rect 35618 7896 35624 7948
rect 35676 7936 35682 7948
rect 37476 7936 37504 7976
rect 39301 7939 39359 7945
rect 39301 7936 39313 7939
rect 35676 7908 37504 7936
rect 37752 7908 39313 7936
rect 35676 7896 35682 7908
rect 37369 7871 37427 7877
rect 37369 7868 37381 7871
rect 35084 7840 37381 7868
rect 37369 7837 37381 7840
rect 37415 7837 37427 7871
rect 37369 7831 37427 7837
rect 22002 7800 22008 7812
rect 19536 7772 22008 7800
rect 22002 7760 22008 7772
rect 22060 7760 22066 7812
rect 30377 7803 30435 7809
rect 30377 7769 30389 7803
rect 30423 7800 30435 7803
rect 30423 7772 32812 7800
rect 30423 7769 30435 7772
rect 30377 7763 30435 7769
rect 16500 7704 18460 7732
rect 18509 7735 18567 7741
rect 18509 7701 18521 7735
rect 18555 7732 18567 7735
rect 19518 7732 19524 7744
rect 18555 7704 19524 7732
rect 18555 7701 18567 7704
rect 18509 7695 18567 7701
rect 19518 7692 19524 7704
rect 19576 7692 19582 7744
rect 20165 7735 20223 7741
rect 20165 7701 20177 7735
rect 20211 7732 20223 7735
rect 20254 7732 20260 7744
rect 20211 7704 20260 7732
rect 20211 7701 20223 7704
rect 20165 7695 20223 7701
rect 20254 7692 20260 7704
rect 20312 7692 20318 7744
rect 22922 7692 22928 7744
rect 22980 7732 22986 7744
rect 23290 7732 23296 7744
rect 22980 7704 23296 7732
rect 22980 7692 22986 7704
rect 23290 7692 23296 7704
rect 23348 7692 23354 7744
rect 30926 7692 30932 7744
rect 30984 7732 30990 7744
rect 31481 7735 31539 7741
rect 31481 7732 31493 7735
rect 30984 7704 31493 7732
rect 30984 7692 30990 7704
rect 31481 7701 31493 7704
rect 31527 7701 31539 7735
rect 32784 7732 32812 7772
rect 32858 7760 32864 7812
rect 32916 7800 32922 7812
rect 35529 7803 35587 7809
rect 35529 7800 35541 7803
rect 32916 7772 35541 7800
rect 32916 7760 32922 7772
rect 35529 7769 35541 7772
rect 35575 7769 35587 7803
rect 35529 7763 35587 7769
rect 36170 7760 36176 7812
rect 36228 7800 36234 7812
rect 37752 7800 37780 7908
rect 39301 7905 39313 7908
rect 39347 7905 39359 7939
rect 39408 7936 39436 7976
rect 40586 7964 40592 8016
rect 40644 7964 40650 8016
rect 40862 7964 40868 8016
rect 40920 7964 40926 8016
rect 41046 7964 41052 8016
rect 41104 7964 41110 8016
rect 41230 7964 41236 8016
rect 41288 7964 41294 8016
rect 41690 7964 41696 8016
rect 41748 7964 41754 8016
rect 41966 7964 41972 8016
rect 42024 7964 42030 8016
rect 42150 7964 42156 8016
rect 42208 7964 42214 8016
rect 43990 7964 43996 8016
rect 44048 7964 44054 8016
rect 42337 7939 42395 7945
rect 42337 7936 42349 7939
rect 39408 7908 42349 7936
rect 39301 7899 39359 7905
rect 42337 7905 42349 7908
rect 42383 7905 42395 7939
rect 42337 7899 42395 7905
rect 37826 7828 37832 7880
rect 37884 7868 37890 7880
rect 37921 7871 37979 7877
rect 37921 7868 37933 7871
rect 37884 7840 37933 7868
rect 37884 7828 37890 7840
rect 37921 7837 37933 7840
rect 37967 7837 37979 7871
rect 37921 7831 37979 7837
rect 38841 7871 38899 7877
rect 38841 7837 38853 7871
rect 38887 7868 38899 7871
rect 40218 7868 40224 7880
rect 38887 7840 40224 7868
rect 38887 7837 38899 7840
rect 38841 7831 38899 7837
rect 40218 7828 40224 7840
rect 40276 7828 40282 7880
rect 41046 7828 41052 7880
rect 41104 7868 41110 7880
rect 41104 7840 42748 7868
rect 41104 7828 41110 7840
rect 36228 7772 37780 7800
rect 38657 7803 38715 7809
rect 36228 7760 36234 7772
rect 38657 7769 38669 7803
rect 38703 7800 38715 7803
rect 39022 7800 39028 7812
rect 38703 7772 39028 7800
rect 38703 7769 38715 7772
rect 38657 7763 38715 7769
rect 39022 7760 39028 7772
rect 39080 7760 39086 7812
rect 40126 7760 40132 7812
rect 40184 7760 40190 7812
rect 40313 7803 40371 7809
rect 40313 7769 40325 7803
rect 40359 7800 40371 7803
rect 42610 7800 42616 7812
rect 40359 7772 42616 7800
rect 40359 7769 40371 7772
rect 40313 7763 40371 7769
rect 42610 7760 42616 7772
rect 42668 7760 42674 7812
rect 34422 7732 34428 7744
rect 32784 7704 34428 7732
rect 31481 7695 31539 7701
rect 34422 7692 34428 7704
rect 34480 7692 34486 7744
rect 37182 7692 37188 7744
rect 37240 7692 37246 7744
rect 38013 7735 38071 7741
rect 38013 7701 38025 7735
rect 38059 7732 38071 7735
rect 39206 7732 39212 7744
rect 38059 7704 39212 7732
rect 38059 7701 38071 7704
rect 38013 7695 38071 7701
rect 39206 7692 39212 7704
rect 39264 7692 39270 7744
rect 41506 7692 41512 7744
rect 41564 7692 41570 7744
rect 42720 7741 42748 7840
rect 42886 7828 42892 7880
rect 42944 7828 42950 7880
rect 43530 7828 43536 7880
rect 43588 7828 43594 7880
rect 44100 7864 44128 8044
rect 44634 8032 44640 8084
rect 44692 8072 44698 8084
rect 44729 8075 44787 8081
rect 44729 8072 44741 8075
rect 44692 8044 44741 8072
rect 44692 8032 44698 8044
rect 44729 8041 44741 8044
rect 44775 8041 44787 8075
rect 44729 8035 44787 8041
rect 45186 8032 45192 8084
rect 45244 8032 45250 8084
rect 45557 8075 45615 8081
rect 45557 8041 45569 8075
rect 45603 8072 45615 8075
rect 47026 8072 47032 8084
rect 45603 8044 47032 8072
rect 45603 8041 45615 8044
rect 45557 8035 45615 8041
rect 47026 8032 47032 8044
rect 47084 8032 47090 8084
rect 44910 7964 44916 8016
rect 44968 8004 44974 8016
rect 47489 8007 47547 8013
rect 47489 8004 47501 8007
rect 44968 7976 47501 8004
rect 44968 7964 44974 7976
rect 47489 7973 47501 7976
rect 47535 7973 47547 8007
rect 47489 7967 47547 7973
rect 44542 7896 44548 7948
rect 44600 7896 44606 7948
rect 45370 7896 45376 7948
rect 45428 7936 45434 7948
rect 49050 7936 49056 7948
rect 45428 7908 49056 7936
rect 45428 7896 45434 7908
rect 46216 7877 46244 7908
rect 49050 7896 49056 7908
rect 49108 7896 49114 7948
rect 49145 7939 49203 7945
rect 49145 7905 49157 7939
rect 49191 7936 49203 7939
rect 49234 7936 49240 7948
rect 49191 7908 49240 7936
rect 49191 7905 49203 7908
rect 49145 7899 49203 7905
rect 49234 7896 49240 7908
rect 49292 7896 49298 7948
rect 44177 7871 44235 7877
rect 44177 7864 44189 7871
rect 44100 7837 44189 7864
rect 44223 7837 44235 7871
rect 44100 7836 44235 7837
rect 44177 7831 44235 7836
rect 45741 7871 45799 7877
rect 45741 7837 45753 7871
rect 45787 7837 45799 7871
rect 45741 7831 45799 7837
rect 46201 7871 46259 7877
rect 46201 7837 46213 7871
rect 46247 7837 46259 7871
rect 46201 7831 46259 7837
rect 46937 7871 46995 7877
rect 46937 7837 46949 7871
rect 46983 7837 46995 7871
rect 46937 7831 46995 7837
rect 42705 7735 42763 7741
rect 42705 7701 42717 7735
rect 42751 7701 42763 7735
rect 42904 7732 42932 7828
rect 43714 7760 43720 7812
rect 43772 7800 43778 7812
rect 45756 7800 45784 7831
rect 43772 7772 45784 7800
rect 46952 7800 46980 7831
rect 47118 7828 47124 7880
rect 47176 7868 47182 7880
rect 47949 7871 48007 7877
rect 47949 7868 47961 7871
rect 47176 7840 47961 7868
rect 47176 7828 47182 7840
rect 47949 7837 47961 7840
rect 47995 7837 48007 7871
rect 47949 7831 48007 7837
rect 48314 7800 48320 7812
rect 46952 7772 48320 7800
rect 43772 7760 43778 7772
rect 48314 7760 48320 7772
rect 48372 7800 48378 7812
rect 49970 7800 49976 7812
rect 48372 7772 49976 7800
rect 48372 7760 48378 7772
rect 49970 7760 49976 7772
rect 50028 7760 50034 7812
rect 43162 7732 43168 7744
rect 42904 7704 43168 7732
rect 42705 7695 42763 7701
rect 43162 7692 43168 7704
rect 43220 7692 43226 7744
rect 43346 7692 43352 7744
rect 43404 7692 43410 7744
rect 44082 7692 44088 7744
rect 44140 7732 44146 7744
rect 45005 7735 45063 7741
rect 45005 7732 45017 7735
rect 44140 7704 45017 7732
rect 44140 7692 44146 7704
rect 45005 7701 45017 7704
rect 45051 7701 45063 7735
rect 45005 7695 45063 7701
rect 46382 7692 46388 7744
rect 46440 7692 46446 7744
rect 46934 7692 46940 7744
rect 46992 7732 46998 7744
rect 47121 7735 47179 7741
rect 47121 7732 47133 7735
rect 46992 7704 47133 7732
rect 46992 7692 46998 7704
rect 47121 7701 47133 7704
rect 47167 7701 47179 7735
rect 47121 7695 47179 7701
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 9214 7488 9220 7540
rect 9272 7528 9278 7540
rect 9769 7531 9827 7537
rect 9769 7528 9781 7531
rect 9272 7500 9781 7528
rect 9272 7488 9278 7500
rect 9769 7497 9781 7500
rect 9815 7497 9827 7531
rect 9769 7491 9827 7497
rect 10321 7531 10379 7537
rect 10321 7497 10333 7531
rect 10367 7528 10379 7531
rect 10413 7531 10471 7537
rect 10413 7528 10425 7531
rect 10367 7500 10425 7528
rect 10367 7497 10379 7500
rect 10321 7491 10379 7497
rect 10413 7497 10425 7500
rect 10459 7528 10471 7531
rect 11238 7528 11244 7540
rect 10459 7500 11244 7528
rect 10459 7497 10471 7500
rect 10413 7491 10471 7497
rect 11238 7488 11244 7500
rect 11296 7488 11302 7540
rect 11330 7488 11336 7540
rect 11388 7488 11394 7540
rect 11793 7531 11851 7537
rect 11793 7497 11805 7531
rect 11839 7497 11851 7531
rect 11793 7491 11851 7497
rect 12437 7531 12495 7537
rect 12437 7497 12449 7531
rect 12483 7528 12495 7531
rect 12526 7528 12532 7540
rect 12483 7500 12532 7528
rect 12483 7497 12495 7500
rect 12437 7491 12495 7497
rect 6086 7420 6092 7472
rect 6144 7460 6150 7472
rect 11808 7460 11836 7491
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 14090 7488 14096 7540
rect 14148 7488 14154 7540
rect 15194 7488 15200 7540
rect 15252 7528 15258 7540
rect 16301 7531 16359 7537
rect 16301 7528 16313 7531
rect 15252 7500 16313 7528
rect 15252 7488 15258 7500
rect 16301 7497 16313 7500
rect 16347 7497 16359 7531
rect 16301 7491 16359 7497
rect 16666 7488 16672 7540
rect 16724 7488 16730 7540
rect 17313 7531 17371 7537
rect 17313 7497 17325 7531
rect 17359 7528 17371 7531
rect 18969 7531 19027 7537
rect 18969 7528 18981 7531
rect 17359 7500 18981 7528
rect 17359 7497 17371 7500
rect 17313 7491 17371 7497
rect 18969 7497 18981 7500
rect 19015 7497 19027 7531
rect 18969 7491 19027 7497
rect 19978 7488 19984 7540
rect 20036 7528 20042 7540
rect 20349 7531 20407 7537
rect 20349 7528 20361 7531
rect 20036 7500 20361 7528
rect 20036 7488 20042 7500
rect 20349 7497 20361 7500
rect 20395 7497 20407 7531
rect 20349 7491 20407 7497
rect 27706 7488 27712 7540
rect 27764 7528 27770 7540
rect 28169 7531 28227 7537
rect 28169 7528 28181 7531
rect 27764 7500 28181 7528
rect 27764 7488 27770 7500
rect 28169 7497 28181 7500
rect 28215 7497 28227 7531
rect 28169 7491 28227 7497
rect 29362 7488 29368 7540
rect 29420 7488 29426 7540
rect 31570 7488 31576 7540
rect 31628 7488 31634 7540
rect 32582 7488 32588 7540
rect 32640 7528 32646 7540
rect 34241 7531 34299 7537
rect 34241 7528 34253 7531
rect 32640 7500 34253 7528
rect 32640 7488 32646 7500
rect 34241 7497 34253 7500
rect 34287 7497 34299 7531
rect 34241 7491 34299 7497
rect 34514 7488 34520 7540
rect 34572 7488 34578 7540
rect 37366 7528 37372 7540
rect 35728 7500 37372 7528
rect 12710 7460 12716 7472
rect 6144 7432 11836 7460
rect 12636 7432 12716 7460
rect 6144 7420 6150 7432
rect 1302 7352 1308 7404
rect 1360 7392 1366 7404
rect 1581 7395 1639 7401
rect 1581 7392 1593 7395
rect 1360 7364 1593 7392
rect 1360 7352 1366 7364
rect 1581 7361 1593 7364
rect 1627 7392 1639 7395
rect 2133 7395 2191 7401
rect 2133 7392 2145 7395
rect 1627 7364 2145 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 2133 7361 2145 7364
rect 2179 7361 2191 7395
rect 2133 7355 2191 7361
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7392 9183 7395
rect 9490 7392 9496 7404
rect 9171 7364 9496 7392
rect 9171 7361 9183 7364
rect 9125 7355 9183 7361
rect 9490 7352 9496 7364
rect 9548 7352 9554 7404
rect 9950 7352 9956 7404
rect 10008 7352 10014 7404
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7392 11207 7395
rect 11974 7392 11980 7404
rect 11195 7364 11980 7392
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 11974 7352 11980 7364
rect 12032 7352 12038 7404
rect 12636 7401 12664 7432
rect 12710 7420 12716 7432
rect 12768 7460 12774 7472
rect 15746 7460 15752 7472
rect 12768 7432 15752 7460
rect 12768 7420 12774 7432
rect 15746 7420 15752 7432
rect 15804 7420 15810 7472
rect 16945 7463 17003 7469
rect 16945 7429 16957 7463
rect 16991 7460 17003 7463
rect 17402 7460 17408 7472
rect 16991 7432 17408 7460
rect 16991 7429 17003 7432
rect 16945 7423 17003 7429
rect 17402 7420 17408 7432
rect 17460 7420 17466 7472
rect 17494 7420 17500 7472
rect 17552 7460 17558 7472
rect 18877 7463 18935 7469
rect 18877 7460 18889 7463
rect 17552 7432 18889 7460
rect 17552 7420 17558 7432
rect 18877 7429 18889 7432
rect 18923 7429 18935 7463
rect 22186 7460 22192 7472
rect 18877 7423 18935 7429
rect 19306 7432 22192 7460
rect 12621 7395 12679 7401
rect 12621 7361 12633 7395
rect 12667 7361 12679 7395
rect 12621 7355 12679 7361
rect 12802 7352 12808 7404
rect 12860 7392 12866 7404
rect 13081 7395 13139 7401
rect 13081 7392 13093 7395
rect 12860 7364 13093 7392
rect 12860 7352 12866 7364
rect 13081 7361 13093 7364
rect 13127 7361 13139 7395
rect 13081 7355 13139 7361
rect 14553 7395 14611 7401
rect 14553 7361 14565 7395
rect 14599 7392 14611 7395
rect 15562 7392 15568 7404
rect 14599 7364 15568 7392
rect 14599 7361 14611 7364
rect 14553 7355 14611 7361
rect 15562 7352 15568 7364
rect 15620 7352 15626 7404
rect 15657 7395 15715 7401
rect 15657 7361 15669 7395
rect 15703 7392 15715 7395
rect 17586 7392 17592 7404
rect 15703 7364 17592 7392
rect 15703 7361 15715 7364
rect 15657 7355 15715 7361
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 17681 7395 17739 7401
rect 17681 7361 17693 7395
rect 17727 7392 17739 7395
rect 18322 7392 18328 7404
rect 17727 7364 18328 7392
rect 17727 7361 17739 7364
rect 17681 7355 17739 7361
rect 18322 7352 18328 7364
rect 18380 7392 18386 7404
rect 19306 7392 19334 7432
rect 22186 7420 22192 7432
rect 22244 7420 22250 7472
rect 33137 7463 33195 7469
rect 33137 7429 33149 7463
rect 33183 7460 33195 7463
rect 35728 7460 35756 7500
rect 37366 7488 37372 7500
rect 37424 7488 37430 7540
rect 39761 7531 39819 7537
rect 39761 7497 39773 7531
rect 39807 7528 39819 7531
rect 39807 7500 44956 7528
rect 39807 7497 39819 7500
rect 39761 7491 39819 7497
rect 33183 7432 35756 7460
rect 33183 7429 33195 7432
rect 33137 7423 33195 7429
rect 35802 7420 35808 7472
rect 35860 7460 35866 7472
rect 35860 7432 39988 7460
rect 35860 7420 35866 7432
rect 18380 7364 19334 7392
rect 18380 7352 18386 7364
rect 19702 7352 19708 7404
rect 19760 7352 19766 7404
rect 20809 7395 20867 7401
rect 20809 7361 20821 7395
rect 20855 7392 20867 7395
rect 22646 7392 22652 7404
rect 20855 7364 22652 7392
rect 20855 7361 20867 7364
rect 20809 7355 20867 7361
rect 22646 7352 22652 7364
rect 22704 7352 22710 7404
rect 22741 7395 22799 7401
rect 22741 7361 22753 7395
rect 22787 7392 22799 7395
rect 22830 7392 22836 7404
rect 22787 7364 22836 7392
rect 22787 7361 22799 7364
rect 22741 7355 22799 7361
rect 22830 7352 22836 7364
rect 22888 7352 22894 7404
rect 23845 7395 23903 7401
rect 23845 7361 23857 7395
rect 23891 7392 23903 7395
rect 24670 7392 24676 7404
rect 23891 7364 24676 7392
rect 23891 7361 23903 7364
rect 23845 7355 23903 7361
rect 24670 7352 24676 7364
rect 24728 7352 24734 7404
rect 24949 7395 25007 7401
rect 24949 7361 24961 7395
rect 24995 7392 25007 7395
rect 25222 7392 25228 7404
rect 24995 7364 25228 7392
rect 24995 7361 25007 7364
rect 24949 7355 25007 7361
rect 25222 7352 25228 7364
rect 25280 7352 25286 7404
rect 27525 7395 27583 7401
rect 27525 7361 27537 7395
rect 27571 7392 27583 7395
rect 28350 7392 28356 7404
rect 27571 7364 28356 7392
rect 27571 7361 27583 7364
rect 27525 7355 27583 7361
rect 28350 7352 28356 7364
rect 28408 7352 28414 7404
rect 28721 7395 28779 7401
rect 28721 7361 28733 7395
rect 28767 7361 28779 7395
rect 28721 7355 28779 7361
rect 29825 7395 29883 7401
rect 29825 7361 29837 7395
rect 29871 7392 29883 7395
rect 29914 7392 29920 7404
rect 29871 7364 29920 7392
rect 29871 7361 29883 7364
rect 29825 7355 29883 7361
rect 10686 7284 10692 7336
rect 10744 7324 10750 7336
rect 13725 7327 13783 7333
rect 13725 7324 13737 7327
rect 10744 7296 13737 7324
rect 10744 7284 10750 7296
rect 13725 7293 13737 7296
rect 13771 7293 13783 7327
rect 13725 7287 13783 7293
rect 14826 7284 14832 7336
rect 14884 7324 14890 7336
rect 15197 7327 15255 7333
rect 15197 7324 15209 7327
rect 14884 7296 15209 7324
rect 14884 7284 14890 7296
rect 15197 7293 15209 7296
rect 15243 7293 15255 7327
rect 15197 7287 15255 7293
rect 16758 7284 16764 7336
rect 16816 7324 16822 7336
rect 17773 7327 17831 7333
rect 17773 7324 17785 7327
rect 16816 7296 17785 7324
rect 16816 7284 16822 7296
rect 17773 7293 17785 7296
rect 17819 7293 17831 7327
rect 17773 7287 17831 7293
rect 17862 7284 17868 7336
rect 17920 7284 17926 7336
rect 18506 7284 18512 7336
rect 18564 7324 18570 7336
rect 19061 7327 19119 7333
rect 19061 7324 19073 7327
rect 18564 7296 19073 7324
rect 18564 7284 18570 7296
rect 19061 7293 19073 7296
rect 19107 7293 19119 7327
rect 19061 7287 19119 7293
rect 22922 7284 22928 7336
rect 22980 7324 22986 7336
rect 28736 7324 28764 7355
rect 29914 7352 29920 7364
rect 29972 7352 29978 7404
rect 30926 7352 30932 7404
rect 30984 7352 30990 7404
rect 32493 7395 32551 7401
rect 32493 7361 32505 7395
rect 32539 7392 32551 7395
rect 32766 7392 32772 7404
rect 32539 7364 32772 7392
rect 32539 7361 32551 7364
rect 32493 7355 32551 7361
rect 32766 7352 32772 7364
rect 32824 7352 32830 7404
rect 33597 7395 33655 7401
rect 33597 7361 33609 7395
rect 33643 7361 33655 7395
rect 33597 7355 33655 7361
rect 34885 7395 34943 7401
rect 34885 7361 34897 7395
rect 34931 7392 34943 7395
rect 35526 7392 35532 7404
rect 34931 7364 35532 7392
rect 34931 7361 34943 7364
rect 34885 7355 34943 7361
rect 30469 7327 30527 7333
rect 30469 7324 30481 7327
rect 22980 7296 26464 7324
rect 28736 7296 30481 7324
rect 22980 7284 22986 7296
rect 9309 7259 9367 7265
rect 9309 7225 9321 7259
rect 9355 7256 9367 7259
rect 17678 7256 17684 7268
rect 9355 7228 17684 7256
rect 9355 7225 9367 7228
rect 9309 7219 9367 7225
rect 17678 7216 17684 7228
rect 17736 7216 17742 7268
rect 26436 7256 26464 7296
rect 30469 7293 30481 7296
rect 30515 7293 30527 7327
rect 33612 7324 33640 7355
rect 35526 7352 35532 7364
rect 35584 7352 35590 7404
rect 35710 7352 35716 7404
rect 35768 7392 35774 7404
rect 35768 7364 37964 7392
rect 35768 7352 35774 7364
rect 37274 7324 37280 7336
rect 33612 7296 37280 7324
rect 30469 7287 30527 7293
rect 37274 7284 37280 7296
rect 37332 7284 37338 7336
rect 37734 7284 37740 7336
rect 37792 7284 37798 7336
rect 37936 7324 37964 7364
rect 38010 7352 38016 7404
rect 38068 7392 38074 7404
rect 39960 7401 39988 7432
rect 40126 7420 40132 7472
rect 40184 7460 40190 7472
rect 40221 7463 40279 7469
rect 40221 7460 40233 7463
rect 40184 7432 40233 7460
rect 40184 7420 40190 7432
rect 40221 7429 40233 7432
rect 40267 7429 40279 7463
rect 40221 7423 40279 7429
rect 40770 7420 40776 7472
rect 40828 7460 40834 7472
rect 43346 7460 43352 7472
rect 40828 7432 43352 7460
rect 40828 7420 40834 7432
rect 43346 7420 43352 7432
rect 43404 7420 43410 7472
rect 43530 7420 43536 7472
rect 43588 7460 43594 7472
rect 44818 7460 44824 7472
rect 43588 7432 44824 7460
rect 43588 7420 43594 7432
rect 44818 7420 44824 7432
rect 44876 7420 44882 7472
rect 44928 7469 44956 7500
rect 45278 7488 45284 7540
rect 45336 7528 45342 7540
rect 45557 7531 45615 7537
rect 45557 7528 45569 7531
rect 45336 7500 45569 7528
rect 45336 7488 45342 7500
rect 45557 7497 45569 7500
rect 45603 7497 45615 7531
rect 45557 7491 45615 7497
rect 46385 7531 46443 7537
rect 46385 7497 46397 7531
rect 46431 7528 46443 7531
rect 50062 7528 50068 7540
rect 46431 7500 50068 7528
rect 46431 7497 46443 7500
rect 46385 7491 46443 7497
rect 50062 7488 50068 7500
rect 50120 7488 50126 7540
rect 44913 7463 44971 7469
rect 44913 7429 44925 7463
rect 44959 7429 44971 7463
rect 44913 7423 44971 7429
rect 45002 7420 45008 7472
rect 45060 7460 45066 7472
rect 47213 7463 47271 7469
rect 47213 7460 47225 7463
rect 45060 7432 47225 7460
rect 45060 7420 45066 7432
rect 47213 7429 47225 7432
rect 47259 7429 47271 7463
rect 47213 7423 47271 7429
rect 49145 7463 49203 7469
rect 49145 7429 49157 7463
rect 49191 7460 49203 7463
rect 49326 7460 49332 7472
rect 49191 7432 49332 7460
rect 49191 7429 49203 7432
rect 49145 7423 49203 7429
rect 49326 7420 49332 7432
rect 49384 7420 49390 7472
rect 38473 7395 38531 7401
rect 38473 7392 38485 7395
rect 38068 7364 38485 7392
rect 38068 7352 38074 7364
rect 38473 7361 38485 7364
rect 38519 7361 38531 7395
rect 39301 7395 39359 7401
rect 39301 7392 39313 7395
rect 38473 7355 38531 7361
rect 38580 7364 39313 7392
rect 38580 7324 38608 7364
rect 39301 7361 39313 7364
rect 39347 7361 39359 7395
rect 39301 7355 39359 7361
rect 39945 7395 40003 7401
rect 39945 7361 39957 7395
rect 39991 7361 40003 7395
rect 39945 7355 40003 7361
rect 42242 7352 42248 7404
rect 42300 7392 42306 7404
rect 43165 7395 43223 7401
rect 43165 7392 43177 7395
rect 42300 7364 43177 7392
rect 42300 7352 42306 7364
rect 43165 7361 43177 7364
rect 43211 7392 43223 7395
rect 43717 7395 43775 7401
rect 43717 7392 43729 7395
rect 43211 7364 43729 7392
rect 43211 7361 43223 7364
rect 43165 7355 43223 7361
rect 43717 7361 43729 7364
rect 43763 7361 43775 7395
rect 43717 7355 43775 7361
rect 44358 7352 44364 7404
rect 44416 7352 44422 7404
rect 45741 7395 45799 7401
rect 45741 7392 45753 7395
rect 44468 7364 45753 7392
rect 37936 7296 38608 7324
rect 38657 7327 38715 7333
rect 38657 7293 38669 7327
rect 38703 7324 38715 7327
rect 40126 7324 40132 7336
rect 38703 7296 40132 7324
rect 38703 7293 38715 7296
rect 38657 7287 38715 7293
rect 40126 7284 40132 7296
rect 40184 7284 40190 7336
rect 42794 7284 42800 7336
rect 42852 7324 42858 7336
rect 44174 7324 44180 7336
rect 42852 7296 43576 7324
rect 42852 7284 42858 7296
rect 35802 7256 35808 7268
rect 26436 7228 35808 7256
rect 35802 7216 35808 7228
rect 35860 7216 35866 7268
rect 43548 7265 43576 7296
rect 43640 7296 44180 7324
rect 39117 7259 39175 7265
rect 39117 7225 39129 7259
rect 39163 7256 39175 7259
rect 43533 7259 43591 7265
rect 39163 7228 43300 7256
rect 39163 7225 39175 7228
rect 39117 7219 39175 7225
rect 1762 7148 1768 7200
rect 1820 7148 1826 7200
rect 18506 7148 18512 7200
rect 18564 7148 18570 7200
rect 21450 7148 21456 7200
rect 21508 7148 21514 7200
rect 21818 7148 21824 7200
rect 21876 7148 21882 7200
rect 23382 7148 23388 7200
rect 23440 7148 23446 7200
rect 24489 7191 24547 7197
rect 24489 7157 24501 7191
rect 24535 7188 24547 7191
rect 24670 7188 24676 7200
rect 24535 7160 24676 7188
rect 24535 7157 24547 7160
rect 24489 7151 24547 7157
rect 24670 7148 24676 7160
rect 24728 7148 24734 7200
rect 25222 7148 25228 7200
rect 25280 7188 25286 7200
rect 25593 7191 25651 7197
rect 25593 7188 25605 7191
rect 25280 7160 25605 7188
rect 25280 7148 25286 7160
rect 25593 7157 25605 7160
rect 25639 7157 25651 7191
rect 25593 7151 25651 7157
rect 34882 7148 34888 7200
rect 34940 7188 34946 7200
rect 35529 7191 35587 7197
rect 35529 7188 35541 7191
rect 34940 7160 35541 7188
rect 34940 7148 34946 7160
rect 35529 7157 35541 7160
rect 35575 7157 35587 7191
rect 35529 7151 35587 7157
rect 42889 7191 42947 7197
rect 42889 7157 42901 7191
rect 42935 7188 42947 7191
rect 42978 7188 42984 7200
rect 42935 7160 42984 7188
rect 42935 7157 42947 7160
rect 42889 7151 42947 7157
rect 42978 7148 42984 7160
rect 43036 7148 43042 7200
rect 43073 7191 43131 7197
rect 43073 7157 43085 7191
rect 43119 7188 43131 7191
rect 43162 7188 43168 7200
rect 43119 7160 43168 7188
rect 43119 7157 43131 7160
rect 43073 7151 43131 7157
rect 43162 7148 43168 7160
rect 43220 7148 43226 7200
rect 43272 7188 43300 7228
rect 43533 7225 43545 7259
rect 43579 7225 43591 7259
rect 43533 7219 43591 7225
rect 43640 7188 43668 7296
rect 44174 7284 44180 7296
rect 44232 7284 44238 7336
rect 44266 7284 44272 7336
rect 44324 7324 44330 7336
rect 44468 7324 44496 7364
rect 45741 7361 45753 7364
rect 45787 7392 45799 7395
rect 45922 7392 45928 7404
rect 45787 7364 45928 7392
rect 45787 7361 45799 7364
rect 45741 7355 45799 7361
rect 45922 7352 45928 7364
rect 45980 7352 45986 7404
rect 46198 7352 46204 7404
rect 46256 7352 46262 7404
rect 46290 7352 46296 7404
rect 46348 7392 46354 7404
rect 47029 7395 47087 7401
rect 47029 7392 47041 7395
rect 46348 7364 47041 7392
rect 46348 7352 46354 7364
rect 47029 7361 47041 7364
rect 47075 7361 47087 7395
rect 47029 7355 47087 7361
rect 47946 7352 47952 7404
rect 48004 7352 48010 7404
rect 44324 7296 44496 7324
rect 44324 7284 44330 7296
rect 44634 7284 44640 7336
rect 44692 7324 44698 7336
rect 46308 7324 46336 7352
rect 44692 7296 46336 7324
rect 44692 7284 44698 7296
rect 47210 7284 47216 7336
rect 47268 7324 47274 7336
rect 47581 7327 47639 7333
rect 47581 7324 47593 7327
rect 47268 7296 47593 7324
rect 47268 7284 47274 7296
rect 47581 7293 47593 7296
rect 47627 7293 47639 7327
rect 47581 7287 47639 7293
rect 50062 7284 50068 7336
rect 50120 7324 50126 7336
rect 50522 7324 50528 7336
rect 50120 7296 50528 7324
rect 50120 7284 50126 7296
rect 50522 7284 50528 7296
rect 50580 7284 50586 7336
rect 45097 7259 45155 7265
rect 45097 7225 45109 7259
rect 45143 7256 45155 7259
rect 47854 7256 47860 7268
rect 45143 7228 47860 7256
rect 45143 7225 45155 7228
rect 45097 7219 45155 7225
rect 47854 7216 47860 7228
rect 47912 7216 47918 7268
rect 43272 7160 43668 7188
rect 44177 7191 44235 7197
rect 44177 7157 44189 7191
rect 44223 7188 44235 7191
rect 44450 7188 44456 7200
rect 44223 7160 44456 7188
rect 44223 7157 44235 7160
rect 44177 7151 44235 7157
rect 44450 7148 44456 7160
rect 44508 7148 44514 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 1762 6944 1768 6996
rect 1820 6984 1826 6996
rect 1820 6956 2774 6984
rect 1820 6944 1826 6956
rect 2746 6916 2774 6956
rect 9490 6944 9496 6996
rect 9548 6944 9554 6996
rect 12710 6944 12716 6996
rect 12768 6984 12774 6996
rect 12805 6987 12863 6993
rect 12805 6984 12817 6987
rect 12768 6956 12817 6984
rect 12768 6944 12774 6956
rect 12805 6953 12817 6956
rect 12851 6953 12863 6987
rect 15102 6984 15108 6996
rect 12805 6947 12863 6953
rect 13556 6956 15108 6984
rect 13556 6916 13584 6956
rect 15102 6944 15108 6956
rect 15160 6944 15166 6996
rect 18414 6944 18420 6996
rect 18472 6984 18478 6996
rect 18601 6987 18659 6993
rect 18601 6984 18613 6987
rect 18472 6956 18613 6984
rect 18472 6944 18478 6956
rect 18601 6953 18613 6956
rect 18647 6953 18659 6987
rect 18601 6947 18659 6953
rect 39298 6944 39304 6996
rect 39356 6984 39362 6996
rect 47946 6984 47952 6996
rect 39356 6956 47952 6984
rect 39356 6944 39362 6956
rect 47946 6944 47952 6956
rect 48004 6944 48010 6996
rect 16390 6916 16396 6928
rect 2746 6888 13584 6916
rect 13648 6888 13860 6916
rect 11057 6851 11115 6857
rect 11057 6817 11069 6851
rect 11103 6848 11115 6851
rect 13648 6848 13676 6888
rect 11103 6820 12434 6848
rect 11103 6817 11115 6820
rect 11057 6811 11115 6817
rect 1210 6740 1216 6792
rect 1268 6780 1274 6792
rect 1581 6783 1639 6789
rect 1581 6780 1593 6783
rect 1268 6752 1593 6780
rect 1268 6740 1274 6752
rect 1581 6749 1593 6752
rect 1627 6749 1639 6783
rect 2501 6783 2559 6789
rect 2501 6780 2513 6783
rect 1581 6743 1639 6749
rect 1780 6752 2513 6780
rect 1302 6672 1308 6724
rect 1360 6712 1366 6724
rect 1780 6712 1808 6752
rect 2501 6749 2513 6752
rect 2547 6780 2559 6783
rect 2777 6783 2835 6789
rect 2777 6780 2789 6783
rect 2547 6752 2789 6780
rect 2547 6749 2559 6752
rect 2501 6743 2559 6749
rect 2777 6749 2789 6752
rect 2823 6749 2835 6783
rect 2777 6743 2835 6749
rect 11330 6740 11336 6792
rect 11388 6740 11394 6792
rect 12406 6780 12434 6820
rect 13372 6820 13676 6848
rect 13372 6780 13400 6820
rect 13722 6808 13728 6860
rect 13780 6808 13786 6860
rect 13832 6848 13860 6888
rect 14384 6888 16396 6916
rect 14384 6848 14412 6888
rect 16390 6876 16396 6888
rect 16448 6876 16454 6928
rect 17589 6919 17647 6925
rect 17589 6885 17601 6919
rect 17635 6885 17647 6919
rect 17589 6879 17647 6885
rect 13832 6820 14412 6848
rect 14476 6820 15424 6848
rect 14476 6785 14504 6820
rect 12406 6752 13400 6780
rect 13464 6752 13676 6780
rect 8754 6712 8760 6724
rect 1360 6684 1808 6712
rect 2332 6684 8760 6712
rect 1360 6672 1366 6684
rect 1762 6604 1768 6656
rect 1820 6604 1826 6656
rect 2332 6653 2360 6684
rect 8754 6672 8760 6684
rect 8812 6672 8818 6724
rect 11790 6672 11796 6724
rect 11848 6712 11854 6724
rect 13464 6712 13492 6752
rect 11848 6684 13492 6712
rect 13541 6715 13599 6721
rect 11848 6672 11854 6684
rect 13541 6681 13553 6715
rect 13587 6681 13599 6715
rect 13648 6712 13676 6752
rect 14461 6779 14519 6785
rect 14461 6745 14473 6779
rect 14507 6745 14519 6779
rect 14461 6739 14519 6745
rect 15286 6740 15292 6792
rect 15344 6740 15350 6792
rect 15396 6780 15424 6820
rect 15562 6808 15568 6860
rect 15620 6848 15626 6860
rect 15933 6851 15991 6857
rect 15933 6848 15945 6851
rect 15620 6820 15945 6848
rect 15620 6808 15626 6820
rect 15933 6817 15945 6820
rect 15979 6817 15991 6851
rect 16850 6848 16856 6860
rect 15933 6811 15991 6817
rect 16040 6820 16856 6848
rect 16040 6780 16068 6820
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 17126 6808 17132 6860
rect 17184 6808 17190 6860
rect 17604 6848 17632 6879
rect 31846 6876 31852 6928
rect 31904 6916 31910 6928
rect 41782 6916 41788 6928
rect 31904 6888 41788 6916
rect 31904 6876 31910 6888
rect 41782 6876 41788 6888
rect 41840 6876 41846 6928
rect 42610 6876 42616 6928
rect 42668 6916 42674 6928
rect 42668 6888 46152 6916
rect 42668 6876 42674 6888
rect 17604 6820 17816 6848
rect 15396 6752 16068 6780
rect 16485 6783 16543 6789
rect 16485 6749 16497 6783
rect 16531 6780 16543 6783
rect 17678 6780 17684 6792
rect 16531 6752 17684 6780
rect 16531 6749 16543 6752
rect 16485 6743 16543 6749
rect 17678 6740 17684 6752
rect 17736 6740 17742 6792
rect 17788 6712 17816 6820
rect 17862 6808 17868 6860
rect 17920 6848 17926 6860
rect 18141 6851 18199 6857
rect 18141 6848 18153 6851
rect 17920 6820 18153 6848
rect 17920 6808 17926 6820
rect 18141 6817 18153 6820
rect 18187 6817 18199 6851
rect 18141 6811 18199 6817
rect 19150 6808 19156 6860
rect 19208 6848 19214 6860
rect 19429 6851 19487 6857
rect 19429 6848 19441 6851
rect 19208 6820 19441 6848
rect 19208 6808 19214 6820
rect 19429 6817 19441 6820
rect 19475 6817 19487 6851
rect 19429 6811 19487 6817
rect 22002 6808 22008 6860
rect 22060 6808 22066 6860
rect 24026 6808 24032 6860
rect 24084 6808 24090 6860
rect 25866 6808 25872 6860
rect 25924 6808 25930 6860
rect 28350 6808 28356 6860
rect 28408 6848 28414 6860
rect 28445 6851 28503 6857
rect 28445 6848 28457 6851
rect 28408 6820 28457 6848
rect 28408 6808 28414 6820
rect 28445 6817 28457 6820
rect 28491 6817 28503 6851
rect 28445 6811 28503 6817
rect 32214 6808 32220 6860
rect 32272 6848 32278 6860
rect 35529 6851 35587 6857
rect 35529 6848 35541 6851
rect 32272 6820 35541 6848
rect 32272 6808 32278 6820
rect 35529 6817 35541 6820
rect 35575 6817 35587 6851
rect 35529 6811 35587 6817
rect 35618 6808 35624 6860
rect 35676 6848 35682 6860
rect 43346 6848 43352 6860
rect 35676 6820 43352 6848
rect 35676 6808 35682 6820
rect 43346 6808 43352 6820
rect 43404 6808 43410 6860
rect 43441 6851 43499 6857
rect 43441 6817 43453 6851
rect 43487 6848 43499 6851
rect 43622 6848 43628 6860
rect 43487 6820 43628 6848
rect 43487 6817 43499 6820
rect 43441 6811 43499 6817
rect 43622 6808 43628 6820
rect 43680 6808 43686 6860
rect 43806 6808 43812 6860
rect 43864 6808 43870 6860
rect 44729 6851 44787 6857
rect 44729 6817 44741 6851
rect 44775 6848 44787 6851
rect 44818 6848 44824 6860
rect 44775 6820 44824 6848
rect 44775 6817 44787 6820
rect 44729 6811 44787 6817
rect 44818 6808 44824 6820
rect 44876 6808 44882 6860
rect 46014 6848 46020 6860
rect 44928 6820 46020 6848
rect 17957 6783 18015 6789
rect 17957 6749 17969 6783
rect 18003 6780 18015 6783
rect 18506 6780 18512 6792
rect 18003 6752 18512 6780
rect 18003 6749 18015 6752
rect 17957 6743 18015 6749
rect 18506 6740 18512 6752
rect 18564 6740 18570 6792
rect 18874 6740 18880 6792
rect 18932 6740 18938 6792
rect 20254 6740 20260 6792
rect 20312 6740 20318 6792
rect 21361 6783 21419 6789
rect 21361 6749 21373 6783
rect 21407 6780 21419 6783
rect 22462 6780 22468 6792
rect 21407 6752 22468 6780
rect 21407 6749 21419 6752
rect 21361 6743 21419 6749
rect 22462 6740 22468 6752
rect 22520 6740 22526 6792
rect 23382 6740 23388 6792
rect 23440 6740 23446 6792
rect 25222 6740 25228 6792
rect 25280 6740 25286 6792
rect 26329 6783 26387 6789
rect 26329 6749 26341 6783
rect 26375 6749 26387 6783
rect 26329 6743 26387 6749
rect 27801 6783 27859 6789
rect 27801 6749 27813 6783
rect 27847 6780 27859 6783
rect 28534 6780 28540 6792
rect 27847 6752 28540 6780
rect 27847 6749 27859 6752
rect 27801 6743 27859 6749
rect 18782 6712 18788 6724
rect 13648 6684 14412 6712
rect 17788 6684 18788 6712
rect 13541 6675 13599 6681
rect 2317 6647 2375 6653
rect 2317 6613 2329 6647
rect 2363 6613 2375 6647
rect 2317 6607 2375 6613
rect 12342 6604 12348 6656
rect 12400 6604 12406 6656
rect 13556 6644 13584 6675
rect 14090 6644 14096 6656
rect 13556 6616 14096 6644
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 14274 6604 14280 6656
rect 14332 6604 14338 6656
rect 14384 6644 14412 6684
rect 18782 6672 18788 6684
rect 18840 6672 18846 6724
rect 19058 6672 19064 6724
rect 19116 6712 19122 6724
rect 20901 6715 20959 6721
rect 20901 6712 20913 6715
rect 19116 6684 20913 6712
rect 19116 6672 19122 6684
rect 20901 6681 20913 6684
rect 20947 6681 20959 6715
rect 20901 6675 20959 6681
rect 21450 6672 21456 6724
rect 21508 6712 21514 6724
rect 26344 6712 26372 6743
rect 28534 6740 28540 6752
rect 28592 6740 28598 6792
rect 29270 6740 29276 6792
rect 29328 6780 29334 6792
rect 29733 6783 29791 6789
rect 29733 6780 29745 6783
rect 29328 6752 29745 6780
rect 29328 6740 29334 6752
rect 29733 6749 29745 6752
rect 29779 6749 29791 6783
rect 29733 6743 29791 6749
rect 30374 6740 30380 6792
rect 30432 6780 30438 6792
rect 30837 6783 30895 6789
rect 30837 6780 30849 6783
rect 30432 6752 30849 6780
rect 30432 6740 30438 6752
rect 30837 6749 30849 6752
rect 30883 6749 30895 6783
rect 30837 6743 30895 6749
rect 32306 6740 32312 6792
rect 32364 6740 32370 6792
rect 33413 6783 33471 6789
rect 33413 6749 33425 6783
rect 33459 6780 33471 6783
rect 33686 6780 33692 6792
rect 33459 6752 33692 6780
rect 33459 6749 33471 6752
rect 33413 6743 33471 6749
rect 33686 6740 33692 6752
rect 33744 6740 33750 6792
rect 34882 6740 34888 6792
rect 34940 6740 34946 6792
rect 43530 6740 43536 6792
rect 43588 6740 43594 6792
rect 43990 6740 43996 6792
rect 44048 6780 44054 6792
rect 44928 6780 44956 6820
rect 46014 6808 46020 6820
rect 46072 6808 46078 6860
rect 44048 6752 44956 6780
rect 44048 6740 44054 6752
rect 45278 6740 45284 6792
rect 45336 6780 45342 6792
rect 45462 6780 45468 6792
rect 45336 6752 45468 6780
rect 45336 6740 45342 6752
rect 45462 6740 45468 6752
rect 45520 6740 45526 6792
rect 45649 6783 45707 6789
rect 45649 6749 45661 6783
rect 45695 6780 45707 6783
rect 45922 6780 45928 6792
rect 45695 6752 45928 6780
rect 45695 6749 45707 6752
rect 45649 6743 45707 6749
rect 45922 6740 45928 6752
rect 45980 6740 45986 6792
rect 46124 6789 46152 6888
rect 46290 6808 46296 6860
rect 46348 6848 46354 6860
rect 46348 6820 48084 6848
rect 46348 6808 46354 6820
rect 46109 6783 46167 6789
rect 46109 6749 46121 6783
rect 46155 6749 46167 6783
rect 46109 6743 46167 6749
rect 47762 6740 47768 6792
rect 47820 6780 47826 6792
rect 47949 6783 48007 6789
rect 47949 6780 47961 6783
rect 47820 6752 47961 6780
rect 47820 6740 47826 6752
rect 47949 6749 47961 6752
rect 47995 6749 48007 6783
rect 48056 6780 48084 6820
rect 49142 6808 49148 6860
rect 49200 6808 49206 6860
rect 50338 6780 50344 6792
rect 48056 6752 50344 6780
rect 47949 6743 48007 6749
rect 50338 6740 50344 6752
rect 50396 6740 50402 6792
rect 21508 6684 26372 6712
rect 21508 6672 21514 6684
rect 30650 6672 30656 6724
rect 30708 6712 30714 6724
rect 32953 6715 33011 6721
rect 32953 6712 32965 6715
rect 30708 6684 32965 6712
rect 30708 6672 30714 6684
rect 32953 6681 32965 6684
rect 32999 6681 33011 6715
rect 32953 6675 33011 6681
rect 34057 6715 34115 6721
rect 34057 6681 34069 6715
rect 34103 6712 34115 6715
rect 36078 6712 36084 6724
rect 34103 6684 36084 6712
rect 34103 6681 34115 6684
rect 34057 6675 34115 6681
rect 36078 6672 36084 6684
rect 36136 6672 36142 6724
rect 37182 6672 37188 6724
rect 37240 6712 37246 6724
rect 44177 6715 44235 6721
rect 44177 6712 44189 6715
rect 37240 6684 44189 6712
rect 37240 6672 37246 6684
rect 44177 6681 44189 6684
rect 44223 6681 44235 6715
rect 44177 6675 44235 6681
rect 44361 6715 44419 6721
rect 44361 6681 44373 6715
rect 44407 6712 44419 6715
rect 47118 6712 47124 6724
rect 44407 6684 47124 6712
rect 44407 6681 44419 6684
rect 44361 6675 44419 6681
rect 47118 6672 47124 6684
rect 47176 6672 47182 6724
rect 47305 6715 47363 6721
rect 47305 6681 47317 6715
rect 47351 6712 47363 6715
rect 48682 6712 48688 6724
rect 47351 6684 48688 6712
rect 47351 6681 47363 6684
rect 47305 6675 47363 6681
rect 48682 6672 48688 6684
rect 48740 6672 48746 6724
rect 14550 6644 14556 6656
rect 14384 6616 14556 6644
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 14642 6604 14648 6656
rect 14700 6644 14706 6656
rect 18049 6647 18107 6653
rect 18049 6644 18061 6647
rect 14700 6616 18061 6644
rect 14700 6604 14706 6616
rect 18049 6613 18061 6616
rect 18095 6613 18107 6647
rect 18049 6607 18107 6613
rect 18322 6604 18328 6656
rect 18380 6644 18386 6656
rect 18969 6647 19027 6653
rect 18969 6644 18981 6647
rect 18380 6616 18981 6644
rect 18380 6604 18386 6616
rect 18969 6613 18981 6616
rect 19015 6613 19027 6647
rect 18969 6607 19027 6613
rect 26970 6604 26976 6656
rect 27028 6604 27034 6656
rect 30282 6604 30288 6656
rect 30340 6644 30346 6656
rect 30377 6647 30435 6653
rect 30377 6644 30389 6647
rect 30340 6616 30389 6644
rect 30340 6604 30346 6616
rect 30377 6613 30389 6616
rect 30423 6613 30435 6647
rect 30377 6607 30435 6613
rect 30466 6604 30472 6656
rect 30524 6644 30530 6656
rect 31481 6647 31539 6653
rect 31481 6644 31493 6647
rect 30524 6616 31493 6644
rect 30524 6604 30530 6616
rect 31481 6613 31493 6616
rect 31527 6613 31539 6647
rect 31481 6607 31539 6613
rect 40310 6604 40316 6656
rect 40368 6644 40374 6656
rect 43254 6644 43260 6656
rect 40368 6616 43260 6644
rect 40368 6604 40374 6616
rect 43254 6604 43260 6616
rect 43312 6604 43318 6656
rect 45002 6604 45008 6656
rect 45060 6604 45066 6656
rect 45462 6604 45468 6656
rect 45520 6604 45526 6656
rect 46014 6604 46020 6656
rect 46072 6644 46078 6656
rect 46842 6644 46848 6656
rect 46072 6616 46848 6644
rect 46072 6604 46078 6616
rect 46842 6604 46848 6616
rect 46900 6604 46906 6656
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 1210 6400 1216 6452
rect 1268 6440 1274 6452
rect 2133 6443 2191 6449
rect 2133 6440 2145 6443
rect 1268 6412 2145 6440
rect 1268 6400 1274 6412
rect 2133 6409 2145 6412
rect 2179 6409 2191 6443
rect 2133 6403 2191 6409
rect 9858 6400 9864 6452
rect 9916 6440 9922 6452
rect 16301 6443 16359 6449
rect 9916 6412 14504 6440
rect 9916 6400 9922 6412
rect 12618 6332 12624 6384
rect 12676 6372 12682 6384
rect 13541 6375 13599 6381
rect 13541 6372 13553 6375
rect 12676 6344 13553 6372
rect 12676 6332 12682 6344
rect 13541 6341 13553 6344
rect 13587 6341 13599 6375
rect 13541 6335 13599 6341
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 14476 6313 14504 6412
rect 16301 6409 16313 6443
rect 16347 6440 16359 6443
rect 16574 6440 16580 6452
rect 16347 6412 16580 6440
rect 16347 6409 16359 6412
rect 16301 6403 16359 6409
rect 16574 6400 16580 6412
rect 16632 6400 16638 6452
rect 17586 6400 17592 6452
rect 17644 6440 17650 6452
rect 18141 6443 18199 6449
rect 18141 6440 18153 6443
rect 17644 6412 18153 6440
rect 17644 6400 17650 6412
rect 18141 6409 18153 6412
rect 18187 6409 18199 6443
rect 18141 6403 18199 6409
rect 19245 6443 19303 6449
rect 19245 6409 19257 6443
rect 19291 6440 19303 6443
rect 19334 6440 19340 6452
rect 19291 6412 19340 6440
rect 19291 6409 19303 6412
rect 19245 6403 19303 6409
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 19702 6400 19708 6452
rect 19760 6440 19766 6452
rect 20349 6443 20407 6449
rect 20349 6440 20361 6443
rect 19760 6412 20361 6440
rect 19760 6400 19766 6412
rect 20349 6409 20361 6412
rect 20395 6409 20407 6443
rect 20349 6403 20407 6409
rect 21910 6400 21916 6452
rect 21968 6440 21974 6452
rect 22649 6443 22707 6449
rect 22649 6440 22661 6443
rect 21968 6412 22661 6440
rect 21968 6400 21974 6412
rect 22649 6409 22661 6412
rect 22695 6409 22707 6443
rect 22649 6403 22707 6409
rect 24210 6400 24216 6452
rect 24268 6400 24274 6452
rect 24946 6400 24952 6452
rect 25004 6440 25010 6452
rect 25317 6443 25375 6449
rect 25317 6440 25329 6443
rect 25004 6412 25329 6440
rect 25004 6400 25010 6412
rect 25317 6409 25329 6412
rect 25363 6409 25375 6443
rect 25317 6403 25375 6409
rect 29270 6400 29276 6452
rect 29328 6400 29334 6452
rect 30469 6443 30527 6449
rect 30469 6409 30481 6443
rect 30515 6440 30527 6443
rect 30558 6440 30564 6452
rect 30515 6412 30564 6440
rect 30515 6409 30527 6412
rect 30469 6403 30527 6409
rect 30558 6400 30564 6412
rect 30616 6400 30622 6452
rect 30834 6400 30840 6452
rect 30892 6440 30898 6452
rect 31573 6443 31631 6449
rect 31573 6440 31585 6443
rect 30892 6412 31585 6440
rect 30892 6400 30898 6412
rect 31573 6409 31585 6412
rect 31619 6409 31631 6443
rect 31573 6403 31631 6409
rect 32306 6400 32312 6452
rect 32364 6440 32370 6452
rect 32953 6443 33011 6449
rect 32953 6440 32965 6443
rect 32364 6412 32965 6440
rect 32364 6400 32370 6412
rect 32953 6409 32965 6412
rect 32999 6409 33011 6443
rect 32953 6403 33011 6409
rect 33413 6443 33471 6449
rect 33413 6409 33425 6443
rect 33459 6440 33471 6443
rect 33502 6440 33508 6452
rect 33459 6412 33508 6440
rect 33459 6409 33471 6412
rect 33413 6403 33471 6409
rect 33502 6400 33508 6412
rect 33560 6400 33566 6452
rect 43990 6400 43996 6452
rect 44048 6400 44054 6452
rect 44177 6443 44235 6449
rect 44177 6409 44189 6443
rect 44223 6440 44235 6443
rect 44266 6440 44272 6452
rect 44223 6412 44272 6440
rect 44223 6409 44235 6412
rect 44177 6403 44235 6409
rect 44266 6400 44272 6412
rect 44324 6400 44330 6452
rect 44358 6400 44364 6452
rect 44416 6400 44422 6452
rect 44450 6400 44456 6452
rect 44508 6440 44514 6452
rect 44637 6443 44695 6449
rect 44637 6440 44649 6443
rect 44508 6412 44649 6440
rect 44508 6400 44514 6412
rect 44637 6409 44649 6412
rect 44683 6409 44695 6443
rect 44637 6403 44695 6409
rect 45097 6443 45155 6449
rect 45097 6409 45109 6443
rect 45143 6440 45155 6443
rect 45646 6440 45652 6452
rect 45143 6412 45652 6440
rect 45143 6409 45155 6412
rect 45097 6403 45155 6409
rect 45646 6400 45652 6412
rect 45704 6400 45710 6452
rect 46014 6400 46020 6452
rect 46072 6400 46078 6452
rect 47210 6400 47216 6452
rect 47268 6400 47274 6452
rect 47397 6443 47455 6449
rect 47397 6409 47409 6443
rect 47443 6440 47455 6443
rect 50890 6440 50896 6452
rect 47443 6412 50896 6440
rect 47443 6409 47455 6412
rect 47397 6403 47455 6409
rect 50890 6400 50896 6412
rect 50948 6400 50954 6452
rect 14918 6332 14924 6384
rect 14976 6372 14982 6384
rect 14976 6344 15792 6372
rect 14976 6332 14982 6344
rect 1581 6307 1639 6313
rect 1581 6304 1593 6307
rect 1360 6276 1593 6304
rect 1360 6264 1366 6276
rect 1581 6273 1593 6276
rect 1627 6304 1639 6307
rect 2317 6307 2375 6313
rect 2317 6304 2329 6307
rect 1627 6276 2329 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 2317 6273 2329 6276
rect 2363 6273 2375 6307
rect 2317 6267 2375 6273
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6273 11851 6307
rect 11793 6267 11851 6273
rect 14461 6307 14519 6313
rect 14461 6273 14473 6307
rect 14507 6273 14519 6307
rect 14461 6267 14519 6273
rect 11808 6236 11836 6267
rect 14550 6264 14556 6316
rect 14608 6304 14614 6316
rect 15197 6307 15255 6313
rect 15197 6304 15209 6307
rect 14608 6276 15209 6304
rect 14608 6264 14614 6276
rect 15197 6273 15209 6276
rect 15243 6273 15255 6307
rect 15197 6267 15255 6273
rect 15657 6307 15715 6313
rect 15657 6273 15669 6307
rect 15703 6273 15715 6307
rect 15657 6267 15715 6273
rect 12342 6236 12348 6248
rect 11808 6208 12348 6236
rect 12342 6196 12348 6208
rect 12400 6196 12406 6248
rect 13630 6196 13636 6248
rect 13688 6236 13694 6248
rect 15672 6236 15700 6267
rect 13688 6208 15700 6236
rect 15764 6236 15792 6344
rect 16482 6332 16488 6384
rect 16540 6372 16546 6384
rect 26970 6372 26976 6384
rect 16540 6344 19748 6372
rect 16540 6332 16546 6344
rect 15930 6264 15936 6316
rect 15988 6304 15994 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 15988 6276 16865 6304
rect 15988 6264 15994 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 17497 6307 17555 6313
rect 17497 6273 17509 6307
rect 17543 6304 17555 6307
rect 18506 6304 18512 6316
rect 17543 6276 18512 6304
rect 17543 6273 17555 6276
rect 17497 6267 17555 6273
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 18601 6307 18659 6313
rect 18601 6273 18613 6307
rect 18647 6304 18659 6307
rect 18874 6304 18880 6316
rect 18647 6276 18880 6304
rect 18647 6273 18659 6276
rect 18601 6267 18659 6273
rect 18874 6264 18880 6276
rect 18932 6264 18938 6316
rect 19720 6313 19748 6344
rect 23584 6344 26976 6372
rect 19705 6307 19763 6313
rect 19705 6273 19717 6307
rect 19751 6273 19763 6307
rect 19705 6267 19763 6273
rect 20809 6307 20867 6313
rect 20809 6273 20821 6307
rect 20855 6304 20867 6307
rect 20990 6304 20996 6316
rect 20855 6276 20996 6304
rect 20855 6273 20867 6276
rect 20809 6267 20867 6273
rect 20990 6264 20996 6276
rect 21048 6264 21054 6316
rect 23584 6313 23612 6344
rect 26970 6332 26976 6344
rect 27028 6332 27034 6384
rect 32858 6372 32864 6384
rect 31726 6344 32864 6372
rect 21453 6307 21511 6313
rect 21453 6273 21465 6307
rect 21499 6304 21511 6307
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21499 6276 22017 6304
rect 21499 6273 21511 6276
rect 21453 6267 21511 6273
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 23569 6307 23627 6313
rect 23569 6273 23581 6307
rect 23615 6273 23627 6307
rect 23569 6267 23627 6273
rect 24670 6264 24676 6316
rect 24728 6264 24734 6316
rect 28629 6307 28687 6313
rect 28629 6273 28641 6307
rect 28675 6304 28687 6307
rect 28902 6304 28908 6316
rect 28675 6276 28908 6304
rect 28675 6273 28687 6276
rect 28629 6267 28687 6273
rect 28902 6264 28908 6276
rect 28960 6264 28966 6316
rect 29825 6307 29883 6313
rect 29825 6273 29837 6307
rect 29871 6304 29883 6307
rect 30466 6304 30472 6316
rect 29871 6276 30472 6304
rect 29871 6273 29883 6276
rect 29825 6267 29883 6273
rect 30466 6264 30472 6276
rect 30524 6264 30530 6316
rect 30929 6307 30987 6313
rect 30929 6273 30941 6307
rect 30975 6304 30987 6307
rect 31726 6304 31754 6344
rect 32858 6332 32864 6344
rect 32916 6332 32922 6384
rect 34330 6332 34336 6384
rect 34388 6372 34394 6384
rect 38197 6375 38255 6381
rect 38197 6372 38209 6375
rect 34388 6344 38209 6372
rect 34388 6332 34394 6344
rect 38197 6341 38209 6344
rect 38243 6372 38255 6375
rect 38657 6375 38715 6381
rect 38657 6372 38669 6375
rect 38243 6344 38669 6372
rect 38243 6341 38255 6344
rect 38197 6335 38255 6341
rect 38657 6341 38669 6344
rect 38703 6341 38715 6375
rect 38657 6335 38715 6341
rect 43254 6332 43260 6384
rect 43312 6372 43318 6384
rect 49145 6375 49203 6381
rect 43312 6344 47992 6372
rect 43312 6332 43318 6344
rect 30975 6276 31754 6304
rect 30975 6273 30987 6276
rect 30929 6267 30987 6273
rect 32030 6264 32036 6316
rect 32088 6304 32094 6316
rect 32309 6307 32367 6313
rect 32309 6304 32321 6307
rect 32088 6276 32321 6304
rect 32088 6264 32094 6276
rect 32309 6273 32321 6276
rect 32355 6273 32367 6307
rect 32309 6267 32367 6273
rect 40034 6264 40040 6316
rect 40092 6304 40098 6316
rect 44453 6307 44511 6313
rect 44453 6304 44465 6307
rect 40092 6276 44465 6304
rect 40092 6264 40098 6276
rect 44453 6273 44465 6276
rect 44499 6273 44511 6307
rect 44453 6267 44511 6273
rect 45462 6264 45468 6316
rect 45520 6308 45526 6316
rect 45557 6308 45615 6313
rect 45520 6307 45615 6308
rect 45520 6280 45569 6307
rect 45520 6264 45526 6280
rect 45557 6273 45569 6280
rect 45603 6273 45615 6307
rect 45557 6267 45615 6273
rect 46201 6307 46259 6313
rect 46201 6273 46213 6307
rect 46247 6304 46259 6307
rect 46290 6304 46296 6316
rect 46247 6276 46296 6304
rect 46247 6273 46259 6276
rect 46201 6267 46259 6273
rect 46290 6264 46296 6276
rect 46348 6264 46354 6316
rect 46842 6264 46848 6316
rect 46900 6264 46906 6316
rect 47670 6264 47676 6316
rect 47728 6264 47734 6316
rect 47964 6313 47992 6344
rect 49145 6341 49157 6375
rect 49191 6372 49203 6375
rect 49234 6372 49240 6384
rect 49191 6344 49240 6372
rect 49191 6341 49203 6344
rect 49145 6335 49203 6341
rect 49234 6332 49240 6344
rect 49292 6332 49298 6384
rect 47949 6307 48007 6313
rect 47949 6273 47961 6307
rect 47995 6273 48007 6307
rect 47949 6267 48007 6273
rect 20898 6236 20904 6248
rect 15764 6208 20904 6236
rect 13688 6196 13694 6208
rect 20898 6196 20904 6208
rect 20956 6196 20962 6248
rect 29086 6196 29092 6248
rect 29144 6236 29150 6248
rect 29144 6208 33364 6236
rect 29144 6196 29150 6208
rect 1765 6171 1823 6177
rect 1765 6137 1777 6171
rect 1811 6168 1823 6171
rect 9306 6168 9312 6180
rect 1811 6140 9312 6168
rect 1811 6137 1823 6140
rect 1765 6131 1823 6137
rect 9306 6128 9312 6140
rect 9364 6128 9370 6180
rect 11977 6171 12035 6177
rect 11977 6137 11989 6171
rect 12023 6168 12035 6171
rect 14277 6171 14335 6177
rect 12023 6140 12434 6168
rect 12023 6137 12035 6140
rect 11977 6131 12035 6137
rect 12406 6100 12434 6140
rect 14277 6137 14289 6171
rect 14323 6168 14335 6171
rect 17770 6168 17776 6180
rect 14323 6140 17776 6168
rect 14323 6137 14335 6140
rect 14277 6131 14335 6137
rect 17770 6128 17776 6140
rect 17828 6128 17834 6180
rect 33336 6168 33364 6208
rect 38378 6196 38384 6248
rect 38436 6196 38442 6248
rect 46934 6236 46940 6248
rect 41386 6208 46940 6236
rect 41386 6168 41414 6208
rect 46934 6196 46940 6208
rect 46992 6196 46998 6248
rect 33336 6140 41414 6168
rect 42518 6128 42524 6180
rect 42576 6168 42582 6180
rect 46382 6168 46388 6180
rect 42576 6140 46388 6168
rect 42576 6128 42582 6140
rect 46382 6128 46388 6140
rect 46440 6128 46446 6180
rect 46658 6128 46664 6180
rect 46716 6128 46722 6180
rect 14918 6100 14924 6112
rect 12406 6072 14924 6100
rect 14918 6060 14924 6072
rect 14976 6060 14982 6112
rect 15013 6103 15071 6109
rect 15013 6069 15025 6103
rect 15059 6100 15071 6103
rect 19610 6100 19616 6112
rect 15059 6072 19616 6100
rect 15059 6069 15071 6072
rect 15013 6063 15071 6069
rect 19610 6060 19616 6072
rect 19668 6060 19674 6112
rect 19702 6060 19708 6112
rect 19760 6100 19766 6112
rect 25314 6100 25320 6112
rect 19760 6072 25320 6100
rect 19760 6060 19766 6072
rect 25314 6060 25320 6072
rect 25372 6060 25378 6112
rect 27522 6060 27528 6112
rect 27580 6100 27586 6112
rect 41874 6100 41880 6112
rect 27580 6072 41880 6100
rect 27580 6060 27586 6072
rect 41874 6060 41880 6072
rect 41932 6060 41938 6112
rect 44913 6103 44971 6109
rect 44913 6069 44925 6103
rect 44959 6100 44971 6103
rect 45094 6100 45100 6112
rect 44959 6072 45100 6100
rect 44959 6069 44971 6072
rect 44913 6063 44971 6069
rect 45094 6060 45100 6072
rect 45152 6060 45158 6112
rect 45278 6060 45284 6112
rect 45336 6100 45342 6112
rect 45373 6103 45431 6109
rect 45373 6100 45385 6103
rect 45336 6072 45385 6100
rect 45336 6060 45342 6072
rect 45373 6069 45385 6072
rect 45419 6069 45431 6103
rect 45373 6063 45431 6069
rect 45462 6060 45468 6112
rect 45520 6100 45526 6112
rect 50246 6100 50252 6112
rect 45520 6072 50252 6100
rect 45520 6060 45526 6072
rect 50246 6060 50252 6072
rect 50304 6060 50310 6112
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 1762 5856 1768 5908
rect 1820 5896 1826 5908
rect 1820 5868 15884 5896
rect 1820 5856 1826 5868
rect 2501 5831 2559 5837
rect 2501 5797 2513 5831
rect 2547 5828 2559 5831
rect 13998 5828 14004 5840
rect 2547 5800 14004 5828
rect 2547 5797 2559 5800
rect 2501 5791 2559 5797
rect 13998 5788 14004 5800
rect 14056 5788 14062 5840
rect 15856 5828 15884 5868
rect 18874 5856 18880 5908
rect 18932 5856 18938 5908
rect 20990 5856 20996 5908
rect 21048 5856 21054 5908
rect 23474 5856 23480 5908
rect 23532 5896 23538 5908
rect 24029 5899 24087 5905
rect 24029 5896 24041 5899
rect 23532 5868 24041 5896
rect 23532 5856 23538 5868
rect 24029 5865 24041 5868
rect 24075 5865 24087 5899
rect 24029 5859 24087 5865
rect 30374 5856 30380 5908
rect 30432 5856 30438 5908
rect 30742 5856 30748 5908
rect 30800 5896 30806 5908
rect 32953 5899 33011 5905
rect 32953 5896 32965 5899
rect 30800 5868 32965 5896
rect 30800 5856 30806 5868
rect 32953 5865 32965 5868
rect 32999 5865 33011 5899
rect 32953 5859 33011 5865
rect 44634 5856 44640 5908
rect 44692 5856 44698 5908
rect 45186 5856 45192 5908
rect 45244 5856 45250 5908
rect 45370 5856 45376 5908
rect 45428 5856 45434 5908
rect 45554 5856 45560 5908
rect 45612 5896 45618 5908
rect 46017 5899 46075 5905
rect 46017 5896 46029 5899
rect 45612 5868 46029 5896
rect 45612 5856 45618 5868
rect 46017 5865 46029 5868
rect 46063 5865 46075 5899
rect 46385 5899 46443 5905
rect 46385 5896 46397 5899
rect 46017 5859 46075 5865
rect 46124 5868 46397 5896
rect 29546 5828 29552 5840
rect 15856 5800 29552 5828
rect 29546 5788 29552 5800
rect 29604 5788 29610 5840
rect 44821 5831 44879 5837
rect 44821 5797 44833 5831
rect 44867 5828 44879 5831
rect 45462 5828 45468 5840
rect 44867 5800 45468 5828
rect 44867 5797 44879 5800
rect 44821 5791 44879 5797
rect 45462 5788 45468 5800
rect 45520 5788 45526 5840
rect 45738 5788 45744 5840
rect 45796 5788 45802 5840
rect 3053 5763 3111 5769
rect 3053 5760 3065 5763
rect 1596 5732 3065 5760
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 1596 5701 1624 5732
rect 3053 5729 3065 5732
rect 3099 5729 3111 5763
rect 3053 5723 3111 5729
rect 15838 5720 15844 5772
rect 15896 5720 15902 5772
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5760 16543 5763
rect 17310 5760 17316 5772
rect 16531 5732 17316 5760
rect 16531 5729 16543 5732
rect 16485 5723 16543 5729
rect 17310 5720 17316 5732
rect 17368 5720 17374 5772
rect 18966 5720 18972 5772
rect 19024 5760 19030 5772
rect 19429 5763 19487 5769
rect 19429 5760 19441 5763
rect 19024 5732 19441 5760
rect 19024 5720 19030 5732
rect 19429 5729 19441 5732
rect 19475 5729 19487 5763
rect 19429 5723 19487 5729
rect 20530 5720 20536 5772
rect 20588 5760 20594 5772
rect 25225 5763 25283 5769
rect 25225 5760 25237 5763
rect 20588 5732 25237 5760
rect 20588 5720 20594 5732
rect 25225 5729 25237 5732
rect 25271 5729 25283 5763
rect 25225 5723 25283 5729
rect 31386 5720 31392 5772
rect 31444 5760 31450 5772
rect 31665 5763 31723 5769
rect 31665 5760 31677 5763
rect 31444 5732 31677 5760
rect 31444 5720 31450 5732
rect 31665 5729 31677 5732
rect 31711 5729 31723 5763
rect 31665 5723 31723 5729
rect 38378 5720 38384 5772
rect 38436 5760 38442 5772
rect 45922 5760 45928 5772
rect 38436 5732 45928 5760
rect 38436 5720 38442 5732
rect 45922 5720 45928 5732
rect 45980 5720 45986 5772
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1360 5664 1593 5692
rect 1360 5652 1366 5664
rect 1581 5661 1593 5664
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5692 2375 5695
rect 2774 5692 2780 5704
rect 2363 5664 2780 5692
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 2774 5652 2780 5664
rect 2832 5692 2838 5704
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 2832 5664 2881 5692
rect 2832 5652 2838 5664
rect 2869 5661 2881 5664
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 17129 5695 17187 5701
rect 17129 5661 17141 5695
rect 17175 5692 17187 5695
rect 17862 5692 17868 5704
rect 17175 5664 17868 5692
rect 17175 5661 17187 5664
rect 17129 5655 17187 5661
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5692 18291 5695
rect 20162 5692 20168 5704
rect 18279 5664 20168 5692
rect 18279 5661 18291 5664
rect 18233 5655 18291 5661
rect 20162 5652 20168 5664
rect 20220 5652 20226 5704
rect 20349 5695 20407 5701
rect 20349 5661 20361 5695
rect 20395 5692 20407 5695
rect 20622 5692 20628 5704
rect 20395 5664 20628 5692
rect 20395 5661 20407 5664
rect 20349 5655 20407 5661
rect 20622 5652 20628 5664
rect 20680 5652 20686 5704
rect 21634 5652 21640 5704
rect 21692 5701 21698 5704
rect 21692 5695 21730 5701
rect 21718 5661 21730 5695
rect 21692 5655 21730 5661
rect 21692 5652 21698 5655
rect 22278 5652 22284 5704
rect 22336 5652 22342 5704
rect 23385 5695 23443 5701
rect 23385 5661 23397 5695
rect 23431 5692 23443 5695
rect 23566 5692 23572 5704
rect 23431 5664 23572 5692
rect 23431 5661 23443 5664
rect 23385 5655 23443 5661
rect 23566 5652 23572 5664
rect 23624 5652 23630 5704
rect 23658 5652 23664 5704
rect 23716 5692 23722 5704
rect 24581 5695 24639 5701
rect 24581 5692 24593 5695
rect 23716 5664 24593 5692
rect 23716 5652 23722 5664
rect 24581 5661 24593 5664
rect 24627 5661 24639 5695
rect 24581 5655 24639 5661
rect 29733 5695 29791 5701
rect 29733 5661 29745 5695
rect 29779 5692 29791 5695
rect 31294 5692 31300 5704
rect 29779 5664 31300 5692
rect 29779 5661 29791 5664
rect 29733 5655 29791 5661
rect 31294 5652 31300 5664
rect 31352 5652 31358 5704
rect 32309 5695 32367 5701
rect 32309 5661 32321 5695
rect 32355 5692 32367 5695
rect 36446 5692 36452 5704
rect 32355 5664 36452 5692
rect 32355 5661 32367 5664
rect 32309 5655 32367 5661
rect 36446 5652 36452 5664
rect 36504 5652 36510 5704
rect 38286 5652 38292 5704
rect 38344 5692 38350 5704
rect 43717 5695 43775 5701
rect 43717 5692 43729 5695
rect 38344 5664 43729 5692
rect 38344 5652 38350 5664
rect 43717 5661 43729 5664
rect 43763 5661 43775 5695
rect 46124 5692 46152 5868
rect 46385 5865 46397 5868
rect 46431 5865 46443 5899
rect 46385 5859 46443 5865
rect 47026 5856 47032 5908
rect 47084 5856 47090 5908
rect 47210 5856 47216 5908
rect 47268 5896 47274 5908
rect 47305 5899 47363 5905
rect 47305 5896 47317 5899
rect 47268 5868 47317 5896
rect 47268 5856 47274 5868
rect 47305 5865 47317 5868
rect 47351 5865 47363 5899
rect 50154 5896 50160 5908
rect 47305 5859 47363 5865
rect 47412 5868 50160 5896
rect 46566 5788 46572 5840
rect 46624 5828 46630 5840
rect 47412 5828 47440 5868
rect 50154 5856 50160 5868
rect 50212 5856 50218 5908
rect 50430 5828 50436 5840
rect 46624 5800 47440 5828
rect 47596 5800 50436 5828
rect 46624 5788 46630 5800
rect 47596 5760 47624 5800
rect 50430 5788 50436 5800
rect 50488 5788 50494 5840
rect 43717 5655 43775 5661
rect 43824 5664 46152 5692
rect 46308 5732 47624 5760
rect 49145 5763 49203 5769
rect 21775 5627 21833 5633
rect 1780 5596 12434 5624
rect 1780 5565 1808 5596
rect 1765 5559 1823 5565
rect 1765 5525 1777 5559
rect 1811 5525 1823 5559
rect 12406 5556 12434 5596
rect 21775 5593 21787 5627
rect 21821 5624 21833 5627
rect 23842 5624 23848 5636
rect 21821 5596 23848 5624
rect 21821 5593 21833 5596
rect 21775 5587 21833 5593
rect 23842 5584 23848 5596
rect 23900 5584 23906 5636
rect 41506 5584 41512 5636
rect 41564 5624 41570 5636
rect 43824 5624 43852 5664
rect 41564 5596 43852 5624
rect 43901 5627 43959 5633
rect 41564 5584 41570 5596
rect 43901 5593 43913 5627
rect 43947 5624 43959 5627
rect 45738 5624 45744 5636
rect 43947 5596 45744 5624
rect 43947 5593 43959 5596
rect 43901 5587 43959 5593
rect 45738 5584 45744 5596
rect 45796 5584 45802 5636
rect 45925 5627 45983 5633
rect 45925 5593 45937 5627
rect 45971 5624 45983 5627
rect 46308 5624 46336 5732
rect 49145 5729 49157 5763
rect 49191 5760 49203 5763
rect 49326 5760 49332 5772
rect 49191 5732 49332 5760
rect 49191 5729 49203 5732
rect 49145 5723 49203 5729
rect 49326 5720 49332 5732
rect 49384 5720 49390 5772
rect 46566 5652 46572 5704
rect 46624 5652 46630 5704
rect 46934 5652 46940 5704
rect 46992 5692 46998 5704
rect 47489 5695 47547 5701
rect 47489 5692 47501 5695
rect 46992 5664 47501 5692
rect 46992 5652 46998 5664
rect 47489 5661 47501 5664
rect 47535 5661 47547 5695
rect 47489 5655 47547 5661
rect 47949 5695 48007 5701
rect 47949 5661 47961 5695
rect 47995 5661 48007 5695
rect 47949 5655 48007 5661
rect 45971 5596 46336 5624
rect 45971 5593 45983 5596
rect 45925 5587 45983 5593
rect 46382 5584 46388 5636
rect 46440 5624 46446 5636
rect 47964 5624 47992 5655
rect 46440 5596 47992 5624
rect 46440 5584 46446 5596
rect 13814 5556 13820 5568
rect 12406 5528 13820 5556
rect 1765 5519 1823 5525
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 17773 5559 17831 5565
rect 17773 5525 17785 5559
rect 17819 5556 17831 5559
rect 18414 5556 18420 5568
rect 17819 5528 18420 5556
rect 17819 5525 17831 5528
rect 17773 5519 17831 5525
rect 18414 5516 18420 5528
rect 18472 5516 18478 5568
rect 18506 5516 18512 5568
rect 18564 5556 18570 5568
rect 22370 5556 22376 5568
rect 18564 5528 22376 5556
rect 18564 5516 18570 5528
rect 22370 5516 22376 5528
rect 22428 5516 22434 5568
rect 22922 5516 22928 5568
rect 22980 5516 22986 5568
rect 45557 5559 45615 5565
rect 45557 5525 45569 5559
rect 45603 5556 45615 5559
rect 48314 5556 48320 5568
rect 45603 5528 48320 5556
rect 45603 5525 45615 5528
rect 45557 5519 45615 5525
rect 48314 5516 48320 5528
rect 48372 5516 48378 5568
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 12158 5312 12164 5364
rect 12216 5352 12222 5364
rect 20165 5355 20223 5361
rect 20165 5352 20177 5355
rect 12216 5324 20177 5352
rect 12216 5312 12222 5324
rect 20165 5321 20177 5324
rect 20211 5321 20223 5355
rect 20165 5315 20223 5321
rect 23566 5312 23572 5364
rect 23624 5312 23630 5364
rect 31478 5312 31484 5364
rect 31536 5352 31542 5364
rect 32309 5355 32367 5361
rect 32309 5352 32321 5355
rect 31536 5324 32321 5352
rect 31536 5312 31542 5324
rect 32309 5321 32321 5324
rect 32355 5321 32367 5355
rect 37642 5352 37648 5364
rect 32309 5315 32367 5321
rect 32600 5324 37648 5352
rect 15010 5244 15016 5296
rect 15068 5284 15074 5296
rect 15068 5256 17632 5284
rect 15068 5244 15074 5256
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5216 1915 5219
rect 8938 5216 8944 5228
rect 1903 5188 8944 5216
rect 1903 5185 1915 5188
rect 1857 5179 1915 5185
rect 8938 5176 8944 5188
rect 8996 5176 9002 5228
rect 16945 5219 17003 5225
rect 16945 5185 16957 5219
rect 16991 5216 17003 5219
rect 17604 5216 17632 5256
rect 17678 5244 17684 5296
rect 17736 5284 17742 5296
rect 19061 5287 19119 5293
rect 19061 5284 19073 5287
rect 17736 5256 19073 5284
rect 17736 5244 17742 5256
rect 19061 5253 19073 5256
rect 19107 5253 19119 5287
rect 19061 5247 19119 5253
rect 26142 5244 26148 5296
rect 26200 5284 26206 5296
rect 32600 5284 32628 5324
rect 37642 5312 37648 5324
rect 37700 5312 37706 5364
rect 45554 5312 45560 5364
rect 45612 5312 45618 5364
rect 45830 5312 45836 5364
rect 45888 5352 45894 5364
rect 46934 5352 46940 5364
rect 45888 5324 46940 5352
rect 45888 5312 45894 5324
rect 46934 5312 46940 5324
rect 46992 5312 46998 5364
rect 47673 5355 47731 5361
rect 47673 5321 47685 5355
rect 47719 5352 47731 5355
rect 49694 5352 49700 5364
rect 47719 5324 49700 5352
rect 47719 5321 47731 5324
rect 47673 5315 47731 5321
rect 49694 5312 49700 5324
rect 49752 5312 49758 5364
rect 26200 5256 32628 5284
rect 26200 5244 26206 5256
rect 32674 5244 32680 5296
rect 32732 5284 32738 5296
rect 39301 5287 39359 5293
rect 39301 5284 39313 5287
rect 32732 5256 39313 5284
rect 32732 5244 32738 5256
rect 39301 5253 39313 5256
rect 39347 5284 39359 5287
rect 39761 5287 39819 5293
rect 39761 5284 39773 5287
rect 39347 5256 39773 5284
rect 39347 5253 39359 5256
rect 39301 5247 39359 5253
rect 39761 5253 39773 5256
rect 39807 5253 39819 5287
rect 39761 5247 39819 5253
rect 49142 5244 49148 5296
rect 49200 5244 49206 5296
rect 17957 5219 18015 5225
rect 17957 5216 17969 5219
rect 16991 5188 17540 5216
rect 17604 5188 17969 5216
rect 16991 5185 17003 5188
rect 16945 5179 17003 5185
rect 1302 5108 1308 5160
rect 1360 5148 1366 5160
rect 1581 5151 1639 5157
rect 1581 5148 1593 5151
rect 1360 5120 1593 5148
rect 1360 5108 1366 5120
rect 1581 5117 1593 5120
rect 1627 5117 1639 5151
rect 1581 5111 1639 5117
rect 17126 5108 17132 5160
rect 17184 5108 17190 5160
rect 17512 5157 17540 5188
rect 17957 5185 17969 5188
rect 18003 5185 18015 5219
rect 17957 5179 18015 5185
rect 18414 5176 18420 5228
rect 18472 5176 18478 5228
rect 19521 5219 19579 5225
rect 19521 5185 19533 5219
rect 19567 5216 19579 5219
rect 20346 5216 20352 5228
rect 19567 5188 20352 5216
rect 19567 5185 19579 5188
rect 19521 5179 19579 5185
rect 20346 5176 20352 5188
rect 20404 5176 20410 5228
rect 20806 5176 20812 5228
rect 20864 5176 20870 5228
rect 22186 5176 22192 5228
rect 22244 5216 22250 5228
rect 22316 5219 22374 5225
rect 22316 5216 22328 5219
rect 22244 5188 22328 5216
rect 22244 5176 22250 5188
rect 22316 5185 22328 5188
rect 22362 5185 22374 5219
rect 22316 5179 22374 5185
rect 22922 5176 22928 5228
rect 22980 5176 22986 5228
rect 23566 5176 23572 5228
rect 23624 5216 23630 5228
rect 24064 5219 24122 5225
rect 24064 5216 24076 5219
rect 23624 5188 24076 5216
rect 23624 5176 23630 5188
rect 24064 5185 24076 5188
rect 24110 5185 24122 5219
rect 24064 5179 24122 5185
rect 24670 5176 24676 5228
rect 24728 5176 24734 5228
rect 38102 5176 38108 5228
rect 38160 5216 38166 5228
rect 38565 5219 38623 5225
rect 38565 5216 38577 5219
rect 38160 5188 38577 5216
rect 38160 5176 38166 5188
rect 38565 5185 38577 5188
rect 38611 5185 38623 5219
rect 38565 5179 38623 5185
rect 40126 5176 40132 5228
rect 40184 5216 40190 5228
rect 45833 5219 45891 5225
rect 45833 5216 45845 5219
rect 40184 5188 45845 5216
rect 40184 5176 40190 5188
rect 45833 5185 45845 5188
rect 45879 5185 45891 5219
rect 45833 5179 45891 5185
rect 47854 5176 47860 5228
rect 47912 5216 47918 5228
rect 47949 5219 48007 5225
rect 47949 5216 47961 5219
rect 47912 5188 47961 5216
rect 47912 5176 47918 5188
rect 47949 5185 47961 5188
rect 47995 5185 48007 5219
rect 47949 5179 48007 5185
rect 17497 5151 17555 5157
rect 17497 5117 17509 5151
rect 17543 5148 17555 5151
rect 22419 5151 22477 5157
rect 17543 5120 22094 5148
rect 17543 5117 17555 5120
rect 17497 5111 17555 5117
rect 17773 5083 17831 5089
rect 17773 5049 17785 5083
rect 17819 5080 17831 5083
rect 19242 5080 19248 5092
rect 17819 5052 19248 5080
rect 17819 5049 17831 5052
rect 17773 5043 17831 5049
rect 19242 5040 19248 5052
rect 19300 5040 19306 5092
rect 22066 5080 22094 5120
rect 22419 5117 22431 5151
rect 22465 5148 22477 5151
rect 24302 5148 24308 5160
rect 22465 5120 24308 5148
rect 22465 5117 22477 5120
rect 22419 5111 22477 5117
rect 24302 5108 24308 5120
rect 24360 5108 24366 5160
rect 39485 5151 39543 5157
rect 39485 5117 39497 5151
rect 39531 5148 39543 5151
rect 40402 5148 40408 5160
rect 39531 5120 40408 5148
rect 39531 5117 39543 5120
rect 39485 5111 39543 5117
rect 40402 5108 40408 5120
rect 40460 5108 40466 5160
rect 46845 5151 46903 5157
rect 46845 5117 46857 5151
rect 46891 5148 46903 5151
rect 48314 5148 48320 5160
rect 46891 5120 48320 5148
rect 46891 5117 46903 5120
rect 46845 5111 46903 5117
rect 48314 5108 48320 5120
rect 48372 5108 48378 5160
rect 35894 5080 35900 5092
rect 22066 5052 35900 5080
rect 35894 5040 35900 5052
rect 35952 5040 35958 5092
rect 38749 5083 38807 5089
rect 38749 5049 38761 5083
rect 38795 5080 38807 5083
rect 44266 5080 44272 5092
rect 38795 5052 44272 5080
rect 38795 5049 38807 5052
rect 38749 5043 38807 5049
rect 44266 5040 44272 5052
rect 44324 5040 44330 5092
rect 21453 5015 21511 5021
rect 21453 4981 21465 5015
rect 21499 5012 21511 5015
rect 22002 5012 22008 5024
rect 21499 4984 22008 5012
rect 21499 4981 21511 4984
rect 21453 4975 21511 4981
rect 22002 4972 22008 4984
rect 22060 4972 22066 5024
rect 24167 5015 24225 5021
rect 24167 4981 24179 5015
rect 24213 5012 24225 5015
rect 24762 5012 24768 5024
rect 24213 4984 24768 5012
rect 24213 4981 24225 4984
rect 24167 4975 24225 4981
rect 24762 4972 24768 4984
rect 24820 4972 24826 5024
rect 24854 4972 24860 5024
rect 24912 5012 24918 5024
rect 25317 5015 25375 5021
rect 25317 5012 25329 5015
rect 24912 4984 25329 5012
rect 24912 4972 24918 4984
rect 25317 4981 25329 4984
rect 25363 4981 25375 5015
rect 25317 4975 25375 4981
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 1302 4768 1308 4820
rect 1360 4808 1366 4820
rect 2133 4811 2191 4817
rect 2133 4808 2145 4811
rect 1360 4780 2145 4808
rect 1360 4768 1366 4780
rect 2133 4777 2145 4780
rect 2179 4777 2191 4811
rect 2133 4771 2191 4777
rect 20162 4768 20168 4820
rect 20220 4768 20226 4820
rect 20714 4768 20720 4820
rect 20772 4808 20778 4820
rect 21082 4808 21088 4820
rect 20772 4780 21088 4808
rect 20772 4768 20778 4780
rect 21082 4768 21088 4780
rect 21140 4808 21146 4820
rect 24029 4811 24087 4817
rect 21140 4780 23980 4808
rect 21140 4768 21146 4780
rect 18693 4743 18751 4749
rect 18693 4709 18705 4743
rect 18739 4740 18751 4743
rect 20898 4740 20904 4752
rect 18739 4712 20904 4740
rect 18739 4709 18751 4712
rect 18693 4703 18751 4709
rect 20898 4700 20904 4712
rect 20956 4700 20962 4752
rect 23952 4740 23980 4780
rect 24029 4777 24041 4811
rect 24075 4808 24087 4811
rect 24670 4808 24676 4820
rect 24075 4780 24676 4808
rect 24075 4777 24087 4780
rect 24029 4771 24087 4777
rect 24670 4768 24676 4780
rect 24728 4768 24734 4820
rect 45830 4768 45836 4820
rect 45888 4768 45894 4820
rect 46198 4768 46204 4820
rect 46256 4808 46262 4820
rect 46477 4811 46535 4817
rect 46477 4808 46489 4811
rect 46256 4780 46489 4808
rect 46256 4768 46262 4780
rect 46477 4777 46489 4780
rect 46523 4777 46535 4811
rect 46477 4771 46535 4777
rect 46750 4768 46756 4820
rect 46808 4768 46814 4820
rect 47029 4811 47087 4817
rect 47029 4777 47041 4811
rect 47075 4808 47087 4811
rect 47302 4808 47308 4820
rect 47075 4780 47308 4808
rect 47075 4777 47087 4780
rect 47029 4771 47087 4777
rect 47302 4768 47308 4780
rect 47360 4768 47366 4820
rect 47394 4768 47400 4820
rect 47452 4808 47458 4820
rect 47581 4811 47639 4817
rect 47581 4808 47593 4811
rect 47452 4780 47593 4808
rect 47452 4768 47458 4780
rect 47581 4777 47593 4780
rect 47627 4777 47639 4811
rect 47581 4771 47639 4777
rect 46109 4743 46167 4749
rect 23952 4712 25728 4740
rect 19150 4632 19156 4684
rect 19208 4672 19214 4684
rect 20714 4672 20720 4684
rect 19208 4644 20720 4672
rect 19208 4632 19214 4644
rect 20714 4632 20720 4644
rect 20772 4632 20778 4684
rect 20993 4675 21051 4681
rect 20993 4641 21005 4675
rect 21039 4672 21051 4675
rect 21818 4672 21824 4684
rect 21039 4644 21824 4672
rect 21039 4641 21051 4644
rect 20993 4635 21051 4641
rect 21818 4632 21824 4644
rect 21876 4672 21882 4684
rect 23017 4675 23075 4681
rect 23017 4672 23029 4675
rect 21876 4644 23029 4672
rect 21876 4632 21882 4644
rect 23017 4641 23029 4644
rect 23063 4672 23075 4675
rect 23290 4672 23296 4684
rect 23063 4644 23296 4672
rect 23063 4641 23075 4644
rect 23017 4635 23075 4641
rect 23290 4632 23296 4644
rect 23348 4632 23354 4684
rect 24762 4632 24768 4684
rect 24820 4672 24826 4684
rect 25700 4681 25728 4712
rect 46109 4709 46121 4743
rect 46155 4740 46167 4743
rect 46566 4740 46572 4752
rect 46155 4712 46572 4740
rect 46155 4709 46167 4712
rect 46109 4703 46167 4709
rect 46566 4700 46572 4712
rect 46624 4700 46630 4752
rect 25409 4675 25467 4681
rect 25409 4672 25421 4675
rect 24820 4644 25421 4672
rect 24820 4632 24826 4644
rect 25409 4641 25421 4644
rect 25455 4641 25467 4675
rect 25409 4635 25467 4641
rect 25685 4675 25743 4681
rect 25685 4641 25697 4675
rect 25731 4641 25743 4675
rect 25685 4635 25743 4641
rect 40218 4632 40224 4684
rect 40276 4672 40282 4684
rect 49145 4675 49203 4681
rect 40276 4644 47992 4672
rect 40276 4632 40282 4644
rect 2317 4607 2375 4613
rect 2317 4604 2329 4607
rect 1688 4576 2329 4604
rect 1302 4496 1308 4548
rect 1360 4536 1366 4548
rect 1688 4545 1716 4576
rect 2317 4573 2329 4576
rect 2363 4573 2375 4607
rect 2317 4567 2375 4573
rect 18782 4564 18788 4616
rect 18840 4604 18846 4616
rect 18877 4607 18935 4613
rect 18877 4604 18889 4607
rect 18840 4576 18889 4604
rect 18840 4564 18846 4576
rect 18877 4573 18889 4576
rect 18923 4573 18935 4607
rect 18877 4567 18935 4573
rect 19521 4607 19579 4613
rect 19521 4573 19533 4607
rect 19567 4604 19579 4607
rect 20438 4604 20444 4616
rect 19567 4576 20444 4604
rect 19567 4573 19579 4576
rect 19521 4567 19579 4573
rect 20438 4564 20444 4576
rect 20496 4564 20502 4616
rect 23385 4607 23443 4613
rect 1673 4539 1731 4545
rect 1673 4536 1685 4539
rect 1360 4508 1685 4536
rect 1360 4496 1366 4508
rect 1673 4505 1685 4508
rect 1719 4505 1731 4539
rect 1673 4499 1731 4505
rect 1857 4539 1915 4545
rect 1857 4505 1869 4539
rect 1903 4536 1915 4539
rect 19702 4536 19708 4548
rect 1903 4508 19708 4536
rect 1903 4505 1915 4508
rect 1857 4499 1915 4505
rect 19702 4496 19708 4508
rect 19760 4496 19766 4548
rect 21266 4496 21272 4548
rect 21324 4496 21330 4548
rect 20717 4471 20775 4477
rect 20717 4437 20729 4471
rect 20763 4468 20775 4471
rect 22094 4468 22100 4480
rect 20763 4440 22100 4468
rect 20763 4437 20775 4440
rect 20717 4431 20775 4437
rect 22094 4428 22100 4440
rect 22152 4468 22158 4480
rect 22388 4468 22416 4590
rect 23385 4573 23397 4607
rect 23431 4604 23443 4607
rect 24026 4604 24032 4616
rect 23431 4576 24032 4604
rect 23431 4573 23443 4576
rect 23385 4567 23443 4573
rect 24026 4564 24032 4576
rect 24084 4564 24090 4616
rect 24616 4607 24674 4613
rect 24616 4604 24628 4607
rect 24136 4576 24628 4604
rect 22830 4496 22836 4548
rect 22888 4536 22894 4548
rect 24136 4536 24164 4576
rect 24616 4573 24628 4576
rect 24662 4573 24674 4607
rect 24616 4567 24674 4573
rect 25222 4564 25228 4616
rect 25280 4564 25286 4616
rect 28626 4564 28632 4616
rect 28684 4604 28690 4616
rect 38105 4607 38163 4613
rect 38105 4604 38117 4607
rect 28684 4576 38117 4604
rect 28684 4564 28690 4576
rect 38105 4573 38117 4576
rect 38151 4604 38163 4607
rect 38565 4607 38623 4613
rect 38565 4604 38577 4607
rect 38151 4576 38577 4604
rect 38151 4573 38163 4576
rect 38105 4567 38163 4573
rect 38565 4573 38577 4576
rect 38611 4573 38623 4607
rect 38565 4567 38623 4573
rect 46290 4564 46296 4616
rect 46348 4564 46354 4616
rect 47964 4613 47992 4644
rect 49145 4641 49157 4675
rect 49191 4672 49203 4675
rect 49418 4672 49424 4684
rect 49191 4644 49424 4672
rect 49191 4641 49203 4644
rect 49145 4635 49203 4641
rect 49418 4632 49424 4644
rect 49476 4632 49482 4684
rect 47213 4607 47271 4613
rect 47213 4573 47225 4607
rect 47259 4573 47271 4607
rect 47213 4567 47271 4573
rect 47949 4607 48007 4613
rect 47949 4573 47961 4607
rect 47995 4573 48007 4607
rect 47949 4567 48007 4573
rect 22888 4508 24164 4536
rect 37369 4539 37427 4545
rect 22888 4496 22894 4508
rect 37369 4505 37381 4539
rect 37415 4505 37427 4539
rect 37369 4499 37427 4505
rect 38289 4539 38347 4545
rect 38289 4505 38301 4539
rect 38335 4536 38347 4539
rect 42794 4536 42800 4548
rect 38335 4508 42800 4536
rect 38335 4505 38347 4508
rect 38289 4499 38347 4505
rect 22152 4440 22416 4468
rect 22152 4428 22158 4440
rect 22738 4428 22744 4480
rect 22796 4428 22802 4480
rect 24719 4471 24777 4477
rect 24719 4437 24731 4471
rect 24765 4468 24777 4471
rect 26142 4468 26148 4480
rect 24765 4440 26148 4468
rect 24765 4437 24777 4440
rect 24719 4431 24777 4437
rect 26142 4428 26148 4440
rect 26200 4428 26206 4480
rect 27154 4428 27160 4480
rect 27212 4468 27218 4480
rect 36909 4471 36967 4477
rect 36909 4468 36921 4471
rect 27212 4440 36921 4468
rect 27212 4428 27218 4440
rect 36909 4437 36921 4440
rect 36955 4468 36967 4471
rect 37384 4468 37412 4499
rect 42794 4496 42800 4508
rect 42852 4496 42858 4548
rect 47228 4536 47256 4567
rect 48958 4536 48964 4548
rect 47228 4508 48964 4536
rect 48958 4496 48964 4508
rect 49016 4496 49022 4548
rect 36955 4440 37412 4468
rect 37461 4471 37519 4477
rect 36955 4437 36967 4440
rect 36909 4431 36967 4437
rect 37461 4437 37473 4471
rect 37507 4468 37519 4471
rect 39390 4468 39396 4480
rect 37507 4440 39396 4468
rect 37507 4437 37519 4440
rect 37461 4431 37519 4437
rect 39390 4428 39396 4440
rect 39448 4428 39454 4480
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 21085 4267 21143 4273
rect 21085 4233 21097 4267
rect 21131 4264 21143 4267
rect 21266 4264 21272 4276
rect 21131 4236 21272 4264
rect 21131 4233 21143 4236
rect 21085 4227 21143 4233
rect 21266 4224 21272 4236
rect 21324 4224 21330 4276
rect 22094 4224 22100 4276
rect 22152 4264 22158 4276
rect 24578 4264 24584 4276
rect 22152 4236 24584 4264
rect 22152 4224 22158 4236
rect 24578 4224 24584 4236
rect 24636 4224 24642 4276
rect 25222 4224 25228 4276
rect 25280 4264 25286 4276
rect 32858 4264 32864 4276
rect 25280 4236 32864 4264
rect 25280 4224 25286 4236
rect 32858 4224 32864 4236
rect 32916 4224 32922 4276
rect 27341 4199 27399 4205
rect 27341 4196 27353 4199
rect 2240 4168 2452 4196
rect 1302 4088 1308 4140
rect 1360 4128 1366 4140
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 1360 4100 1593 4128
rect 1360 4088 1366 4100
rect 1581 4097 1593 4100
rect 1627 4128 1639 4131
rect 2240 4128 2268 4168
rect 1627 4100 2268 4128
rect 2317 4131 2375 4137
rect 1627 4097 1639 4100
rect 1581 4091 1639 4097
rect 2317 4097 2329 4131
rect 2363 4097 2375 4131
rect 2424 4128 2452 4168
rect 27172 4168 27353 4196
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 2424 4100 3065 4128
rect 2317 4091 2375 4097
rect 3053 4097 3065 4100
rect 3099 4097 3111 4131
rect 3053 4091 3111 4097
rect 9677 4131 9735 4137
rect 9677 4097 9689 4131
rect 9723 4128 9735 4131
rect 9858 4128 9864 4140
rect 9723 4100 9864 4128
rect 9723 4097 9735 4100
rect 9677 4091 9735 4097
rect 1210 4020 1216 4072
rect 1268 4060 1274 4072
rect 2332 4060 2360 4091
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 17770 4088 17776 4140
rect 17828 4128 17834 4140
rect 18141 4131 18199 4137
rect 18141 4128 18153 4131
rect 17828 4100 18153 4128
rect 17828 4088 17834 4100
rect 18141 4097 18153 4100
rect 18187 4097 18199 4131
rect 18141 4091 18199 4097
rect 20070 4088 20076 4140
rect 20128 4128 20134 4140
rect 20441 4131 20499 4137
rect 20441 4128 20453 4131
rect 20128 4100 20453 4128
rect 20128 4088 20134 4100
rect 20441 4097 20453 4100
rect 20487 4097 20499 4131
rect 20441 4091 20499 4097
rect 22002 4088 22008 4140
rect 22060 4088 22066 4140
rect 23109 4131 23167 4137
rect 23109 4097 23121 4131
rect 23155 4128 23167 4131
rect 23934 4128 23940 4140
rect 23155 4100 23940 4128
rect 23155 4097 23167 4100
rect 23109 4091 23167 4097
rect 23934 4088 23940 4100
rect 23992 4088 23998 4140
rect 26142 4088 26148 4140
rect 26200 4128 26206 4140
rect 27172 4128 27200 4168
rect 27341 4165 27353 4168
rect 27387 4165 27399 4199
rect 27341 4159 27399 4165
rect 27614 4156 27620 4208
rect 27672 4196 27678 4208
rect 37553 4199 37611 4205
rect 37553 4196 37565 4199
rect 27672 4168 37565 4196
rect 27672 4156 27678 4168
rect 37553 4165 37565 4168
rect 37599 4196 37611 4199
rect 38013 4199 38071 4205
rect 38013 4196 38025 4199
rect 37599 4168 38025 4196
rect 37599 4165 37611 4168
rect 37553 4159 37611 4165
rect 38013 4165 38025 4168
rect 38059 4165 38071 4199
rect 38013 4159 38071 4165
rect 26200 4100 27200 4128
rect 37737 4131 37795 4137
rect 26200 4088 26206 4100
rect 37737 4097 37749 4131
rect 37783 4128 37795 4131
rect 45833 4131 45891 4137
rect 45833 4128 45845 4131
rect 37783 4100 45845 4128
rect 37783 4097 37795 4100
rect 37737 4091 37795 4097
rect 45833 4097 45845 4100
rect 45879 4097 45891 4131
rect 47949 4131 48007 4137
rect 47949 4128 47961 4131
rect 45833 4091 45891 4097
rect 45940 4100 47961 4128
rect 1268 4032 2360 4060
rect 1268 4020 1274 4032
rect 1765 3995 1823 4001
rect 1765 3961 1777 3995
rect 1811 3992 1823 3995
rect 2130 3992 2136 4004
rect 1811 3964 2136 3992
rect 1811 3961 1823 3964
rect 1765 3955 1823 3961
rect 2130 3952 2136 3964
rect 2188 3952 2194 4004
rect 2332 3924 2360 4032
rect 2406 4020 2412 4072
rect 2464 4060 2470 4072
rect 2464 4032 12434 4060
rect 2464 4020 2470 4032
rect 2501 3995 2559 4001
rect 2501 3961 2513 3995
rect 2547 3992 2559 3995
rect 8294 3992 8300 4004
rect 2547 3964 8300 3992
rect 2547 3961 2559 3964
rect 2501 3955 2559 3961
rect 8294 3952 8300 3964
rect 8352 3952 8358 4004
rect 2869 3927 2927 3933
rect 2869 3924 2881 3927
rect 2332 3896 2881 3924
rect 2869 3893 2881 3896
rect 2915 3893 2927 3927
rect 2869 3887 2927 3893
rect 9674 3884 9680 3936
rect 9732 3924 9738 3936
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 9732 3896 10333 3924
rect 9732 3884 9738 3896
rect 10321 3893 10333 3896
rect 10367 3893 10379 3927
rect 12406 3924 12434 4032
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 18325 4063 18383 4069
rect 18325 4060 18337 4063
rect 16264 4032 18337 4060
rect 16264 4020 16270 4032
rect 18325 4029 18337 4032
rect 18371 4029 18383 4063
rect 18325 4023 18383 4029
rect 19981 4063 20039 4069
rect 19981 4029 19993 4063
rect 20027 4060 20039 4063
rect 20162 4060 20168 4072
rect 20027 4032 20168 4060
rect 20027 4029 20039 4032
rect 19981 4023 20039 4029
rect 18340 3992 18368 4023
rect 20162 4020 20168 4032
rect 20220 4020 20226 4072
rect 22649 4063 22707 4069
rect 22649 4029 22661 4063
rect 22695 4060 22707 4063
rect 23658 4060 23664 4072
rect 22695 4032 23664 4060
rect 22695 4029 22707 4032
rect 22649 4023 22707 4029
rect 23658 4020 23664 4032
rect 23716 4020 23722 4072
rect 24121 4063 24179 4069
rect 24121 4029 24133 4063
rect 24167 4060 24179 4063
rect 24167 4032 24256 4060
rect 24167 4029 24179 4032
rect 24121 4023 24179 4029
rect 20714 3992 20720 4004
rect 18340 3964 20720 3992
rect 20714 3952 20720 3964
rect 20772 3952 20778 4004
rect 18506 3924 18512 3936
rect 12406 3896 18512 3924
rect 10321 3887 10379 3893
rect 18506 3884 18512 3896
rect 18564 3884 18570 3936
rect 22738 3884 22744 3936
rect 22796 3924 22802 3936
rect 23201 3927 23259 3933
rect 23201 3924 23213 3927
rect 22796 3896 23213 3924
rect 22796 3884 22802 3896
rect 23201 3893 23213 3896
rect 23247 3924 23259 3927
rect 23382 3924 23388 3936
rect 23247 3896 23388 3924
rect 23247 3893 23259 3896
rect 23201 3887 23259 3893
rect 23382 3884 23388 3896
rect 23440 3884 23446 3936
rect 23566 3884 23572 3936
rect 23624 3884 23630 3936
rect 24228 3924 24256 4032
rect 24302 4020 24308 4072
rect 24360 4020 24366 4072
rect 24946 4020 24952 4072
rect 25004 4020 25010 4072
rect 27157 4063 27215 4069
rect 27157 4029 27169 4063
rect 27203 4029 27215 4063
rect 27157 4023 27215 4029
rect 27172 3992 27200 4023
rect 27614 4020 27620 4072
rect 27672 4020 27678 4072
rect 39206 4020 39212 4072
rect 39264 4060 39270 4072
rect 45940 4060 45968 4100
rect 47949 4097 47961 4100
rect 47995 4097 48007 4131
rect 47949 4091 48007 4097
rect 49145 4131 49203 4137
rect 49145 4097 49157 4131
rect 49191 4128 49203 4131
rect 49234 4128 49240 4140
rect 49191 4100 49240 4128
rect 49191 4097 49203 4100
rect 49145 4091 49203 4097
rect 49234 4088 49240 4100
rect 49292 4088 49298 4140
rect 39264 4032 45968 4060
rect 39264 4020 39270 4032
rect 46658 4020 46664 4072
rect 46716 4020 46722 4072
rect 47673 4063 47731 4069
rect 47673 4029 47685 4063
rect 47719 4060 47731 4063
rect 49786 4060 49792 4072
rect 47719 4032 49792 4060
rect 47719 4029 47731 4032
rect 47673 4023 47731 4029
rect 49786 4020 49792 4032
rect 49844 4020 49850 4072
rect 34422 3992 34428 4004
rect 27172 3964 34428 3992
rect 34422 3952 34428 3964
rect 34480 3952 34486 4004
rect 40494 3952 40500 4004
rect 40552 3992 40558 4004
rect 45554 3992 45560 4004
rect 40552 3964 45560 3992
rect 40552 3952 40558 3964
rect 45554 3952 45560 3964
rect 45612 3952 45618 4004
rect 30834 3924 30840 3936
rect 24228 3896 30840 3924
rect 30834 3884 30840 3896
rect 30892 3884 30898 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 11606 3720 11612 3732
rect 1872 3692 11612 3720
rect 1872 3593 1900 3692
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 20070 3680 20076 3732
rect 20128 3680 20134 3732
rect 24118 3720 24124 3732
rect 20180 3692 24124 3720
rect 3326 3612 3332 3664
rect 3384 3652 3390 3664
rect 19150 3652 19156 3664
rect 3384 3624 19156 3652
rect 3384 3612 3390 3624
rect 19150 3612 19156 3624
rect 19208 3612 19214 3664
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3553 1915 3587
rect 20180 3584 20208 3692
rect 24118 3680 24124 3692
rect 24176 3720 24182 3732
rect 27614 3720 27620 3732
rect 24176 3692 27620 3720
rect 24176 3680 24182 3692
rect 27614 3680 27620 3692
rect 27672 3680 27678 3732
rect 33870 3680 33876 3732
rect 33928 3720 33934 3732
rect 43438 3720 43444 3732
rect 33928 3692 43444 3720
rect 33928 3680 33934 3692
rect 43438 3680 43444 3692
rect 43496 3680 43502 3732
rect 20714 3612 20720 3664
rect 20772 3652 20778 3664
rect 21634 3652 21640 3664
rect 20772 3624 21640 3652
rect 20772 3612 20778 3624
rect 21634 3612 21640 3624
rect 21692 3652 21698 3664
rect 24486 3652 24492 3664
rect 21692 3624 24492 3652
rect 21692 3612 21698 3624
rect 24486 3612 24492 3624
rect 24544 3612 24550 3664
rect 27522 3612 27528 3664
rect 27580 3652 27586 3664
rect 36814 3652 36820 3664
rect 27580 3624 36820 3652
rect 27580 3612 27586 3624
rect 36814 3612 36820 3624
rect 36872 3612 36878 3664
rect 39666 3612 39672 3664
rect 39724 3652 39730 3664
rect 49786 3652 49792 3664
rect 39724 3624 49792 3652
rect 39724 3612 39730 3624
rect 49786 3612 49792 3624
rect 49844 3612 49850 3664
rect 1857 3547 1915 3553
rect 2746 3556 20208 3584
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1581 3519 1639 3525
rect 1581 3516 1593 3519
rect 1360 3488 1593 3516
rect 1360 3476 1366 3488
rect 1581 3485 1593 3488
rect 1627 3485 1639 3519
rect 1581 3479 1639 3485
rect 1026 3408 1032 3460
rect 1084 3448 1090 3460
rect 2746 3448 2774 3556
rect 23290 3544 23296 3596
rect 23348 3584 23354 3596
rect 24581 3587 24639 3593
rect 24581 3584 24593 3587
rect 23348 3556 24593 3584
rect 23348 3544 23354 3556
rect 24581 3553 24593 3556
rect 24627 3553 24639 3587
rect 24581 3547 24639 3553
rect 24854 3544 24860 3596
rect 24912 3544 24918 3596
rect 37090 3544 37096 3596
rect 37148 3584 37154 3596
rect 47670 3584 47676 3596
rect 37148 3556 47676 3584
rect 37148 3544 37154 3556
rect 47670 3544 47676 3556
rect 47728 3544 47734 3596
rect 49142 3544 49148 3596
rect 49200 3544 49206 3596
rect 9582 3476 9588 3528
rect 9640 3476 9646 3528
rect 10042 3476 10048 3528
rect 10100 3476 10106 3528
rect 11146 3476 11152 3528
rect 11204 3476 11210 3528
rect 16206 3476 16212 3528
rect 16264 3476 16270 3528
rect 17129 3519 17187 3525
rect 17129 3485 17141 3519
rect 17175 3485 17187 3519
rect 17129 3479 17187 3485
rect 1084 3420 2774 3448
rect 1084 3408 1090 3420
rect 5350 3340 5356 3392
rect 5408 3380 5414 3392
rect 7466 3380 7472 3392
rect 5408 3352 7472 3380
rect 5408 3340 5414 3352
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 8754 3340 8760 3392
rect 8812 3340 8818 3392
rect 9401 3383 9459 3389
rect 9401 3349 9413 3383
rect 9447 3380 9459 3383
rect 10502 3380 10508 3392
rect 9447 3352 10508 3380
rect 9447 3349 9459 3352
rect 9401 3343 9459 3349
rect 10502 3340 10508 3352
rect 10560 3340 10566 3392
rect 10686 3340 10692 3392
rect 10744 3340 10750 3392
rect 11793 3383 11851 3389
rect 11793 3349 11805 3383
rect 11839 3380 11851 3383
rect 12342 3380 12348 3392
rect 11839 3352 12348 3380
rect 11839 3349 11851 3352
rect 11793 3343 11851 3349
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 12434 3340 12440 3392
rect 12492 3380 12498 3392
rect 16301 3383 16359 3389
rect 16301 3380 16313 3383
rect 12492 3352 16313 3380
rect 12492 3340 12498 3352
rect 16301 3349 16313 3352
rect 16347 3349 16359 3383
rect 16301 3343 16359 3349
rect 16390 3340 16396 3392
rect 16448 3380 16454 3392
rect 16945 3383 17003 3389
rect 16945 3380 16957 3383
rect 16448 3352 16957 3380
rect 16448 3340 16454 3352
rect 16945 3349 16957 3352
rect 16991 3349 17003 3383
rect 17144 3380 17172 3479
rect 17586 3476 17592 3528
rect 17644 3476 17650 3528
rect 18233 3519 18291 3525
rect 18233 3485 18245 3519
rect 18279 3516 18291 3519
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 18279 3488 19441 3516
rect 18279 3485 18291 3488
rect 18233 3479 18291 3485
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 19518 3476 19524 3528
rect 19576 3516 19582 3528
rect 20993 3519 21051 3525
rect 20993 3516 21005 3519
rect 19576 3488 21005 3516
rect 19576 3476 19582 3488
rect 20993 3485 21005 3488
rect 21039 3485 21051 3519
rect 20993 3479 21051 3485
rect 23382 3476 23388 3528
rect 23440 3476 23446 3528
rect 24026 3476 24032 3528
rect 24084 3476 24090 3528
rect 27157 3519 27215 3525
rect 27157 3516 27169 3519
rect 26344 3488 27169 3516
rect 18874 3408 18880 3460
rect 18932 3448 18938 3460
rect 21177 3451 21235 3457
rect 21177 3448 21189 3451
rect 18932 3420 21189 3448
rect 18932 3408 18938 3420
rect 21177 3417 21189 3420
rect 21223 3448 21235 3451
rect 22833 3451 22891 3457
rect 21223 3420 22094 3448
rect 21223 3417 21235 3420
rect 21177 3411 21235 3417
rect 19518 3380 19524 3392
rect 17144 3352 19524 3380
rect 16945 3343 17003 3349
rect 19518 3340 19524 3352
rect 19576 3340 19582 3392
rect 22066 3380 22094 3420
rect 22833 3417 22845 3451
rect 22879 3448 22891 3451
rect 24394 3448 24400 3460
rect 22879 3420 24400 3448
rect 22879 3417 22891 3420
rect 22833 3411 22891 3417
rect 24394 3408 24400 3420
rect 24452 3408 24458 3460
rect 24578 3408 24584 3460
rect 24636 3448 24642 3460
rect 24636 3420 25346 3448
rect 24636 3408 24642 3420
rect 26344 3392 26372 3488
rect 27157 3485 27169 3488
rect 27203 3485 27215 3519
rect 27157 3479 27215 3485
rect 27801 3519 27859 3525
rect 27801 3485 27813 3519
rect 27847 3516 27859 3519
rect 28261 3519 28319 3525
rect 28261 3516 28273 3519
rect 27847 3488 28273 3516
rect 27847 3485 27859 3488
rect 27801 3479 27859 3485
rect 28261 3485 28273 3488
rect 28307 3485 28319 3519
rect 28261 3479 28319 3485
rect 28905 3519 28963 3525
rect 28905 3485 28917 3519
rect 28951 3516 28963 3519
rect 29733 3519 29791 3525
rect 29733 3516 29745 3519
rect 28951 3488 29745 3516
rect 28951 3485 28963 3488
rect 28905 3479 28963 3485
rect 29733 3485 29745 3488
rect 29779 3485 29791 3519
rect 29733 3479 29791 3485
rect 40402 3476 40408 3528
rect 40460 3516 40466 3528
rect 46109 3519 46167 3525
rect 46109 3516 46121 3519
rect 40460 3488 46121 3516
rect 40460 3476 40466 3488
rect 46109 3485 46121 3488
rect 46155 3485 46167 3519
rect 46109 3479 46167 3485
rect 47118 3476 47124 3528
rect 47176 3516 47182 3528
rect 47949 3519 48007 3525
rect 47949 3516 47961 3519
rect 47176 3488 47961 3516
rect 47176 3476 47182 3488
rect 47949 3485 47961 3488
rect 47995 3485 48007 3519
rect 47949 3479 48007 3485
rect 30098 3408 30104 3460
rect 30156 3448 30162 3460
rect 39206 3448 39212 3460
rect 30156 3420 39212 3448
rect 30156 3408 30162 3420
rect 39206 3408 39212 3420
rect 39264 3408 39270 3460
rect 47305 3451 47363 3457
rect 47305 3417 47317 3451
rect 47351 3448 47363 3451
rect 48682 3448 48688 3460
rect 47351 3420 48688 3448
rect 47351 3417 47363 3420
rect 47305 3411 47363 3417
rect 48682 3408 48688 3420
rect 48740 3408 48746 3460
rect 23566 3380 23572 3392
rect 22066 3352 23572 3380
rect 23566 3340 23572 3352
rect 23624 3340 23630 3392
rect 26326 3340 26332 3392
rect 26384 3340 26390 3392
rect 29086 3340 29092 3392
rect 29144 3380 29150 3392
rect 30377 3383 30435 3389
rect 30377 3380 30389 3383
rect 29144 3352 30389 3380
rect 29144 3340 29150 3352
rect 30377 3349 30389 3352
rect 30423 3349 30435 3383
rect 30377 3343 30435 3349
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 1302 3136 1308 3188
rect 1360 3176 1366 3188
rect 2133 3179 2191 3185
rect 2133 3176 2145 3179
rect 1360 3148 2145 3176
rect 1360 3136 1366 3148
rect 2133 3145 2145 3148
rect 2179 3145 2191 3179
rect 2133 3139 2191 3145
rect 9582 3136 9588 3188
rect 9640 3176 9646 3188
rect 10045 3179 10103 3185
rect 10045 3176 10057 3179
rect 9640 3148 10057 3176
rect 9640 3136 9646 3148
rect 10045 3145 10057 3148
rect 10091 3145 10103 3179
rect 10045 3139 10103 3145
rect 11146 3136 11152 3188
rect 11204 3136 11210 3188
rect 16298 3176 16304 3188
rect 14568 3148 16304 3176
rect 10686 3108 10692 3120
rect 9416 3080 10692 3108
rect 1302 3000 1308 3052
rect 1360 3040 1366 3052
rect 9416 3049 9444 3080
rect 10686 3068 10692 3080
rect 10744 3068 10750 3120
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 1360 3012 1593 3040
rect 1360 3000 1366 3012
rect 1581 3009 1593 3012
rect 1627 3040 1639 3043
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 1627 3012 2513 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3009 8355 3043
rect 8297 3003 8355 3009
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 8312 2972 8340 3003
rect 10502 3000 10508 3052
rect 10560 3000 10566 3052
rect 12342 3000 12348 3052
rect 12400 3000 12406 3052
rect 14568 3049 14596 3148
rect 16298 3136 16304 3148
rect 16356 3136 16362 3188
rect 17034 3176 17040 3188
rect 16960 3148 17040 3176
rect 16960 3108 16988 3148
rect 17034 3136 17040 3148
rect 17092 3136 17098 3188
rect 18693 3179 18751 3185
rect 18693 3145 18705 3179
rect 18739 3145 18751 3179
rect 19794 3176 19800 3188
rect 18693 3139 18751 3145
rect 18984 3148 19800 3176
rect 16054 3080 16988 3108
rect 12989 3043 13047 3049
rect 12989 3009 13001 3043
rect 13035 3040 13047 3043
rect 13449 3043 13507 3049
rect 13449 3040 13461 3043
rect 13035 3012 13461 3040
rect 13035 3009 13047 3012
rect 12989 3003 13047 3009
rect 13449 3009 13461 3012
rect 13495 3009 13507 3043
rect 13449 3003 13507 3009
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3040 17095 3043
rect 18708 3040 18736 3139
rect 17083 3012 18736 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 18874 3000 18880 3052
rect 18932 3000 18938 3052
rect 9766 2972 9772 2984
rect 8312 2944 9772 2972
rect 9766 2932 9772 2944
rect 9824 2932 9830 2984
rect 14093 2975 14151 2981
rect 14093 2941 14105 2975
rect 14139 2972 14151 2975
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 14139 2944 14841 2972
rect 14139 2941 14151 2944
rect 14093 2935 14151 2941
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 16482 2932 16488 2984
rect 16540 2972 16546 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 16540 2944 17325 2972
rect 16540 2932 16546 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 1765 2907 1823 2913
rect 1765 2873 1777 2907
rect 1811 2904 1823 2907
rect 1811 2876 7420 2904
rect 1811 2873 1823 2876
rect 1765 2867 1823 2873
rect 2314 2796 2320 2848
rect 2372 2796 2378 2848
rect 2774 2796 2780 2848
rect 2832 2796 2838 2848
rect 7392 2836 7420 2876
rect 7466 2864 7472 2916
rect 7524 2904 7530 2916
rect 18984 2904 19012 3148
rect 19794 3136 19800 3148
rect 19852 3176 19858 3188
rect 19852 3148 22600 3176
rect 19852 3136 19858 3148
rect 19518 3068 19524 3120
rect 19576 3108 19582 3120
rect 22094 3108 22100 3120
rect 19576 3080 22100 3108
rect 19576 3068 19582 3080
rect 22094 3068 22100 3080
rect 22152 3108 22158 3120
rect 22462 3108 22468 3120
rect 22152 3080 22468 3108
rect 22152 3068 22158 3080
rect 22462 3068 22468 3080
rect 22520 3068 22526 3120
rect 22572 3108 22600 3148
rect 22646 3136 22652 3188
rect 22704 3176 22710 3188
rect 22741 3179 22799 3185
rect 22741 3176 22753 3179
rect 22704 3148 22753 3176
rect 22704 3136 22710 3148
rect 22741 3145 22753 3148
rect 22787 3176 22799 3179
rect 22830 3176 22836 3188
rect 22787 3148 22836 3176
rect 22787 3145 22799 3148
rect 22741 3139 22799 3145
rect 22830 3136 22836 3148
rect 22888 3136 22894 3188
rect 23290 3136 23296 3188
rect 23348 3136 23354 3188
rect 23934 3176 23940 3188
rect 23676 3148 23940 3176
rect 23566 3108 23572 3120
rect 22572 3080 23572 3108
rect 23566 3068 23572 3080
rect 23624 3068 23630 3120
rect 22281 3043 22339 3049
rect 22281 3009 22293 3043
rect 22327 3040 22339 3043
rect 23676 3040 23704 3148
rect 23934 3136 23940 3148
rect 23992 3136 23998 3188
rect 24486 3136 24492 3188
rect 24544 3176 24550 3188
rect 27985 3179 28043 3185
rect 27985 3176 27997 3179
rect 24544 3148 27997 3176
rect 24544 3136 24550 3148
rect 27985 3145 27997 3148
rect 28031 3145 28043 3179
rect 27985 3139 28043 3145
rect 23842 3068 23848 3120
rect 23900 3068 23906 3120
rect 29086 3068 29092 3120
rect 29144 3068 29150 3120
rect 29822 3068 29828 3120
rect 29880 3068 29886 3120
rect 49145 3111 49203 3117
rect 49145 3077 49157 3111
rect 49191 3108 49203 3111
rect 49234 3108 49240 3120
rect 49191 3080 49240 3108
rect 49191 3077 49203 3080
rect 49145 3071 49203 3077
rect 49234 3068 49240 3080
rect 49292 3068 49298 3120
rect 22327 3012 23704 3040
rect 22327 3009 22339 3012
rect 22281 3003 22339 3009
rect 27522 3000 27528 3052
rect 27580 3000 27586 3052
rect 28442 3000 28448 3052
rect 28500 3040 28506 3052
rect 28813 3043 28871 3049
rect 28813 3040 28825 3043
rect 28500 3012 28825 3040
rect 28500 3000 28506 3012
rect 28813 3009 28825 3012
rect 28859 3009 28871 3043
rect 28813 3003 28871 3009
rect 39390 3000 39396 3052
rect 39448 3040 39454 3052
rect 43993 3043 44051 3049
rect 43993 3040 44005 3043
rect 39448 3012 44005 3040
rect 39448 3000 39454 3012
rect 43993 3009 44005 3012
rect 44039 3009 44051 3043
rect 43993 3003 44051 3009
rect 45738 3000 45744 3052
rect 45796 3040 45802 3052
rect 45833 3043 45891 3049
rect 45833 3040 45845 3043
rect 45796 3012 45845 3040
rect 45796 3000 45802 3012
rect 45833 3009 45845 3012
rect 45879 3009 45891 3043
rect 45833 3003 45891 3009
rect 45922 3000 45928 3052
rect 45980 3040 45986 3052
rect 47949 3043 48007 3049
rect 47949 3040 47961 3043
rect 45980 3012 47961 3040
rect 45980 3000 45986 3012
rect 47949 3009 47961 3012
rect 47995 3009 48007 3043
rect 47949 3003 48007 3009
rect 19337 2975 19395 2981
rect 19337 2941 19349 2975
rect 19383 2972 19395 2975
rect 19610 2972 19616 2984
rect 19383 2944 19616 2972
rect 19383 2941 19395 2944
rect 19337 2935 19395 2941
rect 19610 2932 19616 2944
rect 19668 2932 19674 2984
rect 21177 2975 21235 2981
rect 21177 2941 21189 2975
rect 21223 2972 21235 2975
rect 23661 2975 23719 2981
rect 21223 2944 22094 2972
rect 21223 2941 21235 2944
rect 21177 2935 21235 2941
rect 7524 2876 12434 2904
rect 7524 2864 7530 2876
rect 8846 2836 8852 2848
rect 7392 2808 8852 2836
rect 8846 2796 8852 2808
rect 8904 2796 8910 2848
rect 8941 2839 8999 2845
rect 8941 2805 8953 2839
rect 8987 2836 8999 2839
rect 10226 2836 10232 2848
rect 8987 2808 10232 2836
rect 8987 2805 8999 2808
rect 8941 2799 8999 2805
rect 10226 2796 10232 2808
rect 10284 2796 10290 2848
rect 12406 2836 12434 2876
rect 16224 2876 19012 2904
rect 22066 2904 22094 2944
rect 23661 2941 23673 2975
rect 23707 2972 23719 2975
rect 23707 2944 23796 2972
rect 23707 2941 23719 2944
rect 23661 2935 23719 2941
rect 22278 2904 22284 2916
rect 22066 2876 22284 2904
rect 16224 2836 16252 2876
rect 22278 2864 22284 2876
rect 22336 2864 22342 2916
rect 23768 2904 23796 2944
rect 23842 2932 23848 2984
rect 23900 2972 23906 2984
rect 24121 2975 24179 2981
rect 24121 2972 24133 2975
rect 23900 2944 24133 2972
rect 23900 2932 23906 2944
rect 24121 2941 24133 2944
rect 24167 2972 24179 2975
rect 26050 2972 26056 2984
rect 24167 2944 26056 2972
rect 24167 2941 24179 2944
rect 24121 2935 24179 2941
rect 26050 2932 26056 2944
rect 26108 2932 26114 2984
rect 30561 2975 30619 2981
rect 30561 2972 30573 2975
rect 27816 2944 30573 2972
rect 24946 2904 24952 2916
rect 23768 2876 24952 2904
rect 24946 2864 24952 2876
rect 25004 2864 25010 2916
rect 12406 2808 16252 2836
rect 16301 2839 16359 2845
rect 16301 2805 16313 2839
rect 16347 2836 16359 2839
rect 17586 2836 17592 2848
rect 16347 2808 17592 2836
rect 16347 2805 16359 2808
rect 16301 2799 16359 2805
rect 17586 2796 17592 2808
rect 17644 2836 17650 2848
rect 27816 2845 27844 2944
rect 30561 2941 30573 2944
rect 30607 2972 30619 2975
rect 45189 2975 45247 2981
rect 30607 2944 31754 2972
rect 30607 2941 30619 2944
rect 30561 2935 30619 2941
rect 22373 2839 22431 2845
rect 22373 2836 22385 2839
rect 17644 2808 22385 2836
rect 17644 2796 17650 2808
rect 22373 2805 22385 2808
rect 22419 2805 22431 2839
rect 22373 2799 22431 2805
rect 27801 2839 27859 2845
rect 27801 2805 27813 2839
rect 27847 2805 27859 2839
rect 31726 2836 31754 2944
rect 45189 2941 45201 2975
rect 45235 2972 45247 2975
rect 46750 2972 46756 2984
rect 45235 2944 46756 2972
rect 45235 2941 45247 2944
rect 45189 2935 45247 2941
rect 46750 2932 46756 2944
rect 46808 2932 46814 2984
rect 46842 2932 46848 2984
rect 46900 2932 46906 2984
rect 38286 2836 38292 2848
rect 31726 2808 38292 2836
rect 27801 2799 27859 2805
rect 38286 2796 38292 2808
rect 38344 2796 38350 2848
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 3053 2635 3111 2641
rect 3053 2601 3065 2635
rect 3099 2632 3111 2635
rect 6362 2632 6368 2644
rect 3099 2604 6368 2632
rect 3099 2601 3111 2604
rect 3053 2595 3111 2601
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 9766 2592 9772 2644
rect 9824 2592 9830 2644
rect 10042 2592 10048 2644
rect 10100 2632 10106 2644
rect 10873 2635 10931 2641
rect 10873 2632 10885 2635
rect 10100 2604 10885 2632
rect 10100 2592 10106 2604
rect 10873 2601 10885 2604
rect 10919 2601 10931 2635
rect 10873 2595 10931 2601
rect 24486 2592 24492 2644
rect 24544 2592 24550 2644
rect 25133 2635 25191 2641
rect 25133 2601 25145 2635
rect 25179 2632 25191 2635
rect 26326 2632 26332 2644
rect 25179 2604 26332 2632
rect 25179 2601 25191 2604
rect 25133 2595 25191 2601
rect 26326 2592 26332 2604
rect 26384 2592 26390 2644
rect 30834 2592 30840 2644
rect 30892 2592 30898 2644
rect 32858 2592 32864 2644
rect 32916 2632 32922 2644
rect 32953 2635 33011 2641
rect 32953 2632 32965 2635
rect 32916 2604 32965 2632
rect 32916 2592 32922 2604
rect 32953 2601 32965 2604
rect 32999 2601 33011 2635
rect 32953 2595 33011 2601
rect 34422 2592 34428 2644
rect 34480 2632 34486 2644
rect 35069 2635 35127 2641
rect 35069 2632 35081 2635
rect 34480 2604 35081 2632
rect 34480 2592 34486 2604
rect 35069 2601 35081 2604
rect 35115 2601 35127 2635
rect 48866 2632 48872 2644
rect 35069 2595 35127 2601
rect 35866 2604 48872 2632
rect 2501 2567 2559 2573
rect 2501 2533 2513 2567
rect 2547 2564 2559 2567
rect 16022 2564 16028 2576
rect 2547 2536 16028 2564
rect 2547 2533 2559 2536
rect 2501 2527 2559 2533
rect 16022 2524 16028 2536
rect 16080 2524 16086 2576
rect 20824 2536 22416 2564
rect 2774 2496 2780 2508
rect 1596 2468 2780 2496
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1596 2437 1624 2468
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 8573 2499 8631 2505
rect 8573 2465 8585 2499
rect 8619 2496 8631 2499
rect 9858 2496 9864 2508
rect 8619 2468 9864 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 9858 2456 9864 2468
rect 9916 2456 9922 2508
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 12253 2499 12311 2505
rect 12253 2496 12265 2499
rect 11756 2468 12265 2496
rect 11756 2456 11762 2468
rect 12253 2465 12265 2468
rect 12299 2465 12311 2499
rect 12253 2459 12311 2465
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 13872 2468 14749 2496
rect 13872 2456 13878 2468
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 14737 2459 14795 2465
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 1360 2400 1593 2428
rect 1360 2388 1366 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 2314 2388 2320 2440
rect 2372 2388 2378 2440
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3513 2431 3571 2437
rect 3513 2428 3525 2431
rect 3292 2400 3525 2428
rect 3292 2388 3298 2400
rect 3513 2397 3525 2400
rect 3559 2397 3571 2431
rect 3513 2391 3571 2397
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2428 7987 2431
rect 8754 2428 8760 2440
rect 7975 2400 8760 2428
rect 7975 2397 7987 2400
rect 7929 2391 7987 2397
rect 8754 2388 8760 2400
rect 8812 2388 8818 2440
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 9674 2428 9680 2440
rect 9171 2400 9680 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 10226 2388 10232 2440
rect 10284 2388 10290 2440
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2428 12035 2431
rect 12434 2428 12440 2440
rect 12023 2400 12440 2428
rect 12023 2397 12035 2400
rect 11977 2391 12035 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2428 14519 2431
rect 16390 2428 16396 2440
rect 14507 2400 16396 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 16390 2388 16396 2400
rect 16448 2388 16454 2440
rect 17681 2431 17739 2437
rect 17681 2397 17693 2431
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 20441 2431 20499 2437
rect 20441 2397 20453 2431
rect 20487 2428 20499 2431
rect 20824 2428 20852 2536
rect 20898 2456 20904 2508
rect 20956 2496 20962 2508
rect 22388 2505 22416 2536
rect 22462 2524 22468 2576
rect 22520 2564 22526 2576
rect 22520 2536 22784 2564
rect 22520 2524 22526 2536
rect 22189 2499 22247 2505
rect 22189 2496 22201 2499
rect 20956 2468 22201 2496
rect 20956 2456 20962 2468
rect 22189 2465 22201 2468
rect 22235 2465 22247 2499
rect 22189 2459 22247 2465
rect 22373 2499 22431 2505
rect 22373 2465 22385 2499
rect 22419 2496 22431 2499
rect 22646 2496 22652 2508
rect 22419 2468 22652 2496
rect 22419 2465 22431 2468
rect 22373 2459 22431 2465
rect 22646 2456 22652 2468
rect 22704 2456 22710 2508
rect 22756 2496 22784 2536
rect 24946 2524 24952 2576
rect 25004 2564 25010 2576
rect 28721 2567 28779 2573
rect 28721 2564 28733 2567
rect 25004 2536 28733 2564
rect 25004 2524 25010 2536
rect 28721 2533 28733 2536
rect 28767 2533 28779 2567
rect 28721 2527 28779 2533
rect 30742 2524 30748 2576
rect 30800 2564 30806 2576
rect 35866 2564 35894 2604
rect 48866 2592 48872 2604
rect 48924 2592 48930 2644
rect 30800 2536 35894 2564
rect 30800 2524 30806 2536
rect 25317 2499 25375 2505
rect 25317 2496 25329 2499
rect 22756 2468 25329 2496
rect 25317 2465 25329 2468
rect 25363 2465 25375 2499
rect 25317 2459 25375 2465
rect 36814 2456 36820 2508
rect 36872 2496 36878 2508
rect 37737 2499 37795 2505
rect 37737 2496 37749 2499
rect 36872 2468 37749 2496
rect 36872 2456 36878 2468
rect 37737 2465 37749 2468
rect 37783 2465 37795 2499
rect 37737 2459 37795 2465
rect 41322 2456 41328 2508
rect 41380 2496 41386 2508
rect 41417 2499 41475 2505
rect 41417 2496 41429 2499
rect 41380 2468 41429 2496
rect 41380 2456 41386 2468
rect 41417 2465 41429 2468
rect 41463 2465 41475 2499
rect 41417 2459 41475 2465
rect 44266 2456 44272 2508
rect 44324 2496 44330 2508
rect 44324 2468 47992 2496
rect 44324 2456 44330 2468
rect 20487 2400 20852 2428
rect 20487 2397 20499 2400
rect 20441 2391 20499 2397
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 2332 2360 2360 2388
rect 1268 2332 2360 2360
rect 1268 2320 1274 2332
rect 6362 2320 6368 2372
rect 6420 2360 6426 2372
rect 6420 2332 12434 2360
rect 6420 2320 6426 2332
rect 1765 2295 1823 2301
rect 1765 2261 1777 2295
rect 1811 2292 1823 2295
rect 6914 2292 6920 2304
rect 1811 2264 6920 2292
rect 1811 2261 1823 2264
rect 1765 2255 1823 2261
rect 6914 2252 6920 2264
rect 6972 2252 6978 2304
rect 12406 2292 12434 2332
rect 14182 2292 14188 2304
rect 12406 2264 14188 2292
rect 14182 2252 14188 2264
rect 14240 2252 14246 2304
rect 17696 2292 17724 2391
rect 23934 2388 23940 2440
rect 23992 2428 23998 2440
rect 24857 2431 24915 2437
rect 24857 2428 24869 2431
rect 23992 2400 24869 2428
rect 23992 2388 23998 2400
rect 24857 2397 24869 2400
rect 24903 2428 24915 2431
rect 27522 2428 27528 2440
rect 24903 2400 27528 2428
rect 24903 2397 24915 2400
rect 24857 2391 24915 2397
rect 27522 2388 27528 2400
rect 27580 2388 27586 2440
rect 28626 2388 28632 2440
rect 28684 2428 28690 2440
rect 28905 2431 28963 2437
rect 28905 2428 28917 2431
rect 28684 2400 28917 2428
rect 28684 2388 28690 2400
rect 28905 2397 28917 2400
rect 28951 2428 28963 2431
rect 29181 2431 29239 2437
rect 29181 2428 29193 2431
rect 28951 2400 29193 2428
rect 28951 2397 28963 2400
rect 28905 2391 28963 2397
rect 29181 2397 29193 2400
rect 29227 2397 29239 2431
rect 29181 2391 29239 2397
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30800 2400 31033 2428
rect 30800 2388 30806 2400
rect 31021 2397 31033 2400
rect 31067 2428 31079 2431
rect 31297 2431 31355 2437
rect 31297 2428 31309 2431
rect 31067 2400 31309 2428
rect 31067 2397 31079 2400
rect 31021 2391 31079 2397
rect 31297 2397 31309 2400
rect 31343 2397 31355 2431
rect 31297 2391 31355 2397
rect 33134 2388 33140 2440
rect 33192 2428 33198 2440
rect 33413 2431 33471 2437
rect 33413 2428 33425 2431
rect 33192 2400 33425 2428
rect 33192 2388 33198 2400
rect 33413 2397 33425 2400
rect 33459 2397 33471 2431
rect 33413 2391 33471 2397
rect 34974 2388 34980 2440
rect 35032 2428 35038 2440
rect 35253 2431 35311 2437
rect 35253 2428 35265 2431
rect 35032 2400 35265 2428
rect 35032 2388 35038 2400
rect 35253 2397 35265 2400
rect 35299 2428 35311 2431
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 35299 2400 35541 2428
rect 35299 2397 35311 2400
rect 35253 2391 35311 2397
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 35529 2391 35587 2397
rect 37108 2400 37473 2428
rect 18322 2320 18328 2372
rect 18380 2360 18386 2372
rect 18417 2363 18475 2369
rect 18417 2360 18429 2363
rect 18380 2332 18429 2360
rect 18380 2320 18386 2332
rect 18417 2329 18429 2332
rect 18463 2329 18475 2363
rect 18417 2323 18475 2329
rect 24029 2363 24087 2369
rect 24029 2329 24041 2363
rect 24075 2360 24087 2363
rect 26510 2360 26516 2372
rect 24075 2332 26516 2360
rect 24075 2329 24087 2332
rect 24029 2323 24087 2329
rect 26510 2320 26516 2332
rect 26568 2320 26574 2372
rect 37108 2304 37136 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 38286 2388 38292 2440
rect 38344 2428 38350 2440
rect 40681 2431 40739 2437
rect 40681 2428 40693 2431
rect 38344 2400 40693 2428
rect 38344 2388 38350 2400
rect 40681 2397 40693 2400
rect 40727 2397 40739 2431
rect 40681 2391 40739 2397
rect 42794 2388 42800 2440
rect 42852 2428 42858 2440
rect 47964 2437 47992 2468
rect 49142 2456 49148 2508
rect 49200 2456 49206 2508
rect 45833 2431 45891 2437
rect 45833 2428 45845 2431
rect 42852 2400 45845 2428
rect 42852 2388 42858 2400
rect 45833 2397 45845 2400
rect 45879 2397 45891 2431
rect 45833 2391 45891 2397
rect 47949 2431 48007 2437
rect 47949 2397 47961 2431
rect 47995 2397 48007 2431
rect 47949 2391 48007 2397
rect 47029 2363 47087 2369
rect 47029 2329 47041 2363
rect 47075 2360 47087 2363
rect 48498 2360 48504 2372
rect 47075 2332 48504 2360
rect 47075 2329 47087 2332
rect 47029 2323 47087 2329
rect 48498 2320 48504 2332
rect 48556 2320 48562 2372
rect 20257 2295 20315 2301
rect 20257 2292 20269 2295
rect 17696 2264 20269 2292
rect 20257 2261 20269 2264
rect 20303 2261 20315 2295
rect 20257 2255 20315 2261
rect 37090 2252 37096 2304
rect 37148 2252 37154 2304
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
rect 8754 1708 8760 1760
rect 8812 1748 8818 1760
rect 9582 1748 9588 1760
rect 8812 1720 9588 1748
rect 8812 1708 8818 1720
rect 9582 1708 9588 1720
rect 9640 1708 9646 1760
<< via1 >>
rect 24216 26324 24268 26376
rect 43812 26324 43864 26376
rect 12256 26256 12308 26308
rect 26332 26256 26384 26308
rect 33508 26188 33560 26240
rect 47216 26188 47268 26240
rect 35808 26120 35860 26172
rect 47492 26120 47544 26172
rect 28356 26052 28408 26104
rect 43352 26052 43404 26104
rect 21180 25984 21232 26036
rect 47124 25984 47176 26036
rect 19708 25916 19760 25968
rect 45560 25916 45612 25968
rect 26884 25848 26936 25900
rect 45192 25848 45244 25900
rect 24308 25780 24360 25832
rect 40868 25780 40920 25832
rect 21732 25712 21784 25764
rect 49240 25712 49292 25764
rect 4344 25644 4396 25696
rect 44180 25644 44232 25696
rect 20352 25576 20404 25628
rect 48780 25576 48832 25628
rect 12072 25508 12124 25560
rect 44456 25508 44508 25560
rect 25136 25440 25188 25492
rect 41880 25440 41932 25492
rect 27252 25372 27304 25424
rect 44364 25372 44416 25424
rect 30564 25304 30616 25356
rect 49056 25304 49108 25356
rect 17316 25236 17368 25288
rect 40316 25236 40368 25288
rect 4068 25168 4120 25220
rect 8852 25168 8904 25220
rect 35900 25168 35952 25220
rect 42524 25168 42576 25220
rect 28264 25100 28316 25152
rect 41420 25100 41472 25152
rect 15016 25032 15068 25084
rect 31760 25032 31812 25084
rect 32220 25032 32272 25084
rect 41972 25032 42024 25084
rect 15200 24964 15252 25016
rect 27068 24964 27120 25016
rect 41328 24964 41380 25016
rect 45836 24964 45888 25016
rect 4712 24896 4764 24948
rect 3424 24828 3476 24880
rect 9864 24828 9916 24880
rect 12716 24896 12768 24948
rect 33508 24896 33560 24948
rect 19892 24828 19944 24880
rect 24584 24828 24636 24880
rect 3700 24760 3752 24812
rect 6276 24760 6328 24812
rect 30932 24760 30984 24812
rect 33968 24760 34020 24812
rect 36820 24828 36872 24880
rect 43444 24828 43496 24880
rect 47768 24760 47820 24812
rect 11796 24692 11848 24744
rect 23388 24692 23440 24744
rect 30012 24692 30064 24744
rect 42800 24692 42852 24744
rect 14188 24624 14240 24676
rect 24860 24624 24912 24676
rect 1768 24556 1820 24608
rect 11336 24556 11388 24608
rect 14832 24556 14884 24608
rect 21364 24556 21416 24608
rect 23664 24556 23716 24608
rect 34152 24624 34204 24676
rect 35532 24624 35584 24676
rect 37556 24624 37608 24676
rect 40684 24624 40736 24676
rect 25964 24556 26016 24608
rect 30840 24556 30892 24608
rect 31300 24556 31352 24608
rect 37464 24556 37516 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 1768 24395 1820 24404
rect 1768 24361 1777 24395
rect 1777 24361 1811 24395
rect 1811 24361 1820 24395
rect 1768 24352 1820 24361
rect 2320 24352 2372 24404
rect 3516 24216 3568 24268
rect 2136 24191 2188 24200
rect 2136 24157 2145 24191
rect 2145 24157 2179 24191
rect 2179 24157 2188 24191
rect 2136 24148 2188 24157
rect 2412 24148 2464 24200
rect 3608 24080 3660 24132
rect 4252 24148 4304 24200
rect 10508 24352 10560 24404
rect 6736 24284 6788 24336
rect 10140 24284 10192 24336
rect 11612 24284 11664 24336
rect 19432 24352 19484 24404
rect 8668 24216 8720 24268
rect 8944 24216 8996 24268
rect 3700 24012 3752 24064
rect 4068 24012 4120 24064
rect 9036 24148 9088 24200
rect 12440 24216 12492 24268
rect 14464 24216 14516 24268
rect 19248 24216 19300 24268
rect 27528 24352 27580 24404
rect 31852 24352 31904 24404
rect 32128 24352 32180 24404
rect 21180 24327 21232 24336
rect 21180 24293 21189 24327
rect 21189 24293 21223 24327
rect 21223 24293 21232 24327
rect 21180 24284 21232 24293
rect 24400 24284 24452 24336
rect 34152 24395 34204 24404
rect 34152 24361 34161 24395
rect 34161 24361 34195 24395
rect 34195 24361 34204 24395
rect 34152 24352 34204 24361
rect 37464 24395 37516 24404
rect 37464 24361 37473 24395
rect 37473 24361 37507 24395
rect 37507 24361 37516 24395
rect 37464 24352 37516 24361
rect 40684 24352 40736 24404
rect 14004 24148 14056 24200
rect 15200 24148 15252 24200
rect 10784 24080 10836 24132
rect 11704 24123 11756 24132
rect 11704 24089 11713 24123
rect 11713 24089 11747 24123
rect 11747 24089 11756 24123
rect 11704 24080 11756 24089
rect 12164 24080 12216 24132
rect 16948 24148 17000 24200
rect 17132 24148 17184 24200
rect 21272 24216 21324 24268
rect 9312 24012 9364 24064
rect 9404 24055 9456 24064
rect 9404 24021 9413 24055
rect 9413 24021 9447 24055
rect 9447 24021 9456 24055
rect 9404 24012 9456 24021
rect 11428 24012 11480 24064
rect 18328 24080 18380 24132
rect 19248 24080 19300 24132
rect 22100 24191 22152 24200
rect 22100 24157 22109 24191
rect 22109 24157 22143 24191
rect 22143 24157 22152 24191
rect 22100 24148 22152 24157
rect 25412 24216 25464 24268
rect 28448 24259 28500 24268
rect 28448 24225 28457 24259
rect 28457 24225 28491 24259
rect 28491 24225 28500 24259
rect 28448 24216 28500 24225
rect 28724 24216 28776 24268
rect 24860 24191 24912 24200
rect 24860 24157 24869 24191
rect 24869 24157 24903 24191
rect 24903 24157 24912 24191
rect 24860 24148 24912 24157
rect 25964 24191 26016 24200
rect 25964 24157 25973 24191
rect 25973 24157 26007 24191
rect 26007 24157 26016 24191
rect 25964 24148 26016 24157
rect 27436 24148 27488 24200
rect 28264 24191 28316 24200
rect 28264 24157 28273 24191
rect 28273 24157 28307 24191
rect 28307 24157 28316 24191
rect 28264 24148 28316 24157
rect 29184 24191 29236 24200
rect 29184 24157 29193 24191
rect 29193 24157 29227 24191
rect 29227 24157 29236 24191
rect 29184 24148 29236 24157
rect 29460 24148 29512 24200
rect 30012 24148 30064 24200
rect 19708 24123 19760 24132
rect 19708 24089 19717 24123
rect 19717 24089 19751 24123
rect 19751 24089 19760 24123
rect 19708 24080 19760 24089
rect 19984 24080 20036 24132
rect 16764 24012 16816 24064
rect 21272 24012 21324 24064
rect 23848 24055 23900 24064
rect 23848 24021 23857 24055
rect 23857 24021 23891 24055
rect 23891 24021 23900 24055
rect 23848 24012 23900 24021
rect 24492 24055 24544 24064
rect 24492 24021 24501 24055
rect 24501 24021 24535 24055
rect 24535 24021 24544 24055
rect 24492 24012 24544 24021
rect 30472 24080 30524 24132
rect 34980 24216 35032 24268
rect 35532 24259 35584 24268
rect 35532 24225 35541 24259
rect 35541 24225 35575 24259
rect 35575 24225 35584 24259
rect 35532 24216 35584 24225
rect 35808 24216 35860 24268
rect 36820 24216 36872 24268
rect 38660 24216 38712 24268
rect 39948 24284 40000 24336
rect 39396 24216 39448 24268
rect 40684 24259 40736 24268
rect 40684 24225 40693 24259
rect 40693 24225 40727 24259
rect 40727 24225 40736 24259
rect 40684 24216 40736 24225
rect 33508 24191 33560 24200
rect 33508 24157 33517 24191
rect 33517 24157 33551 24191
rect 33551 24157 33560 24191
rect 33508 24148 33560 24157
rect 35256 24148 35308 24200
rect 35624 24148 35676 24200
rect 39672 24148 39724 24200
rect 41420 24216 41472 24268
rect 42800 24352 42852 24404
rect 45744 24352 45796 24404
rect 47216 24395 47268 24404
rect 47216 24361 47225 24395
rect 47225 24361 47259 24395
rect 47259 24361 47268 24395
rect 47216 24352 47268 24361
rect 44088 24284 44140 24336
rect 46204 24216 46256 24268
rect 25228 24012 25280 24064
rect 29000 24055 29052 24064
rect 29000 24021 29009 24055
rect 29009 24021 29043 24055
rect 29043 24021 29052 24055
rect 29000 24012 29052 24021
rect 30288 24012 30340 24064
rect 30380 24055 30432 24064
rect 30380 24021 30389 24055
rect 30389 24021 30423 24055
rect 30423 24021 30432 24055
rect 30380 24012 30432 24021
rect 31116 24012 31168 24064
rect 32312 24055 32364 24064
rect 32312 24021 32321 24055
rect 32321 24021 32355 24055
rect 32355 24021 32364 24055
rect 32312 24012 32364 24021
rect 33140 24012 33192 24064
rect 33968 24012 34020 24064
rect 35716 24012 35768 24064
rect 36452 24055 36504 24064
rect 36452 24021 36461 24055
rect 36461 24021 36495 24055
rect 36495 24021 36504 24055
rect 36452 24012 36504 24021
rect 36544 24012 36596 24064
rect 41696 24080 41748 24132
rect 42708 24148 42760 24200
rect 45652 24148 45704 24200
rect 46296 24191 46348 24200
rect 46296 24157 46305 24191
rect 46305 24157 46339 24191
rect 46339 24157 46348 24191
rect 46296 24148 46348 24157
rect 40408 24055 40460 24064
rect 40408 24021 40417 24055
rect 40417 24021 40451 24055
rect 40451 24021 40460 24055
rect 40408 24012 40460 24021
rect 41144 24012 41196 24064
rect 43720 24012 43772 24064
rect 43812 24012 43864 24064
rect 48780 24259 48832 24268
rect 48780 24225 48789 24259
rect 48789 24225 48823 24259
rect 48823 24225 48832 24259
rect 48780 24216 48832 24225
rect 46848 24080 46900 24132
rect 46664 24012 46716 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 2320 23851 2372 23860
rect 2320 23817 2329 23851
rect 2329 23817 2363 23851
rect 2363 23817 2372 23851
rect 2320 23808 2372 23817
rect 3608 23808 3660 23860
rect 4160 23740 4212 23792
rect 6460 23808 6512 23860
rect 18788 23808 18840 23860
rect 8760 23740 8812 23792
rect 9128 23783 9180 23792
rect 9128 23749 9137 23783
rect 9137 23749 9171 23783
rect 9171 23749 9180 23783
rect 9128 23740 9180 23749
rect 10692 23783 10744 23792
rect 10692 23749 10701 23783
rect 10701 23749 10735 23783
rect 10735 23749 10744 23783
rect 10692 23740 10744 23749
rect 15108 23740 15160 23792
rect 17040 23740 17092 23792
rect 3884 23672 3936 23724
rect 4804 23715 4856 23724
rect 4804 23681 4813 23715
rect 4813 23681 4847 23715
rect 4847 23681 4856 23715
rect 4804 23672 4856 23681
rect 6552 23715 6604 23724
rect 6552 23681 6561 23715
rect 6561 23681 6595 23715
rect 6595 23681 6604 23715
rect 6552 23672 6604 23681
rect 9220 23672 9272 23724
rect 4160 23604 4212 23656
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 6920 23604 6972 23656
rect 3700 23536 3752 23588
rect 5632 23536 5684 23588
rect 11796 23715 11848 23724
rect 11796 23681 11805 23715
rect 11805 23681 11839 23715
rect 11839 23681 11848 23715
rect 11796 23672 11848 23681
rect 12072 23715 12124 23724
rect 12072 23681 12081 23715
rect 12081 23681 12115 23715
rect 12115 23681 12124 23715
rect 12072 23672 12124 23681
rect 14648 23672 14700 23724
rect 15016 23715 15068 23724
rect 15016 23681 15025 23715
rect 15025 23681 15059 23715
rect 15059 23681 15068 23715
rect 15016 23672 15068 23681
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 17316 23715 17368 23724
rect 17316 23681 17325 23715
rect 17325 23681 17359 23715
rect 17359 23681 17368 23715
rect 17316 23672 17368 23681
rect 18972 23783 19024 23792
rect 18972 23749 18981 23783
rect 18981 23749 19015 23783
rect 19015 23749 19024 23783
rect 18972 23740 19024 23749
rect 19984 23740 20036 23792
rect 21364 23808 21416 23860
rect 23848 23808 23900 23860
rect 11428 23604 11480 23656
rect 19248 23604 19300 23656
rect 21180 23604 21232 23656
rect 16672 23536 16724 23588
rect 16764 23536 16816 23588
rect 19524 23536 19576 23588
rect 23204 23672 23256 23724
rect 22468 23647 22520 23656
rect 22468 23613 22477 23647
rect 22477 23613 22511 23647
rect 22511 23613 22520 23647
rect 22468 23604 22520 23613
rect 24952 23808 25004 23860
rect 25044 23808 25096 23860
rect 27896 23808 27948 23860
rect 30656 23851 30708 23860
rect 30656 23817 30665 23851
rect 30665 23817 30699 23851
rect 30699 23817 30708 23851
rect 30656 23808 30708 23817
rect 31392 23808 31444 23860
rect 36544 23808 36596 23860
rect 37832 23808 37884 23860
rect 37924 23808 37976 23860
rect 41880 23851 41932 23860
rect 41880 23817 41889 23851
rect 41889 23817 41923 23851
rect 41923 23817 41932 23851
rect 41880 23808 41932 23817
rect 42248 23851 42300 23860
rect 42248 23817 42257 23851
rect 42257 23817 42291 23851
rect 42291 23817 42300 23851
rect 42248 23808 42300 23817
rect 22652 23536 22704 23588
rect 2780 23468 2832 23520
rect 6184 23468 6236 23520
rect 10784 23468 10836 23520
rect 12532 23468 12584 23520
rect 17500 23468 17552 23520
rect 21364 23511 21416 23520
rect 21364 23477 21373 23511
rect 21373 23477 21407 23511
rect 21407 23477 21416 23511
rect 21364 23468 21416 23477
rect 23572 23468 23624 23520
rect 26424 23740 26476 23792
rect 27528 23740 27580 23792
rect 31760 23783 31812 23792
rect 31760 23749 31769 23783
rect 31769 23749 31803 23783
rect 31803 23749 31812 23783
rect 31760 23740 31812 23749
rect 32680 23740 32732 23792
rect 34060 23740 34112 23792
rect 45192 23851 45244 23860
rect 45192 23817 45201 23851
rect 45201 23817 45235 23851
rect 45235 23817 45244 23851
rect 45192 23808 45244 23817
rect 47768 23808 47820 23860
rect 24216 23715 24268 23724
rect 24216 23681 24225 23715
rect 24225 23681 24259 23715
rect 24259 23681 24268 23715
rect 24216 23672 24268 23681
rect 24860 23647 24912 23656
rect 24860 23613 24869 23647
rect 24869 23613 24903 23647
rect 24903 23613 24912 23647
rect 24860 23604 24912 23613
rect 27804 23672 27856 23724
rect 27712 23604 27764 23656
rect 28356 23604 28408 23656
rect 30380 23672 30432 23724
rect 30104 23604 30156 23656
rect 31576 23715 31628 23724
rect 31576 23681 31585 23715
rect 31585 23681 31619 23715
rect 31619 23681 31628 23715
rect 31576 23672 31628 23681
rect 32404 23672 32456 23724
rect 33232 23672 33284 23724
rect 36360 23715 36412 23724
rect 36360 23681 36369 23715
rect 36369 23681 36403 23715
rect 36403 23681 36412 23715
rect 36360 23672 36412 23681
rect 38844 23672 38896 23724
rect 26792 23468 26844 23520
rect 27160 23511 27212 23520
rect 27160 23477 27169 23511
rect 27169 23477 27203 23511
rect 27203 23477 27212 23511
rect 27160 23468 27212 23477
rect 30932 23647 30984 23656
rect 30932 23613 30941 23647
rect 30941 23613 30975 23647
rect 30975 23613 30984 23647
rect 30932 23604 30984 23613
rect 33140 23604 33192 23656
rect 34336 23604 34388 23656
rect 35072 23604 35124 23656
rect 36452 23647 36504 23656
rect 36452 23613 36461 23647
rect 36461 23613 36495 23647
rect 36495 23613 36504 23647
rect 36452 23604 36504 23613
rect 37188 23604 37240 23656
rect 37464 23647 37516 23656
rect 37464 23613 37473 23647
rect 37473 23613 37507 23647
rect 37507 23613 37516 23647
rect 37464 23604 37516 23613
rect 39948 23672 40000 23724
rect 41052 23672 41104 23724
rect 33048 23536 33100 23588
rect 34704 23536 34756 23588
rect 35624 23536 35676 23588
rect 39856 23604 39908 23656
rect 40684 23647 40736 23656
rect 40684 23613 40693 23647
rect 40693 23613 40727 23647
rect 40727 23613 40736 23647
rect 40684 23604 40736 23613
rect 40776 23604 40828 23656
rect 45468 23740 45520 23792
rect 43720 23715 43772 23724
rect 43720 23681 43729 23715
rect 43729 23681 43763 23715
rect 43763 23681 43772 23715
rect 43720 23672 43772 23681
rect 44364 23715 44416 23724
rect 44364 23681 44373 23715
rect 44373 23681 44407 23715
rect 44407 23681 44416 23715
rect 44364 23672 44416 23681
rect 44548 23672 44600 23724
rect 44732 23672 44784 23724
rect 29736 23511 29788 23520
rect 29736 23477 29745 23511
rect 29745 23477 29779 23511
rect 29779 23477 29788 23511
rect 29736 23468 29788 23477
rect 30012 23511 30064 23520
rect 30012 23477 30021 23511
rect 30021 23477 30055 23511
rect 30055 23477 30064 23511
rect 30012 23468 30064 23477
rect 30380 23468 30432 23520
rect 30840 23468 30892 23520
rect 32772 23511 32824 23520
rect 32772 23477 32781 23511
rect 32781 23477 32815 23511
rect 32815 23477 32824 23511
rect 32772 23468 32824 23477
rect 33232 23468 33284 23520
rect 34888 23468 34940 23520
rect 34980 23468 35032 23520
rect 41236 23536 41288 23588
rect 45560 23672 45612 23724
rect 47216 23715 47268 23724
rect 47216 23681 47225 23715
rect 47225 23681 47259 23715
rect 47259 23681 47268 23715
rect 47216 23672 47268 23681
rect 45744 23647 45796 23656
rect 45744 23613 45753 23647
rect 45753 23613 45787 23647
rect 45787 23613 45796 23647
rect 45744 23604 45796 23613
rect 36912 23468 36964 23520
rect 37280 23468 37332 23520
rect 40776 23468 40828 23520
rect 42708 23468 42760 23520
rect 47584 23536 47636 23588
rect 47400 23468 47452 23520
rect 49148 23672 49200 23724
rect 47768 23604 47820 23656
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 14556 23264 14608 23316
rect 14648 23307 14700 23316
rect 14648 23273 14657 23307
rect 14657 23273 14691 23307
rect 14691 23273 14700 23307
rect 14648 23264 14700 23273
rect 14740 23264 14792 23316
rect 17224 23264 17276 23316
rect 17868 23264 17920 23316
rect 3424 23239 3476 23248
rect 3424 23205 3433 23239
rect 3433 23205 3467 23239
rect 3467 23205 3476 23239
rect 3424 23196 3476 23205
rect 4804 23196 4856 23248
rect 2872 23128 2924 23180
rect 4436 23128 4488 23180
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 11244 23171 11296 23180
rect 11244 23137 11253 23171
rect 11253 23137 11287 23171
rect 11287 23137 11296 23171
rect 11244 23128 11296 23137
rect 1768 23103 1820 23112
rect 1768 23069 1777 23103
rect 1777 23069 1811 23103
rect 1811 23069 1820 23103
rect 1768 23060 1820 23069
rect 4252 23103 4304 23112
rect 4252 23069 4261 23103
rect 4261 23069 4295 23103
rect 4295 23069 4304 23103
rect 4252 23060 4304 23069
rect 4344 23060 4396 23112
rect 7472 23060 7524 23112
rect 8300 23060 8352 23112
rect 10508 23103 10560 23112
rect 10508 23069 10517 23103
rect 10517 23069 10551 23103
rect 10551 23069 10560 23103
rect 10508 23060 10560 23069
rect 2780 23035 2832 23044
rect 2780 23001 2789 23035
rect 2789 23001 2823 23035
rect 2823 23001 2832 23035
rect 2780 22992 2832 23001
rect 3240 22992 3292 23044
rect 6736 22992 6788 23044
rect 13360 23171 13412 23180
rect 13360 23137 13369 23171
rect 13369 23137 13403 23171
rect 13403 23137 13412 23171
rect 13360 23128 13412 23137
rect 17040 23196 17092 23248
rect 15752 23128 15804 23180
rect 16396 23171 16448 23180
rect 16396 23137 16405 23171
rect 16405 23137 16439 23171
rect 16439 23137 16448 23171
rect 16396 23128 16448 23137
rect 16764 23128 16816 23180
rect 14556 23060 14608 23112
rect 16580 23060 16632 23112
rect 17132 23103 17184 23112
rect 17132 23069 17141 23103
rect 17141 23069 17175 23103
rect 17175 23069 17184 23103
rect 17132 23060 17184 23069
rect 18512 23060 18564 23112
rect 7748 22924 7800 22976
rect 9680 22924 9732 22976
rect 20260 23264 20312 23316
rect 22468 23264 22520 23316
rect 22652 23264 22704 23316
rect 26056 23264 26108 23316
rect 29276 23264 29328 23316
rect 30932 23264 30984 23316
rect 24124 23196 24176 23248
rect 24492 23196 24544 23248
rect 26700 23196 26752 23248
rect 21180 23128 21232 23180
rect 22376 23128 22428 23180
rect 23940 23128 23992 23180
rect 27252 23128 27304 23180
rect 27620 23196 27672 23248
rect 28816 23196 28868 23248
rect 36820 23264 36872 23316
rect 42340 23264 42392 23316
rect 44180 23264 44232 23316
rect 46296 23264 46348 23316
rect 46388 23264 46440 23316
rect 47308 23264 47360 23316
rect 47860 23264 47912 23316
rect 48780 23264 48832 23316
rect 27896 23128 27948 23180
rect 28448 23128 28500 23180
rect 29092 23171 29144 23180
rect 29092 23137 29101 23171
rect 29101 23137 29135 23171
rect 29135 23137 29144 23171
rect 29092 23128 29144 23137
rect 22928 23060 22980 23112
rect 24768 23060 24820 23112
rect 28080 23103 28132 23112
rect 28080 23069 28089 23103
rect 28089 23069 28123 23103
rect 28123 23069 28132 23103
rect 28080 23060 28132 23069
rect 28540 23060 28592 23112
rect 28632 23060 28684 23112
rect 33416 23128 33468 23180
rect 20812 22992 20864 23044
rect 21088 23035 21140 23044
rect 21088 23001 21097 23035
rect 21097 23001 21131 23035
rect 21131 23001 21140 23035
rect 21088 22992 21140 23001
rect 16764 22924 16816 22976
rect 18328 22924 18380 22976
rect 19984 22924 20036 22976
rect 22744 22992 22796 23044
rect 25320 22992 25372 23044
rect 27344 22992 27396 23044
rect 26516 22924 26568 22976
rect 27160 22967 27212 22976
rect 27160 22933 27169 22967
rect 27169 22933 27203 22967
rect 27203 22933 27212 22967
rect 27160 22924 27212 22933
rect 27620 22967 27672 22976
rect 27620 22933 27629 22967
rect 27629 22933 27663 22967
rect 27663 22933 27672 22967
rect 27620 22924 27672 22933
rect 28908 23035 28960 23044
rect 28908 23001 28917 23035
rect 28917 23001 28951 23035
rect 28951 23001 28960 23035
rect 28908 22992 28960 23001
rect 29644 22967 29696 22976
rect 29644 22933 29653 22967
rect 29653 22933 29687 22967
rect 29687 22933 29696 22967
rect 29644 22924 29696 22933
rect 30196 23035 30248 23044
rect 30196 23001 30205 23035
rect 30205 23001 30239 23035
rect 30239 23001 30248 23035
rect 30196 22992 30248 23001
rect 30840 22924 30892 22976
rect 32680 22992 32732 23044
rect 31760 22924 31812 22976
rect 32772 22924 32824 22976
rect 33324 22924 33376 22976
rect 34060 23196 34112 23248
rect 34152 23196 34204 23248
rect 36268 23196 36320 23248
rect 38660 23196 38712 23248
rect 39764 23196 39816 23248
rect 40408 23196 40460 23248
rect 40960 23196 41012 23248
rect 46940 23239 46992 23248
rect 46940 23205 46949 23239
rect 46949 23205 46983 23239
rect 46983 23205 46992 23239
rect 46940 23196 46992 23205
rect 47124 23196 47176 23248
rect 34612 23128 34664 23180
rect 34888 23171 34940 23180
rect 34888 23137 34897 23171
rect 34897 23137 34931 23171
rect 34931 23137 34940 23171
rect 34888 23128 34940 23137
rect 37464 23128 37516 23180
rect 42616 23128 42668 23180
rect 43444 23128 43496 23180
rect 45100 23128 45152 23180
rect 46664 23128 46716 23180
rect 38844 23060 38896 23112
rect 39488 23103 39540 23112
rect 39488 23069 39497 23103
rect 39497 23069 39531 23103
rect 39531 23069 39540 23103
rect 39488 23060 39540 23069
rect 40040 23103 40092 23112
rect 40040 23069 40049 23103
rect 40049 23069 40083 23103
rect 40083 23069 40092 23103
rect 40040 23060 40092 23069
rect 40316 23103 40368 23112
rect 40316 23069 40325 23103
rect 40325 23069 40359 23103
rect 40359 23069 40368 23103
rect 40316 23060 40368 23069
rect 44456 23060 44508 23112
rect 45192 23103 45244 23112
rect 45192 23069 45201 23103
rect 45201 23069 45235 23103
rect 45235 23069 45244 23103
rect 45192 23060 45244 23069
rect 46848 23060 46900 23112
rect 47124 23060 47176 23112
rect 48872 23060 48924 23112
rect 34520 22992 34572 23044
rect 36544 22992 36596 23044
rect 38660 22992 38712 23044
rect 33692 22924 33744 22976
rect 35532 22924 35584 22976
rect 37096 22924 37148 22976
rect 38384 22924 38436 22976
rect 38936 22924 38988 22976
rect 40960 22924 41012 22976
rect 42064 22924 42116 22976
rect 43260 22992 43312 23044
rect 43720 23035 43772 23044
rect 43720 23001 43729 23035
rect 43729 23001 43763 23035
rect 43763 23001 43772 23035
rect 43720 22992 43772 23001
rect 47032 22992 47084 23044
rect 43996 22924 44048 22976
rect 44824 22967 44876 22976
rect 44824 22933 44833 22967
rect 44833 22933 44867 22967
rect 44867 22933 44876 22967
rect 44824 22924 44876 22933
rect 49424 22967 49476 22976
rect 49424 22933 49433 22967
rect 49433 22933 49467 22967
rect 49467 22933 49476 22967
rect 49424 22924 49476 22933
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 4160 22763 4212 22772
rect 4160 22729 4169 22763
rect 4169 22729 4203 22763
rect 4203 22729 4212 22763
rect 4160 22720 4212 22729
rect 7288 22720 7340 22772
rect 7564 22720 7616 22772
rect 9312 22763 9364 22772
rect 9312 22729 9321 22763
rect 9321 22729 9355 22763
rect 9355 22729 9364 22763
rect 9312 22720 9364 22729
rect 6368 22652 6420 22704
rect 6828 22695 6880 22704
rect 6828 22661 6837 22695
rect 6837 22661 6871 22695
rect 6871 22661 6880 22695
rect 6828 22652 6880 22661
rect 7012 22695 7064 22704
rect 7012 22661 7021 22695
rect 7021 22661 7055 22695
rect 7055 22661 7064 22695
rect 7012 22652 7064 22661
rect 3516 22627 3568 22636
rect 3516 22593 3525 22627
rect 3525 22593 3559 22627
rect 3559 22593 3568 22627
rect 3516 22584 3568 22593
rect 2872 22516 2924 22568
rect 1952 22448 2004 22500
rect 5080 22559 5132 22568
rect 5080 22525 5089 22559
rect 5089 22525 5123 22559
rect 5123 22525 5132 22559
rect 5080 22516 5132 22525
rect 6644 22516 6696 22568
rect 11060 22652 11112 22704
rect 7840 22584 7892 22636
rect 9772 22627 9824 22636
rect 9772 22593 9781 22627
rect 9781 22593 9815 22627
rect 9815 22593 9824 22627
rect 9772 22584 9824 22593
rect 7380 22516 7432 22568
rect 8024 22516 8076 22568
rect 12716 22584 12768 22636
rect 10232 22559 10284 22568
rect 10232 22525 10241 22559
rect 10241 22525 10275 22559
rect 10275 22525 10284 22559
rect 10232 22516 10284 22525
rect 11704 22559 11756 22568
rect 11704 22525 11713 22559
rect 11713 22525 11747 22559
rect 11747 22525 11756 22559
rect 11704 22516 11756 22525
rect 12256 22516 12308 22568
rect 13820 22559 13872 22568
rect 13820 22525 13829 22559
rect 13829 22525 13863 22559
rect 13863 22525 13872 22559
rect 13820 22516 13872 22525
rect 15844 22695 15896 22704
rect 15844 22661 15853 22695
rect 15853 22661 15887 22695
rect 15887 22661 15896 22695
rect 15844 22652 15896 22661
rect 15108 22627 15160 22636
rect 15108 22593 15117 22627
rect 15117 22593 15151 22627
rect 15151 22593 15160 22627
rect 15108 22584 15160 22593
rect 4988 22448 5040 22500
rect 1584 22380 1636 22432
rect 4528 22380 4580 22432
rect 7380 22380 7432 22432
rect 8024 22380 8076 22432
rect 13912 22448 13964 22500
rect 16028 22448 16080 22500
rect 16304 22380 16356 22432
rect 17132 22720 17184 22772
rect 19248 22720 19300 22772
rect 19616 22720 19668 22772
rect 17868 22652 17920 22704
rect 18512 22584 18564 22636
rect 19984 22652 20036 22704
rect 20812 22652 20864 22704
rect 23020 22720 23072 22772
rect 27620 22720 27672 22772
rect 25044 22652 25096 22704
rect 25136 22695 25188 22704
rect 25136 22661 25145 22695
rect 25145 22661 25179 22695
rect 25179 22661 25188 22695
rect 25136 22652 25188 22661
rect 26424 22652 26476 22704
rect 27344 22652 27396 22704
rect 29184 22720 29236 22772
rect 30012 22720 30064 22772
rect 30196 22720 30248 22772
rect 30472 22720 30524 22772
rect 32588 22720 32640 22772
rect 19248 22627 19300 22636
rect 19248 22593 19257 22627
rect 19257 22593 19291 22627
rect 19291 22593 19300 22627
rect 19248 22584 19300 22593
rect 23296 22584 23348 22636
rect 24400 22584 24452 22636
rect 27620 22584 27672 22636
rect 27804 22584 27856 22636
rect 16856 22559 16908 22568
rect 16856 22525 16865 22559
rect 16865 22525 16899 22559
rect 16899 22525 16908 22559
rect 16856 22516 16908 22525
rect 18144 22516 18196 22568
rect 20904 22516 20956 22568
rect 21272 22559 21324 22568
rect 21272 22525 21281 22559
rect 21281 22525 21315 22559
rect 21315 22525 21324 22559
rect 21272 22516 21324 22525
rect 21364 22516 21416 22568
rect 22192 22516 22244 22568
rect 23388 22516 23440 22568
rect 18604 22423 18656 22432
rect 18604 22389 18613 22423
rect 18613 22389 18647 22423
rect 18647 22389 18656 22423
rect 18604 22380 18656 22389
rect 18880 22423 18932 22432
rect 18880 22389 18889 22423
rect 18889 22389 18923 22423
rect 18923 22389 18932 22423
rect 18880 22380 18932 22389
rect 23480 22448 23532 22500
rect 21364 22380 21416 22432
rect 22376 22380 22428 22432
rect 23664 22423 23716 22432
rect 23664 22389 23673 22423
rect 23673 22389 23707 22423
rect 23707 22389 23716 22423
rect 23664 22380 23716 22389
rect 24308 22516 24360 22568
rect 24768 22516 24820 22568
rect 28632 22652 28684 22704
rect 32128 22652 32180 22704
rect 35164 22652 35216 22704
rect 36544 22652 36596 22704
rect 39028 22652 39080 22704
rect 39396 22652 39448 22704
rect 39672 22763 39724 22772
rect 39672 22729 39681 22763
rect 39681 22729 39715 22763
rect 39715 22729 39724 22763
rect 39672 22720 39724 22729
rect 40132 22652 40184 22704
rect 28356 22559 28408 22568
rect 28356 22525 28365 22559
rect 28365 22525 28399 22559
rect 28399 22525 28408 22559
rect 28356 22516 28408 22525
rect 29092 22516 29144 22568
rect 30656 22627 30708 22636
rect 30656 22593 30665 22627
rect 30665 22593 30699 22627
rect 30699 22593 30708 22627
rect 30656 22584 30708 22593
rect 30932 22559 30984 22568
rect 30932 22525 30941 22559
rect 30941 22525 30975 22559
rect 30975 22525 30984 22559
rect 30932 22516 30984 22525
rect 31576 22627 31628 22636
rect 31576 22593 31585 22627
rect 31585 22593 31619 22627
rect 31619 22593 31628 22627
rect 31576 22584 31628 22593
rect 31852 22584 31904 22636
rect 32680 22627 32732 22636
rect 32680 22593 32689 22627
rect 32689 22593 32723 22627
rect 32723 22593 32732 22627
rect 32680 22584 32732 22593
rect 33416 22584 33468 22636
rect 33600 22627 33652 22636
rect 33600 22593 33609 22627
rect 33609 22593 33643 22627
rect 33643 22593 33652 22627
rect 33600 22584 33652 22593
rect 31668 22516 31720 22568
rect 32772 22559 32824 22568
rect 32772 22525 32781 22559
rect 32781 22525 32815 22559
rect 32815 22525 32824 22559
rect 32772 22516 32824 22525
rect 32864 22559 32916 22568
rect 32864 22525 32873 22559
rect 32873 22525 32907 22559
rect 32907 22525 32916 22559
rect 32864 22516 32916 22525
rect 37280 22584 37332 22636
rect 37464 22627 37516 22636
rect 37464 22593 37473 22627
rect 37473 22593 37507 22627
rect 37507 22593 37516 22627
rect 37464 22584 37516 22593
rect 38844 22584 38896 22636
rect 40500 22584 40552 22636
rect 26332 22448 26384 22500
rect 27068 22448 27120 22500
rect 31576 22448 31628 22500
rect 32312 22448 32364 22500
rect 35348 22559 35400 22568
rect 35348 22525 35357 22559
rect 35357 22525 35391 22559
rect 35391 22525 35400 22559
rect 35348 22516 35400 22525
rect 36544 22559 36596 22568
rect 36544 22525 36553 22559
rect 36553 22525 36587 22559
rect 36587 22525 36596 22559
rect 36544 22516 36596 22525
rect 36636 22559 36688 22568
rect 36636 22525 36645 22559
rect 36645 22525 36679 22559
rect 36679 22525 36688 22559
rect 36636 22516 36688 22525
rect 37740 22559 37792 22568
rect 37740 22525 37749 22559
rect 37749 22525 37783 22559
rect 37783 22525 37792 22559
rect 37740 22516 37792 22525
rect 38476 22516 38528 22568
rect 40316 22559 40368 22568
rect 28448 22380 28500 22432
rect 35992 22448 36044 22500
rect 40316 22525 40325 22559
rect 40325 22525 40359 22559
rect 40359 22525 40368 22559
rect 40316 22516 40368 22525
rect 40684 22516 40736 22568
rect 45652 22720 45704 22772
rect 46848 22763 46900 22772
rect 46848 22729 46857 22763
rect 46857 22729 46891 22763
rect 46891 22729 46900 22763
rect 46848 22720 46900 22729
rect 47768 22720 47820 22772
rect 43260 22652 43312 22704
rect 42432 22584 42484 22636
rect 43720 22627 43772 22636
rect 43720 22593 43729 22627
rect 43729 22593 43763 22627
rect 43763 22593 43772 22627
rect 46940 22652 46992 22704
rect 48688 22652 48740 22704
rect 49148 22695 49200 22704
rect 49148 22661 49157 22695
rect 49157 22661 49191 22695
rect 49191 22661 49200 22695
rect 49148 22652 49200 22661
rect 43720 22584 43772 22593
rect 45100 22627 45152 22636
rect 45100 22593 45109 22627
rect 45109 22593 45143 22627
rect 45143 22593 45152 22627
rect 45100 22584 45152 22593
rect 46204 22627 46256 22636
rect 46204 22593 46213 22627
rect 46213 22593 46247 22627
rect 46247 22593 46256 22627
rect 46204 22584 46256 22593
rect 47768 22627 47820 22636
rect 47768 22593 47777 22627
rect 47777 22593 47811 22627
rect 47811 22593 47820 22627
rect 47768 22584 47820 22593
rect 50528 22584 50580 22636
rect 41236 22516 41288 22568
rect 34428 22380 34480 22432
rect 34980 22380 35032 22432
rect 36176 22380 36228 22432
rect 37188 22380 37240 22432
rect 39396 22380 39448 22432
rect 41880 22491 41932 22500
rect 41880 22457 41889 22491
rect 41889 22457 41923 22491
rect 41923 22457 41932 22491
rect 41880 22448 41932 22457
rect 41604 22380 41656 22432
rect 43812 22516 43864 22568
rect 46112 22516 46164 22568
rect 44180 22448 44232 22500
rect 44456 22448 44508 22500
rect 45008 22448 45060 22500
rect 45284 22448 45336 22500
rect 45192 22380 45244 22432
rect 45376 22380 45428 22432
rect 48412 22423 48464 22432
rect 48412 22389 48421 22423
rect 48421 22389 48455 22423
rect 48455 22389 48464 22423
rect 48412 22380 48464 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 2228 22176 2280 22228
rect 4896 22176 4948 22228
rect 6368 22176 6420 22228
rect 9956 22176 10008 22228
rect 10324 22176 10376 22228
rect 14464 22176 14516 22228
rect 15292 22219 15344 22228
rect 15292 22185 15316 22219
rect 15316 22185 15344 22219
rect 15292 22176 15344 22185
rect 16028 22176 16080 22228
rect 18604 22176 18656 22228
rect 3700 22108 3752 22160
rect 1308 22040 1360 22092
rect 3240 22040 3292 22092
rect 6828 22108 6880 22160
rect 11704 22108 11756 22160
rect 11888 22108 11940 22160
rect 3148 21972 3200 22024
rect 5816 22015 5868 22024
rect 5816 21981 5825 22015
rect 5825 21981 5859 22015
rect 5859 21981 5868 22015
rect 5816 21972 5868 21981
rect 6092 21972 6144 22024
rect 7656 21972 7708 22024
rect 9772 22083 9824 22092
rect 9772 22049 9781 22083
rect 9781 22049 9815 22083
rect 9815 22049 9824 22083
rect 9772 22040 9824 22049
rect 12532 22108 12584 22160
rect 3424 21879 3476 21888
rect 3424 21845 3433 21879
rect 3433 21845 3467 21879
rect 3467 21845 3476 21879
rect 3424 21836 3476 21845
rect 11336 21947 11388 21956
rect 11336 21913 11345 21947
rect 11345 21913 11379 21947
rect 11379 21913 11388 21947
rect 11336 21904 11388 21913
rect 5540 21836 5592 21888
rect 7656 21879 7708 21888
rect 7656 21845 7665 21879
rect 7665 21845 7699 21879
rect 7699 21845 7708 21879
rect 7656 21836 7708 21845
rect 9404 21836 9456 21888
rect 9496 21836 9548 21888
rect 15016 22083 15068 22092
rect 15016 22049 15025 22083
rect 15025 22049 15059 22083
rect 15059 22049 15068 22083
rect 16856 22108 16908 22160
rect 17408 22108 17460 22160
rect 19616 22108 19668 22160
rect 15016 22040 15068 22049
rect 12348 21904 12400 21956
rect 12624 21904 12676 21956
rect 14648 21972 14700 22024
rect 16672 21972 16724 22024
rect 16764 21972 16816 22024
rect 17316 21972 17368 22024
rect 17500 22015 17552 22024
rect 17500 21981 17509 22015
rect 17509 21981 17543 22015
rect 17543 21981 17552 22015
rect 17500 21972 17552 21981
rect 17684 22040 17736 22092
rect 21272 22176 21324 22228
rect 21088 22108 21140 22160
rect 23296 22219 23348 22228
rect 23296 22185 23305 22219
rect 23305 22185 23339 22219
rect 23339 22185 23348 22219
rect 23296 22176 23348 22185
rect 23848 22176 23900 22228
rect 24216 22176 24268 22228
rect 24584 22176 24636 22228
rect 27344 22176 27396 22228
rect 28540 22176 28592 22228
rect 28816 22176 28868 22228
rect 17868 21972 17920 22024
rect 19432 21972 19484 22024
rect 22560 22083 22612 22092
rect 22560 22049 22569 22083
rect 22569 22049 22603 22083
rect 22603 22049 22612 22083
rect 22560 22040 22612 22049
rect 23940 22108 23992 22160
rect 23388 22040 23440 22092
rect 23756 22083 23808 22092
rect 23756 22049 23765 22083
rect 23765 22049 23799 22083
rect 23799 22049 23808 22083
rect 23756 22040 23808 22049
rect 23848 22083 23900 22092
rect 23848 22049 23857 22083
rect 23857 22049 23891 22083
rect 23891 22049 23900 22083
rect 23848 22040 23900 22049
rect 26700 22108 26752 22160
rect 28632 22108 28684 22160
rect 26516 22083 26568 22092
rect 26516 22049 26525 22083
rect 26525 22049 26559 22083
rect 26559 22049 26568 22083
rect 26516 22040 26568 22049
rect 14372 21947 14424 21956
rect 13636 21836 13688 21888
rect 13728 21879 13780 21888
rect 13728 21845 13737 21879
rect 13737 21845 13771 21879
rect 13771 21845 13780 21879
rect 13728 21836 13780 21845
rect 13820 21879 13872 21888
rect 13820 21845 13829 21879
rect 13829 21845 13863 21879
rect 13863 21845 13872 21879
rect 13820 21836 13872 21845
rect 14372 21913 14381 21947
rect 14381 21913 14415 21947
rect 14415 21913 14424 21947
rect 14372 21904 14424 21913
rect 15384 21904 15436 21956
rect 17224 21904 17276 21956
rect 22100 21972 22152 22024
rect 25136 22015 25188 22024
rect 25136 21981 25145 22015
rect 25145 21981 25179 22015
rect 25179 21981 25188 22015
rect 29828 22040 29880 22092
rect 30472 22040 30524 22092
rect 31484 22176 31536 22228
rect 34980 22176 35032 22228
rect 35348 22176 35400 22228
rect 32404 22040 32456 22092
rect 32864 22040 32916 22092
rect 25136 21972 25188 21981
rect 27160 22015 27212 22024
rect 27160 21981 27169 22015
rect 27169 21981 27203 22015
rect 27203 21981 27212 22015
rect 27160 21972 27212 21981
rect 27620 21972 27672 22024
rect 21824 21904 21876 21956
rect 22468 21947 22520 21956
rect 22468 21913 22477 21947
rect 22477 21913 22511 21947
rect 22511 21913 22520 21947
rect 22468 21904 22520 21913
rect 24952 21904 25004 21956
rect 25504 21904 25556 21956
rect 25872 21904 25924 21956
rect 28448 21972 28500 22024
rect 30012 21972 30064 22024
rect 30288 21972 30340 22024
rect 34244 22108 34296 22160
rect 34428 22151 34480 22160
rect 34428 22117 34437 22151
rect 34437 22117 34471 22151
rect 34471 22117 34480 22151
rect 34428 22108 34480 22117
rect 38476 22176 38528 22228
rect 39028 22176 39080 22228
rect 36360 22040 36412 22092
rect 36820 22083 36872 22092
rect 36820 22049 36829 22083
rect 36829 22049 36863 22083
rect 36863 22049 36872 22083
rect 36820 22040 36872 22049
rect 34612 21972 34664 22024
rect 34980 21972 35032 22024
rect 29092 21904 29144 21956
rect 31392 21904 31444 21956
rect 31760 21904 31812 21956
rect 32496 21904 32548 21956
rect 38844 22108 38896 22160
rect 39396 22176 39448 22228
rect 39580 22176 39632 22228
rect 44824 22176 44876 22228
rect 38660 22040 38712 22092
rect 39212 22108 39264 22160
rect 39856 22040 39908 22092
rect 48504 22108 48556 22160
rect 42248 22040 42300 22092
rect 41512 21972 41564 22024
rect 41696 22015 41748 22024
rect 41696 21981 41705 22015
rect 41705 21981 41739 22015
rect 41739 21981 41748 22015
rect 41696 21972 41748 21981
rect 41880 21972 41932 22024
rect 43352 22040 43404 22092
rect 42892 21972 42944 22024
rect 43628 21972 43680 22024
rect 44456 22040 44508 22092
rect 44548 22083 44600 22092
rect 44548 22049 44557 22083
rect 44557 22049 44591 22083
rect 44591 22049 44600 22083
rect 44548 22040 44600 22049
rect 46204 22040 46256 22092
rect 44732 21972 44784 22024
rect 45192 22015 45244 22024
rect 45192 21981 45201 22015
rect 45201 21981 45235 22015
rect 45235 21981 45244 22015
rect 45192 21972 45244 21981
rect 46020 21972 46072 22024
rect 14924 21836 14976 21888
rect 17500 21836 17552 21888
rect 19340 21879 19392 21888
rect 19340 21845 19349 21879
rect 19349 21845 19383 21879
rect 19383 21845 19392 21879
rect 19340 21836 19392 21845
rect 19616 21879 19668 21888
rect 19616 21845 19625 21879
rect 19625 21845 19659 21879
rect 19659 21845 19668 21879
rect 19616 21836 19668 21845
rect 19984 21836 20036 21888
rect 20352 21836 20404 21888
rect 20812 21879 20864 21888
rect 20812 21845 20821 21879
rect 20821 21845 20855 21879
rect 20855 21845 20864 21879
rect 20812 21836 20864 21845
rect 21640 21836 21692 21888
rect 22008 21879 22060 21888
rect 22008 21845 22017 21879
rect 22017 21845 22051 21879
rect 22051 21845 22060 21879
rect 22008 21836 22060 21845
rect 24124 21836 24176 21888
rect 24492 21879 24544 21888
rect 24492 21845 24501 21879
rect 24501 21845 24535 21879
rect 24535 21845 24544 21879
rect 24492 21836 24544 21845
rect 24768 21879 24820 21888
rect 24768 21845 24777 21879
rect 24777 21845 24811 21879
rect 24811 21845 24820 21879
rect 24768 21836 24820 21845
rect 25964 21879 26016 21888
rect 25964 21845 25973 21879
rect 25973 21845 26007 21879
rect 26007 21845 26016 21879
rect 25964 21836 26016 21845
rect 26332 21879 26384 21888
rect 26332 21845 26341 21879
rect 26341 21845 26375 21879
rect 26375 21845 26384 21879
rect 26332 21836 26384 21845
rect 28908 21836 28960 21888
rect 33416 21836 33468 21888
rect 33508 21879 33560 21888
rect 33508 21845 33517 21879
rect 33517 21845 33551 21879
rect 33551 21845 33560 21879
rect 33508 21836 33560 21845
rect 33784 21836 33836 21888
rect 33968 21836 34020 21888
rect 34336 21836 34388 21888
rect 35256 21879 35308 21888
rect 35256 21845 35265 21879
rect 35265 21845 35299 21879
rect 35299 21845 35308 21879
rect 35256 21836 35308 21845
rect 37280 21904 37332 21956
rect 40316 21904 40368 21956
rect 40408 21947 40460 21956
rect 40408 21913 40417 21947
rect 40417 21913 40451 21947
rect 40451 21913 40460 21947
rect 40408 21904 40460 21913
rect 40868 21904 40920 21956
rect 41788 21904 41840 21956
rect 44180 21904 44232 21956
rect 46480 21972 46532 22024
rect 48320 21972 48372 22024
rect 48688 21972 48740 22024
rect 49700 21972 49752 22024
rect 47124 21904 47176 21956
rect 47676 21904 47728 21956
rect 36360 21836 36412 21888
rect 36912 21836 36964 21888
rect 37832 21879 37884 21888
rect 37832 21845 37841 21879
rect 37841 21845 37875 21879
rect 37875 21845 37884 21879
rect 37832 21836 37884 21845
rect 37924 21836 37976 21888
rect 38844 21836 38896 21888
rect 39396 21836 39448 21888
rect 40040 21879 40092 21888
rect 40040 21845 40049 21879
rect 40049 21845 40083 21879
rect 40083 21845 40092 21879
rect 40040 21836 40092 21845
rect 40500 21879 40552 21888
rect 40500 21845 40509 21879
rect 40509 21845 40543 21879
rect 40543 21845 40552 21879
rect 40500 21836 40552 21845
rect 41236 21879 41288 21888
rect 41236 21845 41245 21879
rect 41245 21845 41279 21879
rect 41279 21845 41288 21879
rect 41236 21836 41288 21845
rect 42156 21836 42208 21888
rect 43720 21836 43772 21888
rect 44548 21836 44600 21888
rect 45560 21836 45612 21888
rect 47308 21836 47360 21888
rect 48688 21836 48740 21888
rect 49148 21879 49200 21888
rect 49148 21845 49157 21879
rect 49157 21845 49191 21879
rect 49191 21845 49200 21879
rect 49148 21836 49200 21845
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 6000 21675 6052 21684
rect 6000 21641 6009 21675
rect 6009 21641 6043 21675
rect 6043 21641 6052 21675
rect 6000 21632 6052 21641
rect 10140 21675 10192 21684
rect 10140 21641 10149 21675
rect 10149 21641 10183 21675
rect 10183 21641 10192 21675
rect 10140 21632 10192 21641
rect 4344 21607 4396 21616
rect 4344 21573 4353 21607
rect 4353 21573 4387 21607
rect 4387 21573 4396 21607
rect 4344 21564 4396 21573
rect 4436 21564 4488 21616
rect 2596 21496 2648 21548
rect 5908 21496 5960 21548
rect 7932 21564 7984 21616
rect 12716 21632 12768 21684
rect 12808 21675 12860 21684
rect 12808 21641 12817 21675
rect 12817 21641 12851 21675
rect 12851 21641 12860 21675
rect 12808 21632 12860 21641
rect 14188 21632 14240 21684
rect 14280 21632 14332 21684
rect 14464 21632 14516 21684
rect 15016 21632 15068 21684
rect 15108 21632 15160 21684
rect 19616 21632 19668 21684
rect 21640 21632 21692 21684
rect 30656 21632 30708 21684
rect 31576 21632 31628 21684
rect 31760 21632 31812 21684
rect 31852 21632 31904 21684
rect 32496 21632 32548 21684
rect 3332 21428 3384 21480
rect 5632 21428 5684 21480
rect 7564 21360 7616 21412
rect 3148 21292 3200 21344
rect 3976 21292 4028 21344
rect 5632 21292 5684 21344
rect 9036 21496 9088 21548
rect 11704 21564 11756 21616
rect 17224 21564 17276 21616
rect 18144 21607 18196 21616
rect 18144 21573 18153 21607
rect 18153 21573 18187 21607
rect 18187 21573 18196 21607
rect 18144 21564 18196 21573
rect 18604 21564 18656 21616
rect 20352 21564 20404 21616
rect 22008 21564 22060 21616
rect 22284 21607 22336 21616
rect 22284 21573 22293 21607
rect 22293 21573 22327 21607
rect 22327 21573 22336 21607
rect 22284 21564 22336 21573
rect 22376 21564 22428 21616
rect 25872 21564 25924 21616
rect 26148 21564 26200 21616
rect 27344 21564 27396 21616
rect 29000 21564 29052 21616
rect 30380 21564 30432 21616
rect 32036 21564 32088 21616
rect 32956 21564 33008 21616
rect 33416 21675 33468 21684
rect 33416 21641 33425 21675
rect 33425 21641 33459 21675
rect 33459 21641 33468 21675
rect 33416 21632 33468 21641
rect 35808 21632 35860 21684
rect 36544 21632 36596 21684
rect 37832 21632 37884 21684
rect 41236 21632 41288 21684
rect 12256 21539 12308 21548
rect 12256 21505 12265 21539
rect 12265 21505 12299 21539
rect 12299 21505 12308 21539
rect 12256 21496 12308 21505
rect 12532 21496 12584 21548
rect 14740 21539 14792 21548
rect 14740 21505 14749 21539
rect 14749 21505 14783 21539
rect 14783 21505 14792 21539
rect 14740 21496 14792 21505
rect 15568 21496 15620 21548
rect 15844 21496 15896 21548
rect 16672 21496 16724 21548
rect 16948 21539 17000 21548
rect 16948 21505 16957 21539
rect 16957 21505 16991 21539
rect 16991 21505 17000 21539
rect 16948 21496 17000 21505
rect 8852 21471 8904 21480
rect 8852 21437 8861 21471
rect 8861 21437 8895 21471
rect 8895 21437 8904 21471
rect 8852 21428 8904 21437
rect 12072 21428 12124 21480
rect 13912 21428 13964 21480
rect 14924 21471 14976 21480
rect 14924 21437 14933 21471
rect 14933 21437 14967 21471
rect 14967 21437 14976 21471
rect 14924 21428 14976 21437
rect 15384 21428 15436 21480
rect 17316 21428 17368 21480
rect 17684 21428 17736 21480
rect 12256 21360 12308 21412
rect 8852 21292 8904 21344
rect 11060 21292 11112 21344
rect 11612 21335 11664 21344
rect 11612 21301 11621 21335
rect 11621 21301 11655 21335
rect 11655 21301 11664 21335
rect 11612 21292 11664 21301
rect 11704 21292 11756 21344
rect 12624 21292 12676 21344
rect 12716 21292 12768 21344
rect 17592 21360 17644 21412
rect 17868 21471 17920 21480
rect 17868 21437 17877 21471
rect 17877 21437 17911 21471
rect 17911 21437 17920 21471
rect 17868 21428 17920 21437
rect 18236 21428 18288 21480
rect 18788 21428 18840 21480
rect 21088 21496 21140 21548
rect 21916 21496 21968 21548
rect 23756 21496 23808 21548
rect 24124 21496 24176 21548
rect 24308 21539 24360 21548
rect 24308 21505 24317 21539
rect 24317 21505 24351 21539
rect 24351 21505 24360 21539
rect 24308 21496 24360 21505
rect 19156 21360 19208 21412
rect 20536 21471 20588 21480
rect 20536 21437 20545 21471
rect 20545 21437 20579 21471
rect 20579 21437 20588 21471
rect 20536 21428 20588 21437
rect 19800 21360 19852 21412
rect 21272 21428 21324 21480
rect 21640 21360 21692 21412
rect 22284 21428 22336 21480
rect 22652 21428 22704 21480
rect 25136 21428 25188 21480
rect 26332 21428 26384 21480
rect 26884 21428 26936 21480
rect 28816 21496 28868 21548
rect 29736 21496 29788 21548
rect 30932 21496 30984 21548
rect 31576 21496 31628 21548
rect 27804 21428 27856 21480
rect 23388 21360 23440 21412
rect 23664 21360 23716 21412
rect 24308 21360 24360 21412
rect 15660 21292 15712 21344
rect 15752 21292 15804 21344
rect 17224 21292 17276 21344
rect 17316 21292 17368 21344
rect 22100 21292 22152 21344
rect 22744 21292 22796 21344
rect 22928 21292 22980 21344
rect 26424 21360 26476 21412
rect 27620 21360 27672 21412
rect 28908 21360 28960 21412
rect 29276 21428 29328 21480
rect 30012 21428 30064 21480
rect 30380 21428 30432 21480
rect 30656 21428 30708 21480
rect 31392 21471 31444 21480
rect 31392 21437 31401 21471
rect 31401 21437 31435 21471
rect 31435 21437 31444 21471
rect 31392 21428 31444 21437
rect 31484 21471 31536 21480
rect 31484 21437 31493 21471
rect 31493 21437 31527 21471
rect 31527 21437 31536 21471
rect 31484 21428 31536 21437
rect 29460 21360 29512 21412
rect 34060 21607 34112 21616
rect 34060 21573 34069 21607
rect 34069 21573 34103 21607
rect 34103 21573 34112 21607
rect 34060 21564 34112 21573
rect 36268 21564 36320 21616
rect 33600 21496 33652 21548
rect 35164 21496 35216 21548
rect 35624 21496 35676 21548
rect 36360 21496 36412 21548
rect 35256 21428 35308 21480
rect 36268 21428 36320 21480
rect 38476 21564 38528 21616
rect 38568 21607 38620 21616
rect 38568 21573 38577 21607
rect 38577 21573 38611 21607
rect 38611 21573 38620 21607
rect 38568 21564 38620 21573
rect 40040 21564 40092 21616
rect 37648 21539 37700 21548
rect 37648 21505 37657 21539
rect 37657 21505 37691 21539
rect 37691 21505 37700 21539
rect 37648 21496 37700 21505
rect 37832 21539 37884 21548
rect 37832 21505 37841 21539
rect 37841 21505 37875 21539
rect 37875 21505 37884 21539
rect 37832 21496 37884 21505
rect 32404 21360 32456 21412
rect 33600 21360 33652 21412
rect 37280 21428 37332 21480
rect 37464 21428 37516 21480
rect 38568 21428 38620 21480
rect 39028 21428 39080 21480
rect 39120 21428 39172 21480
rect 39948 21496 40000 21548
rect 40408 21496 40460 21548
rect 41604 21564 41656 21616
rect 42524 21632 42576 21684
rect 45468 21632 45520 21684
rect 46480 21632 46532 21684
rect 46572 21675 46624 21684
rect 46572 21641 46581 21675
rect 46581 21641 46615 21675
rect 46615 21641 46624 21675
rect 46572 21632 46624 21641
rect 47032 21675 47084 21684
rect 47032 21641 47041 21675
rect 47041 21641 47075 21675
rect 47075 21641 47084 21675
rect 47032 21632 47084 21641
rect 47400 21632 47452 21684
rect 47676 21632 47728 21684
rect 49056 21675 49108 21684
rect 49056 21641 49065 21675
rect 49065 21641 49099 21675
rect 49099 21641 49108 21675
rect 49056 21632 49108 21641
rect 44456 21564 44508 21616
rect 42524 21496 42576 21548
rect 42800 21496 42852 21548
rect 43720 21539 43772 21548
rect 43720 21505 43729 21539
rect 43729 21505 43763 21539
rect 43763 21505 43772 21539
rect 43720 21496 43772 21505
rect 44824 21539 44876 21548
rect 44824 21505 44833 21539
rect 44833 21505 44867 21539
rect 44867 21505 44876 21539
rect 44824 21496 44876 21505
rect 49148 21564 49200 21616
rect 26332 21335 26384 21344
rect 26332 21301 26341 21335
rect 26341 21301 26375 21335
rect 26375 21301 26384 21335
rect 26332 21292 26384 21301
rect 26608 21292 26660 21344
rect 28172 21292 28224 21344
rect 28356 21292 28408 21344
rect 28632 21292 28684 21344
rect 30380 21292 30432 21344
rect 33784 21292 33836 21344
rect 36820 21360 36872 21412
rect 35532 21335 35584 21344
rect 35532 21301 35541 21335
rect 35541 21301 35575 21335
rect 35575 21301 35584 21335
rect 35532 21292 35584 21301
rect 36360 21292 36412 21344
rect 37188 21292 37240 21344
rect 39948 21360 40000 21412
rect 41512 21428 41564 21480
rect 47492 21496 47544 21548
rect 47952 21428 48004 21480
rect 41236 21360 41288 21412
rect 42156 21360 42208 21412
rect 42524 21360 42576 21412
rect 45192 21360 45244 21412
rect 47768 21360 47820 21412
rect 42064 21292 42116 21344
rect 47400 21292 47452 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 9496 21088 9548 21140
rect 10324 21131 10376 21140
rect 10324 21097 10333 21131
rect 10333 21097 10367 21131
rect 10367 21097 10376 21131
rect 10324 21088 10376 21097
rect 11520 21088 11572 21140
rect 12532 21131 12584 21140
rect 12532 21097 12541 21131
rect 12541 21097 12575 21131
rect 12575 21097 12584 21131
rect 12532 21088 12584 21097
rect 6368 21020 6420 21072
rect 16948 21088 17000 21140
rect 17224 21088 17276 21140
rect 19800 21088 19852 21140
rect 19984 21088 20036 21140
rect 21732 21088 21784 21140
rect 22008 21088 22060 21140
rect 27804 21088 27856 21140
rect 28172 21088 28224 21140
rect 4160 20952 4212 21004
rect 6736 20995 6788 21004
rect 6736 20961 6745 20995
rect 6745 20961 6779 20995
rect 6779 20961 6788 20995
rect 6736 20952 6788 20961
rect 4712 20884 4764 20936
rect 5172 20884 5224 20936
rect 7932 20927 7984 20936
rect 7932 20893 7941 20927
rect 7941 20893 7975 20927
rect 7975 20893 7984 20927
rect 7932 20884 7984 20893
rect 2872 20816 2924 20868
rect 6736 20816 6788 20868
rect 9680 20927 9732 20936
rect 9680 20893 9689 20927
rect 9689 20893 9723 20927
rect 9723 20893 9732 20927
rect 9680 20884 9732 20893
rect 11336 20952 11388 21004
rect 13544 20995 13596 21004
rect 13544 20961 13553 20995
rect 13553 20961 13587 20995
rect 13587 20961 13596 20995
rect 13544 20952 13596 20961
rect 13820 20952 13872 21004
rect 14464 20995 14516 21004
rect 14464 20961 14473 20995
rect 14473 20961 14507 20995
rect 14507 20961 14516 20995
rect 14464 20952 14516 20961
rect 16028 20952 16080 21004
rect 14096 20927 14148 20936
rect 14096 20893 14105 20927
rect 14105 20893 14139 20927
rect 14139 20893 14148 20927
rect 14096 20884 14148 20893
rect 15844 20884 15896 20936
rect 7656 20791 7708 20800
rect 7656 20757 7665 20791
rect 7665 20757 7699 20791
rect 7699 20757 7708 20791
rect 7656 20748 7708 20757
rect 9312 20748 9364 20800
rect 11152 20816 11204 20868
rect 11612 20816 11664 20868
rect 14648 20816 14700 20868
rect 15016 20816 15068 20868
rect 9772 20748 9824 20800
rect 10324 20748 10376 20800
rect 12256 20748 12308 20800
rect 12992 20791 13044 20800
rect 12992 20757 13001 20791
rect 13001 20757 13035 20791
rect 13035 20757 13044 20791
rect 12992 20748 13044 20757
rect 13912 20748 13964 20800
rect 21088 21020 21140 21072
rect 17408 20995 17460 21004
rect 17408 20961 17417 20995
rect 17417 20961 17451 20995
rect 17451 20961 17460 20995
rect 17408 20952 17460 20961
rect 17316 20927 17368 20936
rect 17316 20893 17325 20927
rect 17325 20893 17359 20927
rect 17359 20893 17368 20927
rect 17316 20884 17368 20893
rect 16764 20816 16816 20868
rect 18696 20952 18748 21004
rect 18788 20995 18840 21004
rect 18788 20961 18797 20995
rect 18797 20961 18831 20995
rect 18831 20961 18840 20995
rect 18788 20952 18840 20961
rect 19984 20995 20036 21004
rect 19984 20961 19993 20995
rect 19993 20961 20027 20995
rect 20027 20961 20036 20995
rect 19984 20952 20036 20961
rect 20076 20952 20128 21004
rect 20812 20884 20864 20936
rect 19248 20816 19300 20868
rect 16212 20791 16264 20800
rect 16212 20757 16221 20791
rect 16221 20757 16255 20791
rect 16255 20757 16264 20791
rect 16212 20748 16264 20757
rect 16672 20791 16724 20800
rect 16672 20757 16681 20791
rect 16681 20757 16715 20791
rect 16715 20757 16724 20791
rect 16672 20748 16724 20757
rect 16948 20791 17000 20800
rect 16948 20757 16957 20791
rect 16957 20757 16991 20791
rect 16991 20757 17000 20791
rect 16948 20748 17000 20757
rect 19064 20748 19116 20800
rect 19432 20748 19484 20800
rect 20260 20748 20312 20800
rect 20628 20748 20680 20800
rect 20812 20748 20864 20800
rect 21456 20952 21508 21004
rect 21732 20952 21784 21004
rect 25964 21020 26016 21072
rect 23848 20995 23900 21004
rect 23848 20961 23857 20995
rect 23857 20961 23891 20995
rect 23891 20961 23900 20995
rect 23848 20952 23900 20961
rect 24492 20952 24544 21004
rect 21088 20927 21140 20936
rect 21088 20893 21097 20927
rect 21097 20893 21131 20927
rect 21131 20893 21140 20927
rect 21088 20884 21140 20893
rect 22652 20884 22704 20936
rect 24584 20884 24636 20936
rect 22744 20816 22796 20868
rect 23296 20816 23348 20868
rect 23848 20816 23900 20868
rect 24216 20816 24268 20868
rect 25136 20884 25188 20936
rect 25320 20952 25372 21004
rect 25596 20952 25648 21004
rect 28632 21020 28684 21072
rect 28816 21131 28868 21140
rect 28816 21097 28825 21131
rect 28825 21097 28859 21131
rect 28859 21097 28868 21131
rect 28816 21088 28868 21097
rect 30196 21088 30248 21140
rect 32036 21088 32088 21140
rect 26424 20995 26476 21004
rect 26424 20961 26433 20995
rect 26433 20961 26467 20995
rect 26467 20961 26476 20995
rect 26424 20952 26476 20961
rect 27344 20952 27396 21004
rect 30196 20952 30248 21004
rect 31392 21020 31444 21072
rect 33784 21088 33836 21140
rect 34060 21088 34112 21140
rect 24768 20816 24820 20868
rect 25780 20816 25832 20868
rect 22928 20748 22980 20800
rect 23388 20748 23440 20800
rect 24308 20748 24360 20800
rect 25136 20791 25188 20800
rect 25136 20757 25145 20791
rect 25145 20757 25179 20791
rect 25179 20757 25188 20791
rect 25136 20748 25188 20757
rect 25320 20748 25372 20800
rect 26240 20791 26292 20800
rect 26240 20757 26249 20791
rect 26249 20757 26283 20791
rect 26283 20757 26292 20791
rect 26240 20748 26292 20757
rect 28724 20927 28776 20936
rect 28724 20893 28733 20927
rect 28733 20893 28767 20927
rect 28767 20893 28776 20927
rect 28724 20884 28776 20893
rect 29828 20884 29880 20936
rect 33692 21020 33744 21072
rect 40132 21088 40184 21140
rect 41236 21088 41288 21140
rect 41420 21020 41472 21072
rect 41880 21131 41932 21140
rect 41880 21097 41889 21131
rect 41889 21097 41923 21131
rect 41923 21097 41932 21131
rect 41880 21088 41932 21097
rect 47860 21088 47912 21140
rect 44272 21020 44324 21072
rect 32588 20995 32640 21004
rect 32588 20961 32597 20995
rect 32597 20961 32631 20995
rect 32631 20961 32640 20995
rect 32588 20952 32640 20961
rect 33508 20952 33560 21004
rect 34888 20995 34940 21004
rect 34888 20961 34897 20995
rect 34897 20961 34931 20995
rect 34931 20961 34940 20995
rect 34888 20952 34940 20961
rect 36176 20952 36228 21004
rect 37464 20952 37516 21004
rect 38752 20952 38804 21004
rect 39028 20952 39080 21004
rect 34060 20884 34112 20936
rect 39120 20884 39172 20936
rect 41144 20884 41196 20936
rect 41420 20884 41472 20936
rect 42524 20952 42576 21004
rect 30932 20816 30984 20868
rect 31208 20816 31260 20868
rect 26976 20791 27028 20800
rect 26976 20757 26985 20791
rect 26985 20757 27019 20791
rect 27019 20757 27028 20791
rect 26976 20748 27028 20757
rect 27068 20791 27120 20800
rect 27068 20757 27077 20791
rect 27077 20757 27111 20791
rect 27111 20757 27120 20791
rect 27068 20748 27120 20757
rect 27160 20748 27212 20800
rect 28908 20748 28960 20800
rect 29000 20748 29052 20800
rect 29368 20748 29420 20800
rect 29552 20748 29604 20800
rect 30288 20748 30340 20800
rect 31392 20791 31444 20800
rect 31392 20757 31401 20791
rect 31401 20757 31435 20791
rect 31435 20757 31444 20791
rect 31392 20748 31444 20757
rect 31576 20816 31628 20868
rect 31668 20748 31720 20800
rect 32128 20791 32180 20800
rect 32128 20757 32137 20791
rect 32137 20757 32171 20791
rect 32171 20757 32180 20791
rect 32128 20748 32180 20757
rect 32496 20791 32548 20800
rect 32496 20757 32505 20791
rect 32505 20757 32539 20791
rect 32539 20757 32548 20791
rect 32496 20748 32548 20757
rect 33324 20791 33376 20800
rect 33324 20757 33333 20791
rect 33333 20757 33367 20791
rect 33367 20757 33376 20791
rect 33324 20748 33376 20757
rect 33784 20791 33836 20800
rect 33784 20757 33793 20791
rect 33793 20757 33827 20791
rect 33827 20757 33836 20791
rect 33784 20748 33836 20757
rect 34428 20791 34480 20800
rect 34428 20757 34437 20791
rect 34437 20757 34471 20791
rect 34471 20757 34480 20791
rect 34428 20748 34480 20757
rect 35624 20816 35676 20868
rect 38292 20816 38344 20868
rect 43444 20927 43496 20936
rect 43444 20893 43453 20927
rect 43453 20893 43487 20927
rect 43487 20893 43496 20927
rect 43444 20884 43496 20893
rect 45284 20952 45336 21004
rect 45836 20995 45888 21004
rect 45836 20961 45845 20995
rect 45845 20961 45879 20995
rect 45879 20961 45888 20995
rect 45836 20952 45888 20961
rect 45008 20884 45060 20936
rect 45100 20884 45152 20936
rect 45468 20884 45520 20936
rect 46664 20884 46716 20936
rect 46940 20884 46992 20936
rect 47400 20927 47452 20936
rect 47400 20893 47409 20927
rect 47409 20893 47443 20927
rect 47443 20893 47452 20927
rect 47400 20884 47452 20893
rect 48504 20927 48556 20936
rect 48504 20893 48513 20927
rect 48513 20893 48547 20927
rect 48547 20893 48556 20927
rect 48504 20884 48556 20893
rect 50436 20884 50488 20936
rect 36636 20791 36688 20800
rect 36636 20757 36645 20791
rect 36645 20757 36679 20791
rect 36679 20757 36688 20791
rect 36636 20748 36688 20757
rect 37096 20791 37148 20800
rect 37096 20757 37105 20791
rect 37105 20757 37139 20791
rect 37139 20757 37148 20791
rect 37096 20748 37148 20757
rect 38660 20748 38712 20800
rect 39764 20748 39816 20800
rect 41512 20748 41564 20800
rect 42984 20791 43036 20800
rect 42984 20757 42993 20791
rect 42993 20757 43027 20791
rect 43027 20757 43036 20791
rect 42984 20748 43036 20757
rect 44180 20748 44232 20800
rect 45928 20816 45980 20868
rect 46572 20816 46624 20868
rect 47952 20816 48004 20868
rect 44732 20791 44784 20800
rect 44732 20757 44741 20791
rect 44741 20757 44775 20791
rect 44775 20757 44784 20791
rect 44732 20748 44784 20757
rect 46940 20791 46992 20800
rect 46940 20757 46949 20791
rect 46949 20757 46983 20791
rect 46983 20757 46992 20791
rect 46940 20748 46992 20757
rect 48504 20748 48556 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 50068 20680 50120 20732
rect 50252 20680 50304 20732
rect 3516 20544 3568 20596
rect 4988 20476 5040 20528
rect 9680 20544 9732 20596
rect 3608 20451 3660 20460
rect 3608 20417 3617 20451
rect 3617 20417 3651 20451
rect 3651 20417 3660 20451
rect 3608 20408 3660 20417
rect 6276 20476 6328 20528
rect 2780 20383 2832 20392
rect 2780 20349 2789 20383
rect 2789 20349 2823 20383
rect 2823 20349 2832 20383
rect 2780 20340 2832 20349
rect 3884 20383 3936 20392
rect 3884 20349 3893 20383
rect 3893 20349 3927 20383
rect 3927 20349 3936 20383
rect 3884 20340 3936 20349
rect 2688 20272 2740 20324
rect 8392 20519 8444 20528
rect 8392 20485 8401 20519
rect 8401 20485 8435 20519
rect 8435 20485 8444 20519
rect 8392 20476 8444 20485
rect 8944 20519 8996 20528
rect 8944 20485 8953 20519
rect 8953 20485 8987 20519
rect 8987 20485 8996 20519
rect 8944 20476 8996 20485
rect 9956 20476 10008 20528
rect 8760 20451 8812 20460
rect 8760 20417 8769 20451
rect 8769 20417 8803 20451
rect 8803 20417 8812 20451
rect 8760 20408 8812 20417
rect 9404 20451 9456 20460
rect 9404 20417 9413 20451
rect 9413 20417 9447 20451
rect 9447 20417 9456 20451
rect 9404 20408 9456 20417
rect 11520 20408 11572 20460
rect 11888 20451 11940 20460
rect 11888 20417 11897 20451
rect 11897 20417 11931 20451
rect 11931 20417 11940 20451
rect 11888 20408 11940 20417
rect 13820 20476 13872 20528
rect 15752 20519 15804 20528
rect 15752 20485 15761 20519
rect 15761 20485 15795 20519
rect 15795 20485 15804 20519
rect 15752 20476 15804 20485
rect 16304 20519 16356 20528
rect 16304 20485 16313 20519
rect 16313 20485 16347 20519
rect 16347 20485 16356 20519
rect 16304 20476 16356 20485
rect 9956 20340 10008 20392
rect 15016 20408 15068 20460
rect 15844 20408 15896 20460
rect 16120 20451 16172 20460
rect 16120 20417 16129 20451
rect 16129 20417 16163 20451
rect 16163 20417 16172 20451
rect 16120 20408 16172 20417
rect 16856 20408 16908 20460
rect 18512 20408 18564 20460
rect 13452 20340 13504 20392
rect 13912 20383 13964 20392
rect 13912 20349 13921 20383
rect 13921 20349 13955 20383
rect 13955 20349 13964 20383
rect 13912 20340 13964 20349
rect 7748 20272 7800 20324
rect 9772 20204 9824 20256
rect 10140 20204 10192 20256
rect 13636 20204 13688 20256
rect 20720 20544 20772 20596
rect 20812 20544 20864 20596
rect 22100 20544 22152 20596
rect 22928 20544 22980 20596
rect 22836 20476 22888 20528
rect 15384 20315 15436 20324
rect 15384 20281 15393 20315
rect 15393 20281 15427 20315
rect 15427 20281 15436 20315
rect 15384 20272 15436 20281
rect 18512 20272 18564 20324
rect 17592 20204 17644 20256
rect 18880 20247 18932 20256
rect 18880 20213 18889 20247
rect 18889 20213 18923 20247
rect 18923 20213 18932 20247
rect 18880 20204 18932 20213
rect 19340 20315 19392 20324
rect 19340 20281 19349 20315
rect 19349 20281 19383 20315
rect 19383 20281 19392 20315
rect 19340 20272 19392 20281
rect 22652 20408 22704 20460
rect 24860 20544 24912 20596
rect 23572 20476 23624 20528
rect 24768 20476 24820 20528
rect 22468 20383 22520 20392
rect 22468 20349 22477 20383
rect 22477 20349 22511 20383
rect 22511 20349 22520 20383
rect 22468 20340 22520 20349
rect 22928 20340 22980 20392
rect 21088 20272 21140 20324
rect 24124 20340 24176 20392
rect 26240 20544 26292 20596
rect 28356 20544 28408 20596
rect 28724 20544 28776 20596
rect 28908 20544 28960 20596
rect 30012 20544 30064 20596
rect 30104 20544 30156 20596
rect 30840 20544 30892 20596
rect 37096 20544 37148 20596
rect 37556 20587 37608 20596
rect 37556 20553 37565 20587
rect 37565 20553 37599 20587
rect 37599 20553 37608 20587
rect 37556 20544 37608 20553
rect 24492 20272 24544 20324
rect 25688 20272 25740 20324
rect 26792 20408 26844 20460
rect 26240 20383 26292 20392
rect 26240 20349 26249 20383
rect 26249 20349 26283 20383
rect 26283 20349 26292 20383
rect 26240 20340 26292 20349
rect 26332 20383 26384 20392
rect 26332 20349 26341 20383
rect 26341 20349 26375 20383
rect 26375 20349 26384 20383
rect 26332 20340 26384 20349
rect 27344 20408 27396 20460
rect 29276 20476 29328 20528
rect 32312 20476 32364 20528
rect 33232 20476 33284 20528
rect 34244 20476 34296 20528
rect 34704 20476 34756 20528
rect 36544 20519 36596 20528
rect 36544 20485 36553 20519
rect 36553 20485 36587 20519
rect 36587 20485 36596 20519
rect 36544 20476 36596 20485
rect 36728 20476 36780 20528
rect 41880 20544 41932 20596
rect 41972 20544 42024 20596
rect 43720 20544 43772 20596
rect 45468 20587 45520 20596
rect 45468 20553 45477 20587
rect 45477 20553 45511 20587
rect 45511 20553 45520 20587
rect 45468 20544 45520 20553
rect 45652 20544 45704 20596
rect 38936 20476 38988 20528
rect 40316 20476 40368 20528
rect 42248 20476 42300 20528
rect 28632 20408 28684 20460
rect 29644 20408 29696 20460
rect 27804 20340 27856 20392
rect 31116 20451 31168 20460
rect 31116 20417 31125 20451
rect 31125 20417 31159 20451
rect 31159 20417 31168 20451
rect 31116 20408 31168 20417
rect 35072 20408 35124 20460
rect 35900 20408 35952 20460
rect 37004 20408 37056 20460
rect 37464 20408 37516 20460
rect 37832 20408 37884 20460
rect 39672 20408 39724 20460
rect 40132 20408 40184 20460
rect 27068 20272 27120 20324
rect 28356 20272 28408 20324
rect 30564 20272 30616 20324
rect 32312 20383 32364 20392
rect 32312 20349 32321 20383
rect 32321 20349 32355 20383
rect 32355 20349 32364 20383
rect 32312 20340 32364 20349
rect 34060 20383 34112 20392
rect 34060 20349 34069 20383
rect 34069 20349 34103 20383
rect 34103 20349 34112 20383
rect 34060 20340 34112 20349
rect 35348 20383 35400 20392
rect 35348 20349 35357 20383
rect 35357 20349 35391 20383
rect 35391 20349 35400 20383
rect 35348 20340 35400 20349
rect 35808 20340 35860 20392
rect 21272 20204 21324 20256
rect 22468 20204 22520 20256
rect 23296 20204 23348 20256
rect 23480 20204 23532 20256
rect 25504 20204 25556 20256
rect 29276 20247 29328 20256
rect 29276 20213 29285 20247
rect 29285 20213 29319 20247
rect 29319 20213 29328 20247
rect 29276 20204 29328 20213
rect 29920 20247 29972 20256
rect 29920 20213 29929 20247
rect 29929 20213 29963 20247
rect 29963 20213 29972 20247
rect 29920 20204 29972 20213
rect 30104 20204 30156 20256
rect 34060 20204 34112 20256
rect 36452 20272 36504 20324
rect 34888 20247 34940 20256
rect 34888 20213 34897 20247
rect 34897 20213 34931 20247
rect 34931 20213 34940 20247
rect 34888 20204 34940 20213
rect 35348 20204 35400 20256
rect 36820 20272 36872 20324
rect 40316 20340 40368 20392
rect 40408 20340 40460 20392
rect 40776 20408 40828 20460
rect 41144 20408 41196 20460
rect 42064 20408 42116 20460
rect 42984 20408 43036 20460
rect 47768 20476 47820 20528
rect 49424 20476 49476 20528
rect 45836 20408 45888 20460
rect 39396 20272 39448 20324
rect 44364 20383 44416 20392
rect 44364 20349 44373 20383
rect 44373 20349 44407 20383
rect 44407 20349 44416 20383
rect 44364 20340 44416 20349
rect 44916 20340 44968 20392
rect 45284 20340 45336 20392
rect 46112 20408 46164 20460
rect 49608 20408 49660 20460
rect 46020 20340 46072 20392
rect 49148 20340 49200 20392
rect 46480 20272 46532 20324
rect 37096 20204 37148 20256
rect 37188 20204 37240 20256
rect 37648 20247 37700 20256
rect 37648 20213 37657 20247
rect 37657 20213 37691 20247
rect 37691 20213 37700 20247
rect 37648 20204 37700 20213
rect 37740 20204 37792 20256
rect 40040 20204 40092 20256
rect 40224 20247 40276 20256
rect 40224 20213 40233 20247
rect 40233 20213 40267 20247
rect 40267 20213 40276 20247
rect 40224 20204 40276 20213
rect 40316 20204 40368 20256
rect 40592 20204 40644 20256
rect 42800 20204 42852 20256
rect 44088 20204 44140 20256
rect 44272 20204 44324 20256
rect 45192 20204 45244 20256
rect 46112 20204 46164 20256
rect 47124 20204 47176 20256
rect 49516 20204 49568 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 3516 20000 3568 20052
rect 10968 19932 11020 19984
rect 11152 20000 11204 20052
rect 14188 20000 14240 20052
rect 17868 20000 17920 20052
rect 21088 20000 21140 20052
rect 21180 20000 21232 20052
rect 23296 20000 23348 20052
rect 24768 20000 24820 20052
rect 25596 20000 25648 20052
rect 11428 19932 11480 19984
rect 11520 19975 11572 19984
rect 11520 19941 11529 19975
rect 11529 19941 11563 19975
rect 11563 19941 11572 19975
rect 11520 19932 11572 19941
rect 13636 19932 13688 19984
rect 4896 19907 4948 19916
rect 4896 19873 4905 19907
rect 4905 19873 4939 19907
rect 4939 19873 4948 19907
rect 4896 19864 4948 19873
rect 6184 19864 6236 19916
rect 7288 19864 7340 19916
rect 7840 19864 7892 19916
rect 3332 19796 3384 19848
rect 2872 19728 2924 19780
rect 4896 19728 4948 19780
rect 5724 19728 5776 19780
rect 7196 19796 7248 19848
rect 10140 19864 10192 19916
rect 13728 19864 13780 19916
rect 9772 19839 9824 19848
rect 9772 19805 9781 19839
rect 9781 19805 9815 19839
rect 9815 19805 9824 19839
rect 9772 19796 9824 19805
rect 6276 19728 6328 19780
rect 11980 19839 12032 19848
rect 11980 19805 11989 19839
rect 11989 19805 12023 19839
rect 12023 19805 12032 19839
rect 11980 19796 12032 19805
rect 13544 19796 13596 19848
rect 16304 19864 16356 19916
rect 16856 19864 16908 19916
rect 19248 19932 19300 19984
rect 22560 19932 22612 19984
rect 19984 19864 20036 19916
rect 20168 19907 20220 19916
rect 20168 19873 20177 19907
rect 20177 19873 20211 19907
rect 20211 19873 20220 19907
rect 20168 19864 20220 19873
rect 20720 19907 20772 19916
rect 20720 19873 20729 19907
rect 20729 19873 20763 19907
rect 20763 19873 20772 19907
rect 20720 19864 20772 19873
rect 21640 19864 21692 19916
rect 24308 19932 24360 19984
rect 26240 19932 26292 19984
rect 26976 19932 27028 19984
rect 23756 19907 23808 19916
rect 23756 19873 23765 19907
rect 23765 19873 23799 19907
rect 23799 19873 23808 19907
rect 23756 19864 23808 19873
rect 24860 19864 24912 19916
rect 25228 19907 25280 19916
rect 25228 19873 25237 19907
rect 25237 19873 25271 19907
rect 25271 19873 25280 19907
rect 25228 19864 25280 19873
rect 27436 19907 27488 19916
rect 27436 19873 27445 19907
rect 27445 19873 27479 19907
rect 27479 19873 27488 19907
rect 27436 19864 27488 19873
rect 29736 20043 29788 20052
rect 29736 20009 29745 20043
rect 29745 20009 29779 20043
rect 29779 20009 29788 20043
rect 29736 20000 29788 20009
rect 29276 19932 29328 19984
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 15200 19796 15252 19848
rect 5448 19660 5500 19712
rect 7656 19703 7708 19712
rect 7656 19669 7665 19703
rect 7665 19669 7699 19703
rect 7699 19669 7708 19703
rect 7656 19660 7708 19669
rect 8576 19703 8628 19712
rect 8576 19669 8585 19703
rect 8585 19669 8619 19703
rect 8619 19669 8628 19703
rect 8576 19660 8628 19669
rect 9128 19703 9180 19712
rect 9128 19669 9137 19703
rect 9137 19669 9171 19703
rect 9171 19669 9180 19703
rect 9128 19660 9180 19669
rect 12256 19771 12308 19780
rect 12256 19737 12265 19771
rect 12265 19737 12299 19771
rect 12299 19737 12308 19771
rect 12256 19728 12308 19737
rect 14096 19728 14148 19780
rect 14188 19728 14240 19780
rect 16488 19728 16540 19780
rect 18420 19796 18472 19848
rect 19524 19796 19576 19848
rect 22560 19796 22612 19848
rect 22744 19796 22796 19848
rect 23572 19796 23624 19848
rect 26332 19796 26384 19848
rect 27160 19839 27212 19848
rect 27160 19805 27169 19839
rect 27169 19805 27203 19839
rect 27203 19805 27212 19839
rect 27160 19796 27212 19805
rect 28540 19796 28592 19848
rect 30196 19864 30248 19916
rect 32772 20000 32824 20052
rect 33784 20000 33836 20052
rect 33968 20000 34020 20052
rect 37740 20000 37792 20052
rect 38568 20000 38620 20052
rect 34152 19932 34204 19984
rect 35164 19932 35216 19984
rect 35532 19932 35584 19984
rect 39856 20000 39908 20052
rect 42064 20000 42116 20052
rect 42248 20000 42300 20052
rect 43444 20000 43496 20052
rect 44272 20000 44324 20052
rect 31300 19864 31352 19916
rect 32404 19907 32456 19916
rect 32404 19873 32413 19907
rect 32413 19873 32447 19907
rect 32447 19873 32456 19907
rect 32404 19864 32456 19873
rect 33140 19864 33192 19916
rect 34244 19864 34296 19916
rect 36268 19864 36320 19916
rect 36452 19864 36504 19916
rect 38476 19864 38528 19916
rect 39672 19864 39724 19916
rect 40776 19932 40828 19984
rect 45836 20043 45888 20052
rect 45836 20009 45845 20043
rect 45845 20009 45879 20043
rect 45879 20009 45888 20043
rect 45836 20000 45888 20009
rect 49056 20000 49108 20052
rect 48320 19932 48372 19984
rect 13544 19660 13596 19712
rect 13636 19660 13688 19712
rect 13820 19660 13872 19712
rect 16304 19660 16356 19712
rect 20996 19771 21048 19780
rect 20996 19737 21005 19771
rect 21005 19737 21039 19771
rect 21039 19737 21048 19771
rect 20996 19728 21048 19737
rect 22836 19728 22888 19780
rect 24584 19771 24636 19780
rect 24584 19737 24593 19771
rect 24593 19737 24627 19771
rect 24627 19737 24636 19771
rect 24584 19728 24636 19737
rect 25136 19728 25188 19780
rect 20444 19660 20496 19712
rect 20812 19660 20864 19712
rect 24308 19660 24360 19712
rect 24860 19660 24912 19712
rect 27712 19728 27764 19780
rect 29460 19728 29512 19780
rect 29276 19703 29328 19712
rect 29276 19669 29285 19703
rect 29285 19669 29319 19703
rect 29319 19669 29328 19703
rect 29276 19660 29328 19669
rect 29828 19660 29880 19712
rect 31576 19771 31628 19780
rect 31576 19737 31585 19771
rect 31585 19737 31619 19771
rect 31619 19737 31628 19771
rect 31576 19728 31628 19737
rect 32036 19728 32088 19780
rect 33140 19728 33192 19780
rect 33600 19728 33652 19780
rect 33784 19728 33836 19780
rect 36636 19796 36688 19848
rect 38660 19796 38712 19848
rect 40224 19796 40276 19848
rect 40316 19796 40368 19848
rect 34520 19728 34572 19780
rect 36360 19728 36412 19780
rect 37004 19728 37056 19780
rect 37372 19771 37424 19780
rect 37372 19737 37381 19771
rect 37381 19737 37415 19771
rect 37415 19737 37424 19771
rect 37372 19728 37424 19737
rect 38292 19728 38344 19780
rect 41880 19839 41932 19848
rect 41880 19805 41889 19839
rect 41889 19805 41923 19839
rect 41923 19805 41932 19839
rect 41880 19796 41932 19805
rect 43260 19796 43312 19848
rect 44180 19796 44232 19848
rect 46296 19839 46348 19848
rect 46296 19805 46305 19839
rect 46305 19805 46339 19839
rect 46339 19805 46348 19839
rect 46296 19796 46348 19805
rect 48412 19796 48464 19848
rect 48504 19839 48556 19848
rect 48504 19805 48513 19839
rect 48513 19805 48547 19839
rect 48547 19805 48556 19839
rect 48504 19796 48556 19805
rect 32772 19660 32824 19712
rect 33232 19660 33284 19712
rect 33508 19660 33560 19712
rect 34796 19660 34848 19712
rect 36636 19660 36688 19712
rect 41328 19728 41380 19780
rect 42064 19728 42116 19780
rect 44456 19728 44508 19780
rect 38752 19703 38804 19712
rect 38752 19669 38761 19703
rect 38761 19669 38795 19703
rect 38795 19669 38804 19703
rect 38752 19660 38804 19669
rect 40316 19660 40368 19712
rect 40408 19660 40460 19712
rect 40592 19660 40644 19712
rect 49700 19728 49752 19780
rect 42800 19660 42852 19712
rect 43352 19660 43404 19712
rect 45192 19660 45244 19712
rect 47032 19660 47084 19712
rect 50620 19660 50672 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 4528 19431 4580 19440
rect 4528 19397 4537 19431
rect 4537 19397 4571 19431
rect 4571 19397 4580 19431
rect 4528 19388 4580 19397
rect 7012 19388 7064 19440
rect 6828 19320 6880 19372
rect 9956 19499 10008 19508
rect 9956 19465 9965 19499
rect 9965 19465 9999 19499
rect 9999 19465 10008 19499
rect 9956 19456 10008 19465
rect 10140 19456 10192 19508
rect 11704 19456 11756 19508
rect 15476 19456 15528 19508
rect 15568 19499 15620 19508
rect 15568 19465 15577 19499
rect 15577 19465 15611 19499
rect 15611 19465 15620 19499
rect 15568 19456 15620 19465
rect 19248 19456 19300 19508
rect 10232 19388 10284 19440
rect 7748 19363 7800 19372
rect 7748 19329 7757 19363
rect 7757 19329 7791 19363
rect 7791 19329 7800 19363
rect 7748 19320 7800 19329
rect 8208 19363 8260 19372
rect 8208 19329 8217 19363
rect 8217 19329 8251 19363
rect 8251 19329 8260 19363
rect 8208 19320 8260 19329
rect 8576 19320 8628 19372
rect 10692 19320 10744 19372
rect 2044 19295 2096 19304
rect 2044 19261 2053 19295
rect 2053 19261 2087 19295
rect 2087 19261 2096 19295
rect 2044 19252 2096 19261
rect 5724 19252 5776 19304
rect 11336 19388 11388 19440
rect 11428 19388 11480 19440
rect 13360 19388 13412 19440
rect 14832 19388 14884 19440
rect 18512 19388 18564 19440
rect 12164 19320 12216 19372
rect 14464 19363 14516 19372
rect 14464 19329 14473 19363
rect 14473 19329 14507 19363
rect 14507 19329 14516 19363
rect 14464 19320 14516 19329
rect 14924 19320 14976 19372
rect 15384 19320 15436 19372
rect 16028 19363 16080 19372
rect 16028 19329 16037 19363
rect 16037 19329 16071 19363
rect 16071 19329 16080 19363
rect 16028 19320 16080 19329
rect 16580 19320 16632 19372
rect 17868 19320 17920 19372
rect 19708 19320 19760 19372
rect 21272 19456 21324 19508
rect 25044 19456 25096 19508
rect 25872 19456 25924 19508
rect 28080 19456 28132 19508
rect 28724 19456 28776 19508
rect 28816 19456 28868 19508
rect 29092 19456 29144 19508
rect 30472 19456 30524 19508
rect 32496 19456 32548 19508
rect 21364 19388 21416 19440
rect 21732 19388 21784 19440
rect 22284 19388 22336 19440
rect 24124 19388 24176 19440
rect 24308 19388 24360 19440
rect 2320 19184 2372 19236
rect 4620 19184 4672 19236
rect 5080 19184 5132 19236
rect 7748 19184 7800 19236
rect 7840 19184 7892 19236
rect 10508 19184 10560 19236
rect 11060 19252 11112 19304
rect 12716 19252 12768 19304
rect 13360 19252 13412 19304
rect 14004 19295 14056 19304
rect 14004 19261 14013 19295
rect 14013 19261 14047 19295
rect 14047 19261 14056 19295
rect 14004 19252 14056 19261
rect 14096 19252 14148 19304
rect 14832 19252 14884 19304
rect 15016 19252 15068 19304
rect 15200 19252 15252 19304
rect 16120 19295 16172 19304
rect 16120 19261 16129 19295
rect 16129 19261 16163 19295
rect 16163 19261 16172 19295
rect 16120 19252 16172 19261
rect 6552 19159 6604 19168
rect 6552 19125 6561 19159
rect 6561 19125 6595 19159
rect 6595 19125 6604 19159
rect 6552 19116 6604 19125
rect 7104 19116 7156 19168
rect 7656 19116 7708 19168
rect 7932 19116 7984 19168
rect 8024 19116 8076 19168
rect 9220 19116 9272 19168
rect 9588 19116 9640 19168
rect 12072 19184 12124 19236
rect 11060 19116 11112 19168
rect 11336 19116 11388 19168
rect 12164 19116 12216 19168
rect 12440 19159 12492 19168
rect 12440 19125 12449 19159
rect 12449 19125 12483 19159
rect 12483 19125 12492 19159
rect 12440 19116 12492 19125
rect 13728 19184 13780 19236
rect 21088 19320 21140 19372
rect 21456 19320 21508 19372
rect 22008 19320 22060 19372
rect 21916 19252 21968 19304
rect 23480 19320 23532 19372
rect 24860 19320 24912 19372
rect 17960 19184 18012 19236
rect 19432 19184 19484 19236
rect 21732 19184 21784 19236
rect 22468 19252 22520 19304
rect 23848 19295 23900 19304
rect 17868 19116 17920 19168
rect 20812 19116 20864 19168
rect 21456 19116 21508 19168
rect 22008 19116 22060 19168
rect 22284 19116 22336 19168
rect 23480 19116 23532 19168
rect 23848 19261 23857 19295
rect 23857 19261 23891 19295
rect 23891 19261 23900 19295
rect 23848 19252 23900 19261
rect 23940 19252 23992 19304
rect 24584 19252 24636 19304
rect 25596 19320 25648 19372
rect 25136 19295 25188 19304
rect 25136 19261 25145 19295
rect 25145 19261 25179 19295
rect 25179 19261 25188 19295
rect 26240 19320 26292 19372
rect 25136 19252 25188 19261
rect 27252 19252 27304 19304
rect 27988 19295 28040 19304
rect 25228 19184 25280 19236
rect 25964 19184 26016 19236
rect 26884 19184 26936 19236
rect 27988 19261 27997 19295
rect 27997 19261 28031 19295
rect 28031 19261 28040 19295
rect 27988 19252 28040 19261
rect 29276 19320 29328 19372
rect 29460 19320 29512 19372
rect 31484 19388 31536 19440
rect 33048 19456 33100 19508
rect 33324 19456 33376 19508
rect 34060 19388 34112 19440
rect 34428 19388 34480 19440
rect 40500 19456 40552 19508
rect 40960 19456 41012 19508
rect 41880 19456 41932 19508
rect 42616 19456 42668 19508
rect 43260 19499 43312 19508
rect 43260 19465 43269 19499
rect 43269 19465 43303 19499
rect 43303 19465 43312 19499
rect 43260 19456 43312 19465
rect 43444 19456 43496 19508
rect 28540 19252 28592 19304
rect 27436 19184 27488 19236
rect 29276 19184 29328 19236
rect 31300 19363 31352 19372
rect 31300 19329 31309 19363
rect 31309 19329 31343 19363
rect 31343 19329 31352 19363
rect 31300 19320 31352 19329
rect 31392 19363 31444 19372
rect 31392 19329 31401 19363
rect 31401 19329 31435 19363
rect 31435 19329 31444 19363
rect 31392 19320 31444 19329
rect 34152 19363 34204 19372
rect 34152 19329 34161 19363
rect 34161 19329 34195 19363
rect 34195 19329 34204 19363
rect 34152 19320 34204 19329
rect 34244 19320 34296 19372
rect 32128 19252 32180 19304
rect 32956 19252 33008 19304
rect 30012 19184 30064 19236
rect 26516 19116 26568 19168
rect 28172 19116 28224 19168
rect 29000 19116 29052 19168
rect 30564 19116 30616 19168
rect 33784 19227 33836 19236
rect 33784 19193 33793 19227
rect 33793 19193 33827 19227
rect 33827 19193 33836 19227
rect 33784 19184 33836 19193
rect 34336 19295 34388 19304
rect 34336 19261 34345 19295
rect 34345 19261 34379 19295
rect 34379 19261 34388 19295
rect 34336 19252 34388 19261
rect 34796 19363 34848 19372
rect 34796 19329 34805 19363
rect 34805 19329 34839 19363
rect 34839 19329 34848 19363
rect 34796 19320 34848 19329
rect 36084 19320 36136 19372
rect 36176 19320 36228 19372
rect 39120 19388 39172 19440
rect 41144 19431 41196 19440
rect 41144 19397 41153 19431
rect 41153 19397 41187 19431
rect 41187 19397 41196 19431
rect 41144 19388 41196 19397
rect 41328 19388 41380 19440
rect 37359 19320 37411 19372
rect 37464 19363 37516 19372
rect 37464 19329 37495 19363
rect 37495 19329 37516 19363
rect 37464 19320 37516 19329
rect 37832 19320 37884 19372
rect 40224 19320 40276 19372
rect 40408 19320 40460 19372
rect 35164 19184 35216 19236
rect 35624 19184 35676 19236
rect 30840 19116 30892 19168
rect 32220 19159 32272 19168
rect 32220 19125 32229 19159
rect 32229 19125 32263 19159
rect 32263 19125 32272 19159
rect 32220 19116 32272 19125
rect 34060 19116 34112 19168
rect 36452 19184 36504 19236
rect 40132 19252 40184 19304
rect 40316 19252 40368 19304
rect 40500 19252 40552 19304
rect 35900 19116 35952 19168
rect 38200 19116 38252 19168
rect 40040 19116 40092 19168
rect 40224 19116 40276 19168
rect 41328 19252 41380 19304
rect 41236 19184 41288 19236
rect 41972 19295 42024 19304
rect 41972 19261 41981 19295
rect 41981 19261 42015 19295
rect 42015 19261 42024 19295
rect 41972 19252 42024 19261
rect 42616 19363 42668 19372
rect 42616 19329 42625 19363
rect 42625 19329 42659 19363
rect 42659 19329 42668 19363
rect 42616 19320 42668 19329
rect 44088 19388 44140 19440
rect 42800 19252 42852 19304
rect 45928 19363 45980 19372
rect 45928 19329 45937 19363
rect 45937 19329 45971 19363
rect 45971 19329 45980 19363
rect 45928 19320 45980 19329
rect 46940 19320 46992 19372
rect 49148 19363 49200 19372
rect 49148 19329 49157 19363
rect 49157 19329 49191 19363
rect 49191 19329 49200 19363
rect 49148 19320 49200 19329
rect 50068 19320 50120 19372
rect 50804 19320 50856 19372
rect 44088 19252 44140 19304
rect 44456 19252 44508 19304
rect 42616 19184 42668 19236
rect 45652 19184 45704 19236
rect 41696 19116 41748 19168
rect 41972 19116 42024 19168
rect 42248 19159 42300 19168
rect 42248 19125 42257 19159
rect 42257 19125 42291 19159
rect 42291 19125 42300 19159
rect 42248 19116 42300 19125
rect 46940 19116 46992 19168
rect 47216 19116 47268 19168
rect 47860 19184 47912 19236
rect 48228 19116 48280 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 5448 18912 5500 18964
rect 5540 18912 5592 18964
rect 7012 18912 7064 18964
rect 7748 18912 7800 18964
rect 8024 18912 8076 18964
rect 9036 18955 9088 18964
rect 9036 18921 9045 18955
rect 9045 18921 9079 18955
rect 9079 18921 9088 18955
rect 9036 18912 9088 18921
rect 3516 18844 3568 18896
rect 3424 18776 3476 18828
rect 3884 18708 3936 18760
rect 2780 18683 2832 18692
rect 2780 18649 2789 18683
rect 2789 18649 2823 18683
rect 2823 18649 2832 18683
rect 2780 18640 2832 18649
rect 3424 18640 3476 18692
rect 2872 18572 2924 18624
rect 7104 18776 7156 18828
rect 7656 18844 7708 18896
rect 11060 18912 11112 18964
rect 15108 18912 15160 18964
rect 16672 18912 16724 18964
rect 20168 18955 20220 18964
rect 20168 18921 20177 18955
rect 20177 18921 20211 18955
rect 20211 18921 20220 18955
rect 20168 18912 20220 18921
rect 9220 18844 9272 18896
rect 10324 18844 10376 18896
rect 13728 18844 13780 18896
rect 20996 18912 21048 18964
rect 22284 18912 22336 18964
rect 23480 18912 23532 18964
rect 23664 18912 23716 18964
rect 29000 18955 29052 18964
rect 29000 18921 29009 18955
rect 29009 18921 29043 18955
rect 29043 18921 29052 18955
rect 29000 18912 29052 18921
rect 30104 18912 30156 18964
rect 4988 18708 5040 18760
rect 6552 18708 6604 18760
rect 7840 18708 7892 18760
rect 10048 18776 10100 18828
rect 5540 18640 5592 18692
rect 5724 18640 5776 18692
rect 6184 18683 6236 18692
rect 6184 18649 6193 18683
rect 6193 18649 6227 18683
rect 6227 18649 6236 18683
rect 6184 18640 6236 18649
rect 7748 18640 7800 18692
rect 9496 18751 9548 18760
rect 9496 18717 9505 18751
rect 9505 18717 9539 18751
rect 9539 18717 9548 18751
rect 9496 18708 9548 18717
rect 8484 18640 8536 18692
rect 11152 18640 11204 18692
rect 12164 18640 12216 18692
rect 14280 18819 14332 18828
rect 14280 18785 14289 18819
rect 14289 18785 14323 18819
rect 14323 18785 14332 18819
rect 14280 18776 14332 18785
rect 17960 18776 18012 18828
rect 18880 18776 18932 18828
rect 19984 18776 20036 18828
rect 14188 18640 14240 18692
rect 14556 18683 14608 18692
rect 14556 18649 14565 18683
rect 14565 18649 14599 18683
rect 14599 18649 14608 18683
rect 14556 18640 14608 18649
rect 14832 18640 14884 18692
rect 15016 18640 15068 18692
rect 5816 18615 5868 18624
rect 5816 18581 5825 18615
rect 5825 18581 5859 18615
rect 5859 18581 5868 18615
rect 5816 18572 5868 18581
rect 8576 18615 8628 18624
rect 8576 18581 8585 18615
rect 8585 18581 8619 18615
rect 8619 18581 8628 18615
rect 8576 18572 8628 18581
rect 8944 18572 8996 18624
rect 9588 18572 9640 18624
rect 12808 18615 12860 18624
rect 12808 18581 12817 18615
rect 12817 18581 12851 18615
rect 12851 18581 12860 18615
rect 12808 18572 12860 18581
rect 20352 18708 20404 18760
rect 21732 18844 21784 18896
rect 23940 18776 23992 18828
rect 24860 18887 24912 18896
rect 24860 18853 24869 18887
rect 24869 18853 24903 18887
rect 24903 18853 24912 18887
rect 24860 18844 24912 18853
rect 25320 18776 25372 18828
rect 16488 18683 16540 18692
rect 16488 18649 16497 18683
rect 16497 18649 16531 18683
rect 16531 18649 16540 18683
rect 16488 18640 16540 18649
rect 17500 18640 17552 18692
rect 16120 18572 16172 18624
rect 16948 18572 17000 18624
rect 18880 18640 18932 18692
rect 18328 18572 18380 18624
rect 18972 18615 19024 18624
rect 18972 18581 18981 18615
rect 18981 18581 19015 18615
rect 19015 18581 19024 18615
rect 18972 18572 19024 18581
rect 19524 18683 19576 18692
rect 19524 18649 19533 18683
rect 19533 18649 19567 18683
rect 19567 18649 19576 18683
rect 19524 18640 19576 18649
rect 21180 18708 21232 18760
rect 21364 18751 21416 18760
rect 21364 18717 21373 18751
rect 21373 18717 21407 18751
rect 21407 18717 21416 18751
rect 21364 18708 21416 18717
rect 22744 18708 22796 18760
rect 27068 18844 27120 18896
rect 27712 18844 27764 18896
rect 30380 18912 30432 18964
rect 32220 18912 32272 18964
rect 25964 18776 26016 18828
rect 26516 18776 26568 18828
rect 27344 18819 27396 18828
rect 27344 18785 27353 18819
rect 27353 18785 27387 18819
rect 27387 18785 27396 18819
rect 27344 18776 27396 18785
rect 27436 18708 27488 18760
rect 22836 18640 22888 18692
rect 28724 18776 28776 18828
rect 29368 18776 29420 18828
rect 30564 18844 30616 18896
rect 32588 18844 32640 18896
rect 28908 18708 28960 18760
rect 29276 18751 29328 18760
rect 29276 18717 29285 18751
rect 29285 18717 29319 18751
rect 29319 18717 29328 18751
rect 29276 18708 29328 18717
rect 29736 18708 29788 18760
rect 32312 18776 32364 18828
rect 22284 18572 22336 18624
rect 22744 18615 22796 18624
rect 22744 18581 22753 18615
rect 22753 18581 22787 18615
rect 22787 18581 22796 18615
rect 22744 18572 22796 18581
rect 23480 18615 23532 18624
rect 23480 18581 23489 18615
rect 23489 18581 23523 18615
rect 23523 18581 23532 18615
rect 23480 18572 23532 18581
rect 23756 18572 23808 18624
rect 24308 18572 24360 18624
rect 25872 18572 25924 18624
rect 26332 18572 26384 18624
rect 28172 18640 28224 18692
rect 29828 18640 29880 18692
rect 31116 18640 31168 18692
rect 31576 18708 31628 18760
rect 32128 18708 32180 18760
rect 33600 18776 33652 18828
rect 33876 18776 33928 18828
rect 34244 18776 34296 18828
rect 34612 18776 34664 18828
rect 36084 18776 36136 18828
rect 36268 18819 36320 18828
rect 36268 18785 36277 18819
rect 36277 18785 36311 18819
rect 36311 18785 36320 18819
rect 36268 18776 36320 18785
rect 38568 18844 38620 18896
rect 39580 18887 39632 18896
rect 39580 18853 39589 18887
rect 39589 18853 39623 18887
rect 39623 18853 39632 18887
rect 39580 18844 39632 18853
rect 39672 18844 39724 18896
rect 44180 18912 44232 18964
rect 46296 18912 46348 18964
rect 47400 18955 47452 18964
rect 47400 18921 47409 18955
rect 47409 18921 47443 18955
rect 47443 18921 47452 18955
rect 47400 18912 47452 18921
rect 48412 18955 48464 18964
rect 48412 18921 48421 18955
rect 48421 18921 48455 18955
rect 48455 18921 48464 18955
rect 48412 18912 48464 18921
rect 48964 18912 49016 18964
rect 38752 18776 38804 18828
rect 39856 18776 39908 18828
rect 41604 18776 41656 18828
rect 42616 18776 42668 18828
rect 32220 18640 32272 18692
rect 32404 18640 32456 18692
rect 36176 18708 36228 18760
rect 38660 18708 38712 18760
rect 39764 18708 39816 18760
rect 40040 18751 40092 18760
rect 40040 18717 40049 18751
rect 40049 18717 40083 18751
rect 40083 18717 40092 18751
rect 40040 18708 40092 18717
rect 34060 18640 34112 18692
rect 34336 18640 34388 18692
rect 28080 18572 28132 18624
rect 29368 18572 29420 18624
rect 29460 18572 29512 18624
rect 29644 18572 29696 18624
rect 33324 18572 33376 18624
rect 34796 18572 34848 18624
rect 35256 18683 35308 18692
rect 35256 18649 35265 18683
rect 35265 18649 35299 18683
rect 35299 18649 35308 18683
rect 35256 18640 35308 18649
rect 35440 18640 35492 18692
rect 36820 18640 36872 18692
rect 37832 18640 37884 18692
rect 39948 18640 40000 18692
rect 40316 18683 40368 18692
rect 40316 18649 40346 18683
rect 40346 18649 40368 18683
rect 40316 18640 40368 18649
rect 42156 18708 42208 18760
rect 42248 18751 42300 18760
rect 42248 18717 42257 18751
rect 42257 18717 42291 18751
rect 42291 18717 42300 18751
rect 42248 18708 42300 18717
rect 47124 18844 47176 18896
rect 43720 18776 43772 18828
rect 44824 18776 44876 18828
rect 43904 18708 43956 18760
rect 46296 18751 46348 18760
rect 46296 18717 46305 18751
rect 46305 18717 46339 18751
rect 46339 18717 46348 18751
rect 46296 18708 46348 18717
rect 36728 18572 36780 18624
rect 38752 18572 38804 18624
rect 38844 18615 38896 18624
rect 38844 18581 38853 18615
rect 38853 18581 38887 18615
rect 38887 18581 38896 18615
rect 38844 18572 38896 18581
rect 38936 18615 38988 18624
rect 38936 18581 38945 18615
rect 38945 18581 38979 18615
rect 38979 18581 38988 18615
rect 38936 18572 38988 18581
rect 40592 18572 40644 18624
rect 41604 18572 41656 18624
rect 41696 18572 41748 18624
rect 49700 18640 49752 18692
rect 42616 18572 42668 18624
rect 43720 18572 43772 18624
rect 44272 18572 44324 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 3516 18368 3568 18420
rect 3608 18411 3660 18420
rect 3608 18377 3617 18411
rect 3617 18377 3651 18411
rect 3651 18377 3660 18411
rect 3608 18368 3660 18377
rect 12164 18368 12216 18420
rect 12624 18368 12676 18420
rect 6552 18300 6604 18352
rect 8852 18300 8904 18352
rect 10048 18300 10100 18352
rect 10876 18343 10928 18352
rect 10876 18309 10885 18343
rect 10885 18309 10919 18343
rect 10919 18309 10928 18343
rect 10876 18300 10928 18309
rect 11060 18300 11112 18352
rect 14648 18368 14700 18420
rect 17316 18411 17368 18420
rect 17316 18377 17325 18411
rect 17325 18377 17359 18411
rect 17359 18377 17368 18411
rect 17316 18368 17368 18377
rect 18696 18368 18748 18420
rect 13360 18300 13412 18352
rect 14188 18300 14240 18352
rect 22192 18411 22244 18420
rect 22192 18377 22201 18411
rect 22201 18377 22235 18411
rect 22235 18377 22244 18411
rect 22192 18368 22244 18377
rect 23480 18368 23532 18420
rect 25780 18368 25832 18420
rect 24768 18300 24820 18352
rect 3608 18232 3660 18284
rect 2044 18207 2096 18216
rect 2044 18173 2053 18207
rect 2053 18173 2087 18207
rect 2087 18173 2096 18207
rect 2044 18164 2096 18173
rect 6000 18232 6052 18284
rect 7012 18232 7064 18284
rect 7380 18275 7432 18284
rect 7380 18241 7389 18275
rect 7389 18241 7423 18275
rect 7423 18241 7432 18275
rect 7380 18232 7432 18241
rect 8484 18275 8536 18284
rect 8484 18241 8493 18275
rect 8493 18241 8527 18275
rect 8527 18241 8536 18275
rect 8484 18232 8536 18241
rect 11796 18275 11848 18284
rect 11796 18241 11805 18275
rect 11805 18241 11839 18275
rect 11839 18241 11848 18275
rect 11796 18232 11848 18241
rect 15568 18232 15620 18284
rect 7104 18164 7156 18216
rect 8852 18164 8904 18216
rect 3884 18096 3936 18148
rect 5724 18028 5776 18080
rect 5908 18028 5960 18080
rect 7840 18096 7892 18148
rect 8300 18096 8352 18148
rect 10232 18207 10284 18216
rect 10232 18173 10241 18207
rect 10241 18173 10275 18207
rect 10275 18173 10284 18207
rect 10232 18164 10284 18173
rect 11980 18164 12032 18216
rect 12164 18096 12216 18148
rect 12532 18096 12584 18148
rect 9404 18028 9456 18080
rect 11244 18028 11296 18080
rect 12900 18164 12952 18216
rect 15292 18207 15344 18216
rect 15292 18173 15301 18207
rect 15301 18173 15335 18207
rect 15335 18173 15344 18207
rect 15292 18164 15344 18173
rect 15844 18164 15896 18216
rect 14648 18096 14700 18148
rect 16304 18232 16356 18284
rect 17868 18232 17920 18284
rect 19156 18232 19208 18284
rect 19432 18232 19484 18284
rect 16212 18164 16264 18216
rect 17500 18164 17552 18216
rect 20996 18232 21048 18284
rect 22008 18232 22060 18284
rect 22284 18232 22336 18284
rect 25136 18232 25188 18284
rect 26608 18368 26660 18420
rect 27068 18368 27120 18420
rect 27252 18368 27304 18420
rect 30840 18368 30892 18420
rect 31576 18368 31628 18420
rect 31760 18368 31812 18420
rect 34428 18368 34480 18420
rect 36176 18411 36228 18420
rect 36176 18377 36185 18411
rect 36185 18377 36219 18411
rect 36219 18377 36228 18411
rect 36176 18368 36228 18377
rect 36636 18368 36688 18420
rect 36728 18368 36780 18420
rect 38660 18368 38712 18420
rect 38936 18368 38988 18420
rect 26424 18300 26476 18352
rect 28816 18300 28868 18352
rect 33324 18300 33376 18352
rect 33600 18300 33652 18352
rect 27068 18232 27120 18284
rect 27160 18275 27212 18284
rect 27160 18241 27169 18275
rect 27169 18241 27203 18275
rect 27203 18241 27212 18275
rect 27160 18232 27212 18241
rect 28724 18232 28776 18284
rect 22836 18207 22888 18216
rect 22836 18173 22845 18207
rect 22845 18173 22879 18207
rect 22879 18173 22888 18207
rect 22836 18164 22888 18173
rect 24584 18207 24636 18216
rect 24584 18173 24593 18207
rect 24593 18173 24627 18207
rect 24627 18173 24636 18207
rect 24584 18164 24636 18173
rect 14280 18028 14332 18080
rect 14832 18071 14884 18080
rect 14832 18037 14841 18071
rect 14841 18037 14875 18071
rect 14875 18037 14884 18071
rect 14832 18028 14884 18037
rect 16396 18028 16448 18080
rect 17960 18028 18012 18080
rect 19156 18028 19208 18080
rect 26148 18207 26200 18216
rect 26148 18173 26157 18207
rect 26157 18173 26191 18207
rect 26191 18173 26200 18207
rect 26148 18164 26200 18173
rect 27528 18164 27580 18216
rect 25044 18096 25096 18148
rect 26608 18096 26660 18148
rect 20904 18028 20956 18080
rect 21456 18028 21508 18080
rect 24952 18071 25004 18080
rect 24952 18037 24961 18071
rect 24961 18037 24995 18071
rect 24995 18037 25004 18071
rect 24952 18028 25004 18037
rect 25964 18028 26016 18080
rect 30564 18232 30616 18284
rect 30840 18232 30892 18284
rect 30932 18275 30984 18284
rect 30932 18241 30941 18275
rect 30941 18241 30975 18275
rect 30975 18241 30984 18275
rect 30932 18232 30984 18241
rect 31392 18164 31444 18216
rect 32220 18275 32272 18284
rect 32220 18241 32229 18275
rect 32229 18241 32263 18275
rect 32263 18241 32272 18275
rect 32220 18232 32272 18241
rect 34336 18300 34388 18352
rect 34704 18343 34756 18352
rect 34704 18309 34713 18343
rect 34713 18309 34747 18343
rect 34747 18309 34756 18343
rect 34704 18300 34756 18309
rect 37832 18300 37884 18352
rect 32128 18164 32180 18216
rect 32680 18164 32732 18216
rect 30380 18096 30432 18148
rect 33232 18207 33284 18216
rect 33232 18173 33241 18207
rect 33241 18173 33275 18207
rect 33275 18173 33284 18207
rect 33232 18164 33284 18173
rect 33324 18164 33376 18216
rect 33416 18164 33468 18216
rect 34060 18164 34112 18216
rect 36728 18275 36780 18284
rect 36728 18241 36737 18275
rect 36737 18241 36771 18275
rect 36771 18241 36780 18275
rect 36728 18232 36780 18241
rect 37280 18232 37332 18284
rect 34428 18207 34480 18216
rect 34428 18173 34437 18207
rect 34437 18173 34471 18207
rect 34471 18173 34480 18207
rect 34428 18164 34480 18173
rect 39120 18300 39172 18352
rect 40132 18300 40184 18352
rect 39948 18232 40000 18284
rect 40592 18368 40644 18420
rect 38292 18164 38344 18216
rect 40316 18232 40368 18284
rect 40592 18232 40644 18284
rect 30564 18071 30616 18080
rect 30564 18037 30573 18071
rect 30573 18037 30607 18071
rect 30607 18037 30616 18071
rect 30564 18028 30616 18037
rect 30748 18028 30800 18080
rect 31668 18028 31720 18080
rect 32680 18071 32732 18080
rect 32680 18037 32689 18071
rect 32689 18037 32723 18071
rect 32723 18037 32732 18071
rect 32680 18028 32732 18037
rect 33968 18028 34020 18080
rect 36176 18096 36228 18148
rect 36820 18096 36872 18148
rect 35992 18028 36044 18080
rect 37464 18028 37516 18080
rect 40776 18164 40828 18216
rect 41236 18343 41288 18352
rect 41236 18309 41245 18343
rect 41245 18309 41279 18343
rect 41279 18309 41288 18343
rect 41236 18300 41288 18309
rect 42800 18368 42852 18420
rect 44916 18368 44968 18420
rect 49240 18411 49292 18420
rect 49240 18377 49249 18411
rect 49249 18377 49283 18411
rect 49283 18377 49292 18411
rect 49240 18368 49292 18377
rect 42156 18300 42208 18352
rect 42708 18300 42760 18352
rect 46480 18300 46532 18352
rect 46940 18300 46992 18352
rect 47860 18300 47912 18352
rect 42616 18275 42668 18284
rect 42616 18241 42625 18275
rect 42625 18241 42659 18275
rect 42659 18241 42668 18275
rect 42616 18232 42668 18241
rect 43720 18275 43772 18284
rect 43720 18241 43729 18275
rect 43729 18241 43763 18275
rect 43763 18241 43772 18275
rect 43720 18232 43772 18241
rect 44364 18275 44416 18284
rect 44364 18241 44373 18275
rect 44373 18241 44407 18275
rect 44407 18241 44416 18275
rect 44364 18232 44416 18241
rect 44548 18232 44600 18284
rect 47032 18232 47084 18284
rect 47124 18232 47176 18284
rect 50068 18232 50120 18284
rect 41420 18207 41472 18216
rect 41420 18173 41429 18207
rect 41429 18173 41463 18207
rect 41463 18173 41472 18207
rect 41420 18164 41472 18173
rect 41512 18164 41564 18216
rect 41604 18164 41656 18216
rect 40316 18139 40368 18148
rect 40316 18105 40325 18139
rect 40325 18105 40359 18139
rect 40359 18105 40368 18139
rect 46296 18164 46348 18216
rect 47584 18164 47636 18216
rect 48872 18164 48924 18216
rect 40316 18096 40368 18105
rect 43996 18096 44048 18148
rect 47124 18096 47176 18148
rect 40040 18028 40092 18080
rect 40132 18028 40184 18080
rect 40960 18028 41012 18080
rect 41144 18028 41196 18080
rect 42340 18028 42392 18080
rect 42800 18028 42852 18080
rect 45376 18028 45428 18080
rect 46664 18028 46716 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 2872 17824 2924 17876
rect 6644 17824 6696 17876
rect 9496 17824 9548 17876
rect 1216 17688 1268 17740
rect 4160 17688 4212 17740
rect 10968 17756 11020 17808
rect 9772 17688 9824 17740
rect 3424 17663 3476 17672
rect 3424 17629 3433 17663
rect 3433 17629 3467 17663
rect 3467 17629 3476 17663
rect 3424 17620 3476 17629
rect 4620 17663 4672 17672
rect 4620 17629 4629 17663
rect 4629 17629 4663 17663
rect 4663 17629 4672 17663
rect 4620 17620 4672 17629
rect 5724 17663 5776 17672
rect 5724 17629 5733 17663
rect 5733 17629 5767 17663
rect 5767 17629 5776 17663
rect 5724 17620 5776 17629
rect 6828 17663 6880 17672
rect 6828 17629 6837 17663
rect 6837 17629 6871 17663
rect 6871 17629 6880 17663
rect 6828 17620 6880 17629
rect 9956 17620 10008 17672
rect 14740 17824 14792 17876
rect 14924 17824 14976 17876
rect 19616 17824 19668 17876
rect 11152 17731 11204 17740
rect 11152 17697 11161 17731
rect 11161 17697 11195 17731
rect 11195 17697 11204 17731
rect 11152 17688 11204 17697
rect 11980 17688 12032 17740
rect 12164 17688 12216 17740
rect 13268 17756 13320 17808
rect 13452 17756 13504 17808
rect 20904 17824 20956 17876
rect 24216 17824 24268 17876
rect 12808 17688 12860 17740
rect 22652 17756 22704 17808
rect 17040 17688 17092 17740
rect 17960 17688 18012 17740
rect 19248 17688 19300 17740
rect 12532 17620 12584 17672
rect 8944 17527 8996 17536
rect 8944 17493 8953 17527
rect 8953 17493 8987 17527
rect 8987 17493 8996 17527
rect 8944 17484 8996 17493
rect 9220 17552 9272 17604
rect 9588 17552 9640 17604
rect 10508 17484 10560 17536
rect 10876 17552 10928 17604
rect 13544 17595 13596 17604
rect 13544 17561 13553 17595
rect 13553 17561 13587 17595
rect 13587 17561 13596 17595
rect 13544 17552 13596 17561
rect 14280 17663 14332 17672
rect 14280 17629 14289 17663
rect 14289 17629 14323 17663
rect 14323 17629 14332 17663
rect 14280 17620 14332 17629
rect 15016 17552 15068 17604
rect 13360 17484 13412 17536
rect 14740 17484 14792 17536
rect 17132 17552 17184 17604
rect 19432 17620 19484 17672
rect 22008 17688 22060 17740
rect 26240 17688 26292 17740
rect 26976 17824 27028 17876
rect 27436 17824 27488 17876
rect 27620 17867 27672 17876
rect 27620 17833 27629 17867
rect 27629 17833 27663 17867
rect 27663 17833 27672 17867
rect 27620 17824 27672 17833
rect 28080 17824 28132 17876
rect 30196 17824 30248 17876
rect 30656 17824 30708 17876
rect 27252 17756 27304 17808
rect 28080 17731 28132 17740
rect 28080 17697 28089 17731
rect 28089 17697 28123 17731
rect 28123 17697 28132 17731
rect 28080 17688 28132 17697
rect 28632 17688 28684 17740
rect 29460 17688 29512 17740
rect 32588 17756 32640 17808
rect 33416 17756 33468 17808
rect 34152 17824 34204 17876
rect 34980 17824 35032 17876
rect 35992 17867 36044 17876
rect 35992 17833 36001 17867
rect 36001 17833 36035 17867
rect 36035 17833 36044 17867
rect 35992 17824 36044 17833
rect 35900 17756 35952 17808
rect 36452 17756 36504 17808
rect 37924 17824 37976 17876
rect 44456 17824 44508 17876
rect 46480 17824 46532 17876
rect 38476 17756 38528 17808
rect 38568 17756 38620 17808
rect 39672 17756 39724 17808
rect 41512 17756 41564 17808
rect 46020 17756 46072 17808
rect 32312 17688 32364 17740
rect 33600 17688 33652 17740
rect 34152 17731 34204 17740
rect 34152 17697 34161 17731
rect 34161 17697 34195 17731
rect 34195 17697 34204 17731
rect 34152 17688 34204 17697
rect 15936 17484 15988 17536
rect 16672 17527 16724 17536
rect 16672 17493 16681 17527
rect 16681 17493 16715 17527
rect 16715 17493 16724 17527
rect 16672 17484 16724 17493
rect 17316 17527 17368 17536
rect 17316 17493 17325 17527
rect 17325 17493 17359 17527
rect 17359 17493 17368 17527
rect 17316 17484 17368 17493
rect 17684 17527 17736 17536
rect 17684 17493 17693 17527
rect 17693 17493 17727 17527
rect 17727 17493 17736 17527
rect 17684 17484 17736 17493
rect 18328 17552 18380 17604
rect 18788 17552 18840 17604
rect 19156 17552 19208 17604
rect 19800 17596 19852 17648
rect 22836 17620 22888 17672
rect 23112 17620 23164 17672
rect 20812 17552 20864 17604
rect 21272 17552 21324 17604
rect 23664 17552 23716 17604
rect 23756 17595 23808 17604
rect 23756 17561 23765 17595
rect 23765 17561 23799 17595
rect 23799 17561 23808 17595
rect 23756 17552 23808 17561
rect 24768 17552 24820 17604
rect 19800 17484 19852 17536
rect 21364 17484 21416 17536
rect 21916 17484 21968 17536
rect 23480 17484 23532 17536
rect 23848 17527 23900 17536
rect 23848 17493 23857 17527
rect 23857 17493 23891 17527
rect 23891 17493 23900 17527
rect 23848 17484 23900 17493
rect 24124 17484 24176 17536
rect 26424 17552 26476 17604
rect 28356 17620 28408 17672
rect 32588 17620 32640 17672
rect 34520 17688 34572 17740
rect 34704 17688 34756 17740
rect 35532 17731 35584 17740
rect 35532 17697 35541 17731
rect 35541 17697 35575 17731
rect 35575 17697 35584 17731
rect 35532 17688 35584 17697
rect 35808 17688 35860 17740
rect 35992 17688 36044 17740
rect 34428 17620 34480 17672
rect 38292 17688 38344 17740
rect 38384 17688 38436 17740
rect 38016 17620 38068 17672
rect 39856 17688 39908 17740
rect 40040 17731 40092 17740
rect 40040 17697 40049 17731
rect 40049 17697 40083 17731
rect 40083 17697 40092 17731
rect 40040 17688 40092 17697
rect 43996 17688 44048 17740
rect 44456 17731 44508 17740
rect 44456 17697 44465 17731
rect 44465 17697 44499 17731
rect 44499 17697 44508 17731
rect 44456 17688 44508 17697
rect 27896 17552 27948 17604
rect 27068 17484 27120 17536
rect 27436 17484 27488 17536
rect 28448 17527 28500 17536
rect 28448 17493 28457 17527
rect 28457 17493 28491 17527
rect 28491 17493 28500 17527
rect 28448 17484 28500 17493
rect 28540 17484 28592 17536
rect 29000 17484 29052 17536
rect 29736 17527 29788 17536
rect 29736 17493 29745 17527
rect 29745 17493 29779 17527
rect 29779 17493 29788 17527
rect 29736 17484 29788 17493
rect 30104 17527 30156 17536
rect 30104 17493 30113 17527
rect 30113 17493 30147 17527
rect 30147 17493 30156 17527
rect 30104 17484 30156 17493
rect 30196 17527 30248 17536
rect 30196 17493 30205 17527
rect 30205 17493 30239 17527
rect 30239 17493 30248 17527
rect 30196 17484 30248 17493
rect 30932 17484 30984 17536
rect 35808 17552 35860 17604
rect 34060 17484 34112 17536
rect 36820 17552 36872 17604
rect 36176 17484 36228 17536
rect 38476 17484 38528 17536
rect 39396 17552 39448 17604
rect 39120 17527 39172 17536
rect 39120 17493 39129 17527
rect 39129 17493 39163 17527
rect 39163 17493 39172 17527
rect 39120 17484 39172 17493
rect 39212 17484 39264 17536
rect 39488 17484 39540 17536
rect 42248 17663 42300 17672
rect 42248 17629 42257 17663
rect 42257 17629 42291 17663
rect 42291 17629 42300 17663
rect 42248 17620 42300 17629
rect 40776 17552 40828 17604
rect 44732 17552 44784 17604
rect 46020 17620 46072 17672
rect 48412 17620 48464 17672
rect 48504 17663 48556 17672
rect 48504 17629 48513 17663
rect 48513 17629 48547 17663
rect 48547 17629 48556 17663
rect 48504 17620 48556 17629
rect 47584 17552 47636 17604
rect 42616 17484 42668 17536
rect 43352 17484 43404 17536
rect 45836 17527 45888 17536
rect 45836 17493 45845 17527
rect 45845 17493 45879 17527
rect 45879 17493 45888 17527
rect 45836 17484 45888 17493
rect 45928 17484 45980 17536
rect 47124 17484 47176 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 49976 17348 50028 17400
rect 50712 17348 50764 17400
rect 1768 17280 1820 17332
rect 4620 17280 4672 17332
rect 6368 17280 6420 17332
rect 7380 17280 7432 17332
rect 4804 17212 4856 17264
rect 1860 17144 1912 17196
rect 2780 17144 2832 17196
rect 1308 17076 1360 17128
rect 4344 17144 4396 17196
rect 5448 17144 5500 17196
rect 8116 17212 8168 17264
rect 6736 17144 6788 17196
rect 12072 17280 12124 17332
rect 12440 17323 12492 17332
rect 12440 17289 12449 17323
rect 12449 17289 12483 17323
rect 12483 17289 12492 17323
rect 12440 17280 12492 17289
rect 7012 17076 7064 17128
rect 8484 17076 8536 17128
rect 7748 17008 7800 17060
rect 9956 17255 10008 17264
rect 9956 17221 9965 17255
rect 9965 17221 9999 17255
rect 9999 17221 10008 17255
rect 9956 17212 10008 17221
rect 13820 17280 13872 17332
rect 14464 17280 14516 17332
rect 15476 17280 15528 17332
rect 13268 17212 13320 17264
rect 10232 17144 10284 17196
rect 10968 17144 11020 17196
rect 13912 17212 13964 17264
rect 17040 17212 17092 17264
rect 10048 17076 10100 17128
rect 10600 17076 10652 17128
rect 12624 17119 12676 17128
rect 12624 17085 12633 17119
rect 12633 17085 12667 17119
rect 12667 17085 12676 17119
rect 12624 17076 12676 17085
rect 15016 17144 15068 17196
rect 15476 17144 15528 17196
rect 17500 17212 17552 17264
rect 17960 17212 18012 17264
rect 19616 17255 19668 17264
rect 19616 17221 19625 17255
rect 19625 17221 19659 17255
rect 19659 17221 19668 17255
rect 19616 17212 19668 17221
rect 18696 17144 18748 17196
rect 15752 17076 15804 17128
rect 16028 17119 16080 17128
rect 16028 17085 16037 17119
rect 16037 17085 16071 17119
rect 16071 17085 16080 17119
rect 16028 17076 16080 17085
rect 16120 17119 16172 17128
rect 16120 17085 16129 17119
rect 16129 17085 16163 17119
rect 16163 17085 16172 17119
rect 16120 17076 16172 17085
rect 16304 17076 16356 17128
rect 19248 17144 19300 17196
rect 20996 17144 21048 17196
rect 24860 17280 24912 17332
rect 25412 17280 25464 17332
rect 26792 17280 26844 17332
rect 30104 17280 30156 17332
rect 31944 17280 31996 17332
rect 32036 17280 32088 17332
rect 32680 17280 32732 17332
rect 24124 17212 24176 17264
rect 26424 17212 26476 17264
rect 27436 17212 27488 17264
rect 28816 17212 28868 17264
rect 30472 17212 30524 17264
rect 31208 17212 31260 17264
rect 23112 17187 23164 17196
rect 23112 17153 23121 17187
rect 23121 17153 23155 17187
rect 23155 17153 23164 17187
rect 23112 17144 23164 17153
rect 25412 17144 25464 17196
rect 26148 17144 26200 17196
rect 26240 17144 26292 17196
rect 27252 17144 27304 17196
rect 30748 17144 30800 17196
rect 21272 17076 21324 17128
rect 22376 17076 22428 17128
rect 25504 17076 25556 17128
rect 25596 17076 25648 17128
rect 26608 17076 26660 17128
rect 26700 17119 26752 17128
rect 26700 17085 26709 17119
rect 26709 17085 26743 17119
rect 26743 17085 26752 17119
rect 26700 17076 26752 17085
rect 30012 17076 30064 17128
rect 31576 17144 31628 17196
rect 31852 17144 31904 17196
rect 2044 16940 2096 16992
rect 3608 16940 3660 16992
rect 9128 16940 9180 16992
rect 10048 16940 10100 16992
rect 10416 16983 10468 16992
rect 10416 16949 10425 16983
rect 10425 16949 10459 16983
rect 10459 16949 10468 16983
rect 10416 16940 10468 16949
rect 11796 17051 11848 17060
rect 11796 17017 11805 17051
rect 11805 17017 11839 17051
rect 11839 17017 11848 17051
rect 11796 17008 11848 17017
rect 16212 17008 16264 17060
rect 18512 17008 18564 17060
rect 18696 17008 18748 17060
rect 20720 17008 20772 17060
rect 20904 17008 20956 17060
rect 22008 17008 22060 17060
rect 12072 16983 12124 16992
rect 12072 16949 12081 16983
rect 12081 16949 12115 16983
rect 12115 16949 12124 16983
rect 12072 16940 12124 16949
rect 15108 16983 15160 16992
rect 15108 16949 15117 16983
rect 15117 16949 15151 16983
rect 15151 16949 15160 16983
rect 15108 16940 15160 16949
rect 17960 16940 18012 16992
rect 18052 16940 18104 16992
rect 19156 16940 19208 16992
rect 20352 16940 20404 16992
rect 22192 16940 22244 16992
rect 24492 17008 24544 17060
rect 27712 17008 27764 17060
rect 29552 17008 29604 17060
rect 30380 17008 30432 17060
rect 30748 17008 30800 17060
rect 31668 17076 31720 17128
rect 32864 17255 32916 17264
rect 32864 17221 32873 17255
rect 32873 17221 32907 17255
rect 32907 17221 32916 17255
rect 32864 17212 32916 17221
rect 34888 17280 34940 17332
rect 35532 17280 35584 17332
rect 32312 17144 32364 17196
rect 34520 17144 34572 17196
rect 32128 17076 32180 17128
rect 33324 17076 33376 17128
rect 37280 17212 37332 17264
rect 37556 17280 37608 17332
rect 38200 17280 38252 17332
rect 38844 17280 38896 17332
rect 39028 17280 39080 17332
rect 39120 17280 39172 17332
rect 40960 17280 41012 17332
rect 48412 17323 48464 17332
rect 48412 17289 48421 17323
rect 48421 17289 48455 17323
rect 48455 17289 48464 17323
rect 48412 17280 48464 17289
rect 49056 17280 49108 17332
rect 40776 17212 40828 17264
rect 41144 17212 41196 17264
rect 35532 17144 35584 17196
rect 36544 17144 36596 17196
rect 35716 17076 35768 17128
rect 31484 17008 31536 17060
rect 32588 17008 32640 17060
rect 33876 17008 33928 17060
rect 36636 17119 36688 17128
rect 36636 17085 36645 17119
rect 36645 17085 36679 17119
rect 36679 17085 36688 17119
rect 36636 17076 36688 17085
rect 36820 17076 36872 17128
rect 37464 17187 37516 17196
rect 37464 17153 37473 17187
rect 37473 17153 37507 17187
rect 37507 17153 37516 17187
rect 37464 17144 37516 17153
rect 38292 17144 38344 17196
rect 41236 17187 41288 17196
rect 41236 17153 41245 17187
rect 41245 17153 41279 17187
rect 41279 17153 41288 17187
rect 41236 17144 41288 17153
rect 45836 17212 45888 17264
rect 47124 17212 47176 17264
rect 38384 17076 38436 17128
rect 42156 17187 42208 17196
rect 42156 17153 42165 17187
rect 42165 17153 42199 17187
rect 42199 17153 42208 17187
rect 42156 17144 42208 17153
rect 42616 17187 42668 17196
rect 42616 17153 42625 17187
rect 42625 17153 42659 17187
rect 42659 17153 42668 17187
rect 42616 17144 42668 17153
rect 43720 17187 43772 17196
rect 43720 17153 43729 17187
rect 43729 17153 43763 17187
rect 43763 17153 43772 17187
rect 43720 17144 43772 17153
rect 45468 17144 45520 17196
rect 45928 17187 45980 17196
rect 45928 17153 45937 17187
rect 45937 17153 45971 17187
rect 45971 17153 45980 17187
rect 45928 17144 45980 17153
rect 41512 17119 41564 17128
rect 41512 17085 41521 17119
rect 41521 17085 41555 17119
rect 41555 17085 41564 17119
rect 41512 17076 41564 17085
rect 43260 17119 43312 17128
rect 43260 17085 43269 17119
rect 43269 17085 43303 17119
rect 43303 17085 43312 17119
rect 43260 17076 43312 17085
rect 44088 17076 44140 17128
rect 47124 17076 47176 17128
rect 49148 17212 49200 17264
rect 48780 17144 48832 17196
rect 49056 17144 49108 17196
rect 49884 17076 49936 17128
rect 28356 16940 28408 16992
rect 29184 16940 29236 16992
rect 29644 16940 29696 16992
rect 30012 16983 30064 16992
rect 30012 16949 30021 16983
rect 30021 16949 30055 16983
rect 30055 16949 30064 16983
rect 30012 16940 30064 16949
rect 31208 16940 31260 16992
rect 31852 16983 31904 16992
rect 31852 16949 31861 16983
rect 31861 16949 31895 16983
rect 31895 16949 31904 16983
rect 31852 16940 31904 16949
rect 32864 16940 32916 16992
rect 34336 16983 34388 16992
rect 34336 16949 34345 16983
rect 34345 16949 34379 16983
rect 34379 16949 34388 16983
rect 34336 16940 34388 16949
rect 35900 16940 35952 16992
rect 37648 17008 37700 17060
rect 38200 16940 38252 16992
rect 44732 17008 44784 17060
rect 46480 17008 46532 17060
rect 46756 17008 46808 17060
rect 47768 17008 47820 17060
rect 40960 16940 41012 16992
rect 41420 16940 41472 16992
rect 44088 16940 44140 16992
rect 44272 16940 44324 16992
rect 45560 16940 45612 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 2872 16736 2924 16788
rect 5356 16668 5408 16720
rect 7196 16668 7248 16720
rect 3884 16532 3936 16584
rect 5264 16532 5316 16584
rect 1308 16464 1360 16516
rect 5448 16532 5500 16584
rect 8300 16736 8352 16788
rect 8944 16736 8996 16788
rect 10048 16736 10100 16788
rect 10968 16736 11020 16788
rect 11060 16736 11112 16788
rect 12164 16668 12216 16720
rect 12624 16736 12676 16788
rect 13636 16736 13688 16788
rect 13820 16779 13872 16788
rect 13820 16745 13829 16779
rect 13829 16745 13863 16779
rect 13863 16745 13872 16779
rect 13820 16736 13872 16745
rect 16028 16736 16080 16788
rect 17776 16736 17828 16788
rect 17868 16779 17920 16788
rect 17868 16745 17877 16779
rect 17877 16745 17911 16779
rect 17911 16745 17920 16779
rect 17868 16736 17920 16745
rect 17960 16736 18012 16788
rect 18972 16779 19024 16788
rect 18972 16745 18981 16779
rect 18981 16745 19015 16779
rect 19015 16745 19024 16779
rect 18972 16736 19024 16745
rect 20996 16736 21048 16788
rect 16120 16668 16172 16720
rect 16212 16668 16264 16720
rect 18052 16668 18104 16720
rect 8116 16643 8168 16652
rect 8116 16609 8125 16643
rect 8125 16609 8159 16643
rect 8159 16609 8168 16643
rect 8116 16600 8168 16609
rect 8944 16600 8996 16652
rect 6368 16464 6420 16516
rect 9128 16532 9180 16584
rect 9220 16575 9272 16584
rect 9220 16541 9229 16575
rect 9229 16541 9263 16575
rect 9263 16541 9272 16575
rect 9220 16532 9272 16541
rect 10968 16575 11020 16584
rect 10968 16541 10977 16575
rect 10977 16541 11011 16575
rect 11011 16541 11020 16575
rect 10968 16532 11020 16541
rect 11612 16600 11664 16652
rect 13268 16643 13320 16652
rect 13268 16609 13277 16643
rect 13277 16609 13311 16643
rect 13311 16609 13320 16643
rect 13268 16600 13320 16609
rect 13820 16600 13872 16652
rect 11060 16464 11112 16516
rect 11152 16464 11204 16516
rect 13544 16532 13596 16584
rect 14648 16575 14700 16584
rect 14648 16541 14657 16575
rect 14657 16541 14691 16575
rect 14691 16541 14700 16575
rect 14648 16532 14700 16541
rect 14740 16575 14792 16584
rect 14740 16541 14749 16575
rect 14749 16541 14783 16575
rect 14783 16541 14792 16575
rect 14740 16532 14792 16541
rect 15752 16600 15804 16652
rect 17960 16600 18012 16652
rect 15108 16532 15160 16584
rect 3608 16396 3660 16448
rect 5908 16396 5960 16448
rect 6828 16396 6880 16448
rect 7196 16396 7248 16448
rect 9036 16396 9088 16448
rect 9220 16396 9272 16448
rect 10876 16396 10928 16448
rect 11796 16439 11848 16448
rect 11796 16405 11805 16439
rect 11805 16405 11839 16439
rect 11839 16405 11848 16439
rect 11796 16396 11848 16405
rect 11888 16439 11940 16448
rect 11888 16405 11897 16439
rect 11897 16405 11931 16439
rect 11931 16405 11940 16439
rect 11888 16396 11940 16405
rect 12348 16396 12400 16448
rect 12440 16396 12492 16448
rect 12992 16439 13044 16448
rect 12992 16405 13001 16439
rect 13001 16405 13035 16439
rect 13035 16405 13044 16439
rect 12992 16396 13044 16405
rect 13544 16396 13596 16448
rect 13820 16464 13872 16516
rect 16580 16532 16632 16584
rect 16764 16575 16816 16584
rect 16764 16541 16773 16575
rect 16773 16541 16807 16575
rect 16807 16541 16816 16575
rect 16764 16532 16816 16541
rect 19156 16668 19208 16720
rect 21732 16736 21784 16788
rect 21916 16736 21968 16788
rect 23756 16736 23808 16788
rect 24308 16736 24360 16788
rect 26608 16736 26660 16788
rect 26700 16736 26752 16788
rect 27988 16736 28040 16788
rect 29552 16779 29604 16788
rect 18972 16600 19024 16652
rect 19708 16600 19760 16652
rect 20352 16600 20404 16652
rect 16396 16464 16448 16516
rect 14464 16396 14516 16448
rect 15016 16396 15068 16448
rect 17868 16464 17920 16516
rect 16856 16396 16908 16448
rect 27528 16668 27580 16720
rect 29552 16745 29561 16779
rect 29561 16745 29595 16779
rect 29595 16745 29604 16779
rect 29552 16736 29604 16745
rect 29644 16736 29696 16788
rect 30012 16736 30064 16788
rect 30196 16736 30248 16788
rect 33324 16736 33376 16788
rect 33692 16736 33744 16788
rect 34244 16736 34296 16788
rect 34704 16736 34756 16788
rect 35532 16736 35584 16788
rect 20720 16643 20772 16652
rect 20720 16609 20729 16643
rect 20729 16609 20763 16643
rect 20763 16609 20772 16643
rect 20720 16600 20772 16609
rect 20812 16600 20864 16652
rect 22836 16600 22888 16652
rect 24768 16600 24820 16652
rect 25964 16600 26016 16652
rect 27344 16600 27396 16652
rect 29828 16668 29880 16720
rect 27988 16643 28040 16652
rect 27988 16609 27997 16643
rect 27997 16609 28031 16643
rect 28031 16609 28040 16643
rect 27988 16600 28040 16609
rect 28540 16600 28592 16652
rect 28816 16600 28868 16652
rect 30012 16600 30064 16652
rect 30104 16643 30156 16652
rect 30104 16609 30113 16643
rect 30113 16609 30147 16643
rect 30147 16609 30156 16643
rect 30104 16600 30156 16609
rect 33324 16600 33376 16652
rect 33416 16600 33468 16652
rect 22376 16532 22428 16584
rect 23388 16532 23440 16584
rect 24124 16532 24176 16584
rect 18236 16439 18288 16448
rect 18236 16405 18245 16439
rect 18245 16405 18279 16439
rect 18279 16405 18288 16439
rect 18236 16396 18288 16405
rect 18604 16396 18656 16448
rect 19432 16439 19484 16448
rect 19432 16405 19441 16439
rect 19441 16405 19475 16439
rect 19475 16405 19484 16439
rect 19432 16396 19484 16405
rect 19800 16439 19852 16448
rect 19800 16405 19809 16439
rect 19809 16405 19843 16439
rect 19843 16405 19852 16439
rect 19800 16396 19852 16405
rect 19892 16396 19944 16448
rect 23848 16464 23900 16516
rect 27896 16575 27948 16584
rect 27896 16541 27905 16575
rect 27905 16541 27939 16575
rect 27939 16541 27948 16575
rect 27896 16532 27948 16541
rect 29276 16532 29328 16584
rect 29552 16532 29604 16584
rect 31484 16532 31536 16584
rect 31944 16532 31996 16584
rect 23296 16439 23348 16448
rect 23296 16405 23305 16439
rect 23305 16405 23339 16439
rect 23339 16405 23348 16439
rect 23296 16396 23348 16405
rect 23664 16439 23716 16448
rect 23664 16405 23673 16439
rect 23673 16405 23707 16439
rect 23707 16405 23716 16439
rect 23664 16396 23716 16405
rect 24492 16396 24544 16448
rect 26148 16396 26200 16448
rect 26700 16439 26752 16448
rect 26700 16405 26709 16439
rect 26709 16405 26743 16439
rect 26743 16405 26752 16439
rect 26700 16396 26752 16405
rect 27620 16464 27672 16516
rect 28724 16464 28776 16516
rect 30656 16464 30708 16516
rect 34428 16600 34480 16652
rect 38108 16736 38160 16788
rect 38752 16736 38804 16788
rect 38200 16668 38252 16720
rect 38568 16668 38620 16720
rect 41328 16736 41380 16788
rect 42248 16736 42300 16788
rect 43720 16736 43772 16788
rect 44824 16736 44876 16788
rect 38844 16600 38896 16652
rect 39304 16600 39356 16652
rect 39488 16643 39540 16652
rect 39488 16609 39497 16643
rect 39497 16609 39531 16643
rect 39531 16609 39540 16643
rect 39488 16600 39540 16609
rect 40224 16600 40276 16652
rect 40500 16643 40552 16652
rect 40500 16609 40509 16643
rect 40509 16609 40543 16643
rect 40543 16609 40552 16643
rect 40500 16600 40552 16609
rect 40960 16600 41012 16652
rect 44548 16668 44600 16720
rect 45192 16668 45244 16720
rect 45836 16668 45888 16720
rect 47216 16668 47268 16720
rect 41972 16600 42024 16652
rect 44272 16600 44324 16652
rect 48412 16600 48464 16652
rect 48964 16600 49016 16652
rect 34888 16575 34940 16584
rect 34888 16541 34897 16575
rect 34897 16541 34931 16575
rect 34931 16541 34940 16575
rect 34888 16532 34940 16541
rect 27712 16396 27764 16448
rect 28908 16439 28960 16448
rect 28908 16405 28917 16439
rect 28917 16405 28951 16439
rect 28951 16405 28960 16439
rect 28908 16396 28960 16405
rect 33324 16396 33376 16448
rect 33600 16396 33652 16448
rect 33692 16396 33744 16448
rect 35808 16464 35860 16516
rect 43352 16532 43404 16584
rect 44364 16532 44416 16584
rect 44456 16532 44508 16584
rect 45192 16575 45244 16584
rect 45192 16541 45201 16575
rect 45201 16541 45235 16575
rect 45235 16541 45244 16575
rect 45192 16532 45244 16541
rect 45468 16532 45520 16584
rect 37740 16464 37792 16516
rect 36636 16439 36688 16448
rect 36636 16405 36645 16439
rect 36645 16405 36679 16439
rect 36679 16405 36688 16439
rect 36636 16396 36688 16405
rect 39488 16464 39540 16516
rect 41880 16464 41932 16516
rect 45376 16464 45428 16516
rect 47216 16532 47268 16584
rect 48780 16532 48832 16584
rect 49240 16464 49292 16516
rect 38384 16396 38436 16448
rect 38660 16439 38712 16448
rect 38660 16405 38669 16439
rect 38669 16405 38703 16439
rect 38703 16405 38712 16439
rect 38660 16396 38712 16405
rect 38752 16439 38804 16448
rect 38752 16405 38761 16439
rect 38761 16405 38795 16439
rect 38795 16405 38804 16439
rect 38752 16396 38804 16405
rect 39672 16396 39724 16448
rect 40040 16439 40092 16448
rect 40040 16405 40049 16439
rect 40049 16405 40083 16439
rect 40083 16405 40092 16439
rect 40040 16396 40092 16405
rect 42248 16396 42300 16448
rect 45468 16396 45520 16448
rect 45928 16396 45980 16448
rect 47032 16396 47084 16448
rect 47400 16396 47452 16448
rect 48504 16396 48556 16448
rect 48964 16396 49016 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 6000 16235 6052 16244
rect 6000 16201 6009 16235
rect 6009 16201 6043 16235
rect 6043 16201 6052 16235
rect 6000 16192 6052 16201
rect 6368 16192 6420 16244
rect 7748 16192 7800 16244
rect 7840 16192 7892 16244
rect 3976 16124 4028 16176
rect 7104 16124 7156 16176
rect 1768 16099 1820 16108
rect 1768 16065 1777 16099
rect 1777 16065 1811 16099
rect 1811 16065 1820 16099
rect 1768 16056 1820 16065
rect 3608 16099 3660 16108
rect 3608 16065 3617 16099
rect 3617 16065 3651 16099
rect 3651 16065 3660 16099
rect 3608 16056 3660 16065
rect 5264 16056 5316 16108
rect 1308 15988 1360 16040
rect 3884 15988 3936 16040
rect 6460 16056 6512 16108
rect 8116 16099 8168 16108
rect 8116 16065 8125 16099
rect 8125 16065 8159 16099
rect 8159 16065 8168 16099
rect 8116 16056 8168 16065
rect 8852 16192 8904 16244
rect 8668 16124 8720 16176
rect 10784 16124 10836 16176
rect 11888 16192 11940 16244
rect 12440 16235 12492 16244
rect 12440 16201 12449 16235
rect 12449 16201 12483 16235
rect 12483 16201 12492 16235
rect 12440 16192 12492 16201
rect 12164 16124 12216 16176
rect 13452 16192 13504 16244
rect 14832 16235 14884 16244
rect 14832 16201 14841 16235
rect 14841 16201 14875 16235
rect 14875 16201 14884 16235
rect 14832 16192 14884 16201
rect 15384 16192 15436 16244
rect 15568 16192 15620 16244
rect 16028 16235 16080 16244
rect 16028 16201 16037 16235
rect 16037 16201 16071 16235
rect 16071 16201 16080 16235
rect 16028 16192 16080 16201
rect 16396 16192 16448 16244
rect 20904 16192 20956 16244
rect 21180 16192 21232 16244
rect 23296 16192 23348 16244
rect 24308 16192 24360 16244
rect 24860 16192 24912 16244
rect 25872 16192 25924 16244
rect 26700 16192 26752 16244
rect 27344 16192 27396 16244
rect 28908 16192 28960 16244
rect 30656 16192 30708 16244
rect 30840 16192 30892 16244
rect 31576 16192 31628 16244
rect 31852 16192 31904 16244
rect 31944 16235 31996 16244
rect 31944 16201 31953 16235
rect 31953 16201 31987 16235
rect 31987 16201 31996 16235
rect 31944 16192 31996 16201
rect 32220 16192 32272 16244
rect 32404 16192 32456 16244
rect 32864 16192 32916 16244
rect 34704 16192 34756 16244
rect 4804 15852 4856 15904
rect 5816 15988 5868 16040
rect 8576 16056 8628 16108
rect 10508 16099 10560 16108
rect 10508 16065 10517 16099
rect 10517 16065 10551 16099
rect 10551 16065 10560 16099
rect 10508 16056 10560 16065
rect 14556 16124 14608 16176
rect 9036 15988 9088 16040
rect 7748 15963 7800 15972
rect 7748 15929 7757 15963
rect 7757 15929 7791 15963
rect 7791 15929 7800 15963
rect 7748 15920 7800 15929
rect 7932 15920 7984 15972
rect 13544 16056 13596 16108
rect 13912 16056 13964 16108
rect 14740 16099 14792 16108
rect 14740 16065 14749 16099
rect 14749 16065 14783 16099
rect 14783 16065 14792 16099
rect 14740 16056 14792 16065
rect 13268 15988 13320 16040
rect 13728 16031 13780 16040
rect 13728 15997 13737 16031
rect 13737 15997 13771 16031
rect 13771 15997 13780 16031
rect 13728 15988 13780 15997
rect 15108 15988 15160 16040
rect 16120 16031 16172 16040
rect 16120 15997 16129 16031
rect 16129 15997 16163 16031
rect 16163 15997 16172 16031
rect 16120 15988 16172 15997
rect 16304 15988 16356 16040
rect 16856 16167 16908 16176
rect 16856 16133 16865 16167
rect 16865 16133 16899 16167
rect 16899 16133 16908 16167
rect 16856 16124 16908 16133
rect 17776 16124 17828 16176
rect 17960 16124 18012 16176
rect 20720 16124 20772 16176
rect 17408 15988 17460 16040
rect 18604 16056 18656 16108
rect 18696 16099 18748 16108
rect 18696 16065 18705 16099
rect 18705 16065 18739 16099
rect 18739 16065 18748 16099
rect 18696 16056 18748 16065
rect 19156 16099 19208 16108
rect 19156 16065 19165 16099
rect 19165 16065 19199 16099
rect 19199 16065 19208 16099
rect 19156 16056 19208 16065
rect 20996 16056 21048 16108
rect 21088 16056 21140 16108
rect 21640 16056 21692 16108
rect 9312 15920 9364 15972
rect 11060 15920 11112 15972
rect 16580 15920 16632 15972
rect 18788 15988 18840 16040
rect 17868 15920 17920 15972
rect 18512 15920 18564 15972
rect 8300 15852 8352 15904
rect 8852 15895 8904 15904
rect 8852 15861 8861 15895
rect 8861 15861 8895 15895
rect 8895 15861 8904 15895
rect 8852 15852 8904 15861
rect 8944 15852 8996 15904
rect 10600 15852 10652 15904
rect 11888 15852 11940 15904
rect 12164 15852 12216 15904
rect 13912 15852 13964 15904
rect 14740 15852 14792 15904
rect 16304 15852 16356 15904
rect 17224 15895 17276 15904
rect 17224 15861 17233 15895
rect 17233 15861 17267 15895
rect 17267 15861 17276 15895
rect 17224 15852 17276 15861
rect 17592 15852 17644 15904
rect 17960 15852 18012 15904
rect 18788 15852 18840 15904
rect 19616 15852 19668 15904
rect 20904 15988 20956 16040
rect 23848 16056 23900 16108
rect 24768 16056 24820 16108
rect 25320 16056 25372 16108
rect 25780 16056 25832 16108
rect 26700 16099 26752 16108
rect 22468 16031 22520 16040
rect 22468 15997 22477 16031
rect 22477 15997 22511 16031
rect 22511 15997 22520 16031
rect 22468 15988 22520 15997
rect 20628 15920 20680 15972
rect 20996 15852 21048 15904
rect 21364 15852 21416 15904
rect 21640 15852 21692 15904
rect 22836 15988 22888 16040
rect 24400 15988 24452 16040
rect 25044 16031 25096 16040
rect 25044 15997 25053 16031
rect 25053 15997 25087 16031
rect 25087 15997 25096 16031
rect 25044 15988 25096 15997
rect 25872 15988 25924 16040
rect 26700 16065 26709 16099
rect 26709 16065 26743 16099
rect 26743 16065 26752 16099
rect 26700 16056 26752 16065
rect 26884 16124 26936 16176
rect 27344 16056 27396 16108
rect 23572 15920 23624 15972
rect 25780 15920 25832 15972
rect 27620 15988 27672 16040
rect 28356 16099 28408 16108
rect 28356 16065 28365 16099
rect 28365 16065 28399 16099
rect 28399 16065 28408 16099
rect 28356 16056 28408 16065
rect 29276 15988 29328 16040
rect 27252 15920 27304 15972
rect 33692 16124 33744 16176
rect 34796 16124 34848 16176
rect 35164 16124 35216 16176
rect 35808 16124 35860 16176
rect 29644 16056 29696 16108
rect 23296 15852 23348 15904
rect 24492 15852 24544 15904
rect 26792 15852 26844 15904
rect 27344 15852 27396 15904
rect 27712 15852 27764 15904
rect 30196 16031 30248 16040
rect 30196 15997 30205 16031
rect 30205 15997 30239 16031
rect 30239 15997 30248 16031
rect 30196 15988 30248 15997
rect 30564 16056 30616 16108
rect 32404 16056 32456 16108
rect 34152 16056 34204 16108
rect 34888 16056 34940 16108
rect 30380 15920 30432 15972
rect 32128 15988 32180 16040
rect 32312 15920 32364 15972
rect 33968 16031 34020 16040
rect 33968 15997 33977 16031
rect 33977 15997 34011 16031
rect 34011 15997 34020 16031
rect 33968 15988 34020 15997
rect 34336 15988 34388 16040
rect 38476 16124 38528 16176
rect 38568 16167 38620 16176
rect 38568 16133 38577 16167
rect 38577 16133 38611 16167
rect 38611 16133 38620 16167
rect 38568 16124 38620 16133
rect 40040 16192 40092 16244
rect 41328 16192 41380 16244
rect 42708 16124 42760 16176
rect 44364 16235 44416 16244
rect 44364 16201 44373 16235
rect 44373 16201 44407 16235
rect 44407 16201 44416 16235
rect 44364 16192 44416 16201
rect 44548 16192 44600 16244
rect 48780 16235 48832 16244
rect 48780 16201 48789 16235
rect 48789 16201 48823 16235
rect 48823 16201 48832 16235
rect 48780 16192 48832 16201
rect 45560 16124 45612 16176
rect 36820 16056 36872 16108
rect 38292 16099 38344 16108
rect 38292 16065 38301 16099
rect 38301 16065 38335 16099
rect 38335 16065 38344 16099
rect 38292 16056 38344 16065
rect 39672 16056 39724 16108
rect 40408 16099 40460 16108
rect 40408 16065 40417 16099
rect 40417 16065 40451 16099
rect 40451 16065 40460 16099
rect 40408 16056 40460 16065
rect 41144 16099 41196 16108
rect 41144 16065 41153 16099
rect 41153 16065 41187 16099
rect 41187 16065 41196 16099
rect 41144 16056 41196 16065
rect 36636 15988 36688 16040
rect 41328 16031 41380 16040
rect 41328 15997 41337 16031
rect 41337 15997 41371 16031
rect 41371 15997 41380 16031
rect 41328 15988 41380 15997
rect 42064 15988 42116 16040
rect 42340 15988 42392 16040
rect 42616 16099 42668 16108
rect 42616 16065 42625 16099
rect 42625 16065 42659 16099
rect 42659 16065 42668 16099
rect 42616 16056 42668 16065
rect 44824 16099 44876 16108
rect 44824 16065 44833 16099
rect 44833 16065 44867 16099
rect 44867 16065 44876 16099
rect 44824 16056 44876 16065
rect 46572 16124 46624 16176
rect 44364 15988 44416 16040
rect 45928 16099 45980 16108
rect 45928 16065 45937 16099
rect 45937 16065 45971 16099
rect 45971 16065 45980 16099
rect 45928 16056 45980 16065
rect 47400 16124 47452 16176
rect 48320 16124 48372 16176
rect 45468 15988 45520 16040
rect 49240 16056 49292 16108
rect 36820 15920 36872 15972
rect 37004 15920 37056 15972
rect 30288 15852 30340 15904
rect 30564 15852 30616 15904
rect 30840 15895 30892 15904
rect 30840 15861 30849 15895
rect 30849 15861 30883 15895
rect 30883 15861 30892 15895
rect 30840 15852 30892 15861
rect 31944 15852 31996 15904
rect 33508 15852 33560 15904
rect 34704 15852 34756 15904
rect 35624 15852 35676 15904
rect 35808 15852 35860 15904
rect 37740 15895 37792 15904
rect 37740 15861 37749 15895
rect 37749 15861 37783 15895
rect 37783 15861 37792 15895
rect 37740 15852 37792 15861
rect 39856 15852 39908 15904
rect 45192 15920 45244 15972
rect 40960 15852 41012 15904
rect 41420 15852 41472 15904
rect 41880 15852 41932 15904
rect 42524 15852 42576 15904
rect 42800 15852 42852 15904
rect 45468 15895 45520 15904
rect 45468 15861 45477 15895
rect 45477 15861 45511 15895
rect 45511 15861 45520 15895
rect 45468 15852 45520 15861
rect 46572 15895 46624 15904
rect 46572 15861 46581 15895
rect 46581 15861 46615 15895
rect 46615 15861 46624 15895
rect 46572 15852 46624 15861
rect 47032 15852 47084 15904
rect 48780 15852 48832 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 3884 15648 3936 15700
rect 4068 15648 4120 15700
rect 5356 15648 5408 15700
rect 7380 15648 7432 15700
rect 7932 15648 7984 15700
rect 1308 15512 1360 15564
rect 7380 15512 7432 15564
rect 8116 15512 8168 15564
rect 3608 15444 3660 15496
rect 3424 15376 3476 15428
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 4620 15444 4672 15453
rect 5724 15487 5776 15496
rect 5724 15453 5733 15487
rect 5733 15453 5767 15487
rect 5767 15453 5776 15487
rect 5724 15444 5776 15453
rect 6828 15487 6880 15496
rect 6828 15453 6837 15487
rect 6837 15453 6871 15487
rect 6871 15453 6880 15487
rect 6828 15444 6880 15453
rect 8484 15580 8536 15632
rect 8300 15512 8352 15564
rect 9220 15580 9272 15632
rect 10048 15512 10100 15564
rect 10784 15512 10836 15564
rect 11704 15648 11756 15700
rect 12440 15648 12492 15700
rect 13452 15648 13504 15700
rect 11796 15580 11848 15632
rect 15292 15648 15344 15700
rect 12808 15555 12860 15564
rect 12808 15521 12817 15555
rect 12817 15521 12851 15555
rect 12851 15521 12860 15555
rect 12808 15512 12860 15521
rect 12992 15555 13044 15564
rect 12992 15521 13001 15555
rect 13001 15521 13035 15555
rect 13035 15521 13044 15555
rect 12992 15512 13044 15521
rect 13360 15512 13412 15564
rect 13912 15512 13964 15564
rect 14740 15555 14792 15564
rect 14740 15521 14749 15555
rect 14749 15521 14783 15555
rect 14783 15521 14792 15555
rect 14740 15512 14792 15521
rect 14924 15555 14976 15564
rect 14924 15521 14933 15555
rect 14933 15521 14967 15555
rect 14967 15521 14976 15555
rect 14924 15512 14976 15521
rect 15752 15580 15804 15632
rect 16120 15580 16172 15632
rect 19524 15648 19576 15700
rect 19892 15648 19944 15700
rect 20444 15648 20496 15700
rect 20996 15648 21048 15700
rect 24124 15648 24176 15700
rect 24768 15648 24820 15700
rect 26240 15648 26292 15700
rect 26608 15691 26660 15700
rect 26608 15657 26617 15691
rect 26617 15657 26651 15691
rect 26651 15657 26660 15691
rect 26608 15648 26660 15657
rect 16028 15555 16080 15564
rect 16028 15521 16037 15555
rect 16037 15521 16071 15555
rect 16071 15521 16080 15555
rect 16028 15512 16080 15521
rect 16856 15512 16908 15564
rect 18696 15580 18748 15632
rect 5356 15376 5408 15428
rect 9496 15419 9548 15428
rect 9496 15385 9505 15419
rect 9505 15385 9539 15419
rect 9539 15385 9548 15419
rect 9496 15376 9548 15385
rect 16396 15444 16448 15496
rect 17408 15512 17460 15564
rect 20720 15512 20772 15564
rect 20812 15512 20864 15564
rect 21824 15580 21876 15632
rect 22284 15580 22336 15632
rect 21456 15555 21508 15564
rect 21456 15521 21465 15555
rect 21465 15521 21499 15555
rect 21499 15521 21508 15555
rect 21456 15512 21508 15521
rect 18420 15444 18472 15496
rect 22192 15444 22244 15496
rect 22652 15444 22704 15496
rect 12440 15376 12492 15428
rect 6644 15308 6696 15360
rect 9312 15308 9364 15360
rect 9588 15351 9640 15360
rect 9588 15317 9597 15351
rect 9597 15317 9631 15351
rect 9631 15317 9640 15351
rect 9588 15308 9640 15317
rect 11704 15308 11756 15360
rect 12164 15308 12216 15360
rect 12716 15351 12768 15360
rect 12716 15317 12725 15351
rect 12725 15317 12759 15351
rect 12759 15317 12768 15351
rect 12716 15308 12768 15317
rect 13636 15308 13688 15360
rect 15200 15308 15252 15360
rect 15752 15308 15804 15360
rect 16672 15308 16724 15360
rect 17132 15351 17184 15360
rect 17132 15317 17141 15351
rect 17141 15317 17175 15351
rect 17175 15317 17184 15351
rect 17132 15308 17184 15317
rect 17224 15308 17276 15360
rect 17408 15308 17460 15360
rect 21272 15419 21324 15428
rect 21272 15385 21281 15419
rect 21281 15385 21315 15419
rect 21315 15385 21324 15419
rect 21272 15376 21324 15385
rect 18420 15351 18472 15360
rect 18420 15317 18429 15351
rect 18429 15317 18463 15351
rect 18463 15317 18472 15351
rect 18420 15308 18472 15317
rect 19616 15308 19668 15360
rect 20260 15308 20312 15360
rect 21640 15376 21692 15428
rect 23572 15512 23624 15564
rect 24400 15512 24452 15564
rect 23296 15487 23348 15496
rect 23296 15453 23305 15487
rect 23305 15453 23339 15487
rect 23339 15453 23348 15487
rect 23296 15444 23348 15453
rect 26332 15512 26384 15564
rect 24952 15444 25004 15496
rect 25596 15444 25648 15496
rect 26148 15444 26200 15496
rect 24400 15376 24452 15428
rect 24676 15376 24728 15428
rect 25228 15376 25280 15428
rect 27528 15580 27580 15632
rect 29644 15580 29696 15632
rect 30196 15580 30248 15632
rect 27620 15555 27672 15564
rect 27620 15521 27629 15555
rect 27629 15521 27663 15555
rect 27663 15521 27672 15555
rect 27620 15512 27672 15521
rect 27712 15512 27764 15564
rect 28356 15512 28408 15564
rect 28908 15512 28960 15564
rect 29920 15512 29972 15564
rect 29736 15444 29788 15496
rect 30288 15555 30340 15564
rect 30288 15521 30297 15555
rect 30297 15521 30331 15555
rect 30331 15521 30340 15555
rect 30288 15512 30340 15521
rect 30564 15580 30616 15632
rect 32312 15580 32364 15632
rect 31944 15512 31996 15564
rect 32588 15512 32640 15564
rect 30380 15444 30432 15496
rect 30564 15444 30616 15496
rect 30840 15444 30892 15496
rect 32772 15444 32824 15496
rect 27528 15419 27580 15428
rect 27528 15385 27537 15419
rect 27537 15385 27571 15419
rect 27571 15385 27580 15419
rect 27528 15376 27580 15385
rect 22560 15308 22612 15360
rect 23480 15308 23532 15360
rect 23756 15308 23808 15360
rect 23848 15308 23900 15360
rect 24124 15308 24176 15360
rect 25044 15308 25096 15360
rect 27896 15376 27948 15428
rect 30840 15351 30892 15360
rect 30840 15317 30849 15351
rect 30849 15317 30883 15351
rect 30883 15317 30892 15351
rect 30840 15308 30892 15317
rect 32496 15376 32548 15428
rect 33416 15555 33468 15564
rect 33416 15521 33425 15555
rect 33425 15521 33459 15555
rect 33459 15521 33468 15555
rect 33416 15512 33468 15521
rect 34704 15648 34756 15700
rect 34152 15555 34204 15564
rect 34152 15521 34161 15555
rect 34161 15521 34195 15555
rect 34195 15521 34204 15555
rect 34152 15512 34204 15521
rect 34336 15512 34388 15564
rect 37096 15580 37148 15632
rect 35808 15555 35860 15564
rect 35808 15521 35817 15555
rect 35817 15521 35851 15555
rect 35851 15521 35860 15555
rect 35808 15512 35860 15521
rect 36360 15487 36412 15496
rect 36360 15453 36369 15487
rect 36369 15453 36403 15487
rect 36403 15453 36412 15487
rect 36360 15444 36412 15453
rect 37280 15376 37332 15428
rect 32956 15351 33008 15360
rect 32956 15317 32965 15351
rect 32965 15317 32999 15351
rect 32999 15317 33008 15351
rect 32956 15308 33008 15317
rect 34060 15308 34112 15360
rect 34612 15308 34664 15360
rect 35532 15351 35584 15360
rect 35532 15317 35541 15351
rect 35541 15317 35575 15351
rect 35575 15317 35584 15351
rect 35532 15308 35584 15317
rect 36820 15308 36872 15360
rect 37004 15351 37056 15360
rect 37004 15317 37013 15351
rect 37013 15317 37047 15351
rect 37047 15317 37056 15351
rect 37004 15308 37056 15317
rect 45468 15648 45520 15700
rect 39488 15623 39540 15632
rect 39488 15589 39497 15623
rect 39497 15589 39531 15623
rect 39531 15589 39540 15623
rect 39488 15580 39540 15589
rect 41328 15580 41380 15632
rect 42708 15580 42760 15632
rect 46572 15580 46624 15632
rect 44272 15512 44324 15564
rect 45008 15512 45060 15564
rect 45468 15555 45520 15564
rect 45468 15521 45477 15555
rect 45477 15521 45511 15555
rect 45511 15521 45520 15555
rect 45468 15512 45520 15521
rect 49884 15512 49936 15564
rect 37464 15487 37516 15496
rect 37464 15453 37473 15487
rect 37473 15453 37507 15487
rect 37507 15453 37516 15487
rect 37464 15444 37516 15453
rect 38844 15444 38896 15496
rect 39120 15444 39172 15496
rect 39396 15444 39448 15496
rect 42248 15487 42300 15496
rect 42248 15453 42257 15487
rect 42257 15453 42291 15487
rect 42291 15453 42300 15487
rect 42248 15444 42300 15453
rect 41696 15376 41748 15428
rect 44640 15487 44692 15496
rect 44640 15453 44649 15487
rect 44649 15453 44683 15487
rect 44683 15453 44692 15487
rect 44640 15444 44692 15453
rect 39120 15308 39172 15360
rect 39304 15308 39356 15360
rect 39764 15308 39816 15360
rect 43444 15376 43496 15428
rect 49332 15444 49384 15496
rect 48320 15376 48372 15428
rect 50436 15376 50488 15428
rect 43996 15351 44048 15360
rect 43996 15317 44005 15351
rect 44005 15317 44039 15351
rect 44039 15317 44048 15351
rect 43996 15308 44048 15317
rect 44456 15351 44508 15360
rect 44456 15317 44465 15351
rect 44465 15317 44499 15351
rect 44499 15317 44508 15351
rect 44456 15308 44508 15317
rect 46848 15308 46900 15360
rect 47768 15351 47820 15360
rect 47768 15317 47777 15351
rect 47777 15317 47811 15351
rect 47811 15317 47820 15351
rect 47768 15308 47820 15317
rect 48596 15308 48648 15360
rect 49608 15308 49660 15360
rect 49792 15308 49844 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 7012 15104 7064 15156
rect 7748 15104 7800 15156
rect 9680 15104 9732 15156
rect 3424 15036 3476 15088
rect 6736 15036 6788 15088
rect 7840 15036 7892 15088
rect 9128 15036 9180 15088
rect 10876 15079 10928 15088
rect 10876 15045 10885 15079
rect 10885 15045 10919 15079
rect 10919 15045 10928 15079
rect 10876 15036 10928 15045
rect 1308 14900 1360 14952
rect 6828 14968 6880 15020
rect 7932 14968 7984 15020
rect 8024 15011 8076 15020
rect 8024 14977 8033 15011
rect 8033 14977 8067 15011
rect 8067 14977 8076 15011
rect 8024 14968 8076 14977
rect 8484 14968 8536 15020
rect 11704 14968 11756 15020
rect 6184 14900 6236 14952
rect 9496 14900 9548 14952
rect 9864 14900 9916 14952
rect 10324 14900 10376 14952
rect 7104 14832 7156 14884
rect 7564 14832 7616 14884
rect 7748 14832 7800 14884
rect 7840 14832 7892 14884
rect 12900 15104 12952 15156
rect 13268 15104 13320 15156
rect 14740 15104 14792 15156
rect 16396 15104 16448 15156
rect 18328 15104 18380 15156
rect 18880 15104 18932 15156
rect 19616 15104 19668 15156
rect 19800 15104 19852 15156
rect 21456 15147 21508 15156
rect 21456 15113 21465 15147
rect 21465 15113 21499 15147
rect 21499 15113 21508 15147
rect 21456 15104 21508 15113
rect 21824 15104 21876 15156
rect 22008 15104 22060 15156
rect 23756 15104 23808 15156
rect 25412 15147 25464 15156
rect 25412 15113 25421 15147
rect 25421 15113 25455 15147
rect 25455 15113 25464 15147
rect 25412 15104 25464 15113
rect 27252 15104 27304 15156
rect 14004 15036 14056 15088
rect 12164 14968 12216 15020
rect 12256 14900 12308 14952
rect 12532 14968 12584 15020
rect 13544 15011 13596 15020
rect 13544 14977 13553 15011
rect 13553 14977 13587 15011
rect 13587 14977 13596 15011
rect 13544 14968 13596 14977
rect 6000 14807 6052 14816
rect 6000 14773 6009 14807
rect 6009 14773 6043 14807
rect 6043 14773 6052 14807
rect 6000 14764 6052 14773
rect 8300 14764 8352 14816
rect 9772 14764 9824 14816
rect 9956 14764 10008 14816
rect 13268 14900 13320 14952
rect 12808 14832 12860 14884
rect 13820 14900 13872 14952
rect 16212 15036 16264 15088
rect 16028 14968 16080 15020
rect 16396 15011 16448 15020
rect 16396 14977 16405 15011
rect 16405 14977 16439 15011
rect 16439 14977 16448 15011
rect 16396 14968 16448 14977
rect 16672 14968 16724 15020
rect 17040 14968 17092 15020
rect 17776 15036 17828 15088
rect 19524 15036 19576 15088
rect 14280 14943 14332 14952
rect 14280 14909 14289 14943
rect 14289 14909 14323 14943
rect 14323 14909 14332 14943
rect 14280 14900 14332 14909
rect 15844 14900 15896 14952
rect 16120 14900 16172 14952
rect 18512 14968 18564 15020
rect 18696 14968 18748 15020
rect 20812 15036 20864 15088
rect 22836 15036 22888 15088
rect 19800 14968 19852 15020
rect 20168 14968 20220 15020
rect 20628 15011 20680 15020
rect 20628 14977 20637 15011
rect 20637 14977 20671 15011
rect 20671 14977 20680 15011
rect 20628 14968 20680 14977
rect 21548 14968 21600 15020
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 23572 14968 23624 15020
rect 12624 14764 12676 14816
rect 13544 14764 13596 14816
rect 19524 14943 19576 14952
rect 19524 14909 19533 14943
rect 19533 14909 19567 14943
rect 19567 14909 19576 14943
rect 19524 14900 19576 14909
rect 19892 14900 19944 14952
rect 20720 14943 20772 14952
rect 20720 14909 20729 14943
rect 20729 14909 20763 14943
rect 20763 14909 20772 14943
rect 20720 14900 20772 14909
rect 15660 14764 15712 14816
rect 18696 14764 18748 14816
rect 19064 14807 19116 14816
rect 19064 14773 19073 14807
rect 19073 14773 19107 14807
rect 19107 14773 19116 14807
rect 19064 14764 19116 14773
rect 19708 14832 19760 14884
rect 22468 14900 22520 14952
rect 23112 14900 23164 14952
rect 24032 14968 24084 15020
rect 22192 14832 22244 14884
rect 23204 14764 23256 14816
rect 23480 14807 23532 14816
rect 23480 14773 23489 14807
rect 23489 14773 23523 14807
rect 23523 14773 23532 14807
rect 23480 14764 23532 14773
rect 23756 14900 23808 14952
rect 24676 14943 24728 14952
rect 24676 14909 24685 14943
rect 24685 14909 24719 14943
rect 24719 14909 24728 14943
rect 24676 14900 24728 14909
rect 25872 15036 25924 15088
rect 26976 15036 27028 15088
rect 27988 15104 28040 15156
rect 28448 15104 28500 15156
rect 28724 15147 28776 15156
rect 28724 15113 28733 15147
rect 28733 15113 28767 15147
rect 28767 15113 28776 15147
rect 28724 15104 28776 15113
rect 28816 15147 28868 15156
rect 28816 15113 28825 15147
rect 28825 15113 28859 15147
rect 28859 15113 28868 15147
rect 28816 15104 28868 15113
rect 28908 15104 28960 15156
rect 29828 15104 29880 15156
rect 32220 15104 32272 15156
rect 27804 15036 27856 15088
rect 24860 14900 24912 14952
rect 26240 14900 26292 14952
rect 26424 14943 26476 14952
rect 26424 14909 26433 14943
rect 26433 14909 26467 14943
rect 26467 14909 26476 14943
rect 26424 14900 26476 14909
rect 26608 14943 26660 14952
rect 26608 14909 26617 14943
rect 26617 14909 26651 14943
rect 26651 14909 26660 14943
rect 26608 14900 26660 14909
rect 27160 14900 27212 14952
rect 28264 14968 28316 15020
rect 28724 14968 28776 15020
rect 29092 14968 29144 15020
rect 27896 14900 27948 14952
rect 28724 14832 28776 14884
rect 29276 15036 29328 15088
rect 29736 15036 29788 15088
rect 30656 14968 30708 15020
rect 30840 14968 30892 15020
rect 33232 15104 33284 15156
rect 35348 15147 35400 15156
rect 35348 15113 35357 15147
rect 35357 15113 35391 15147
rect 35391 15113 35400 15147
rect 35348 15104 35400 15113
rect 35992 15104 36044 15156
rect 37372 15104 37424 15156
rect 40868 15104 40920 15156
rect 37832 15036 37884 15088
rect 38752 15036 38804 15088
rect 40776 15036 40828 15088
rect 32496 14968 32548 15020
rect 30380 14900 30432 14952
rect 31392 14943 31444 14952
rect 31392 14909 31401 14943
rect 31401 14909 31435 14943
rect 31435 14909 31444 14943
rect 31392 14900 31444 14909
rect 33416 14968 33468 15020
rect 33692 14968 33744 15020
rect 34888 14968 34940 15020
rect 36452 15011 36504 15020
rect 36452 14977 36461 15011
rect 36461 14977 36495 15011
rect 36495 14977 36504 15011
rect 36452 14968 36504 14977
rect 37096 14968 37148 15020
rect 37464 14968 37516 15020
rect 39948 14968 40000 15020
rect 42800 15036 42852 15088
rect 33508 14900 33560 14952
rect 34336 14900 34388 14952
rect 35532 14943 35584 14952
rect 35532 14909 35541 14943
rect 35541 14909 35575 14943
rect 35575 14909 35584 14943
rect 35532 14900 35584 14909
rect 35624 14900 35676 14952
rect 32220 14832 32272 14884
rect 36360 14832 36412 14884
rect 28448 14764 28500 14816
rect 28540 14764 28592 14816
rect 29092 14764 29144 14816
rect 29368 14764 29420 14816
rect 30656 14764 30708 14816
rect 31576 14764 31628 14816
rect 32864 14764 32916 14816
rect 33232 14764 33284 14816
rect 34336 14764 34388 14816
rect 35900 14764 35952 14816
rect 36268 14764 36320 14816
rect 36820 14900 36872 14952
rect 37556 14900 37608 14952
rect 38292 14943 38344 14952
rect 38292 14909 38301 14943
rect 38301 14909 38335 14943
rect 38335 14909 38344 14943
rect 38292 14900 38344 14909
rect 38384 14900 38436 14952
rect 37832 14764 37884 14816
rect 39304 14832 39356 14884
rect 44824 15104 44876 15156
rect 47676 15104 47728 15156
rect 49240 15147 49292 15156
rect 49240 15113 49249 15147
rect 49249 15113 49283 15147
rect 49283 15113 49292 15147
rect 49240 15104 49292 15113
rect 44364 15036 44416 15088
rect 44640 15036 44692 15088
rect 43996 14968 44048 15020
rect 45652 14968 45704 15020
rect 45928 14968 45980 15020
rect 48688 15036 48740 15088
rect 47676 14968 47728 15020
rect 47860 14968 47912 15020
rect 48596 15011 48648 15020
rect 48596 14977 48605 15011
rect 48605 14977 48639 15011
rect 48639 14977 48648 15011
rect 48596 14968 48648 14977
rect 47032 14900 47084 14952
rect 39764 14807 39816 14816
rect 39764 14773 39773 14807
rect 39773 14773 39807 14807
rect 39807 14773 39816 14807
rect 39764 14764 39816 14773
rect 39856 14764 39908 14816
rect 41972 14764 42024 14816
rect 42064 14807 42116 14816
rect 42064 14773 42073 14807
rect 42073 14773 42107 14807
rect 42107 14773 42116 14807
rect 42064 14764 42116 14773
rect 42432 14764 42484 14816
rect 44180 14764 44232 14816
rect 45192 14764 45244 14816
rect 45468 14764 45520 14816
rect 45652 14764 45704 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 50896 14628 50948 14680
rect 3516 14603 3568 14612
rect 3516 14569 3525 14603
rect 3525 14569 3559 14603
rect 3559 14569 3568 14603
rect 3516 14560 3568 14569
rect 5724 14560 5776 14612
rect 7932 14560 7984 14612
rect 8668 14560 8720 14612
rect 9404 14560 9456 14612
rect 9956 14560 10008 14612
rect 13820 14560 13872 14612
rect 13912 14603 13964 14612
rect 13912 14569 13921 14603
rect 13921 14569 13955 14603
rect 13955 14569 13964 14603
rect 13912 14560 13964 14569
rect 14004 14560 14056 14612
rect 14556 14560 14608 14612
rect 14648 14560 14700 14612
rect 16028 14560 16080 14612
rect 16856 14560 16908 14612
rect 17684 14560 17736 14612
rect 1952 14492 2004 14544
rect 2228 14492 2280 14544
rect 3976 14535 4028 14544
rect 3976 14501 3985 14535
rect 3985 14501 4019 14535
rect 4019 14501 4028 14535
rect 3976 14492 4028 14501
rect 5264 14492 5316 14544
rect 6736 14492 6788 14544
rect 11152 14492 11204 14544
rect 17868 14492 17920 14544
rect 19708 14560 19760 14612
rect 18696 14492 18748 14544
rect 18880 14492 18932 14544
rect 19248 14492 19300 14544
rect 1308 14424 1360 14476
rect 1952 14356 2004 14408
rect 7012 14424 7064 14476
rect 7564 14424 7616 14476
rect 11244 14424 11296 14476
rect 12440 14424 12492 14476
rect 4896 14356 4948 14408
rect 6000 14356 6052 14408
rect 4804 14288 4856 14340
rect 8760 14356 8812 14408
rect 8944 14356 8996 14408
rect 10048 14356 10100 14408
rect 10508 14399 10560 14408
rect 10508 14365 10517 14399
rect 10517 14365 10551 14399
rect 10551 14365 10560 14399
rect 10508 14356 10560 14365
rect 10784 14356 10836 14408
rect 14648 14424 14700 14476
rect 14832 14467 14884 14476
rect 14832 14433 14841 14467
rect 14841 14433 14875 14467
rect 14875 14433 14884 14467
rect 14832 14424 14884 14433
rect 13360 14356 13412 14408
rect 16764 14424 16816 14476
rect 18788 14467 18840 14476
rect 18788 14433 18797 14467
rect 18797 14433 18831 14467
rect 18831 14433 18840 14467
rect 18788 14424 18840 14433
rect 21456 14424 21508 14476
rect 21824 14424 21876 14476
rect 25136 14560 25188 14612
rect 27712 14560 27764 14612
rect 27896 14560 27948 14612
rect 28264 14603 28316 14612
rect 28264 14569 28273 14603
rect 28273 14569 28307 14603
rect 28307 14569 28316 14603
rect 28264 14560 28316 14569
rect 24308 14492 24360 14544
rect 24768 14492 24820 14544
rect 28080 14492 28132 14544
rect 29552 14492 29604 14544
rect 31576 14492 31628 14544
rect 32220 14492 32272 14544
rect 32312 14492 32364 14544
rect 33324 14560 33376 14612
rect 33968 14560 34020 14612
rect 42064 14560 42116 14612
rect 42800 14560 42852 14612
rect 47492 14560 47544 14612
rect 49332 14603 49384 14612
rect 49332 14569 49341 14603
rect 49341 14569 49375 14603
rect 49375 14569 49384 14603
rect 49332 14560 49384 14569
rect 24584 14424 24636 14476
rect 28724 14424 28776 14476
rect 29644 14424 29696 14476
rect 1768 14220 1820 14272
rect 7564 14220 7616 14272
rect 8300 14220 8352 14272
rect 11704 14220 11756 14272
rect 11888 14331 11940 14340
rect 11888 14297 11897 14331
rect 11897 14297 11931 14331
rect 11931 14297 11940 14331
rect 11888 14288 11940 14297
rect 14004 14288 14056 14340
rect 15292 14288 15344 14340
rect 16212 14356 16264 14408
rect 16856 14356 16908 14408
rect 17040 14399 17092 14408
rect 17040 14365 17049 14399
rect 17049 14365 17083 14399
rect 17083 14365 17092 14399
rect 17040 14356 17092 14365
rect 20536 14356 20588 14408
rect 20812 14399 20864 14408
rect 20812 14365 20821 14399
rect 20821 14365 20855 14399
rect 20855 14365 20864 14399
rect 20812 14356 20864 14365
rect 22192 14356 22244 14408
rect 24492 14356 24544 14408
rect 25596 14356 25648 14408
rect 25780 14356 25832 14408
rect 25964 14399 26016 14408
rect 25964 14365 25973 14399
rect 25973 14365 26007 14399
rect 26007 14365 26016 14399
rect 25964 14356 26016 14365
rect 27344 14356 27396 14408
rect 29368 14356 29420 14408
rect 30104 14424 30156 14476
rect 30656 14424 30708 14476
rect 38384 14492 38436 14544
rect 32588 14467 32640 14476
rect 32588 14433 32597 14467
rect 32597 14433 32631 14467
rect 32631 14433 32640 14467
rect 32588 14424 32640 14433
rect 32772 14424 32824 14476
rect 35716 14424 35768 14476
rect 33784 14356 33836 14408
rect 34060 14356 34112 14408
rect 13636 14220 13688 14272
rect 13912 14220 13964 14272
rect 14648 14263 14700 14272
rect 14648 14229 14657 14263
rect 14657 14229 14691 14263
rect 14691 14229 14700 14263
rect 14648 14220 14700 14229
rect 15476 14263 15528 14272
rect 15476 14229 15485 14263
rect 15485 14229 15519 14263
rect 15519 14229 15528 14263
rect 15476 14220 15528 14229
rect 16764 14288 16816 14340
rect 17684 14288 17736 14340
rect 21088 14331 21140 14340
rect 21088 14297 21097 14331
rect 21097 14297 21131 14331
rect 21131 14297 21140 14331
rect 21088 14288 21140 14297
rect 25228 14288 25280 14340
rect 29552 14288 29604 14340
rect 30012 14331 30064 14340
rect 30012 14297 30021 14331
rect 30021 14297 30055 14331
rect 30055 14297 30064 14331
rect 30012 14288 30064 14297
rect 15752 14220 15804 14272
rect 17592 14220 17644 14272
rect 18420 14220 18472 14272
rect 18880 14220 18932 14272
rect 19524 14220 19576 14272
rect 19984 14263 20036 14272
rect 19984 14229 19993 14263
rect 19993 14229 20027 14263
rect 20027 14229 20036 14263
rect 19984 14220 20036 14229
rect 22560 14220 22612 14272
rect 25780 14220 25832 14272
rect 26516 14220 26568 14272
rect 27712 14263 27764 14272
rect 27712 14229 27721 14263
rect 27721 14229 27755 14263
rect 27755 14229 27764 14263
rect 27712 14220 27764 14229
rect 28264 14220 28316 14272
rect 28908 14263 28960 14272
rect 28908 14229 28917 14263
rect 28917 14229 28951 14263
rect 28951 14229 28960 14263
rect 28908 14220 28960 14229
rect 30748 14220 30800 14272
rect 31484 14288 31536 14340
rect 32680 14288 32732 14340
rect 34796 14288 34848 14340
rect 35624 14288 35676 14340
rect 34336 14220 34388 14272
rect 34612 14220 34664 14272
rect 36820 14424 36872 14476
rect 37464 14424 37516 14476
rect 39212 14492 39264 14544
rect 39304 14535 39356 14544
rect 39304 14501 39313 14535
rect 39313 14501 39347 14535
rect 39347 14501 39356 14535
rect 39304 14492 39356 14501
rect 39396 14492 39448 14544
rect 39856 14492 39908 14544
rect 40224 14492 40276 14544
rect 44088 14492 44140 14544
rect 39764 14424 39816 14476
rect 37372 14331 37424 14340
rect 37372 14297 37381 14331
rect 37381 14297 37415 14331
rect 37415 14297 37424 14331
rect 37372 14288 37424 14297
rect 38844 14356 38896 14408
rect 38936 14356 38988 14408
rect 43168 14424 43220 14476
rect 41512 14356 41564 14408
rect 43260 14356 43312 14408
rect 39120 14288 39172 14340
rect 39212 14288 39264 14340
rect 39856 14288 39908 14340
rect 40132 14288 40184 14340
rect 38936 14220 38988 14272
rect 41972 14220 42024 14272
rect 44364 14356 44416 14408
rect 45376 14356 45428 14408
rect 47308 14356 47360 14408
rect 47768 14356 47820 14408
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 3608 14059 3660 14068
rect 3608 14025 3617 14059
rect 3617 14025 3651 14059
rect 3651 14025 3660 14059
rect 3608 14016 3660 14025
rect 4896 14059 4948 14068
rect 4896 14025 4905 14059
rect 4905 14025 4939 14059
rect 4939 14025 4948 14059
rect 4896 14016 4948 14025
rect 6000 14059 6052 14068
rect 6000 14025 6009 14059
rect 6009 14025 6043 14059
rect 6043 14025 6052 14059
rect 6000 14016 6052 14025
rect 6368 14016 6420 14068
rect 6828 14016 6880 14068
rect 10048 14059 10100 14068
rect 10048 14025 10057 14059
rect 10057 14025 10091 14059
rect 10091 14025 10100 14059
rect 10048 14016 10100 14025
rect 10508 14016 10560 14068
rect 13728 14016 13780 14068
rect 14464 14059 14516 14068
rect 14464 14025 14473 14059
rect 14473 14025 14507 14059
rect 14507 14025 14516 14059
rect 14464 14016 14516 14025
rect 14556 14016 14608 14068
rect 15476 14016 15528 14068
rect 15660 14059 15712 14068
rect 15660 14025 15669 14059
rect 15669 14025 15703 14059
rect 15703 14025 15712 14059
rect 15660 14016 15712 14025
rect 15936 14016 15988 14068
rect 16212 14059 16264 14068
rect 16212 14025 16221 14059
rect 16221 14025 16255 14059
rect 16255 14025 16264 14059
rect 16212 14016 16264 14025
rect 16396 14016 16448 14068
rect 19064 14016 19116 14068
rect 5908 13948 5960 14000
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 2780 13880 2832 13932
rect 2872 13880 2924 13932
rect 3608 13880 3660 13932
rect 4068 13880 4120 13932
rect 940 13812 992 13864
rect 6000 13812 6052 13864
rect 6644 13880 6696 13932
rect 9956 13948 10008 14000
rect 12440 13948 12492 14000
rect 15752 13948 15804 14000
rect 16304 13948 16356 14000
rect 18328 13991 18380 14000
rect 18328 13957 18337 13991
rect 18337 13957 18371 13991
rect 18371 13957 18380 13991
rect 18328 13948 18380 13957
rect 20812 14016 20864 14068
rect 21456 14059 21508 14068
rect 21456 14025 21465 14059
rect 21465 14025 21499 14059
rect 21499 14025 21508 14059
rect 21456 14016 21508 14025
rect 22008 14059 22060 14068
rect 22008 14025 22017 14059
rect 22017 14025 22051 14059
rect 22051 14025 22060 14059
rect 22008 14016 22060 14025
rect 22836 14016 22888 14068
rect 23664 14016 23716 14068
rect 7840 13812 7892 13864
rect 11244 13880 11296 13932
rect 11704 13923 11756 13932
rect 11704 13889 11713 13923
rect 11713 13889 11747 13923
rect 11747 13889 11756 13923
rect 11704 13880 11756 13889
rect 13544 13880 13596 13932
rect 15200 13880 15252 13932
rect 15660 13880 15712 13932
rect 17132 13880 17184 13932
rect 18512 13880 18564 13932
rect 22192 13948 22244 14000
rect 22744 13948 22796 14000
rect 12808 13812 12860 13864
rect 9220 13744 9272 13796
rect 9312 13744 9364 13796
rect 6552 13676 6604 13728
rect 6828 13676 6880 13728
rect 7564 13676 7616 13728
rect 9864 13676 9916 13728
rect 12164 13676 12216 13728
rect 12348 13676 12400 13728
rect 12716 13676 12768 13728
rect 12808 13719 12860 13728
rect 12808 13685 12817 13719
rect 12817 13685 12851 13719
rect 12851 13685 12860 13719
rect 12808 13676 12860 13685
rect 13544 13744 13596 13796
rect 15016 13812 15068 13864
rect 17040 13812 17092 13864
rect 19524 13812 19576 13864
rect 22100 13880 22152 13932
rect 14464 13676 14516 13728
rect 17868 13744 17920 13796
rect 22100 13744 22152 13796
rect 22652 13880 22704 13932
rect 24492 13948 24544 14000
rect 25964 14016 26016 14068
rect 26516 14016 26568 14068
rect 24676 13880 24728 13932
rect 27344 13948 27396 14000
rect 31760 14016 31812 14068
rect 32772 14059 32824 14068
rect 32772 14025 32781 14059
rect 32781 14025 32815 14059
rect 32815 14025 32824 14059
rect 32772 14016 32824 14025
rect 33508 14016 33560 14068
rect 27160 13923 27212 13932
rect 27160 13889 27169 13923
rect 27169 13889 27203 13923
rect 27203 13889 27212 13923
rect 27160 13880 27212 13889
rect 31300 13948 31352 14000
rect 32680 13948 32732 14000
rect 35348 14059 35400 14068
rect 35348 14025 35357 14059
rect 35357 14025 35391 14059
rect 35391 14025 35400 14059
rect 35348 14016 35400 14025
rect 35992 13991 36044 14000
rect 35992 13957 36001 13991
rect 36001 13957 36035 13991
rect 36035 13957 36044 13991
rect 35992 13948 36044 13957
rect 36820 13991 36872 14000
rect 36820 13957 36829 13991
rect 36829 13957 36863 13991
rect 36863 13957 36872 13991
rect 36820 13948 36872 13957
rect 38476 14016 38528 14068
rect 41512 14016 41564 14068
rect 43260 14059 43312 14068
rect 43260 14025 43269 14059
rect 43269 14025 43303 14059
rect 43303 14025 43312 14059
rect 43260 14016 43312 14025
rect 44364 14059 44416 14068
rect 44364 14025 44373 14059
rect 44373 14025 44407 14059
rect 44407 14025 44416 14059
rect 44364 14016 44416 14025
rect 44548 14016 44600 14068
rect 45560 14016 45612 14068
rect 45744 14016 45796 14068
rect 47032 14016 47084 14068
rect 47400 14016 47452 14068
rect 47768 14016 47820 14068
rect 48320 14016 48372 14068
rect 29368 13923 29420 13932
rect 29368 13889 29377 13923
rect 29377 13889 29411 13923
rect 29411 13889 29420 13923
rect 29368 13880 29420 13889
rect 30748 13880 30800 13932
rect 31024 13880 31076 13932
rect 22652 13744 22704 13796
rect 24124 13744 24176 13796
rect 29736 13812 29788 13864
rect 30196 13812 30248 13864
rect 31668 13812 31720 13864
rect 33140 13923 33192 13932
rect 33140 13889 33149 13923
rect 33149 13889 33183 13923
rect 33183 13889 33192 13923
rect 33140 13880 33192 13889
rect 36176 13880 36228 13932
rect 34704 13812 34756 13864
rect 35900 13812 35952 13864
rect 37096 13812 37148 13864
rect 16580 13676 16632 13728
rect 19248 13719 19300 13728
rect 19248 13685 19257 13719
rect 19257 13685 19291 13719
rect 19291 13685 19300 13719
rect 19248 13676 19300 13685
rect 21364 13676 21416 13728
rect 22376 13676 22428 13728
rect 22836 13676 22888 13728
rect 23480 13676 23532 13728
rect 24952 13676 25004 13728
rect 32864 13744 32916 13796
rect 35348 13744 35400 13796
rect 39764 13880 39816 13932
rect 39856 13923 39908 13932
rect 39856 13889 39865 13923
rect 39865 13889 39899 13923
rect 39899 13889 39908 13923
rect 39856 13880 39908 13889
rect 39948 13880 40000 13932
rect 43352 13948 43404 14000
rect 43904 13948 43956 14000
rect 37280 13744 37332 13796
rect 38016 13744 38068 13796
rect 38292 13812 38344 13864
rect 38200 13744 38252 13796
rect 40500 13855 40552 13864
rect 40500 13821 40509 13855
rect 40509 13821 40543 13855
rect 40543 13821 40552 13855
rect 40500 13812 40552 13821
rect 42708 13880 42760 13932
rect 45284 13880 45336 13932
rect 41696 13812 41748 13864
rect 44640 13812 44692 13864
rect 42616 13744 42668 13796
rect 34428 13676 34480 13728
rect 34612 13676 34664 13728
rect 38292 13676 38344 13728
rect 38568 13676 38620 13728
rect 40592 13676 40644 13728
rect 42524 13676 42576 13728
rect 50620 13948 50672 14000
rect 46296 13923 46348 13932
rect 46296 13889 46305 13923
rect 46305 13889 46339 13923
rect 46339 13889 46348 13923
rect 46296 13880 46348 13889
rect 46388 13880 46440 13932
rect 47860 13880 47912 13932
rect 48596 13880 48648 13932
rect 49148 13880 49200 13932
rect 47492 13676 47544 13728
rect 47768 13676 47820 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 3424 13515 3476 13524
rect 3424 13481 3433 13515
rect 3433 13481 3467 13515
rect 3467 13481 3476 13515
rect 3424 13472 3476 13481
rect 7472 13515 7524 13524
rect 7472 13481 7481 13515
rect 7481 13481 7515 13515
rect 7515 13481 7524 13515
rect 7472 13472 7524 13481
rect 11888 13472 11940 13524
rect 12440 13472 12492 13524
rect 12716 13472 12768 13524
rect 16028 13472 16080 13524
rect 17868 13515 17920 13524
rect 17868 13481 17877 13515
rect 17877 13481 17911 13515
rect 17911 13481 17920 13515
rect 17868 13472 17920 13481
rect 18328 13515 18380 13524
rect 18328 13481 18337 13515
rect 18337 13481 18371 13515
rect 18371 13481 18380 13515
rect 18328 13472 18380 13481
rect 18788 13472 18840 13524
rect 19524 13472 19576 13524
rect 19984 13472 20036 13524
rect 2136 13404 2188 13456
rect 4528 13404 4580 13456
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 2780 13336 2832 13345
rect 3976 13243 4028 13252
rect 3976 13209 3985 13243
rect 3985 13209 4019 13243
rect 4019 13209 4028 13243
rect 3976 13200 4028 13209
rect 5080 13268 5132 13320
rect 8484 13404 8536 13456
rect 8760 13404 8812 13456
rect 9128 13404 9180 13456
rect 9956 13447 10008 13456
rect 9956 13413 9965 13447
rect 9965 13413 9999 13447
rect 9999 13413 10008 13447
rect 9956 13404 10008 13413
rect 13084 13404 13136 13456
rect 13452 13404 13504 13456
rect 15384 13404 15436 13456
rect 20168 13404 20220 13456
rect 9588 13336 9640 13388
rect 10324 13336 10376 13388
rect 10784 13336 10836 13388
rect 11152 13336 11204 13388
rect 11888 13336 11940 13388
rect 12440 13336 12492 13388
rect 12992 13336 13044 13388
rect 13176 13379 13228 13388
rect 13176 13345 13185 13379
rect 13185 13345 13219 13379
rect 13219 13345 13228 13379
rect 13176 13336 13228 13345
rect 13544 13336 13596 13388
rect 7840 13268 7892 13320
rect 8852 13268 8904 13320
rect 9864 13268 9916 13320
rect 12072 13268 12124 13320
rect 6460 13200 6512 13252
rect 11704 13200 11756 13252
rect 18696 13379 18748 13388
rect 18696 13345 18705 13379
rect 18705 13345 18739 13379
rect 18739 13345 18748 13379
rect 18696 13336 18748 13345
rect 18880 13379 18932 13388
rect 18880 13345 18889 13379
rect 18889 13345 18923 13379
rect 18923 13345 18932 13379
rect 18880 13336 18932 13345
rect 20076 13336 20128 13388
rect 21640 13472 21692 13524
rect 24584 13472 24636 13524
rect 27160 13472 27212 13524
rect 30104 13515 30156 13524
rect 30104 13481 30113 13515
rect 30113 13481 30147 13515
rect 30147 13481 30156 13515
rect 30104 13472 30156 13481
rect 14280 13268 14332 13320
rect 19616 13268 19668 13320
rect 20812 13336 20864 13388
rect 21548 13336 21600 13388
rect 21640 13336 21692 13388
rect 23020 13379 23072 13388
rect 23020 13345 23029 13379
rect 23029 13345 23063 13379
rect 23063 13345 23072 13379
rect 23020 13336 23072 13345
rect 23480 13268 23532 13320
rect 6092 13132 6144 13184
rect 8484 13132 8536 13184
rect 10600 13132 10652 13184
rect 14372 13243 14424 13252
rect 14372 13209 14381 13243
rect 14381 13209 14415 13243
rect 14415 13209 14424 13243
rect 14372 13200 14424 13209
rect 14832 13200 14884 13252
rect 16488 13200 16540 13252
rect 18696 13200 18748 13252
rect 18880 13200 18932 13252
rect 19800 13200 19852 13252
rect 20904 13200 20956 13252
rect 21180 13243 21232 13252
rect 21180 13209 21189 13243
rect 21189 13209 21223 13243
rect 21223 13209 21232 13243
rect 21180 13200 21232 13209
rect 24492 13336 24544 13388
rect 25964 13404 26016 13456
rect 26792 13336 26844 13388
rect 28908 13404 28960 13456
rect 29368 13336 29420 13388
rect 29552 13447 29604 13456
rect 29552 13413 29561 13447
rect 29561 13413 29595 13447
rect 29595 13413 29604 13447
rect 29552 13404 29604 13413
rect 29644 13404 29696 13456
rect 32588 13472 32640 13524
rect 33324 13472 33376 13524
rect 34060 13472 34112 13524
rect 34888 13515 34940 13524
rect 34888 13481 34897 13515
rect 34897 13481 34931 13515
rect 34931 13481 34940 13515
rect 34888 13472 34940 13481
rect 30380 13447 30432 13456
rect 30380 13413 30389 13447
rect 30389 13413 30423 13447
rect 30423 13413 30432 13447
rect 30380 13404 30432 13413
rect 32680 13404 32732 13456
rect 36360 13404 36412 13456
rect 38200 13515 38252 13524
rect 38200 13481 38209 13515
rect 38209 13481 38243 13515
rect 38243 13481 38252 13515
rect 38200 13472 38252 13481
rect 39672 13515 39724 13524
rect 39672 13481 39681 13515
rect 39681 13481 39715 13515
rect 39715 13481 39724 13515
rect 39672 13472 39724 13481
rect 39856 13472 39908 13524
rect 42800 13472 42852 13524
rect 45008 13515 45060 13524
rect 45008 13481 45017 13515
rect 45017 13481 45051 13515
rect 45051 13481 45060 13515
rect 45008 13472 45060 13481
rect 48412 13472 48464 13524
rect 33508 13336 33560 13388
rect 33692 13336 33744 13388
rect 34244 13336 34296 13388
rect 34428 13336 34480 13388
rect 35624 13336 35676 13388
rect 36176 13336 36228 13388
rect 36820 13336 36872 13388
rect 37280 13336 37332 13388
rect 38476 13336 38528 13388
rect 43812 13404 43864 13456
rect 28448 13268 28500 13320
rect 32312 13268 32364 13320
rect 34060 13268 34112 13320
rect 35164 13268 35216 13320
rect 38936 13268 38988 13320
rect 12164 13175 12216 13184
rect 12164 13141 12173 13175
rect 12173 13141 12207 13175
rect 12207 13141 12216 13175
rect 12164 13132 12216 13141
rect 12348 13132 12400 13184
rect 12716 13175 12768 13184
rect 12716 13141 12725 13175
rect 12725 13141 12759 13175
rect 12759 13141 12768 13175
rect 12716 13132 12768 13141
rect 13176 13132 13228 13184
rect 14096 13132 14148 13184
rect 15200 13132 15252 13184
rect 19432 13132 19484 13184
rect 20168 13175 20220 13184
rect 20168 13141 20177 13175
rect 20177 13141 20211 13175
rect 20211 13141 20220 13175
rect 20168 13132 20220 13141
rect 20260 13132 20312 13184
rect 21272 13132 21324 13184
rect 21364 13132 21416 13184
rect 23296 13175 23348 13184
rect 23296 13141 23305 13175
rect 23305 13141 23339 13175
rect 23339 13141 23348 13175
rect 23296 13132 23348 13141
rect 23664 13175 23716 13184
rect 23664 13141 23673 13175
rect 23673 13141 23707 13175
rect 23707 13141 23716 13175
rect 23664 13132 23716 13141
rect 24768 13200 24820 13252
rect 24308 13132 24360 13184
rect 24952 13200 25004 13252
rect 27436 13200 27488 13252
rect 28540 13200 28592 13252
rect 29000 13200 29052 13252
rect 29460 13200 29512 13252
rect 31024 13243 31076 13252
rect 31024 13209 31033 13243
rect 31033 13209 31067 13243
rect 31067 13209 31076 13243
rect 31024 13200 31076 13209
rect 31484 13200 31536 13252
rect 32772 13200 32824 13252
rect 34520 13200 34572 13252
rect 35440 13200 35492 13252
rect 39672 13268 39724 13320
rect 40040 13311 40092 13320
rect 40040 13277 40049 13311
rect 40049 13277 40083 13311
rect 40083 13277 40092 13311
rect 40040 13268 40092 13277
rect 41696 13268 41748 13320
rect 44180 13336 44232 13388
rect 44916 13404 44968 13456
rect 44548 13336 44600 13388
rect 43260 13268 43312 13320
rect 44916 13268 44968 13320
rect 46940 13404 46992 13456
rect 47492 13447 47544 13456
rect 47492 13413 47501 13447
rect 47501 13413 47535 13447
rect 47535 13413 47544 13447
rect 47492 13404 47544 13413
rect 48320 13336 48372 13388
rect 48412 13336 48464 13388
rect 48688 13336 48740 13388
rect 46940 13268 46992 13320
rect 49148 13311 49200 13320
rect 49148 13277 49157 13311
rect 49157 13277 49191 13311
rect 49191 13277 49200 13311
rect 49148 13268 49200 13277
rect 25688 13132 25740 13184
rect 28816 13132 28868 13184
rect 29828 13175 29880 13184
rect 29828 13141 29837 13175
rect 29837 13141 29871 13175
rect 29871 13141 29880 13175
rect 29828 13132 29880 13141
rect 30288 13132 30340 13184
rect 32680 13132 32732 13184
rect 36176 13132 36228 13184
rect 40316 13200 40368 13252
rect 41420 13200 41472 13252
rect 39304 13175 39356 13184
rect 39304 13141 39313 13175
rect 39313 13141 39347 13175
rect 39347 13141 39356 13175
rect 39304 13132 39356 13141
rect 39948 13132 40000 13184
rect 43720 13132 43772 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 3884 12928 3936 12980
rect 4988 12928 5040 12980
rect 6000 12971 6052 12980
rect 6000 12937 6009 12971
rect 6009 12937 6043 12971
rect 6043 12937 6052 12971
rect 6000 12928 6052 12937
rect 6368 12928 6420 12980
rect 6828 12971 6880 12980
rect 6828 12937 6837 12971
rect 6837 12937 6871 12971
rect 6871 12937 6880 12971
rect 6828 12928 6880 12937
rect 8852 12971 8904 12980
rect 8852 12937 8861 12971
rect 8861 12937 8895 12971
rect 8895 12937 8904 12971
rect 8852 12928 8904 12937
rect 9772 12928 9824 12980
rect 3056 12860 3108 12912
rect 4620 12860 4672 12912
rect 11152 12860 11204 12912
rect 13452 12971 13504 12980
rect 13452 12937 13461 12971
rect 13461 12937 13495 12971
rect 13495 12937 13504 12971
rect 13452 12928 13504 12937
rect 13820 12928 13872 12980
rect 15108 12928 15160 12980
rect 15844 12928 15896 12980
rect 16764 12928 16816 12980
rect 18880 12928 18932 12980
rect 19432 12928 19484 12980
rect 20352 12928 20404 12980
rect 13084 12860 13136 12912
rect 18696 12903 18748 12912
rect 1308 12792 1360 12844
rect 2044 12792 2096 12844
rect 2780 12724 2832 12776
rect 4804 12724 4856 12776
rect 5540 12792 5592 12844
rect 7104 12835 7156 12844
rect 7104 12801 7113 12835
rect 7113 12801 7147 12835
rect 7147 12801 7156 12835
rect 7104 12792 7156 12801
rect 6460 12724 6512 12776
rect 6736 12724 6788 12776
rect 9312 12835 9364 12844
rect 9312 12801 9321 12835
rect 9321 12801 9355 12835
rect 9355 12801 9364 12835
rect 9312 12792 9364 12801
rect 9680 12724 9732 12776
rect 10232 12724 10284 12776
rect 10968 12767 11020 12776
rect 10968 12733 10977 12767
rect 10977 12733 11011 12767
rect 11011 12733 11020 12767
rect 10968 12724 11020 12733
rect 11888 12724 11940 12776
rect 12164 12767 12216 12776
rect 12164 12733 12173 12767
rect 12173 12733 12207 12767
rect 12207 12733 12216 12767
rect 12164 12724 12216 12733
rect 5816 12588 5868 12640
rect 6184 12588 6236 12640
rect 7104 12588 7156 12640
rect 7748 12588 7800 12640
rect 11612 12656 11664 12708
rect 12072 12656 12124 12708
rect 12348 12767 12400 12776
rect 12348 12733 12357 12767
rect 12357 12733 12391 12767
rect 12391 12733 12400 12767
rect 12348 12724 12400 12733
rect 12992 12792 13044 12844
rect 13452 12792 13504 12844
rect 14280 12792 14332 12844
rect 16120 12792 16172 12844
rect 13728 12724 13780 12776
rect 15844 12724 15896 12776
rect 18696 12869 18705 12903
rect 18705 12869 18739 12903
rect 18739 12869 18748 12903
rect 18696 12860 18748 12869
rect 19248 12860 19300 12912
rect 22192 12903 22244 12912
rect 22192 12869 22201 12903
rect 22201 12869 22235 12903
rect 22235 12869 22244 12903
rect 22192 12860 22244 12869
rect 23020 12860 23072 12912
rect 23480 12860 23532 12912
rect 24400 12928 24452 12980
rect 24676 12928 24728 12980
rect 26148 12928 26200 12980
rect 17500 12792 17552 12844
rect 17684 12792 17736 12844
rect 19432 12792 19484 12844
rect 19524 12792 19576 12844
rect 22008 12792 22060 12844
rect 23572 12792 23624 12844
rect 28356 12860 28408 12912
rect 28540 12860 28592 12912
rect 29276 12928 29328 12980
rect 30472 12928 30524 12980
rect 31300 12860 31352 12912
rect 31760 12860 31812 12912
rect 25412 12792 25464 12844
rect 13636 12656 13688 12708
rect 16028 12656 16080 12708
rect 19064 12724 19116 12776
rect 20536 12724 20588 12776
rect 9588 12588 9640 12640
rect 9956 12631 10008 12640
rect 9956 12597 9965 12631
rect 9965 12597 9999 12631
rect 9999 12597 10008 12631
rect 9956 12588 10008 12597
rect 10416 12631 10468 12640
rect 10416 12597 10425 12631
rect 10425 12597 10459 12631
rect 10459 12597 10468 12631
rect 10416 12588 10468 12597
rect 11520 12588 11572 12640
rect 13452 12588 13504 12640
rect 17684 12588 17736 12640
rect 18880 12588 18932 12640
rect 19340 12699 19392 12708
rect 19340 12665 19349 12699
rect 19349 12665 19383 12699
rect 19383 12665 19392 12699
rect 19340 12656 19392 12665
rect 20444 12699 20496 12708
rect 20444 12665 20453 12699
rect 20453 12665 20487 12699
rect 20487 12665 20496 12699
rect 20444 12656 20496 12665
rect 21088 12656 21140 12708
rect 20812 12588 20864 12640
rect 21364 12767 21416 12776
rect 21364 12733 21373 12767
rect 21373 12733 21407 12767
rect 21407 12733 21416 12767
rect 21364 12724 21416 12733
rect 22744 12724 22796 12776
rect 26516 12792 26568 12844
rect 26240 12767 26292 12776
rect 26240 12733 26249 12767
rect 26249 12733 26283 12767
rect 26283 12733 26292 12767
rect 26240 12724 26292 12733
rect 26332 12724 26384 12776
rect 27620 12724 27672 12776
rect 32220 12792 32272 12844
rect 32312 12835 32364 12844
rect 32312 12801 32321 12835
rect 32321 12801 32355 12835
rect 32355 12801 32364 12835
rect 32312 12792 32364 12801
rect 37832 12928 37884 12980
rect 35072 12860 35124 12912
rect 35992 12860 36044 12912
rect 36912 12860 36964 12912
rect 38752 12860 38804 12912
rect 36820 12792 36872 12844
rect 40592 12971 40644 12980
rect 40592 12937 40601 12971
rect 40601 12937 40635 12971
rect 40635 12937 40644 12971
rect 40592 12928 40644 12937
rect 41696 12971 41748 12980
rect 41696 12937 41705 12971
rect 41705 12937 41739 12971
rect 41739 12937 41748 12971
rect 41696 12928 41748 12937
rect 43260 12971 43312 12980
rect 43260 12937 43269 12971
rect 43269 12937 43303 12971
rect 43303 12937 43312 12971
rect 43260 12928 43312 12937
rect 44916 12971 44968 12980
rect 44916 12937 44925 12971
rect 44925 12937 44959 12971
rect 44959 12937 44968 12971
rect 44916 12928 44968 12937
rect 46940 12928 46992 12980
rect 47032 12928 47084 12980
rect 40040 12860 40092 12912
rect 22376 12656 22428 12708
rect 23756 12656 23808 12708
rect 25320 12656 25372 12708
rect 26884 12656 26936 12708
rect 22192 12588 22244 12640
rect 25688 12588 25740 12640
rect 30472 12724 30524 12776
rect 31300 12767 31352 12776
rect 31300 12733 31309 12767
rect 31309 12733 31343 12767
rect 31343 12733 31352 12767
rect 31300 12724 31352 12733
rect 34244 12724 34296 12776
rect 34612 12724 34664 12776
rect 35256 12724 35308 12776
rect 35716 12724 35768 12776
rect 36728 12724 36780 12776
rect 37372 12656 37424 12708
rect 29920 12588 29972 12640
rect 30840 12588 30892 12640
rect 33324 12588 33376 12640
rect 35348 12588 35400 12640
rect 36544 12588 36596 12640
rect 39580 12724 39632 12776
rect 39948 12835 40000 12844
rect 39948 12801 39957 12835
rect 39957 12801 39991 12835
rect 39991 12801 40000 12835
rect 39948 12792 40000 12801
rect 41144 12792 41196 12844
rect 44732 12860 44784 12912
rect 45560 12860 45612 12912
rect 46756 12860 46808 12912
rect 42616 12835 42668 12844
rect 42616 12801 42625 12835
rect 42625 12801 42659 12835
rect 42659 12801 42668 12835
rect 42616 12792 42668 12801
rect 43720 12835 43772 12844
rect 43720 12801 43729 12835
rect 43729 12801 43763 12835
rect 43763 12801 43772 12835
rect 43720 12792 43772 12801
rect 41880 12724 41932 12776
rect 45376 12792 45428 12844
rect 46572 12835 46624 12844
rect 46572 12801 46581 12835
rect 46581 12801 46615 12835
rect 46615 12801 46624 12835
rect 46572 12792 46624 12801
rect 44732 12656 44784 12708
rect 45192 12656 45244 12708
rect 47676 12792 47728 12844
rect 49148 12835 49200 12844
rect 49148 12801 49157 12835
rect 49157 12801 49191 12835
rect 49191 12801 49200 12835
rect 49148 12792 49200 12801
rect 37832 12588 37884 12640
rect 39580 12588 39632 12640
rect 41144 12588 41196 12640
rect 44640 12631 44692 12640
rect 44640 12597 44649 12631
rect 44649 12597 44683 12631
rect 44683 12597 44692 12631
rect 44640 12588 44692 12597
rect 47676 12588 47728 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 2320 12427 2372 12436
rect 2320 12393 2329 12427
rect 2329 12393 2363 12427
rect 2363 12393 2372 12427
rect 2320 12384 2372 12393
rect 2780 12427 2832 12436
rect 2780 12393 2789 12427
rect 2789 12393 2823 12427
rect 2823 12393 2832 12427
rect 2780 12384 2832 12393
rect 6368 12427 6420 12436
rect 6368 12393 6377 12427
rect 6377 12393 6411 12427
rect 6411 12393 6420 12427
rect 6368 12384 6420 12393
rect 7656 12384 7708 12436
rect 9864 12427 9916 12436
rect 9864 12393 9873 12427
rect 9873 12393 9907 12427
rect 9907 12393 9916 12427
rect 9864 12384 9916 12393
rect 10048 12384 10100 12436
rect 10968 12384 11020 12436
rect 11888 12384 11940 12436
rect 11980 12384 12032 12436
rect 9680 12316 9732 12368
rect 11612 12316 11664 12368
rect 12072 12316 12124 12368
rect 13084 12316 13136 12368
rect 14648 12384 14700 12436
rect 14740 12384 14792 12436
rect 18604 12384 18656 12436
rect 20168 12384 20220 12436
rect 20444 12384 20496 12436
rect 23940 12384 23992 12436
rect 3424 12291 3476 12300
rect 3424 12257 3433 12291
rect 3433 12257 3467 12291
rect 3467 12257 3476 12291
rect 3424 12248 3476 12257
rect 6368 12248 6420 12300
rect 7196 12248 7248 12300
rect 7472 12248 7524 12300
rect 7564 12248 7616 12300
rect 3700 12180 3752 12232
rect 3884 12180 3936 12232
rect 4068 12180 4120 12232
rect 4620 12223 4672 12232
rect 4620 12189 4629 12223
rect 4629 12189 4663 12223
rect 4663 12189 4672 12223
rect 4620 12180 4672 12189
rect 7840 12180 7892 12232
rect 10324 12291 10376 12300
rect 10324 12257 10333 12291
rect 10333 12257 10367 12291
rect 10367 12257 10376 12291
rect 10324 12248 10376 12257
rect 12992 12248 13044 12300
rect 14004 12316 14056 12368
rect 16120 12316 16172 12368
rect 17040 12316 17092 12368
rect 18696 12316 18748 12368
rect 13544 12291 13596 12300
rect 13544 12257 13553 12291
rect 13553 12257 13587 12291
rect 13587 12257 13596 12291
rect 13544 12248 13596 12257
rect 14556 12248 14608 12300
rect 15292 12248 15344 12300
rect 14280 12223 14332 12232
rect 8852 12112 8904 12164
rect 4068 12044 4120 12096
rect 4620 12044 4672 12096
rect 7564 12044 7616 12096
rect 8576 12087 8628 12096
rect 8576 12053 8585 12087
rect 8585 12053 8619 12087
rect 8619 12053 8628 12087
rect 8576 12044 8628 12053
rect 10600 12155 10652 12164
rect 10600 12121 10609 12155
rect 10609 12121 10643 12155
rect 10643 12121 10652 12155
rect 10600 12112 10652 12121
rect 12348 12112 12400 12164
rect 12992 12112 13044 12164
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 16856 12248 16908 12300
rect 18420 12248 18472 12300
rect 18788 12248 18840 12300
rect 20260 12248 20312 12300
rect 23480 12248 23532 12300
rect 27068 12384 27120 12436
rect 24400 12248 24452 12300
rect 29000 12384 29052 12436
rect 30288 12384 30340 12436
rect 27804 12316 27856 12368
rect 30564 12316 30616 12368
rect 42156 12384 42208 12436
rect 42432 12384 42484 12436
rect 45376 12384 45428 12436
rect 37188 12316 37240 12368
rect 15844 12180 15896 12232
rect 16488 12180 16540 12232
rect 20076 12180 20128 12232
rect 22284 12223 22336 12232
rect 22284 12189 22293 12223
rect 22293 12189 22327 12223
rect 22327 12189 22336 12223
rect 22284 12180 22336 12189
rect 23940 12180 23992 12232
rect 24584 12223 24636 12232
rect 24584 12189 24593 12223
rect 24593 12189 24627 12223
rect 24627 12189 24636 12223
rect 24584 12180 24636 12189
rect 27620 12248 27672 12300
rect 28080 12248 28132 12300
rect 28816 12248 28868 12300
rect 29460 12248 29512 12300
rect 30196 12248 30248 12300
rect 29552 12180 29604 12232
rect 29644 12180 29696 12232
rect 30380 12180 30432 12232
rect 32312 12248 32364 12300
rect 34612 12248 34664 12300
rect 33508 12180 33560 12232
rect 35716 12248 35768 12300
rect 35808 12248 35860 12300
rect 37556 12248 37608 12300
rect 38568 12248 38620 12300
rect 36452 12180 36504 12232
rect 13912 12112 13964 12164
rect 14004 12112 14056 12164
rect 10968 12044 11020 12096
rect 11888 12044 11940 12096
rect 16304 12112 16356 12164
rect 18328 12155 18380 12164
rect 18328 12121 18337 12155
rect 18337 12121 18371 12155
rect 18371 12121 18380 12155
rect 18328 12112 18380 12121
rect 18512 12112 18564 12164
rect 19064 12112 19116 12164
rect 19984 12155 20036 12164
rect 19984 12121 19993 12155
rect 19993 12121 20027 12155
rect 20027 12121 20036 12155
rect 19984 12112 20036 12121
rect 20720 12112 20772 12164
rect 20996 12112 21048 12164
rect 21640 12155 21692 12164
rect 21640 12121 21649 12155
rect 21649 12121 21683 12155
rect 21683 12121 21692 12155
rect 21640 12112 21692 12121
rect 24216 12112 24268 12164
rect 25320 12112 25372 12164
rect 17408 12044 17460 12096
rect 17500 12044 17552 12096
rect 18696 12044 18748 12096
rect 18788 12044 18840 12096
rect 19248 12044 19300 12096
rect 20260 12044 20312 12096
rect 22560 12044 22612 12096
rect 23296 12044 23348 12096
rect 24860 12044 24912 12096
rect 29092 12112 29144 12164
rect 29276 12112 29328 12164
rect 29368 12112 29420 12164
rect 30196 12112 30248 12164
rect 31484 12112 31536 12164
rect 33784 12112 33836 12164
rect 35440 12112 35492 12164
rect 27068 12044 27120 12096
rect 27252 12087 27304 12096
rect 27252 12053 27261 12087
rect 27261 12053 27295 12087
rect 27295 12053 27304 12087
rect 27252 12044 27304 12053
rect 27712 12044 27764 12096
rect 28080 12044 28132 12096
rect 28448 12087 28500 12096
rect 28448 12053 28457 12087
rect 28457 12053 28491 12087
rect 28491 12053 28500 12087
rect 28448 12044 28500 12053
rect 29644 12044 29696 12096
rect 32404 12087 32456 12096
rect 32404 12053 32413 12087
rect 32413 12053 32447 12087
rect 32447 12053 32456 12087
rect 32404 12044 32456 12053
rect 32864 12087 32916 12096
rect 32864 12053 32873 12087
rect 32873 12053 32907 12087
rect 32907 12053 32916 12087
rect 32864 12044 32916 12053
rect 33968 12087 34020 12096
rect 33968 12053 33977 12087
rect 33977 12053 34011 12087
rect 34011 12053 34020 12087
rect 33968 12044 34020 12053
rect 34060 12044 34112 12096
rect 34336 12044 34388 12096
rect 34980 12044 35032 12096
rect 35348 12044 35400 12096
rect 35808 12044 35860 12096
rect 35992 12044 36044 12096
rect 36544 12112 36596 12164
rect 41420 12316 41472 12368
rect 43076 12316 43128 12368
rect 39212 12248 39264 12300
rect 45652 12316 45704 12368
rect 47308 12316 47360 12368
rect 39672 12180 39724 12232
rect 39856 12180 39908 12232
rect 40132 12180 40184 12232
rect 41144 12223 41196 12232
rect 41144 12189 41153 12223
rect 41153 12189 41187 12223
rect 41187 12189 41196 12223
rect 41144 12180 41196 12189
rect 41420 12180 41472 12232
rect 46756 12291 46808 12300
rect 46756 12257 46765 12291
rect 46765 12257 46799 12291
rect 46799 12257 46808 12291
rect 46756 12248 46808 12257
rect 49148 12291 49200 12300
rect 49148 12257 49157 12291
rect 49157 12257 49191 12291
rect 49191 12257 49200 12291
rect 49148 12248 49200 12257
rect 37740 12112 37792 12164
rect 37464 12044 37516 12096
rect 38476 12044 38528 12096
rect 38660 12087 38712 12096
rect 38660 12053 38669 12087
rect 38669 12053 38703 12087
rect 38703 12053 38712 12087
rect 38660 12044 38712 12053
rect 39488 12087 39540 12096
rect 39488 12053 39497 12087
rect 39497 12053 39531 12087
rect 39531 12053 39540 12087
rect 39488 12044 39540 12053
rect 39672 12044 39724 12096
rect 42984 12044 43036 12096
rect 45284 12180 45336 12232
rect 46388 12180 46440 12232
rect 46848 12180 46900 12232
rect 44180 12112 44232 12164
rect 45008 12112 45060 12164
rect 50712 12112 50764 12164
rect 43996 12087 44048 12096
rect 43996 12053 44005 12087
rect 44005 12053 44039 12087
rect 44039 12053 44048 12087
rect 43996 12044 44048 12053
rect 45468 12044 45520 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 1768 11883 1820 11892
rect 1768 11849 1777 11883
rect 1777 11849 1811 11883
rect 1811 11849 1820 11883
rect 1768 11840 1820 11849
rect 2596 11883 2648 11892
rect 2596 11849 2605 11883
rect 2605 11849 2639 11883
rect 2639 11849 2648 11883
rect 2596 11840 2648 11849
rect 3608 11840 3660 11892
rect 2872 11772 2924 11824
rect 4344 11840 4396 11892
rect 4804 11840 4856 11892
rect 5448 11883 5500 11892
rect 5448 11849 5457 11883
rect 5457 11849 5491 11883
rect 5491 11849 5500 11883
rect 5448 11840 5500 11849
rect 1308 11704 1360 11756
rect 1860 11704 1912 11756
rect 4068 11772 4120 11824
rect 10232 11840 10284 11892
rect 6092 11772 6144 11824
rect 2872 11636 2924 11688
rect 3700 11704 3752 11756
rect 5264 11704 5316 11756
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 7196 11747 7248 11756
rect 7196 11713 7205 11747
rect 7205 11713 7239 11747
rect 7239 11713 7248 11747
rect 7196 11704 7248 11713
rect 7748 11772 7800 11824
rect 6092 11636 6144 11688
rect 7840 11679 7892 11688
rect 7840 11645 7849 11679
rect 7849 11645 7883 11679
rect 7883 11645 7892 11679
rect 7840 11636 7892 11645
rect 4620 11568 4672 11620
rect 5264 11611 5316 11620
rect 5264 11577 5273 11611
rect 5273 11577 5307 11611
rect 5307 11577 5316 11611
rect 5264 11568 5316 11577
rect 5540 11568 5592 11620
rect 9864 11704 9916 11756
rect 13912 11840 13964 11892
rect 14464 11840 14516 11892
rect 16028 11840 16080 11892
rect 10968 11772 11020 11824
rect 11980 11815 12032 11824
rect 11980 11781 11989 11815
rect 11989 11781 12023 11815
rect 12023 11781 12032 11815
rect 11980 11772 12032 11781
rect 12072 11772 12124 11824
rect 12256 11772 12308 11824
rect 13728 11815 13780 11824
rect 13728 11781 13737 11815
rect 13737 11781 13771 11815
rect 13771 11781 13780 11815
rect 13728 11772 13780 11781
rect 15292 11772 15344 11824
rect 14280 11704 14332 11756
rect 14924 11704 14976 11756
rect 21088 11840 21140 11892
rect 18236 11772 18288 11824
rect 25228 11840 25280 11892
rect 25780 11883 25832 11892
rect 25780 11849 25789 11883
rect 25789 11849 25823 11883
rect 25823 11849 25832 11883
rect 25780 11840 25832 11849
rect 25872 11840 25924 11892
rect 29368 11840 29420 11892
rect 30196 11840 30248 11892
rect 30748 11840 30800 11892
rect 22284 11772 22336 11824
rect 23756 11772 23808 11824
rect 23940 11772 23992 11824
rect 26056 11772 26108 11824
rect 27252 11772 27304 11824
rect 28356 11772 28408 11824
rect 29092 11772 29144 11824
rect 32772 11840 32824 11892
rect 32864 11840 32916 11892
rect 36912 11840 36964 11892
rect 35992 11772 36044 11824
rect 37740 11815 37792 11824
rect 37740 11781 37749 11815
rect 37749 11781 37783 11815
rect 37783 11781 37792 11815
rect 37740 11772 37792 11781
rect 39212 11883 39264 11892
rect 39212 11849 39221 11883
rect 39221 11849 39255 11883
rect 39255 11849 39264 11883
rect 39212 11840 39264 11849
rect 40316 11883 40368 11892
rect 40316 11849 40325 11883
rect 40325 11849 40359 11883
rect 40359 11849 40368 11883
rect 40316 11840 40368 11849
rect 41420 11883 41472 11892
rect 41420 11849 41429 11883
rect 41429 11849 41463 11883
rect 41463 11849 41472 11883
rect 41420 11840 41472 11849
rect 41880 11883 41932 11892
rect 41880 11849 41889 11883
rect 41889 11849 41923 11883
rect 41923 11849 41932 11883
rect 41880 11840 41932 11849
rect 42432 11840 42484 11892
rect 44272 11840 44324 11892
rect 44364 11883 44416 11892
rect 44364 11849 44373 11883
rect 44373 11849 44407 11883
rect 44407 11849 44416 11883
rect 44364 11840 44416 11849
rect 44732 11840 44784 11892
rect 47124 11883 47176 11892
rect 47124 11849 47133 11883
rect 47133 11849 47167 11883
rect 47167 11849 47176 11883
rect 47124 11840 47176 11849
rect 39856 11772 39908 11824
rect 10324 11636 10376 11688
rect 10784 11568 10836 11620
rect 10968 11568 11020 11620
rect 13360 11636 13412 11688
rect 15016 11679 15068 11688
rect 15016 11645 15025 11679
rect 15025 11645 15059 11679
rect 15059 11645 15068 11679
rect 15016 11636 15068 11645
rect 15568 11636 15620 11688
rect 16212 11679 16264 11688
rect 16212 11645 16221 11679
rect 16221 11645 16255 11679
rect 16255 11645 16264 11679
rect 16212 11636 16264 11645
rect 14188 11568 14240 11620
rect 17500 11704 17552 11756
rect 20720 11704 20772 11756
rect 21088 11747 21140 11756
rect 21088 11713 21097 11747
rect 21097 11713 21131 11747
rect 21131 11713 21140 11747
rect 21088 11704 21140 11713
rect 21824 11704 21876 11756
rect 24400 11704 24452 11756
rect 19248 11636 19300 11688
rect 21272 11636 21324 11688
rect 21364 11679 21416 11688
rect 21364 11645 21373 11679
rect 21373 11645 21407 11679
rect 21407 11645 21416 11679
rect 21364 11636 21416 11645
rect 21640 11636 21692 11688
rect 23940 11636 23992 11688
rect 25044 11636 25096 11688
rect 25412 11636 25464 11688
rect 25596 11704 25648 11756
rect 3884 11543 3936 11552
rect 3884 11509 3893 11543
rect 3893 11509 3927 11543
rect 3927 11509 3936 11543
rect 3884 11500 3936 11509
rect 4344 11500 4396 11552
rect 7380 11500 7432 11552
rect 9404 11500 9456 11552
rect 11060 11500 11112 11552
rect 11336 11500 11388 11552
rect 12440 11500 12492 11552
rect 13084 11500 13136 11552
rect 13360 11500 13412 11552
rect 19064 11568 19116 11620
rect 16672 11500 16724 11552
rect 16764 11543 16816 11552
rect 16764 11509 16773 11543
rect 16773 11509 16807 11543
rect 16807 11509 16816 11543
rect 16764 11500 16816 11509
rect 17224 11500 17276 11552
rect 17776 11500 17828 11552
rect 17960 11500 18012 11552
rect 20444 11568 20496 11620
rect 20996 11568 21048 11620
rect 23664 11568 23716 11620
rect 26424 11568 26476 11620
rect 27344 11568 27396 11620
rect 29920 11704 29972 11756
rect 32680 11747 32732 11756
rect 32680 11713 32689 11747
rect 32689 11713 32723 11747
rect 32723 11713 32732 11747
rect 32680 11704 32732 11713
rect 35808 11704 35860 11756
rect 38844 11704 38896 11756
rect 40224 11704 40276 11756
rect 40592 11704 40644 11756
rect 41512 11704 41564 11756
rect 42156 11704 42208 11756
rect 27620 11679 27672 11688
rect 27620 11645 27629 11679
rect 27629 11645 27663 11679
rect 27663 11645 27672 11679
rect 27620 11636 27672 11645
rect 27804 11679 27856 11688
rect 27804 11645 27813 11679
rect 27813 11645 27847 11679
rect 27847 11645 27856 11679
rect 27804 11636 27856 11645
rect 27712 11568 27764 11620
rect 19340 11500 19392 11552
rect 19616 11500 19668 11552
rect 19892 11500 19944 11552
rect 22284 11500 22336 11552
rect 22468 11500 22520 11552
rect 24952 11500 25004 11552
rect 27068 11500 27120 11552
rect 27160 11543 27212 11552
rect 27160 11509 27169 11543
rect 27169 11509 27203 11543
rect 27203 11509 27212 11543
rect 27160 11500 27212 11509
rect 27252 11500 27304 11552
rect 28632 11636 28684 11688
rect 30196 11636 30248 11688
rect 31852 11636 31904 11688
rect 29920 11568 29972 11620
rect 33508 11679 33560 11688
rect 33508 11645 33517 11679
rect 33517 11645 33551 11679
rect 33551 11645 33560 11679
rect 33508 11636 33560 11645
rect 33784 11679 33836 11688
rect 33784 11645 33793 11679
rect 33793 11645 33827 11679
rect 33827 11645 33836 11679
rect 33784 11636 33836 11645
rect 34520 11636 34572 11688
rect 35900 11636 35952 11688
rect 36544 11636 36596 11688
rect 37188 11636 37240 11688
rect 35716 11568 35768 11620
rect 37740 11636 37792 11688
rect 42984 11636 43036 11688
rect 44180 11747 44232 11756
rect 44180 11713 44189 11747
rect 44189 11713 44223 11747
rect 44223 11713 44232 11747
rect 44180 11704 44232 11713
rect 44916 11747 44968 11756
rect 44916 11713 44925 11747
rect 44925 11713 44959 11747
rect 44959 11713 44968 11747
rect 44916 11704 44968 11713
rect 45376 11704 45428 11756
rect 46112 11772 46164 11824
rect 49148 11815 49200 11824
rect 49148 11781 49157 11815
rect 49157 11781 49191 11815
rect 49191 11781 49200 11815
rect 49148 11772 49200 11781
rect 46848 11704 46900 11756
rect 46940 11747 46992 11756
rect 46940 11713 46949 11747
rect 46949 11713 46983 11747
rect 46983 11713 46992 11747
rect 46940 11704 46992 11713
rect 47032 11704 47084 11756
rect 45192 11636 45244 11688
rect 41696 11568 41748 11620
rect 43076 11568 43128 11620
rect 29736 11500 29788 11552
rect 30932 11500 30984 11552
rect 31116 11500 31168 11552
rect 35624 11500 35676 11552
rect 39764 11500 39816 11552
rect 42432 11500 42484 11552
rect 45468 11568 45520 11620
rect 44272 11500 44324 11552
rect 50804 11636 50856 11688
rect 47124 11500 47176 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 2688 11271 2740 11280
rect 2688 11237 2697 11271
rect 2697 11237 2731 11271
rect 2731 11237 2740 11271
rect 2688 11228 2740 11237
rect 3332 11339 3384 11348
rect 3332 11305 3341 11339
rect 3341 11305 3375 11339
rect 3375 11305 3384 11339
rect 3332 11296 3384 11305
rect 3700 11296 3752 11348
rect 4436 11339 4488 11348
rect 4436 11305 4445 11339
rect 4445 11305 4479 11339
rect 4479 11305 4488 11339
rect 4436 11296 4488 11305
rect 5172 11339 5224 11348
rect 5172 11305 5181 11339
rect 5181 11305 5215 11339
rect 5215 11305 5224 11339
rect 5172 11296 5224 11305
rect 5724 11339 5776 11348
rect 5724 11305 5733 11339
rect 5733 11305 5767 11339
rect 5767 11305 5776 11339
rect 5724 11296 5776 11305
rect 6276 11339 6328 11348
rect 6276 11305 6285 11339
rect 6285 11305 6319 11339
rect 6319 11305 6328 11339
rect 6276 11296 6328 11305
rect 8944 11339 8996 11348
rect 8944 11305 8953 11339
rect 8953 11305 8987 11339
rect 8987 11305 8996 11339
rect 8944 11296 8996 11305
rect 9312 11339 9364 11348
rect 9312 11305 9321 11339
rect 9321 11305 9355 11339
rect 9355 11305 9364 11339
rect 9312 11296 9364 11305
rect 14004 11296 14056 11348
rect 14464 11296 14516 11348
rect 14832 11296 14884 11348
rect 18512 11296 18564 11348
rect 18604 11296 18656 11348
rect 5540 11228 5592 11280
rect 1584 11135 1636 11144
rect 1584 11101 1593 11135
rect 1593 11101 1627 11135
rect 1627 11101 1636 11135
rect 1584 11092 1636 11101
rect 4344 11135 4396 11144
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 2780 11024 2832 11076
rect 9864 11228 9916 11280
rect 14924 11228 14976 11280
rect 15200 11228 15252 11280
rect 6460 11092 6512 11144
rect 8944 11160 8996 11212
rect 9128 11203 9180 11212
rect 9128 11169 9137 11203
rect 9137 11169 9171 11203
rect 9171 11169 9180 11203
rect 9128 11160 9180 11169
rect 10048 11160 10100 11212
rect 12256 11160 12308 11212
rect 12716 11160 12768 11212
rect 13728 11160 13780 11212
rect 14648 11160 14700 11212
rect 15476 11160 15528 11212
rect 16856 11228 16908 11280
rect 18420 11228 18472 11280
rect 18512 11160 18564 11212
rect 18604 11203 18656 11212
rect 18604 11169 18613 11203
rect 18613 11169 18647 11203
rect 18647 11169 18656 11203
rect 18604 11160 18656 11169
rect 18788 11296 18840 11348
rect 19432 11296 19484 11348
rect 19892 11339 19944 11348
rect 19892 11305 19901 11339
rect 19901 11305 19935 11339
rect 19935 11305 19944 11339
rect 19892 11296 19944 11305
rect 20076 11339 20128 11348
rect 20076 11305 20085 11339
rect 20085 11305 20119 11339
rect 20119 11305 20128 11339
rect 20076 11296 20128 11305
rect 20628 11296 20680 11348
rect 24952 11296 25004 11348
rect 25228 11296 25280 11348
rect 26332 11339 26384 11348
rect 26332 11305 26341 11339
rect 26341 11305 26375 11339
rect 26375 11305 26384 11339
rect 26332 11296 26384 11305
rect 27712 11296 27764 11348
rect 29552 11296 29604 11348
rect 23388 11271 23440 11280
rect 23388 11237 23397 11271
rect 23397 11237 23431 11271
rect 23431 11237 23440 11271
rect 23388 11228 23440 11237
rect 29920 11228 29972 11280
rect 10232 11092 10284 11144
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 12808 11092 12860 11144
rect 16396 11092 16448 11144
rect 7380 11024 7432 11076
rect 12348 11024 12400 11076
rect 13912 11024 13964 11076
rect 14188 11024 14240 11076
rect 1952 10956 2004 11008
rect 5264 10956 5316 11008
rect 6920 10956 6972 11008
rect 12440 10956 12492 11008
rect 14648 10956 14700 11008
rect 15752 10999 15804 11008
rect 15752 10965 15761 10999
rect 15761 10965 15795 10999
rect 15795 10965 15804 10999
rect 15752 10956 15804 10965
rect 16120 11067 16172 11076
rect 16120 11033 16129 11067
rect 16129 11033 16163 11067
rect 16163 11033 16172 11067
rect 16120 11024 16172 11033
rect 17960 11092 18012 11144
rect 21364 11160 21416 11212
rect 22652 11160 22704 11212
rect 24584 11203 24636 11212
rect 24584 11169 24593 11203
rect 24593 11169 24627 11203
rect 24627 11169 24636 11203
rect 24584 11160 24636 11169
rect 26792 11160 26844 11212
rect 27252 11160 27304 11212
rect 29092 11160 29144 11212
rect 29276 11160 29328 11212
rect 32772 11296 32824 11348
rect 32220 11228 32272 11280
rect 34888 11296 34940 11348
rect 35072 11339 35124 11348
rect 35072 11305 35081 11339
rect 35081 11305 35115 11339
rect 35115 11305 35124 11339
rect 35072 11296 35124 11305
rect 35164 11296 35216 11348
rect 35992 11296 36044 11348
rect 34060 11228 34112 11280
rect 32128 11160 32180 11212
rect 34980 11228 35032 11280
rect 38568 11296 38620 11348
rect 39120 11339 39172 11348
rect 39120 11305 39129 11339
rect 39129 11305 39163 11339
rect 39163 11305 39172 11339
rect 39120 11296 39172 11305
rect 39856 11296 39908 11348
rect 37556 11228 37608 11280
rect 40592 11296 40644 11348
rect 41788 11296 41840 11348
rect 42708 11296 42760 11348
rect 43444 11296 43496 11348
rect 41880 11228 41932 11280
rect 44548 11296 44600 11348
rect 44732 11228 44784 11280
rect 45284 11296 45336 11348
rect 46572 11296 46624 11348
rect 47400 11339 47452 11348
rect 47400 11305 47409 11339
rect 47409 11305 47443 11339
rect 47443 11305 47452 11339
rect 47400 11296 47452 11305
rect 45192 11228 45244 11280
rect 48504 11228 48556 11280
rect 17316 11067 17368 11076
rect 17316 11033 17325 11067
rect 17325 11033 17359 11067
rect 17359 11033 17368 11067
rect 17316 11024 17368 11033
rect 16948 10956 17000 11008
rect 17684 10956 17736 11008
rect 18972 11092 19024 11144
rect 19432 11092 19484 11144
rect 19708 11092 19760 11144
rect 21640 11135 21692 11144
rect 21640 11101 21649 11135
rect 21649 11101 21683 11135
rect 21683 11101 21692 11135
rect 21640 11092 21692 11101
rect 28632 11092 28684 11144
rect 18236 11024 18288 11076
rect 21824 11024 21876 11076
rect 21916 11067 21968 11076
rect 21916 11033 21925 11067
rect 21925 11033 21959 11067
rect 21959 11033 21968 11067
rect 21916 11024 21968 11033
rect 19248 10956 19300 11008
rect 20720 10956 20772 11008
rect 22376 11024 22428 11076
rect 25136 11024 25188 11076
rect 25412 11024 25464 11076
rect 29828 11092 29880 11144
rect 30288 11092 30340 11144
rect 33416 11135 33468 11144
rect 33416 11101 33425 11135
rect 33425 11101 33459 11135
rect 33459 11101 33468 11135
rect 33416 11092 33468 11101
rect 30748 11024 30800 11076
rect 31760 11024 31812 11076
rect 35256 11160 35308 11212
rect 35716 11160 35768 11212
rect 41972 11160 42024 11212
rect 44180 11160 44232 11212
rect 46848 11160 46900 11212
rect 34152 11135 34204 11144
rect 34152 11101 34161 11135
rect 34161 11101 34195 11135
rect 34195 11101 34204 11135
rect 34152 11092 34204 11101
rect 35164 11092 35216 11144
rect 35808 11092 35860 11144
rect 37280 11092 37332 11144
rect 24952 10956 25004 11008
rect 29000 10956 29052 11008
rect 32588 10999 32640 11008
rect 32588 10965 32597 10999
rect 32597 10965 32631 10999
rect 32631 10965 32640 10999
rect 37648 11024 37700 11076
rect 38292 11092 38344 11144
rect 38568 11092 38620 11144
rect 39672 11135 39724 11144
rect 39672 11101 39681 11135
rect 39681 11101 39715 11135
rect 39715 11101 39724 11135
rect 39672 11092 39724 11101
rect 32588 10956 32640 10965
rect 36176 10956 36228 11008
rect 36544 10956 36596 11008
rect 38844 11024 38896 11076
rect 40132 11092 40184 11144
rect 41144 11135 41196 11144
rect 41144 11101 41153 11135
rect 41153 11101 41187 11135
rect 41187 11101 41196 11135
rect 41144 11092 41196 11101
rect 42064 11092 42116 11144
rect 43352 11092 43404 11144
rect 43444 11092 43496 11144
rect 44548 11092 44600 11144
rect 45468 11092 45520 11144
rect 46112 11092 46164 11144
rect 47400 11092 47452 11144
rect 49148 11203 49200 11212
rect 49148 11169 49157 11203
rect 49157 11169 49191 11203
rect 49191 11169 49200 11203
rect 49148 11160 49200 11169
rect 41604 11024 41656 11076
rect 42708 11024 42760 11076
rect 43260 11024 43312 11076
rect 45284 11024 45336 11076
rect 49424 11024 49476 11076
rect 39028 10956 39080 11008
rect 44548 10956 44600 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 2872 10795 2924 10804
rect 2872 10761 2881 10795
rect 2881 10761 2915 10795
rect 2915 10761 2924 10795
rect 2872 10752 2924 10761
rect 4068 10752 4120 10804
rect 4528 10752 4580 10804
rect 1216 10616 1268 10668
rect 3332 10684 3384 10736
rect 5264 10684 5316 10736
rect 8852 10752 8904 10804
rect 9312 10752 9364 10804
rect 11612 10795 11664 10804
rect 11612 10761 11621 10795
rect 11621 10761 11655 10795
rect 11655 10761 11664 10795
rect 11612 10752 11664 10761
rect 11704 10752 11756 10804
rect 12716 10752 12768 10804
rect 15568 10752 15620 10804
rect 7104 10727 7156 10736
rect 7104 10693 7113 10727
rect 7113 10693 7147 10727
rect 7147 10693 7156 10727
rect 7104 10684 7156 10693
rect 10784 10684 10836 10736
rect 1308 10548 1360 10600
rect 3700 10659 3752 10668
rect 3700 10625 3709 10659
rect 3709 10625 3743 10659
rect 3743 10625 3752 10659
rect 3700 10616 3752 10625
rect 3792 10616 3844 10668
rect 6184 10616 6236 10668
rect 6920 10659 6972 10668
rect 6920 10625 6929 10659
rect 6929 10625 6963 10659
rect 6963 10625 6972 10659
rect 6920 10616 6972 10625
rect 2412 10548 2464 10600
rect 4344 10548 4396 10600
rect 6000 10548 6052 10600
rect 8300 10659 8352 10668
rect 8300 10625 8309 10659
rect 8309 10625 8343 10659
rect 8343 10625 8352 10659
rect 8300 10616 8352 10625
rect 9036 10616 9088 10668
rect 9404 10659 9456 10668
rect 9404 10625 9413 10659
rect 9413 10625 9447 10659
rect 9447 10625 9456 10659
rect 9404 10616 9456 10625
rect 9956 10616 10008 10668
rect 11428 10616 11480 10668
rect 12164 10616 12216 10668
rect 12256 10616 12308 10668
rect 13360 10684 13412 10736
rect 15292 10684 15344 10736
rect 17316 10752 17368 10804
rect 17776 10752 17828 10804
rect 18512 10752 18564 10804
rect 19340 10752 19392 10804
rect 19432 10795 19484 10804
rect 19432 10761 19441 10795
rect 19441 10761 19475 10795
rect 19475 10761 19484 10795
rect 19432 10752 19484 10761
rect 15108 10616 15160 10668
rect 10968 10548 11020 10600
rect 12532 10591 12584 10600
rect 12532 10557 12541 10591
rect 12541 10557 12575 10591
rect 12575 10557 12584 10591
rect 12532 10548 12584 10557
rect 12808 10548 12860 10600
rect 14464 10548 14516 10600
rect 15200 10591 15252 10600
rect 15200 10557 15209 10591
rect 15209 10557 15243 10591
rect 15243 10557 15252 10591
rect 15200 10548 15252 10557
rect 1768 10523 1820 10532
rect 1768 10489 1777 10523
rect 1777 10489 1811 10523
rect 1811 10489 1820 10523
rect 1768 10480 1820 10489
rect 8024 10480 8076 10532
rect 5724 10412 5776 10464
rect 6000 10412 6052 10464
rect 10692 10480 10744 10532
rect 17316 10659 17368 10668
rect 17316 10625 17325 10659
rect 17325 10625 17359 10659
rect 17359 10625 17368 10659
rect 17316 10616 17368 10625
rect 16580 10548 16632 10600
rect 17776 10616 17828 10668
rect 19616 10684 19668 10736
rect 18972 10616 19024 10668
rect 21640 10752 21692 10804
rect 24032 10752 24084 10804
rect 20720 10684 20772 10736
rect 21824 10684 21876 10736
rect 17868 10548 17920 10600
rect 11244 10412 11296 10464
rect 12164 10412 12216 10464
rect 18512 10480 18564 10532
rect 18696 10591 18748 10600
rect 18696 10557 18705 10591
rect 18705 10557 18739 10591
rect 18739 10557 18748 10591
rect 18696 10548 18748 10557
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 19984 10591 20036 10600
rect 19984 10557 19993 10591
rect 19993 10557 20027 10591
rect 20027 10557 20036 10591
rect 19984 10548 20036 10557
rect 20628 10548 20680 10600
rect 26240 10752 26292 10804
rect 26516 10795 26568 10804
rect 26516 10761 26525 10795
rect 26525 10761 26559 10795
rect 26559 10761 26568 10795
rect 26516 10752 26568 10761
rect 27804 10752 27856 10804
rect 28724 10752 28776 10804
rect 24400 10684 24452 10736
rect 27160 10684 27212 10736
rect 31668 10752 31720 10804
rect 23480 10616 23532 10668
rect 24216 10659 24268 10668
rect 24216 10625 24225 10659
rect 24225 10625 24259 10659
rect 24259 10625 24268 10659
rect 24216 10616 24268 10625
rect 28080 10616 28132 10668
rect 29184 10616 29236 10668
rect 31484 10616 31536 10668
rect 32404 10616 32456 10668
rect 32864 10616 32916 10668
rect 35072 10752 35124 10804
rect 35532 10795 35584 10804
rect 35532 10761 35541 10795
rect 35541 10761 35575 10795
rect 35575 10761 35584 10795
rect 35532 10752 35584 10761
rect 36636 10752 36688 10804
rect 37004 10752 37056 10804
rect 37096 10795 37148 10804
rect 37096 10761 37105 10795
rect 37105 10761 37139 10795
rect 37139 10761 37148 10795
rect 37096 10752 37148 10761
rect 37556 10752 37608 10804
rect 38016 10752 38068 10804
rect 42064 10795 42116 10804
rect 42064 10761 42073 10795
rect 42073 10761 42107 10795
rect 42107 10761 42116 10795
rect 42064 10752 42116 10761
rect 43444 10752 43496 10804
rect 47676 10795 47728 10804
rect 47676 10761 47685 10795
rect 47685 10761 47719 10795
rect 47719 10761 47728 10795
rect 47676 10752 47728 10761
rect 35440 10684 35492 10736
rect 36176 10616 36228 10668
rect 22744 10591 22796 10600
rect 22744 10557 22753 10591
rect 22753 10557 22787 10591
rect 22787 10557 22796 10591
rect 22744 10548 22796 10557
rect 23296 10591 23348 10600
rect 23296 10557 23305 10591
rect 23305 10557 23339 10591
rect 23339 10557 23348 10591
rect 23296 10548 23348 10557
rect 25872 10548 25924 10600
rect 26056 10548 26108 10600
rect 26976 10548 27028 10600
rect 27804 10548 27856 10600
rect 28540 10548 28592 10600
rect 29736 10548 29788 10600
rect 30656 10548 30708 10600
rect 15200 10412 15252 10464
rect 17132 10412 17184 10464
rect 17960 10412 18012 10464
rect 19156 10455 19208 10464
rect 19156 10421 19165 10455
rect 19165 10421 19199 10455
rect 19199 10421 19208 10455
rect 19156 10412 19208 10421
rect 23572 10480 23624 10532
rect 21364 10412 21416 10464
rect 23664 10412 23716 10464
rect 24032 10412 24084 10464
rect 24308 10412 24360 10464
rect 24676 10412 24728 10464
rect 29552 10455 29604 10464
rect 29552 10421 29561 10455
rect 29561 10421 29595 10455
rect 29595 10421 29604 10455
rect 29552 10412 29604 10421
rect 32680 10548 32732 10600
rect 32772 10548 32824 10600
rect 31392 10480 31444 10532
rect 31944 10480 31996 10532
rect 33508 10480 33560 10532
rect 36268 10548 36320 10600
rect 36544 10548 36596 10600
rect 36636 10591 36688 10600
rect 36636 10557 36645 10591
rect 36645 10557 36679 10591
rect 36679 10557 36688 10591
rect 36636 10548 36688 10557
rect 37464 10684 37516 10736
rect 36912 10616 36964 10668
rect 37648 10616 37700 10668
rect 37832 10659 37884 10668
rect 37832 10625 37841 10659
rect 37841 10625 37875 10659
rect 37875 10625 37884 10659
rect 37832 10616 37884 10625
rect 38568 10616 38620 10668
rect 39580 10616 39632 10668
rect 43628 10684 43680 10736
rect 45560 10684 45612 10736
rect 35348 10480 35400 10532
rect 32036 10412 32088 10464
rect 33324 10412 33376 10464
rect 36912 10412 36964 10464
rect 38108 10548 38160 10600
rect 38292 10548 38344 10600
rect 40960 10616 41012 10668
rect 44088 10616 44140 10668
rect 44548 10659 44600 10668
rect 44548 10625 44557 10659
rect 44557 10625 44591 10659
rect 44591 10625 44600 10659
rect 44548 10616 44600 10625
rect 46204 10684 46256 10736
rect 48596 10684 48648 10736
rect 49332 10684 49384 10736
rect 46112 10659 46164 10668
rect 46112 10625 46121 10659
rect 46121 10625 46155 10659
rect 46155 10625 46164 10659
rect 46112 10616 46164 10625
rect 39856 10548 39908 10600
rect 41880 10548 41932 10600
rect 42156 10591 42208 10600
rect 42156 10557 42165 10591
rect 42165 10557 42199 10591
rect 42199 10557 42208 10591
rect 42156 10548 42208 10557
rect 42616 10548 42668 10600
rect 43720 10548 43772 10600
rect 44732 10548 44784 10600
rect 38568 10480 38620 10532
rect 40408 10455 40460 10464
rect 40408 10421 40417 10455
rect 40417 10421 40451 10455
rect 40451 10421 40460 10455
rect 40408 10412 40460 10421
rect 40684 10412 40736 10464
rect 43996 10480 44048 10532
rect 45376 10480 45428 10532
rect 48872 10548 48924 10600
rect 44088 10412 44140 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 1584 10208 1636 10260
rect 3700 10208 3752 10260
rect 5172 10251 5224 10260
rect 5172 10217 5181 10251
rect 5181 10217 5215 10251
rect 5215 10217 5224 10251
rect 5172 10208 5224 10217
rect 5908 10251 5960 10260
rect 5908 10217 5917 10251
rect 5917 10217 5951 10251
rect 5951 10217 5960 10251
rect 5908 10208 5960 10217
rect 7380 10251 7432 10260
rect 7380 10217 7389 10251
rect 7389 10217 7423 10251
rect 7423 10217 7432 10251
rect 7380 10208 7432 10217
rect 4252 10115 4304 10124
rect 4252 10081 4261 10115
rect 4261 10081 4295 10115
rect 4295 10081 4304 10115
rect 4252 10072 4304 10081
rect 5816 10140 5868 10192
rect 8668 10208 8720 10260
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 9588 10208 9640 10260
rect 12808 10208 12860 10260
rect 13912 10208 13964 10260
rect 15292 10208 15344 10260
rect 16212 10208 16264 10260
rect 16580 10208 16632 10260
rect 16948 10251 17000 10260
rect 16948 10217 16957 10251
rect 16957 10217 16991 10251
rect 16991 10217 17000 10251
rect 16948 10208 17000 10217
rect 8392 10140 8444 10192
rect 10876 10140 10928 10192
rect 12072 10140 12124 10192
rect 15568 10140 15620 10192
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 5540 10004 5592 10056
rect 5632 9936 5684 9988
rect 6368 9936 6420 9988
rect 10416 10072 10468 10124
rect 12348 10115 12400 10124
rect 12348 10081 12357 10115
rect 12357 10081 12391 10115
rect 12391 10081 12400 10115
rect 12348 10072 12400 10081
rect 13452 10115 13504 10124
rect 13452 10081 13461 10115
rect 13461 10081 13495 10115
rect 13495 10081 13504 10115
rect 13452 10072 13504 10081
rect 13636 10115 13688 10124
rect 13636 10081 13645 10115
rect 13645 10081 13679 10115
rect 13679 10081 13688 10115
rect 13636 10072 13688 10081
rect 6000 9868 6052 9920
rect 8024 10004 8076 10056
rect 8392 10004 8444 10056
rect 8484 10004 8536 10056
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 12164 10047 12216 10056
rect 12164 10013 12173 10047
rect 12173 10013 12207 10047
rect 12207 10013 12216 10047
rect 12164 10004 12216 10013
rect 9680 9936 9732 9988
rect 13268 10004 13320 10056
rect 16304 10072 16356 10124
rect 16120 10004 16172 10056
rect 17408 10208 17460 10260
rect 18052 10208 18104 10260
rect 18604 10208 18656 10260
rect 23756 10208 23808 10260
rect 24216 10208 24268 10260
rect 25964 10208 26016 10260
rect 17500 10072 17552 10124
rect 18512 10072 18564 10124
rect 22100 10140 22152 10192
rect 13176 9936 13228 9988
rect 14464 9936 14516 9988
rect 14832 9936 14884 9988
rect 15292 9936 15344 9988
rect 17776 10004 17828 10056
rect 17960 9936 18012 9988
rect 11796 9911 11848 9920
rect 11796 9877 11805 9911
rect 11805 9877 11839 9911
rect 11839 9877 11848 9911
rect 11796 9868 11848 9877
rect 13360 9911 13412 9920
rect 13360 9877 13369 9911
rect 13369 9877 13403 9911
rect 13403 9877 13412 9911
rect 13360 9868 13412 9877
rect 13820 9868 13872 9920
rect 18052 9868 18104 9920
rect 18144 9911 18196 9920
rect 18144 9877 18153 9911
rect 18153 9877 18187 9911
rect 18187 9877 18196 9911
rect 18144 9868 18196 9877
rect 19156 9868 19208 9920
rect 19708 10072 19760 10124
rect 20352 10072 20404 10124
rect 22008 10072 22060 10124
rect 22652 10072 22704 10124
rect 23388 10115 23440 10124
rect 23388 10081 23397 10115
rect 23397 10081 23431 10115
rect 23431 10081 23440 10115
rect 23388 10072 23440 10081
rect 23296 10004 23348 10056
rect 19340 9936 19392 9988
rect 20720 9936 20772 9988
rect 21272 9936 21324 9988
rect 22008 9936 22060 9988
rect 22652 9936 22704 9988
rect 23572 10072 23624 10124
rect 24768 10140 24820 10192
rect 25228 10115 25280 10124
rect 25228 10081 25237 10115
rect 25237 10081 25271 10115
rect 25271 10081 25280 10115
rect 25228 10072 25280 10081
rect 24952 10047 25004 10056
rect 24952 10013 24961 10047
rect 24961 10013 24995 10047
rect 24995 10013 25004 10047
rect 24952 10004 25004 10013
rect 25320 10004 25372 10056
rect 25964 10072 26016 10124
rect 24400 9936 24452 9988
rect 25412 9936 25464 9988
rect 20076 9868 20128 9920
rect 22192 9911 22244 9920
rect 22192 9877 22201 9911
rect 22201 9877 22235 9911
rect 22235 9877 22244 9911
rect 22192 9868 22244 9877
rect 22928 9868 22980 9920
rect 26792 10115 26844 10124
rect 26792 10081 26801 10115
rect 26801 10081 26835 10115
rect 26835 10081 26844 10115
rect 26792 10072 26844 10081
rect 28908 10208 28960 10260
rect 30932 10208 30984 10260
rect 28448 10140 28500 10192
rect 29184 10072 29236 10124
rect 29552 10072 29604 10124
rect 30380 10115 30432 10124
rect 30380 10081 30389 10115
rect 30389 10081 30423 10115
rect 30423 10081 30432 10115
rect 30380 10072 30432 10081
rect 31392 10072 31444 10124
rect 33784 10208 33836 10260
rect 36452 10208 36504 10260
rect 36636 10208 36688 10260
rect 38660 10208 38712 10260
rect 41144 10208 41196 10260
rect 43720 10251 43772 10260
rect 43720 10217 43729 10251
rect 43729 10217 43763 10251
rect 43763 10217 43772 10251
rect 43720 10208 43772 10217
rect 45192 10208 45244 10260
rect 48412 10208 48464 10260
rect 34520 10140 34572 10192
rect 33508 10072 33560 10124
rect 40408 10140 40460 10192
rect 36912 10072 36964 10124
rect 38016 10115 38068 10124
rect 38016 10081 38025 10115
rect 38025 10081 38059 10115
rect 38059 10081 38068 10115
rect 38016 10072 38068 10081
rect 28632 9936 28684 9988
rect 29276 9936 29328 9988
rect 27804 9868 27856 9920
rect 28080 9868 28132 9920
rect 36452 10004 36504 10056
rect 39396 10072 39448 10124
rect 38660 10047 38712 10056
rect 38660 10013 38669 10047
rect 38669 10013 38703 10047
rect 38703 10013 38712 10047
rect 38660 10004 38712 10013
rect 40684 10004 40736 10056
rect 42064 10072 42116 10124
rect 30656 9868 30708 9920
rect 30840 9868 30892 9920
rect 31116 9868 31168 9920
rect 31300 9868 31352 9920
rect 32404 9936 32456 9988
rect 36176 9936 36228 9988
rect 34152 9868 34204 9920
rect 34980 9868 35032 9920
rect 36636 9911 36688 9920
rect 36636 9877 36645 9911
rect 36645 9877 36679 9911
rect 36679 9877 36688 9911
rect 36636 9868 36688 9877
rect 37096 9911 37148 9920
rect 37096 9877 37105 9911
rect 37105 9877 37139 9911
rect 37139 9877 37148 9911
rect 37096 9868 37148 9877
rect 37188 9868 37240 9920
rect 38108 9868 38160 9920
rect 39856 9936 39908 9988
rect 42616 10047 42668 10056
rect 42616 10013 42625 10047
rect 42625 10013 42659 10047
rect 42659 10013 42668 10047
rect 42616 10004 42668 10013
rect 43812 10004 43864 10056
rect 44456 10047 44508 10056
rect 44456 10013 44465 10047
rect 44465 10013 44499 10047
rect 44499 10013 44508 10047
rect 44456 10004 44508 10013
rect 45560 10004 45612 10056
rect 46204 10140 46256 10192
rect 47676 10140 47728 10192
rect 46848 10115 46900 10124
rect 46848 10081 46857 10115
rect 46857 10081 46891 10115
rect 46891 10081 46900 10115
rect 46848 10072 46900 10081
rect 49148 10115 49200 10124
rect 49148 10081 49157 10115
rect 49157 10081 49191 10115
rect 49191 10081 49200 10115
rect 49148 10072 49200 10081
rect 41972 9868 42024 9920
rect 42064 9911 42116 9920
rect 42064 9877 42073 9911
rect 42073 9877 42107 9911
rect 42107 9877 42116 9911
rect 42064 9868 42116 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 2412 9707 2464 9716
rect 2412 9673 2421 9707
rect 2421 9673 2455 9707
rect 2455 9673 2464 9707
rect 2412 9664 2464 9673
rect 3608 9664 3660 9716
rect 1216 9528 1268 9580
rect 2136 9528 2188 9580
rect 3516 9528 3568 9580
rect 3608 9571 3660 9580
rect 3608 9537 3617 9571
rect 3617 9537 3651 9571
rect 3651 9537 3660 9571
rect 3608 9528 3660 9537
rect 3976 9528 4028 9580
rect 8300 9664 8352 9716
rect 13176 9664 13228 9716
rect 13452 9664 13504 9716
rect 15752 9664 15804 9716
rect 16212 9664 16264 9716
rect 16948 9664 17000 9716
rect 17132 9664 17184 9716
rect 17500 9664 17552 9716
rect 17776 9664 17828 9716
rect 18144 9664 18196 9716
rect 18420 9664 18472 9716
rect 18512 9664 18564 9716
rect 20444 9664 20496 9716
rect 21364 9664 21416 9716
rect 23388 9664 23440 9716
rect 4712 9639 4764 9648
rect 4712 9605 4721 9639
rect 4721 9605 4755 9639
rect 4755 9605 4764 9639
rect 4712 9596 4764 9605
rect 5724 9596 5776 9648
rect 11060 9596 11112 9648
rect 11244 9596 11296 9648
rect 14004 9596 14056 9648
rect 4160 9528 4212 9580
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 6000 9571 6052 9580
rect 6000 9537 6009 9571
rect 6009 9537 6043 9571
rect 6043 9537 6052 9571
rect 6000 9528 6052 9537
rect 9220 9528 9272 9580
rect 10324 9528 10376 9580
rect 10508 9571 10560 9580
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 12164 9571 12216 9580
rect 12164 9537 12173 9571
rect 12173 9537 12207 9571
rect 12207 9537 12216 9571
rect 12164 9528 12216 9537
rect 13268 9571 13320 9580
rect 13268 9537 13277 9571
rect 13277 9537 13311 9571
rect 13311 9537 13320 9571
rect 13268 9528 13320 9537
rect 15016 9528 15068 9580
rect 15476 9528 15528 9580
rect 16396 9528 16448 9580
rect 16764 9528 16816 9580
rect 6184 9460 6236 9512
rect 1768 9435 1820 9444
rect 1768 9401 1777 9435
rect 1777 9401 1811 9435
rect 1811 9401 1820 9435
rect 1768 9392 1820 9401
rect 2780 9435 2832 9444
rect 2780 9401 2789 9435
rect 2789 9401 2823 9435
rect 2823 9401 2832 9435
rect 2780 9392 2832 9401
rect 6920 9460 6972 9512
rect 9956 9460 10008 9512
rect 11980 9460 12032 9512
rect 13544 9460 13596 9512
rect 2504 9324 2556 9376
rect 7196 9392 7248 9444
rect 5540 9324 5592 9376
rect 7748 9324 7800 9376
rect 8024 9367 8076 9376
rect 8024 9333 8033 9367
rect 8033 9333 8067 9367
rect 8067 9333 8076 9367
rect 8024 9324 8076 9333
rect 9956 9324 10008 9376
rect 13268 9392 13320 9444
rect 16212 9460 16264 9512
rect 18788 9596 18840 9648
rect 19708 9596 19760 9648
rect 21548 9639 21600 9648
rect 21548 9605 21557 9639
rect 21557 9605 21591 9639
rect 21591 9605 21600 9639
rect 21548 9596 21600 9605
rect 22100 9596 22152 9648
rect 20720 9528 20772 9580
rect 22192 9528 22244 9580
rect 24400 9596 24452 9648
rect 23296 9528 23348 9580
rect 23480 9571 23532 9580
rect 23480 9537 23489 9571
rect 23489 9537 23523 9571
rect 23523 9537 23532 9571
rect 23480 9528 23532 9537
rect 25964 9528 26016 9580
rect 17132 9503 17184 9512
rect 17132 9469 17141 9503
rect 17141 9469 17175 9503
rect 17175 9469 17184 9503
rect 17132 9460 17184 9469
rect 18420 9460 18472 9512
rect 18512 9460 18564 9512
rect 19248 9460 19300 9512
rect 18328 9392 18380 9444
rect 20076 9460 20128 9512
rect 22284 9460 22336 9512
rect 21824 9392 21876 9444
rect 22008 9392 22060 9444
rect 23756 9503 23808 9512
rect 23756 9469 23765 9503
rect 23765 9469 23799 9503
rect 23799 9469 23808 9503
rect 23756 9460 23808 9469
rect 24308 9460 24360 9512
rect 28448 9596 28500 9648
rect 29276 9528 29328 9580
rect 30012 9664 30064 9716
rect 32404 9664 32456 9716
rect 32864 9664 32916 9716
rect 34244 9664 34296 9716
rect 29644 9596 29696 9648
rect 30472 9528 30524 9580
rect 26608 9460 26660 9512
rect 27252 9503 27304 9512
rect 27252 9469 27261 9503
rect 27261 9469 27295 9503
rect 27295 9469 27304 9503
rect 27252 9460 27304 9469
rect 30564 9460 30616 9512
rect 31392 9571 31444 9580
rect 31392 9537 31401 9571
rect 31401 9537 31435 9571
rect 31435 9537 31444 9571
rect 31392 9528 31444 9537
rect 31760 9460 31812 9512
rect 32588 9639 32640 9648
rect 32588 9605 32597 9639
rect 32597 9605 32631 9639
rect 32631 9605 32640 9639
rect 32588 9596 32640 9605
rect 33324 9596 33376 9648
rect 34796 9596 34848 9648
rect 35072 9596 35124 9648
rect 36452 9639 36504 9648
rect 36452 9605 36461 9639
rect 36461 9605 36495 9639
rect 36495 9605 36504 9639
rect 36452 9596 36504 9605
rect 37004 9664 37056 9716
rect 37832 9664 37884 9716
rect 38660 9664 38712 9716
rect 32312 9571 32364 9580
rect 32312 9537 32321 9571
rect 32321 9537 32355 9571
rect 32355 9537 32364 9571
rect 32312 9528 32364 9537
rect 33876 9528 33928 9580
rect 33784 9460 33836 9512
rect 29276 9392 29328 9444
rect 29828 9392 29880 9444
rect 11704 9367 11756 9376
rect 11704 9333 11713 9367
rect 11713 9333 11747 9367
rect 11747 9333 11756 9367
rect 11704 9324 11756 9333
rect 14556 9324 14608 9376
rect 15292 9324 15344 9376
rect 15384 9324 15436 9376
rect 17776 9324 17828 9376
rect 18236 9324 18288 9376
rect 19708 9324 19760 9376
rect 22100 9324 22152 9376
rect 22376 9324 22428 9376
rect 22652 9324 22704 9376
rect 28724 9324 28776 9376
rect 28816 9324 28868 9376
rect 33968 9324 34020 9376
rect 34244 9324 34296 9376
rect 34888 9571 34940 9580
rect 34888 9537 34897 9571
rect 34897 9537 34931 9571
rect 34931 9537 34940 9571
rect 34888 9528 34940 9537
rect 34428 9460 34480 9512
rect 35900 9528 35952 9580
rect 36360 9571 36412 9580
rect 36360 9537 36369 9571
rect 36369 9537 36403 9571
rect 36403 9537 36412 9571
rect 36360 9528 36412 9537
rect 35072 9503 35124 9512
rect 35072 9469 35081 9503
rect 35081 9469 35115 9503
rect 35115 9469 35124 9503
rect 35072 9460 35124 9469
rect 35532 9503 35584 9512
rect 35532 9469 35541 9503
rect 35541 9469 35575 9503
rect 35575 9469 35584 9503
rect 35532 9460 35584 9469
rect 36636 9528 36688 9580
rect 37188 9596 37240 9648
rect 39120 9596 39172 9648
rect 37280 9528 37332 9580
rect 37832 9528 37884 9580
rect 38568 9571 38620 9580
rect 38568 9537 38577 9571
rect 38577 9537 38611 9571
rect 38611 9537 38620 9571
rect 38568 9528 38620 9537
rect 38936 9528 38988 9580
rect 40132 9664 40184 9716
rect 39856 9596 39908 9648
rect 39764 9571 39816 9580
rect 39764 9537 39773 9571
rect 39773 9537 39807 9571
rect 39807 9537 39816 9571
rect 39764 9528 39816 9537
rect 40592 9571 40644 9580
rect 35716 9392 35768 9444
rect 37556 9392 37608 9444
rect 35992 9367 36044 9376
rect 35992 9333 36001 9367
rect 36001 9333 36035 9367
rect 36035 9333 36044 9367
rect 35992 9324 36044 9333
rect 37004 9367 37056 9376
rect 37004 9333 37013 9367
rect 37013 9333 37047 9367
rect 37047 9333 37056 9367
rect 37004 9324 37056 9333
rect 37280 9324 37332 9376
rect 38476 9392 38528 9444
rect 38660 9392 38712 9444
rect 40592 9537 40601 9571
rect 40601 9537 40635 9571
rect 40635 9537 40644 9571
rect 40592 9528 40644 9537
rect 39948 9460 40000 9512
rect 41236 9503 41288 9512
rect 41236 9469 41245 9503
rect 41245 9469 41279 9503
rect 41279 9469 41288 9503
rect 41236 9460 41288 9469
rect 41420 9528 41472 9580
rect 42892 9571 42944 9580
rect 42892 9537 42901 9571
rect 42901 9537 42935 9571
rect 42935 9537 42944 9571
rect 42892 9528 42944 9537
rect 43260 9528 43312 9580
rect 43720 9528 43772 9580
rect 44548 9596 44600 9648
rect 47216 9596 47268 9648
rect 47860 9596 47912 9648
rect 49424 9596 49476 9648
rect 45100 9528 45152 9580
rect 45744 9528 45796 9580
rect 46480 9528 46532 9580
rect 42524 9460 42576 9512
rect 42616 9503 42668 9512
rect 42616 9469 42625 9503
rect 42625 9469 42659 9503
rect 42659 9469 42668 9503
rect 42616 9460 42668 9469
rect 42708 9460 42760 9512
rect 43904 9503 43956 9512
rect 43904 9469 43913 9503
rect 43913 9469 43947 9503
rect 43947 9469 43956 9503
rect 43904 9460 43956 9469
rect 45192 9503 45244 9512
rect 45192 9469 45201 9503
rect 45201 9469 45235 9503
rect 45235 9469 45244 9503
rect 45192 9460 45244 9469
rect 47492 9392 47544 9444
rect 38936 9324 38988 9376
rect 39856 9367 39908 9376
rect 39856 9333 39865 9367
rect 39865 9333 39899 9367
rect 39899 9333 39908 9367
rect 39856 9324 39908 9333
rect 47124 9324 47176 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 3608 9163 3660 9172
rect 3608 9129 3617 9163
rect 3617 9129 3651 9163
rect 3651 9129 3660 9163
rect 3608 9120 3660 9129
rect 8484 9120 8536 9172
rect 10324 9163 10376 9172
rect 10324 9129 10333 9163
rect 10333 9129 10367 9163
rect 10367 9129 10376 9163
rect 10324 9120 10376 9129
rect 10600 9120 10652 9172
rect 12256 9120 12308 9172
rect 13728 9120 13780 9172
rect 15292 9120 15344 9172
rect 15476 9120 15528 9172
rect 2228 8984 2280 9036
rect 8024 9052 8076 9104
rect 7288 8984 7340 9036
rect 7748 9027 7800 9036
rect 7748 8993 7757 9027
rect 7757 8993 7791 9027
rect 7791 8993 7800 9027
rect 7748 8984 7800 8993
rect 1308 8916 1360 8968
rect 1216 8848 1268 8900
rect 3424 8916 3476 8968
rect 7656 8916 7708 8968
rect 8392 8848 8444 8900
rect 1768 8823 1820 8832
rect 1768 8789 1777 8823
rect 1777 8789 1811 8823
rect 1811 8789 1820 8823
rect 1768 8780 1820 8789
rect 4344 8780 4396 8832
rect 5356 8780 5408 8832
rect 16028 9052 16080 9104
rect 8576 8984 8628 9036
rect 9680 8959 9732 8968
rect 9680 8925 9689 8959
rect 9689 8925 9723 8959
rect 9723 8925 9732 8959
rect 9680 8916 9732 8925
rect 13452 9027 13504 9036
rect 13452 8993 13461 9027
rect 13461 8993 13495 9027
rect 13495 8993 13504 9027
rect 13452 8984 13504 8993
rect 13636 9027 13688 9036
rect 13636 8993 13645 9027
rect 13645 8993 13679 9027
rect 13679 8993 13688 9027
rect 13636 8984 13688 8993
rect 14924 8984 14976 9036
rect 15568 9027 15620 9036
rect 15568 8993 15577 9027
rect 15577 8993 15611 9027
rect 15611 8993 15620 9027
rect 15568 8984 15620 8993
rect 16212 9027 16264 9036
rect 16212 8993 16221 9027
rect 16221 8993 16255 9027
rect 16255 8993 16264 9027
rect 16212 8984 16264 8993
rect 17684 9120 17736 9172
rect 19432 9120 19484 9172
rect 18696 9095 18748 9104
rect 18696 9061 18705 9095
rect 18705 9061 18739 9095
rect 18739 9061 18748 9095
rect 18696 9052 18748 9061
rect 20812 9120 20864 9172
rect 22284 9120 22336 9172
rect 25136 9120 25188 9172
rect 34888 9120 34940 9172
rect 13268 8916 13320 8968
rect 15108 8916 15160 8968
rect 15384 8959 15436 8968
rect 15384 8925 15393 8959
rect 15393 8925 15427 8959
rect 15427 8925 15436 8959
rect 15384 8916 15436 8925
rect 8852 8848 8904 8900
rect 11704 8848 11756 8900
rect 8576 8780 8628 8832
rect 11612 8780 11664 8832
rect 13636 8848 13688 8900
rect 15200 8848 15252 8900
rect 16948 8848 17000 8900
rect 13176 8780 13228 8832
rect 13452 8780 13504 8832
rect 14924 8780 14976 8832
rect 15016 8823 15068 8832
rect 15016 8789 15025 8823
rect 15025 8789 15059 8823
rect 15059 8789 15068 8823
rect 15016 8780 15068 8789
rect 18512 8916 18564 8968
rect 18696 8916 18748 8968
rect 25964 9052 26016 9104
rect 28540 9052 28592 9104
rect 28816 9052 28868 9104
rect 31300 9052 31352 9104
rect 19248 8984 19300 9036
rect 21824 8984 21876 9036
rect 23480 8984 23532 9036
rect 27620 8984 27672 9036
rect 28724 9027 28776 9036
rect 28724 8993 28733 9027
rect 28733 8993 28767 9027
rect 28767 8993 28776 9027
rect 28724 8984 28776 8993
rect 28908 9027 28960 9036
rect 28908 8993 28917 9027
rect 28917 8993 28951 9027
rect 28951 8993 28960 9027
rect 28908 8984 28960 8993
rect 30748 8984 30800 9036
rect 19708 8959 19760 8968
rect 19708 8925 19717 8959
rect 19717 8925 19751 8959
rect 19751 8925 19760 8959
rect 19708 8916 19760 8925
rect 24492 8916 24544 8968
rect 25044 8916 25096 8968
rect 27068 8959 27120 8968
rect 27068 8925 27077 8959
rect 27077 8925 27111 8959
rect 27111 8925 27120 8959
rect 27068 8916 27120 8925
rect 28448 8916 28500 8968
rect 29736 8959 29788 8968
rect 29736 8925 29745 8959
rect 29745 8925 29779 8959
rect 29779 8925 29788 8959
rect 29736 8916 29788 8925
rect 31484 8916 31536 8968
rect 31944 9027 31996 9036
rect 31944 8993 31953 9027
rect 31953 8993 31987 9027
rect 31987 8993 31996 9027
rect 31944 8984 31996 8993
rect 33692 9095 33744 9104
rect 33692 9061 33701 9095
rect 33701 9061 33735 9095
rect 33735 9061 33744 9095
rect 33692 9052 33744 9061
rect 34704 9052 34756 9104
rect 35256 9052 35308 9104
rect 34152 9027 34204 9036
rect 34152 8993 34161 9027
rect 34161 8993 34195 9027
rect 34195 8993 34204 9027
rect 34152 8984 34204 8993
rect 35164 8984 35216 9036
rect 36544 9120 36596 9172
rect 37188 9120 37240 9172
rect 38568 9120 38620 9172
rect 38844 9120 38896 9172
rect 39764 9120 39816 9172
rect 43812 9163 43864 9172
rect 43812 9129 43821 9163
rect 43821 9129 43855 9163
rect 43855 9129 43864 9163
rect 43812 9120 43864 9129
rect 45008 9120 45060 9172
rect 45928 9120 45980 9172
rect 47584 9120 47636 9172
rect 35624 9052 35676 9104
rect 36636 9052 36688 9104
rect 37372 9052 37424 9104
rect 38384 9052 38436 9104
rect 38936 9052 38988 9104
rect 39856 9052 39908 9104
rect 35532 8984 35584 9036
rect 39120 8984 39172 9036
rect 40868 8984 40920 9036
rect 42432 8984 42484 9036
rect 33324 8916 33376 8968
rect 33508 8916 33560 8968
rect 35624 8916 35676 8968
rect 35808 8916 35860 8968
rect 36084 8959 36136 8968
rect 36084 8925 36093 8959
rect 36093 8925 36127 8959
rect 36127 8925 36136 8959
rect 36084 8916 36136 8925
rect 36452 8916 36504 8968
rect 18604 8848 18656 8900
rect 18512 8780 18564 8832
rect 20536 8848 20588 8900
rect 20720 8848 20772 8900
rect 22928 8848 22980 8900
rect 27252 8848 27304 8900
rect 32220 8891 32272 8900
rect 32220 8857 32229 8891
rect 32229 8857 32263 8891
rect 32263 8857 32272 8891
rect 32220 8848 32272 8857
rect 34244 8848 34296 8900
rect 37556 8916 37608 8968
rect 41972 8916 42024 8968
rect 43536 8959 43588 8968
rect 43536 8925 43545 8959
rect 43545 8925 43579 8959
rect 43579 8925 43588 8959
rect 43536 8916 43588 8925
rect 44088 8916 44140 8968
rect 44548 8984 44600 9036
rect 46756 8916 46808 8968
rect 49240 8984 49292 9036
rect 24216 8780 24268 8832
rect 24492 8780 24544 8832
rect 25964 8780 26016 8832
rect 34980 8780 35032 8832
rect 35256 8780 35308 8832
rect 37648 8780 37700 8832
rect 38476 8823 38528 8832
rect 38476 8789 38485 8823
rect 38485 8789 38519 8823
rect 38519 8789 38528 8823
rect 38476 8780 38528 8789
rect 38936 8848 38988 8900
rect 39304 8891 39356 8900
rect 39304 8857 39313 8891
rect 39313 8857 39347 8891
rect 39347 8857 39356 8891
rect 39304 8848 39356 8857
rect 39580 8848 39632 8900
rect 40316 8891 40368 8900
rect 40316 8857 40325 8891
rect 40325 8857 40359 8891
rect 40359 8857 40368 8891
rect 40316 8848 40368 8857
rect 47860 8848 47912 8900
rect 41972 8780 42024 8832
rect 43720 8780 43772 8832
rect 43904 8780 43956 8832
rect 48320 8780 48372 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 1308 8576 1360 8628
rect 5632 8576 5684 8628
rect 7564 8576 7616 8628
rect 1216 8508 1268 8560
rect 6000 8508 6052 8560
rect 1584 8415 1636 8424
rect 1584 8381 1593 8415
rect 1593 8381 1627 8415
rect 1627 8381 1636 8415
rect 1584 8372 1636 8381
rect 2872 8372 2924 8424
rect 3148 8483 3200 8492
rect 3148 8449 3157 8483
rect 3157 8449 3191 8483
rect 3191 8449 3200 8483
rect 3148 8440 3200 8449
rect 10140 8508 10192 8560
rect 8576 8372 8628 8424
rect 9404 8483 9456 8492
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 9404 8440 9456 8449
rect 13544 8576 13596 8628
rect 14004 8576 14056 8628
rect 14188 8576 14240 8628
rect 14372 8576 14424 8628
rect 15568 8576 15620 8628
rect 16396 8576 16448 8628
rect 18144 8576 18196 8628
rect 18236 8576 18288 8628
rect 18788 8576 18840 8628
rect 18328 8508 18380 8560
rect 19892 8576 19944 8628
rect 20904 8576 20956 8628
rect 2780 8347 2832 8356
rect 2780 8313 2789 8347
rect 2789 8313 2823 8347
rect 2823 8313 2832 8347
rect 2780 8304 2832 8313
rect 3332 8304 3384 8356
rect 11520 8372 11572 8424
rect 11612 8415 11664 8424
rect 11612 8381 11621 8415
rect 11621 8381 11655 8415
rect 11655 8381 11664 8415
rect 11612 8372 11664 8381
rect 12716 8372 12768 8424
rect 13728 8372 13780 8424
rect 14556 8483 14608 8492
rect 14556 8449 14565 8483
rect 14565 8449 14599 8483
rect 14599 8449 14608 8483
rect 14556 8440 14608 8449
rect 15568 8372 15620 8424
rect 15844 8440 15896 8492
rect 18052 8440 18104 8492
rect 20720 8508 20772 8560
rect 22928 8576 22980 8628
rect 24400 8576 24452 8628
rect 24768 8576 24820 8628
rect 29000 8576 29052 8628
rect 23848 8508 23900 8560
rect 32496 8576 32548 8628
rect 32864 8576 32916 8628
rect 33968 8619 34020 8628
rect 33968 8585 33977 8619
rect 33977 8585 34011 8619
rect 34011 8585 34020 8619
rect 33968 8576 34020 8585
rect 34060 8619 34112 8628
rect 34060 8585 34069 8619
rect 34069 8585 34103 8619
rect 34103 8585 34112 8619
rect 34060 8576 34112 8585
rect 36360 8576 36412 8628
rect 38292 8576 38344 8628
rect 38384 8576 38436 8628
rect 39028 8619 39080 8628
rect 39028 8585 39037 8619
rect 39037 8585 39071 8619
rect 39071 8585 39080 8619
rect 39028 8576 39080 8585
rect 39580 8576 39632 8628
rect 23572 8440 23624 8492
rect 24400 8440 24452 8492
rect 24492 8483 24544 8492
rect 24492 8449 24501 8483
rect 24501 8449 24535 8483
rect 24535 8449 24544 8483
rect 24492 8440 24544 8449
rect 25964 8483 26016 8492
rect 25964 8449 25973 8483
rect 25973 8449 26007 8483
rect 26007 8449 26016 8483
rect 25964 8440 26016 8449
rect 26608 8440 26660 8492
rect 29828 8440 29880 8492
rect 31392 8483 31444 8492
rect 31392 8449 31401 8483
rect 31401 8449 31435 8483
rect 31435 8449 31444 8483
rect 31392 8440 31444 8449
rect 35348 8551 35400 8560
rect 35348 8517 35357 8551
rect 35357 8517 35391 8551
rect 35391 8517 35400 8551
rect 35348 8508 35400 8517
rect 36636 8508 36688 8560
rect 38016 8508 38068 8560
rect 38936 8508 38988 8560
rect 32680 8440 32732 8492
rect 11980 8304 12032 8356
rect 13176 8304 13228 8356
rect 12808 8236 12860 8288
rect 16488 8304 16540 8356
rect 17592 8415 17644 8424
rect 17592 8381 17601 8415
rect 17601 8381 17635 8415
rect 17635 8381 17644 8415
rect 17592 8372 17644 8381
rect 17960 8372 18012 8424
rect 18236 8304 18288 8356
rect 17408 8236 17460 8288
rect 17776 8236 17828 8288
rect 18420 8236 18472 8288
rect 19248 8372 19300 8424
rect 20444 8372 20496 8424
rect 21824 8372 21876 8424
rect 20812 8304 20864 8356
rect 28448 8415 28500 8424
rect 28448 8381 28457 8415
rect 28457 8381 28491 8415
rect 28491 8381 28500 8415
rect 28448 8372 28500 8381
rect 30288 8372 30340 8424
rect 31760 8372 31812 8424
rect 32128 8372 32180 8424
rect 32864 8415 32916 8424
rect 32864 8381 32873 8415
rect 32873 8381 32907 8415
rect 32907 8381 32916 8415
rect 32864 8372 32916 8381
rect 33048 8415 33100 8424
rect 33048 8381 33057 8415
rect 33057 8381 33091 8415
rect 33091 8381 33100 8415
rect 33048 8372 33100 8381
rect 34244 8415 34296 8424
rect 34244 8381 34253 8415
rect 34253 8381 34287 8415
rect 34287 8381 34296 8415
rect 34244 8372 34296 8381
rect 35440 8372 35492 8424
rect 36268 8440 36320 8492
rect 37464 8483 37516 8492
rect 37464 8449 37473 8483
rect 37473 8449 37507 8483
rect 37507 8449 37516 8483
rect 37464 8440 37516 8449
rect 40040 8508 40092 8560
rect 41236 8508 41288 8560
rect 42340 8576 42392 8628
rect 44180 8576 44232 8628
rect 43812 8508 43864 8560
rect 43996 8508 44048 8560
rect 45376 8551 45428 8560
rect 45376 8517 45385 8551
rect 45385 8517 45419 8551
rect 45419 8517 45428 8551
rect 45376 8508 45428 8517
rect 22008 8236 22060 8288
rect 23480 8236 23532 8288
rect 27988 8279 28040 8288
rect 27988 8245 27997 8279
rect 27997 8245 28031 8279
rect 28031 8245 28040 8279
rect 27988 8236 28040 8245
rect 35808 8304 35860 8356
rect 37832 8372 37884 8424
rect 37464 8304 37516 8356
rect 38016 8304 38068 8356
rect 39120 8372 39172 8424
rect 39488 8372 39540 8424
rect 40868 8372 40920 8424
rect 42156 8440 42208 8492
rect 44180 8483 44232 8492
rect 44180 8449 44189 8483
rect 44189 8449 44223 8483
rect 44223 8449 44232 8483
rect 44180 8440 44232 8449
rect 47768 8508 47820 8560
rect 49148 8551 49200 8560
rect 49148 8517 49157 8551
rect 49157 8517 49191 8551
rect 49191 8517 49200 8551
rect 49148 8508 49200 8517
rect 42524 8372 42576 8424
rect 42708 8372 42760 8424
rect 43444 8415 43496 8424
rect 43444 8381 43453 8415
rect 43453 8381 43487 8415
rect 43487 8381 43496 8415
rect 43444 8372 43496 8381
rect 38936 8304 38988 8356
rect 41328 8304 41380 8356
rect 42064 8304 42116 8356
rect 47860 8440 47912 8492
rect 46848 8415 46900 8424
rect 46848 8381 46857 8415
rect 46857 8381 46891 8415
rect 46891 8381 46900 8415
rect 46848 8372 46900 8381
rect 34888 8236 34940 8288
rect 35900 8236 35952 8288
rect 39948 8236 40000 8288
rect 41420 8236 41472 8288
rect 46388 8304 46440 8356
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 2136 8075 2188 8084
rect 2136 8041 2145 8075
rect 2145 8041 2179 8075
rect 2179 8041 2188 8075
rect 2136 8032 2188 8041
rect 8392 8075 8444 8084
rect 8392 8041 8401 8075
rect 8401 8041 8435 8075
rect 8435 8041 8444 8075
rect 8392 8032 8444 8041
rect 9772 8032 9824 8084
rect 11428 8032 11480 8084
rect 10048 7939 10100 7948
rect 10048 7905 10057 7939
rect 10057 7905 10091 7939
rect 10091 7905 10100 7939
rect 10048 7896 10100 7905
rect 11152 7896 11204 7948
rect 14740 8032 14792 8084
rect 17960 8032 18012 8084
rect 18420 8032 18472 8084
rect 19248 8032 19300 8084
rect 21456 8032 21508 8084
rect 22192 8032 22244 8084
rect 1308 7828 1360 7880
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 10232 7828 10284 7880
rect 11336 7828 11388 7880
rect 15200 7964 15252 8016
rect 17776 7964 17828 8016
rect 21180 7964 21232 8016
rect 23756 8032 23808 8084
rect 24400 8075 24452 8084
rect 24400 8041 24409 8075
rect 24409 8041 24443 8075
rect 24443 8041 24452 8075
rect 24400 8032 24452 8041
rect 27068 8032 27120 8084
rect 27804 8032 27856 8084
rect 28356 8032 28408 8084
rect 35900 8032 35952 8084
rect 35992 8032 36044 8084
rect 23848 7964 23900 8016
rect 27436 7964 27488 8016
rect 31116 7964 31168 8016
rect 12072 7896 12124 7948
rect 11980 7871 12032 7880
rect 11980 7837 11989 7871
rect 11989 7837 12023 7871
rect 12023 7837 12032 7871
rect 11980 7828 12032 7837
rect 22560 7896 22612 7948
rect 31760 7896 31812 7948
rect 15200 7871 15252 7880
rect 15200 7837 15209 7871
rect 15209 7837 15243 7871
rect 15243 7837 15252 7871
rect 15200 7828 15252 7837
rect 16304 7871 16356 7880
rect 16304 7837 16313 7871
rect 16313 7837 16347 7871
rect 16347 7837 16356 7871
rect 16304 7828 16356 7837
rect 7472 7692 7524 7744
rect 14188 7735 14240 7744
rect 14188 7701 14197 7735
rect 14197 7701 14231 7735
rect 14231 7701 14240 7735
rect 14188 7692 14240 7701
rect 16580 7803 16632 7812
rect 16580 7769 16589 7803
rect 16589 7769 16623 7803
rect 16623 7769 16632 7803
rect 16580 7760 16632 7769
rect 17040 7760 17092 7812
rect 18696 7760 18748 7812
rect 19616 7828 19668 7880
rect 21732 7871 21784 7880
rect 21732 7837 21741 7871
rect 21741 7837 21775 7871
rect 21775 7837 21784 7871
rect 21732 7828 21784 7837
rect 24952 7828 25004 7880
rect 25044 7871 25096 7880
rect 25044 7837 25053 7871
rect 25053 7837 25087 7871
rect 25087 7837 25096 7871
rect 25044 7828 25096 7837
rect 27988 7828 28040 7880
rect 29368 7828 29420 7880
rect 29460 7828 29512 7880
rect 30932 7828 30984 7880
rect 31576 7828 31628 7880
rect 32956 7828 33008 7880
rect 33324 7871 33376 7880
rect 33324 7837 33333 7871
rect 33333 7837 33367 7871
rect 33367 7837 33376 7871
rect 33324 7828 33376 7837
rect 34520 7828 34572 7880
rect 34888 7871 34940 7880
rect 34888 7837 34897 7871
rect 34897 7837 34931 7871
rect 34931 7837 34940 7871
rect 34888 7828 34940 7837
rect 35624 7896 35676 7948
rect 22008 7760 22060 7812
rect 19524 7692 19576 7744
rect 20260 7692 20312 7744
rect 22928 7735 22980 7744
rect 22928 7701 22937 7735
rect 22937 7701 22971 7735
rect 22971 7701 22980 7735
rect 22928 7692 22980 7701
rect 23296 7692 23348 7744
rect 30932 7692 30984 7744
rect 32864 7760 32916 7812
rect 36176 7760 36228 7812
rect 40592 8007 40644 8016
rect 40592 7973 40601 8007
rect 40601 7973 40635 8007
rect 40635 7973 40644 8007
rect 40592 7964 40644 7973
rect 40868 8007 40920 8016
rect 40868 7973 40877 8007
rect 40877 7973 40911 8007
rect 40911 7973 40920 8007
rect 40868 7964 40920 7973
rect 41052 8007 41104 8016
rect 41052 7973 41061 8007
rect 41061 7973 41095 8007
rect 41095 7973 41104 8007
rect 41052 7964 41104 7973
rect 41236 8007 41288 8016
rect 41236 7973 41245 8007
rect 41245 7973 41279 8007
rect 41279 7973 41288 8007
rect 41236 7964 41288 7973
rect 41696 8007 41748 8016
rect 41696 7973 41705 8007
rect 41705 7973 41739 8007
rect 41739 7973 41748 8007
rect 41696 7964 41748 7973
rect 41972 8007 42024 8016
rect 41972 7973 41981 8007
rect 41981 7973 42015 8007
rect 42015 7973 42024 8007
rect 41972 7964 42024 7973
rect 42156 8007 42208 8016
rect 42156 7973 42165 8007
rect 42165 7973 42199 8007
rect 42199 7973 42208 8007
rect 42156 7964 42208 7973
rect 43996 8007 44048 8016
rect 43996 7973 44005 8007
rect 44005 7973 44039 8007
rect 44039 7973 44048 8007
rect 43996 7964 44048 7973
rect 37832 7828 37884 7880
rect 40224 7828 40276 7880
rect 41052 7828 41104 7880
rect 39028 7760 39080 7812
rect 40132 7803 40184 7812
rect 40132 7769 40141 7803
rect 40141 7769 40175 7803
rect 40175 7769 40184 7803
rect 40132 7760 40184 7769
rect 42616 7760 42668 7812
rect 34428 7692 34480 7744
rect 37188 7735 37240 7744
rect 37188 7701 37197 7735
rect 37197 7701 37231 7735
rect 37231 7701 37240 7735
rect 37188 7692 37240 7701
rect 39212 7692 39264 7744
rect 41512 7735 41564 7744
rect 41512 7701 41521 7735
rect 41521 7701 41555 7735
rect 41555 7701 41564 7735
rect 41512 7692 41564 7701
rect 42892 7871 42944 7880
rect 42892 7837 42901 7871
rect 42901 7837 42935 7871
rect 42935 7837 42944 7871
rect 42892 7828 42944 7837
rect 43536 7871 43588 7880
rect 43536 7837 43545 7871
rect 43545 7837 43579 7871
rect 43579 7837 43588 7871
rect 43536 7828 43588 7837
rect 44640 8032 44692 8084
rect 45192 8075 45244 8084
rect 45192 8041 45201 8075
rect 45201 8041 45235 8075
rect 45235 8041 45244 8075
rect 45192 8032 45244 8041
rect 47032 8032 47084 8084
rect 44916 7964 44968 8016
rect 44548 7939 44600 7948
rect 44548 7905 44557 7939
rect 44557 7905 44591 7939
rect 44591 7905 44600 7939
rect 44548 7896 44600 7905
rect 45376 7896 45428 7948
rect 49056 7896 49108 7948
rect 49240 7896 49292 7948
rect 43720 7760 43772 7812
rect 47124 7828 47176 7880
rect 48320 7760 48372 7812
rect 49976 7760 50028 7812
rect 43168 7692 43220 7744
rect 43352 7735 43404 7744
rect 43352 7701 43361 7735
rect 43361 7701 43395 7735
rect 43395 7701 43404 7735
rect 43352 7692 43404 7701
rect 44088 7692 44140 7744
rect 46388 7735 46440 7744
rect 46388 7701 46397 7735
rect 46397 7701 46431 7735
rect 46431 7701 46440 7735
rect 46388 7692 46440 7701
rect 46940 7692 46992 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 9220 7488 9272 7540
rect 11244 7488 11296 7540
rect 11336 7531 11388 7540
rect 11336 7497 11345 7531
rect 11345 7497 11379 7531
rect 11379 7497 11388 7531
rect 11336 7488 11388 7497
rect 6092 7420 6144 7472
rect 12532 7488 12584 7540
rect 14096 7531 14148 7540
rect 14096 7497 14105 7531
rect 14105 7497 14139 7531
rect 14139 7497 14148 7531
rect 14096 7488 14148 7497
rect 15200 7488 15252 7540
rect 16672 7531 16724 7540
rect 16672 7497 16681 7531
rect 16681 7497 16715 7531
rect 16715 7497 16724 7531
rect 16672 7488 16724 7497
rect 19984 7488 20036 7540
rect 27712 7488 27764 7540
rect 29368 7531 29420 7540
rect 29368 7497 29377 7531
rect 29377 7497 29411 7531
rect 29411 7497 29420 7531
rect 29368 7488 29420 7497
rect 31576 7531 31628 7540
rect 31576 7497 31585 7531
rect 31585 7497 31619 7531
rect 31619 7497 31628 7531
rect 31576 7488 31628 7497
rect 32588 7488 32640 7540
rect 34520 7531 34572 7540
rect 34520 7497 34529 7531
rect 34529 7497 34563 7531
rect 34563 7497 34572 7531
rect 34520 7488 34572 7497
rect 1308 7352 1360 7404
rect 9496 7352 9548 7404
rect 9956 7395 10008 7404
rect 9956 7361 9965 7395
rect 9965 7361 9999 7395
rect 9999 7361 10008 7395
rect 9956 7352 10008 7361
rect 11980 7395 12032 7404
rect 11980 7361 11989 7395
rect 11989 7361 12023 7395
rect 12023 7361 12032 7395
rect 11980 7352 12032 7361
rect 12716 7420 12768 7472
rect 15752 7420 15804 7472
rect 17408 7420 17460 7472
rect 17500 7420 17552 7472
rect 12808 7352 12860 7404
rect 15568 7352 15620 7404
rect 17592 7352 17644 7404
rect 18328 7352 18380 7404
rect 22192 7420 22244 7472
rect 37372 7488 37424 7540
rect 35808 7420 35860 7472
rect 19708 7395 19760 7404
rect 19708 7361 19717 7395
rect 19717 7361 19751 7395
rect 19751 7361 19760 7395
rect 19708 7352 19760 7361
rect 22652 7352 22704 7404
rect 22836 7352 22888 7404
rect 24676 7352 24728 7404
rect 25228 7352 25280 7404
rect 28356 7352 28408 7404
rect 10692 7284 10744 7336
rect 14832 7284 14884 7336
rect 16764 7284 16816 7336
rect 17868 7327 17920 7336
rect 17868 7293 17877 7327
rect 17877 7293 17911 7327
rect 17911 7293 17920 7327
rect 17868 7284 17920 7293
rect 18512 7284 18564 7336
rect 22928 7284 22980 7336
rect 29920 7352 29972 7404
rect 30932 7395 30984 7404
rect 30932 7361 30941 7395
rect 30941 7361 30975 7395
rect 30975 7361 30984 7395
rect 30932 7352 30984 7361
rect 32772 7352 32824 7404
rect 17684 7216 17736 7268
rect 35532 7352 35584 7404
rect 35716 7352 35768 7404
rect 37280 7284 37332 7336
rect 37740 7327 37792 7336
rect 37740 7293 37749 7327
rect 37749 7293 37783 7327
rect 37783 7293 37792 7327
rect 37740 7284 37792 7293
rect 38016 7395 38068 7404
rect 38016 7361 38025 7395
rect 38025 7361 38059 7395
rect 38059 7361 38068 7395
rect 40132 7420 40184 7472
rect 40776 7420 40828 7472
rect 43352 7420 43404 7472
rect 43536 7420 43588 7472
rect 44824 7420 44876 7472
rect 45284 7488 45336 7540
rect 50068 7488 50120 7540
rect 45008 7420 45060 7472
rect 49332 7420 49384 7472
rect 38016 7352 38068 7361
rect 42248 7352 42300 7404
rect 44364 7395 44416 7404
rect 44364 7361 44373 7395
rect 44373 7361 44407 7395
rect 44407 7361 44416 7395
rect 44364 7352 44416 7361
rect 40132 7284 40184 7336
rect 42800 7284 42852 7336
rect 35808 7216 35860 7268
rect 1768 7191 1820 7200
rect 1768 7157 1777 7191
rect 1777 7157 1811 7191
rect 1811 7157 1820 7191
rect 1768 7148 1820 7157
rect 18512 7191 18564 7200
rect 18512 7157 18521 7191
rect 18521 7157 18555 7191
rect 18555 7157 18564 7191
rect 18512 7148 18564 7157
rect 21456 7191 21508 7200
rect 21456 7157 21465 7191
rect 21465 7157 21499 7191
rect 21499 7157 21508 7191
rect 21456 7148 21508 7157
rect 21824 7191 21876 7200
rect 21824 7157 21833 7191
rect 21833 7157 21867 7191
rect 21867 7157 21876 7191
rect 21824 7148 21876 7157
rect 23388 7191 23440 7200
rect 23388 7157 23397 7191
rect 23397 7157 23431 7191
rect 23431 7157 23440 7191
rect 23388 7148 23440 7157
rect 24676 7148 24728 7200
rect 25228 7148 25280 7200
rect 34888 7148 34940 7200
rect 42984 7148 43036 7200
rect 43168 7148 43220 7200
rect 44180 7284 44232 7336
rect 44272 7284 44324 7336
rect 45928 7352 45980 7404
rect 46204 7395 46256 7404
rect 46204 7361 46213 7395
rect 46213 7361 46247 7395
rect 46247 7361 46256 7395
rect 46204 7352 46256 7361
rect 46296 7352 46348 7404
rect 47952 7395 48004 7404
rect 47952 7361 47961 7395
rect 47961 7361 47995 7395
rect 47995 7361 48004 7395
rect 47952 7352 48004 7361
rect 44640 7284 44692 7336
rect 47216 7284 47268 7336
rect 50068 7284 50120 7336
rect 50528 7284 50580 7336
rect 47860 7216 47912 7268
rect 44456 7148 44508 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 1768 6944 1820 6996
rect 9496 6987 9548 6996
rect 9496 6953 9505 6987
rect 9505 6953 9539 6987
rect 9539 6953 9548 6987
rect 9496 6944 9548 6953
rect 12716 6944 12768 6996
rect 15108 6944 15160 6996
rect 18420 6944 18472 6996
rect 39304 6944 39356 6996
rect 47952 6944 48004 6996
rect 1216 6740 1268 6792
rect 1308 6672 1360 6724
rect 11336 6783 11388 6792
rect 11336 6749 11345 6783
rect 11345 6749 11379 6783
rect 11379 6749 11388 6783
rect 11336 6740 11388 6749
rect 13728 6851 13780 6860
rect 13728 6817 13737 6851
rect 13737 6817 13771 6851
rect 13771 6817 13780 6851
rect 13728 6808 13780 6817
rect 16396 6876 16448 6928
rect 1768 6647 1820 6656
rect 1768 6613 1777 6647
rect 1777 6613 1811 6647
rect 1811 6613 1820 6647
rect 1768 6604 1820 6613
rect 8760 6672 8812 6724
rect 11796 6672 11848 6724
rect 15292 6783 15344 6792
rect 15292 6749 15301 6783
rect 15301 6749 15335 6783
rect 15335 6749 15344 6783
rect 15292 6740 15344 6749
rect 15568 6808 15620 6860
rect 16856 6808 16908 6860
rect 17132 6851 17184 6860
rect 17132 6817 17141 6851
rect 17141 6817 17175 6851
rect 17175 6817 17184 6851
rect 17132 6808 17184 6817
rect 31852 6876 31904 6928
rect 41788 6876 41840 6928
rect 42616 6876 42668 6928
rect 17684 6740 17736 6792
rect 17868 6808 17920 6860
rect 19156 6808 19208 6860
rect 22008 6851 22060 6860
rect 22008 6817 22017 6851
rect 22017 6817 22051 6851
rect 22051 6817 22060 6851
rect 22008 6808 22060 6817
rect 24032 6851 24084 6860
rect 24032 6817 24041 6851
rect 24041 6817 24075 6851
rect 24075 6817 24084 6851
rect 24032 6808 24084 6817
rect 25872 6851 25924 6860
rect 25872 6817 25881 6851
rect 25881 6817 25915 6851
rect 25915 6817 25924 6851
rect 25872 6808 25924 6817
rect 28356 6808 28408 6860
rect 32220 6808 32272 6860
rect 35624 6808 35676 6860
rect 43352 6808 43404 6860
rect 43628 6808 43680 6860
rect 43812 6851 43864 6860
rect 43812 6817 43821 6851
rect 43821 6817 43855 6851
rect 43855 6817 43864 6851
rect 43812 6808 43864 6817
rect 44824 6808 44876 6860
rect 18512 6740 18564 6792
rect 18880 6783 18932 6792
rect 18880 6749 18889 6783
rect 18889 6749 18923 6783
rect 18923 6749 18932 6783
rect 18880 6740 18932 6749
rect 20260 6783 20312 6792
rect 20260 6749 20269 6783
rect 20269 6749 20303 6783
rect 20303 6749 20312 6783
rect 20260 6740 20312 6749
rect 22468 6740 22520 6792
rect 23388 6783 23440 6792
rect 23388 6749 23397 6783
rect 23397 6749 23431 6783
rect 23431 6749 23440 6783
rect 23388 6740 23440 6749
rect 25228 6783 25280 6792
rect 25228 6749 25237 6783
rect 25237 6749 25271 6783
rect 25271 6749 25280 6783
rect 25228 6740 25280 6749
rect 12348 6647 12400 6656
rect 12348 6613 12357 6647
rect 12357 6613 12391 6647
rect 12391 6613 12400 6647
rect 12348 6604 12400 6613
rect 14096 6604 14148 6656
rect 14280 6647 14332 6656
rect 14280 6613 14289 6647
rect 14289 6613 14323 6647
rect 14323 6613 14332 6647
rect 14280 6604 14332 6613
rect 18788 6672 18840 6724
rect 19064 6672 19116 6724
rect 21456 6672 21508 6724
rect 28540 6740 28592 6792
rect 29276 6740 29328 6792
rect 30380 6740 30432 6792
rect 32312 6783 32364 6792
rect 32312 6749 32321 6783
rect 32321 6749 32355 6783
rect 32355 6749 32364 6783
rect 32312 6740 32364 6749
rect 33692 6740 33744 6792
rect 34888 6783 34940 6792
rect 34888 6749 34897 6783
rect 34897 6749 34931 6783
rect 34931 6749 34940 6783
rect 34888 6740 34940 6749
rect 43536 6783 43588 6792
rect 43536 6749 43545 6783
rect 43545 6749 43579 6783
rect 43579 6749 43588 6783
rect 43536 6740 43588 6749
rect 43996 6740 44048 6792
rect 46020 6808 46072 6860
rect 45284 6740 45336 6792
rect 45468 6740 45520 6792
rect 45928 6740 45980 6792
rect 46296 6808 46348 6860
rect 47768 6740 47820 6792
rect 49148 6851 49200 6860
rect 49148 6817 49157 6851
rect 49157 6817 49191 6851
rect 49191 6817 49200 6851
rect 49148 6808 49200 6817
rect 50344 6740 50396 6792
rect 30656 6672 30708 6724
rect 36084 6672 36136 6724
rect 37188 6672 37240 6724
rect 47124 6672 47176 6724
rect 48688 6672 48740 6724
rect 14556 6604 14608 6656
rect 14648 6604 14700 6656
rect 18328 6604 18380 6656
rect 26976 6647 27028 6656
rect 26976 6613 26985 6647
rect 26985 6613 27019 6647
rect 27019 6613 27028 6647
rect 26976 6604 27028 6613
rect 30288 6604 30340 6656
rect 30472 6604 30524 6656
rect 40316 6604 40368 6656
rect 43260 6604 43312 6656
rect 45008 6647 45060 6656
rect 45008 6613 45017 6647
rect 45017 6613 45051 6647
rect 45051 6613 45060 6647
rect 45008 6604 45060 6613
rect 45468 6647 45520 6656
rect 45468 6613 45477 6647
rect 45477 6613 45511 6647
rect 45511 6613 45520 6647
rect 45468 6604 45520 6613
rect 46020 6604 46072 6656
rect 46848 6604 46900 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 1216 6400 1268 6452
rect 9864 6400 9916 6452
rect 12624 6332 12676 6384
rect 1308 6264 1360 6316
rect 16580 6400 16632 6452
rect 17592 6400 17644 6452
rect 19340 6400 19392 6452
rect 19708 6400 19760 6452
rect 21916 6400 21968 6452
rect 24216 6443 24268 6452
rect 24216 6409 24225 6443
rect 24225 6409 24259 6443
rect 24259 6409 24268 6443
rect 24216 6400 24268 6409
rect 24952 6400 25004 6452
rect 29276 6443 29328 6452
rect 29276 6409 29285 6443
rect 29285 6409 29319 6443
rect 29319 6409 29328 6443
rect 29276 6400 29328 6409
rect 30564 6400 30616 6452
rect 30840 6400 30892 6452
rect 32312 6400 32364 6452
rect 33508 6400 33560 6452
rect 43996 6443 44048 6452
rect 43996 6409 44005 6443
rect 44005 6409 44039 6443
rect 44039 6409 44048 6443
rect 43996 6400 44048 6409
rect 44272 6400 44324 6452
rect 44364 6443 44416 6452
rect 44364 6409 44373 6443
rect 44373 6409 44407 6443
rect 44407 6409 44416 6443
rect 44364 6400 44416 6409
rect 44456 6400 44508 6452
rect 45652 6400 45704 6452
rect 46020 6443 46072 6452
rect 46020 6409 46029 6443
rect 46029 6409 46063 6443
rect 46063 6409 46072 6443
rect 46020 6400 46072 6409
rect 47216 6443 47268 6452
rect 47216 6409 47225 6443
rect 47225 6409 47259 6443
rect 47259 6409 47268 6443
rect 47216 6400 47268 6409
rect 50896 6400 50948 6452
rect 14924 6332 14976 6384
rect 14556 6264 14608 6316
rect 12348 6239 12400 6248
rect 12348 6205 12357 6239
rect 12357 6205 12391 6239
rect 12391 6205 12400 6239
rect 12348 6196 12400 6205
rect 13636 6196 13688 6248
rect 16488 6332 16540 6384
rect 15936 6264 15988 6316
rect 18512 6264 18564 6316
rect 18880 6264 18932 6316
rect 20996 6264 21048 6316
rect 26976 6332 27028 6384
rect 24676 6307 24728 6316
rect 24676 6273 24685 6307
rect 24685 6273 24719 6307
rect 24719 6273 24728 6307
rect 24676 6264 24728 6273
rect 28908 6264 28960 6316
rect 30472 6264 30524 6316
rect 32864 6332 32916 6384
rect 34336 6332 34388 6384
rect 43260 6332 43312 6384
rect 32036 6264 32088 6316
rect 40040 6264 40092 6316
rect 45468 6264 45520 6316
rect 46296 6264 46348 6316
rect 46848 6307 46900 6316
rect 46848 6273 46857 6307
rect 46857 6273 46891 6307
rect 46891 6273 46900 6307
rect 46848 6264 46900 6273
rect 47676 6307 47728 6316
rect 47676 6273 47685 6307
rect 47685 6273 47719 6307
rect 47719 6273 47728 6307
rect 47676 6264 47728 6273
rect 49240 6332 49292 6384
rect 20904 6196 20956 6248
rect 29092 6196 29144 6248
rect 9312 6128 9364 6180
rect 17776 6128 17828 6180
rect 38384 6239 38436 6248
rect 38384 6205 38393 6239
rect 38393 6205 38427 6239
rect 38427 6205 38436 6239
rect 38384 6196 38436 6205
rect 46940 6196 46992 6248
rect 42524 6128 42576 6180
rect 46388 6128 46440 6180
rect 46664 6171 46716 6180
rect 46664 6137 46673 6171
rect 46673 6137 46707 6171
rect 46707 6137 46716 6171
rect 46664 6128 46716 6137
rect 14924 6060 14976 6112
rect 19616 6060 19668 6112
rect 19708 6060 19760 6112
rect 25320 6060 25372 6112
rect 27528 6060 27580 6112
rect 41880 6060 41932 6112
rect 45100 6060 45152 6112
rect 45284 6060 45336 6112
rect 45468 6060 45520 6112
rect 50252 6060 50304 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 1768 5856 1820 5908
rect 14004 5788 14056 5840
rect 18880 5899 18932 5908
rect 18880 5865 18889 5899
rect 18889 5865 18923 5899
rect 18923 5865 18932 5899
rect 18880 5856 18932 5865
rect 20996 5899 21048 5908
rect 20996 5865 21005 5899
rect 21005 5865 21039 5899
rect 21039 5865 21048 5899
rect 20996 5856 21048 5865
rect 23480 5856 23532 5908
rect 30380 5899 30432 5908
rect 30380 5865 30389 5899
rect 30389 5865 30423 5899
rect 30423 5865 30432 5899
rect 30380 5856 30432 5865
rect 30748 5856 30800 5908
rect 44640 5899 44692 5908
rect 44640 5865 44649 5899
rect 44649 5865 44683 5899
rect 44683 5865 44692 5899
rect 44640 5856 44692 5865
rect 45192 5899 45244 5908
rect 45192 5865 45201 5899
rect 45201 5865 45235 5899
rect 45235 5865 45244 5899
rect 45192 5856 45244 5865
rect 45376 5899 45428 5908
rect 45376 5865 45385 5899
rect 45385 5865 45419 5899
rect 45419 5865 45428 5899
rect 45376 5856 45428 5865
rect 45560 5856 45612 5908
rect 29552 5788 29604 5840
rect 45468 5788 45520 5840
rect 45744 5831 45796 5840
rect 45744 5797 45753 5831
rect 45753 5797 45787 5831
rect 45787 5797 45796 5831
rect 45744 5788 45796 5797
rect 1308 5652 1360 5704
rect 15844 5763 15896 5772
rect 15844 5729 15853 5763
rect 15853 5729 15887 5763
rect 15887 5729 15896 5763
rect 15844 5720 15896 5729
rect 17316 5720 17368 5772
rect 18972 5720 19024 5772
rect 20536 5720 20588 5772
rect 31392 5720 31444 5772
rect 38384 5720 38436 5772
rect 45928 5720 45980 5772
rect 2780 5652 2832 5704
rect 17868 5652 17920 5704
rect 20168 5652 20220 5704
rect 20628 5652 20680 5704
rect 21640 5695 21692 5704
rect 21640 5661 21684 5695
rect 21684 5661 21692 5695
rect 21640 5652 21692 5661
rect 22284 5695 22336 5704
rect 22284 5661 22293 5695
rect 22293 5661 22327 5695
rect 22327 5661 22336 5695
rect 22284 5652 22336 5661
rect 23572 5652 23624 5704
rect 23664 5652 23716 5704
rect 31300 5652 31352 5704
rect 36452 5652 36504 5704
rect 38292 5652 38344 5704
rect 47032 5899 47084 5908
rect 47032 5865 47041 5899
rect 47041 5865 47075 5899
rect 47075 5865 47084 5899
rect 47032 5856 47084 5865
rect 47216 5856 47268 5908
rect 46572 5788 46624 5840
rect 50160 5856 50212 5908
rect 50436 5788 50488 5840
rect 23848 5584 23900 5636
rect 41512 5584 41564 5636
rect 45744 5584 45796 5636
rect 49332 5720 49384 5772
rect 46572 5695 46624 5704
rect 46572 5661 46581 5695
rect 46581 5661 46615 5695
rect 46615 5661 46624 5695
rect 46572 5652 46624 5661
rect 46940 5652 46992 5704
rect 46388 5584 46440 5636
rect 13820 5516 13872 5568
rect 18420 5516 18472 5568
rect 18512 5516 18564 5568
rect 22376 5516 22428 5568
rect 22928 5559 22980 5568
rect 22928 5525 22937 5559
rect 22937 5525 22971 5559
rect 22971 5525 22980 5559
rect 22928 5516 22980 5525
rect 48320 5516 48372 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 12164 5312 12216 5364
rect 23572 5355 23624 5364
rect 23572 5321 23581 5355
rect 23581 5321 23615 5355
rect 23615 5321 23624 5355
rect 23572 5312 23624 5321
rect 31484 5312 31536 5364
rect 15016 5244 15068 5296
rect 8944 5176 8996 5228
rect 17684 5244 17736 5296
rect 26148 5244 26200 5296
rect 37648 5312 37700 5364
rect 45560 5355 45612 5364
rect 45560 5321 45569 5355
rect 45569 5321 45603 5355
rect 45603 5321 45612 5355
rect 45560 5312 45612 5321
rect 45836 5312 45888 5364
rect 46940 5312 46992 5364
rect 49700 5312 49752 5364
rect 32680 5244 32732 5296
rect 49148 5287 49200 5296
rect 49148 5253 49157 5287
rect 49157 5253 49191 5287
rect 49191 5253 49200 5287
rect 49148 5244 49200 5253
rect 1308 5108 1360 5160
rect 17132 5151 17184 5160
rect 17132 5117 17141 5151
rect 17141 5117 17175 5151
rect 17175 5117 17184 5151
rect 17132 5108 17184 5117
rect 18420 5219 18472 5228
rect 18420 5185 18429 5219
rect 18429 5185 18463 5219
rect 18463 5185 18472 5219
rect 18420 5176 18472 5185
rect 20352 5176 20404 5228
rect 20812 5219 20864 5228
rect 20812 5185 20821 5219
rect 20821 5185 20855 5219
rect 20855 5185 20864 5219
rect 20812 5176 20864 5185
rect 22192 5176 22244 5228
rect 22928 5219 22980 5228
rect 22928 5185 22937 5219
rect 22937 5185 22971 5219
rect 22971 5185 22980 5219
rect 22928 5176 22980 5185
rect 23572 5176 23624 5228
rect 24676 5219 24728 5228
rect 24676 5185 24685 5219
rect 24685 5185 24719 5219
rect 24719 5185 24728 5219
rect 24676 5176 24728 5185
rect 38108 5219 38160 5228
rect 38108 5185 38117 5219
rect 38117 5185 38151 5219
rect 38151 5185 38160 5219
rect 38108 5176 38160 5185
rect 40132 5176 40184 5228
rect 47860 5176 47912 5228
rect 19248 5040 19300 5092
rect 24308 5108 24360 5160
rect 40408 5108 40460 5160
rect 48320 5108 48372 5160
rect 35900 5040 35952 5092
rect 44272 5040 44324 5092
rect 22008 4972 22060 5024
rect 24768 4972 24820 5024
rect 24860 4972 24912 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 1308 4768 1360 4820
rect 20168 4811 20220 4820
rect 20168 4777 20177 4811
rect 20177 4777 20211 4811
rect 20211 4777 20220 4811
rect 20168 4768 20220 4777
rect 20720 4768 20772 4820
rect 21088 4768 21140 4820
rect 20904 4700 20956 4752
rect 24676 4768 24728 4820
rect 45836 4811 45888 4820
rect 45836 4777 45845 4811
rect 45845 4777 45879 4811
rect 45879 4777 45888 4811
rect 45836 4768 45888 4777
rect 46204 4768 46256 4820
rect 46756 4811 46808 4820
rect 46756 4777 46765 4811
rect 46765 4777 46799 4811
rect 46799 4777 46808 4811
rect 46756 4768 46808 4777
rect 47308 4768 47360 4820
rect 47400 4768 47452 4820
rect 19156 4632 19208 4684
rect 20720 4632 20772 4684
rect 21824 4632 21876 4684
rect 23296 4632 23348 4684
rect 24768 4632 24820 4684
rect 46572 4700 46624 4752
rect 40224 4632 40276 4684
rect 1308 4496 1360 4548
rect 18788 4564 18840 4616
rect 20444 4564 20496 4616
rect 19708 4496 19760 4548
rect 21272 4539 21324 4548
rect 21272 4505 21281 4539
rect 21281 4505 21315 4539
rect 21315 4505 21324 4539
rect 21272 4496 21324 4505
rect 22100 4428 22152 4480
rect 24032 4564 24084 4616
rect 22836 4496 22888 4548
rect 25228 4607 25280 4616
rect 25228 4573 25237 4607
rect 25237 4573 25271 4607
rect 25271 4573 25280 4607
rect 25228 4564 25280 4573
rect 28632 4564 28684 4616
rect 46296 4607 46348 4616
rect 46296 4573 46305 4607
rect 46305 4573 46339 4607
rect 46339 4573 46348 4607
rect 46296 4564 46348 4573
rect 49424 4632 49476 4684
rect 22744 4471 22796 4480
rect 22744 4437 22753 4471
rect 22753 4437 22787 4471
rect 22787 4437 22796 4471
rect 22744 4428 22796 4437
rect 26148 4428 26200 4480
rect 27160 4428 27212 4480
rect 42800 4496 42852 4548
rect 48964 4496 49016 4548
rect 39396 4428 39448 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 21272 4224 21324 4276
rect 22100 4224 22152 4276
rect 24584 4224 24636 4276
rect 25228 4224 25280 4276
rect 32864 4224 32916 4276
rect 1308 4088 1360 4140
rect 1216 4020 1268 4072
rect 9864 4088 9916 4140
rect 17776 4088 17828 4140
rect 20076 4088 20128 4140
rect 22008 4131 22060 4140
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22008 4088 22060 4097
rect 23940 4088 23992 4140
rect 26148 4088 26200 4140
rect 27620 4156 27672 4208
rect 2136 3952 2188 4004
rect 2412 4020 2464 4072
rect 8300 3952 8352 4004
rect 9680 3884 9732 3936
rect 16212 4020 16264 4072
rect 20168 4020 20220 4072
rect 23664 4020 23716 4072
rect 20720 3952 20772 4004
rect 18512 3884 18564 3936
rect 22744 3884 22796 3936
rect 23388 3884 23440 3936
rect 23572 3927 23624 3936
rect 23572 3893 23581 3927
rect 23581 3893 23615 3927
rect 23615 3893 23624 3927
rect 23572 3884 23624 3893
rect 24308 4063 24360 4072
rect 24308 4029 24317 4063
rect 24317 4029 24351 4063
rect 24351 4029 24360 4063
rect 24308 4020 24360 4029
rect 24952 4063 25004 4072
rect 24952 4029 24961 4063
rect 24961 4029 24995 4063
rect 24995 4029 25004 4063
rect 24952 4020 25004 4029
rect 27620 4063 27672 4072
rect 27620 4029 27629 4063
rect 27629 4029 27663 4063
rect 27663 4029 27672 4063
rect 27620 4020 27672 4029
rect 39212 4020 39264 4072
rect 49240 4088 49292 4140
rect 46664 4063 46716 4072
rect 46664 4029 46673 4063
rect 46673 4029 46707 4063
rect 46707 4029 46716 4063
rect 46664 4020 46716 4029
rect 49792 4020 49844 4072
rect 34428 3952 34480 4004
rect 40500 3952 40552 4004
rect 45560 3952 45612 4004
rect 30840 3884 30892 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 11612 3680 11664 3732
rect 20076 3723 20128 3732
rect 20076 3689 20085 3723
rect 20085 3689 20119 3723
rect 20119 3689 20128 3723
rect 20076 3680 20128 3689
rect 3332 3612 3384 3664
rect 19156 3612 19208 3664
rect 24124 3680 24176 3732
rect 27620 3680 27672 3732
rect 33876 3680 33928 3732
rect 43444 3680 43496 3732
rect 20720 3612 20772 3664
rect 21640 3612 21692 3664
rect 24492 3612 24544 3664
rect 27528 3612 27580 3664
rect 36820 3612 36872 3664
rect 39672 3612 39724 3664
rect 49792 3612 49844 3664
rect 1308 3476 1360 3528
rect 1032 3408 1084 3460
rect 23296 3544 23348 3596
rect 24860 3587 24912 3596
rect 24860 3553 24869 3587
rect 24869 3553 24903 3587
rect 24903 3553 24912 3587
rect 24860 3544 24912 3553
rect 37096 3544 37148 3596
rect 47676 3544 47728 3596
rect 49148 3587 49200 3596
rect 49148 3553 49157 3587
rect 49157 3553 49191 3587
rect 49191 3553 49200 3587
rect 49148 3544 49200 3553
rect 9588 3519 9640 3528
rect 9588 3485 9597 3519
rect 9597 3485 9631 3519
rect 9631 3485 9640 3519
rect 9588 3476 9640 3485
rect 10048 3519 10100 3528
rect 10048 3485 10057 3519
rect 10057 3485 10091 3519
rect 10091 3485 10100 3519
rect 10048 3476 10100 3485
rect 11152 3519 11204 3528
rect 11152 3485 11161 3519
rect 11161 3485 11195 3519
rect 11195 3485 11204 3519
rect 11152 3476 11204 3485
rect 16212 3519 16264 3528
rect 16212 3485 16221 3519
rect 16221 3485 16255 3519
rect 16255 3485 16264 3519
rect 16212 3476 16264 3485
rect 5356 3340 5408 3392
rect 7472 3340 7524 3392
rect 8760 3383 8812 3392
rect 8760 3349 8769 3383
rect 8769 3349 8803 3383
rect 8803 3349 8812 3383
rect 8760 3340 8812 3349
rect 10508 3340 10560 3392
rect 10692 3383 10744 3392
rect 10692 3349 10701 3383
rect 10701 3349 10735 3383
rect 10735 3349 10744 3383
rect 10692 3340 10744 3349
rect 12348 3340 12400 3392
rect 12440 3340 12492 3392
rect 16396 3340 16448 3392
rect 17592 3519 17644 3528
rect 17592 3485 17601 3519
rect 17601 3485 17635 3519
rect 17635 3485 17644 3519
rect 17592 3476 17644 3485
rect 19524 3476 19576 3528
rect 23388 3519 23440 3528
rect 23388 3485 23397 3519
rect 23397 3485 23431 3519
rect 23431 3485 23440 3519
rect 23388 3476 23440 3485
rect 24032 3519 24084 3528
rect 24032 3485 24041 3519
rect 24041 3485 24075 3519
rect 24075 3485 24084 3519
rect 24032 3476 24084 3485
rect 18880 3408 18932 3460
rect 19524 3340 19576 3392
rect 24400 3408 24452 3460
rect 24584 3408 24636 3460
rect 40408 3476 40460 3528
rect 47124 3476 47176 3528
rect 30104 3408 30156 3460
rect 39212 3408 39264 3460
rect 48688 3408 48740 3460
rect 23572 3340 23624 3392
rect 26332 3383 26384 3392
rect 26332 3349 26341 3383
rect 26341 3349 26375 3383
rect 26375 3349 26384 3383
rect 26332 3340 26384 3349
rect 29092 3340 29144 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 1308 3136 1360 3188
rect 9588 3136 9640 3188
rect 11152 3179 11204 3188
rect 11152 3145 11161 3179
rect 11161 3145 11195 3179
rect 11195 3145 11204 3179
rect 11152 3136 11204 3145
rect 1308 3000 1360 3052
rect 10692 3068 10744 3120
rect 10508 3043 10560 3052
rect 10508 3009 10517 3043
rect 10517 3009 10551 3043
rect 10551 3009 10560 3043
rect 10508 3000 10560 3009
rect 12348 3043 12400 3052
rect 12348 3009 12357 3043
rect 12357 3009 12391 3043
rect 12391 3009 12400 3043
rect 12348 3000 12400 3009
rect 16304 3136 16356 3188
rect 17040 3136 17092 3188
rect 18880 3043 18932 3052
rect 18880 3009 18889 3043
rect 18889 3009 18923 3043
rect 18923 3009 18932 3043
rect 18880 3000 18932 3009
rect 9772 2932 9824 2984
rect 16488 2932 16540 2984
rect 2320 2839 2372 2848
rect 2320 2805 2329 2839
rect 2329 2805 2363 2839
rect 2363 2805 2372 2839
rect 2320 2796 2372 2805
rect 2780 2839 2832 2848
rect 2780 2805 2789 2839
rect 2789 2805 2823 2839
rect 2823 2805 2832 2839
rect 2780 2796 2832 2805
rect 7472 2864 7524 2916
rect 19800 3136 19852 3188
rect 19524 3111 19576 3120
rect 19524 3077 19533 3111
rect 19533 3077 19567 3111
rect 19567 3077 19576 3111
rect 19524 3068 19576 3077
rect 22100 3068 22152 3120
rect 22468 3068 22520 3120
rect 22652 3136 22704 3188
rect 22836 3136 22888 3188
rect 23296 3179 23348 3188
rect 23296 3145 23305 3179
rect 23305 3145 23339 3179
rect 23339 3145 23348 3179
rect 23296 3136 23348 3145
rect 23572 3068 23624 3120
rect 23940 3136 23992 3188
rect 24492 3136 24544 3188
rect 23848 3111 23900 3120
rect 23848 3077 23857 3111
rect 23857 3077 23891 3111
rect 23891 3077 23900 3111
rect 23848 3068 23900 3077
rect 29092 3111 29144 3120
rect 29092 3077 29101 3111
rect 29101 3077 29135 3111
rect 29135 3077 29144 3111
rect 29092 3068 29144 3077
rect 29828 3068 29880 3120
rect 49240 3068 49292 3120
rect 27528 3043 27580 3052
rect 27528 3009 27537 3043
rect 27537 3009 27571 3043
rect 27571 3009 27580 3043
rect 27528 3000 27580 3009
rect 28448 3000 28500 3052
rect 39396 3000 39448 3052
rect 45744 3000 45796 3052
rect 45928 3000 45980 3052
rect 19616 2932 19668 2984
rect 8852 2796 8904 2848
rect 10232 2796 10284 2848
rect 22284 2864 22336 2916
rect 23848 2932 23900 2984
rect 26056 2932 26108 2984
rect 24952 2864 25004 2916
rect 17592 2796 17644 2848
rect 46756 2932 46808 2984
rect 46848 2975 46900 2984
rect 46848 2941 46857 2975
rect 46857 2941 46891 2975
rect 46891 2941 46900 2975
rect 46848 2932 46900 2941
rect 38292 2796 38344 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 6368 2592 6420 2644
rect 9772 2635 9824 2644
rect 9772 2601 9781 2635
rect 9781 2601 9815 2635
rect 9815 2601 9824 2635
rect 9772 2592 9824 2601
rect 10048 2592 10100 2644
rect 24492 2635 24544 2644
rect 24492 2601 24501 2635
rect 24501 2601 24535 2635
rect 24535 2601 24544 2635
rect 24492 2592 24544 2601
rect 26332 2592 26384 2644
rect 30840 2635 30892 2644
rect 30840 2601 30849 2635
rect 30849 2601 30883 2635
rect 30883 2601 30892 2635
rect 30840 2592 30892 2601
rect 32864 2592 32916 2644
rect 34428 2592 34480 2644
rect 16028 2524 16080 2576
rect 1308 2388 1360 2440
rect 2780 2456 2832 2508
rect 9864 2456 9916 2508
rect 11704 2456 11756 2508
rect 13820 2456 13872 2508
rect 2320 2431 2372 2440
rect 2320 2397 2329 2431
rect 2329 2397 2363 2431
rect 2363 2397 2372 2431
rect 2320 2388 2372 2397
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 8760 2388 8812 2440
rect 9680 2388 9732 2440
rect 10232 2431 10284 2440
rect 10232 2397 10241 2431
rect 10241 2397 10275 2431
rect 10275 2397 10284 2431
rect 10232 2388 10284 2397
rect 12440 2388 12492 2440
rect 16396 2388 16448 2440
rect 20904 2456 20956 2508
rect 22468 2524 22520 2576
rect 22652 2456 22704 2508
rect 24952 2524 25004 2576
rect 30748 2524 30800 2576
rect 48872 2592 48924 2644
rect 36820 2456 36872 2508
rect 41328 2456 41380 2508
rect 44272 2456 44324 2508
rect 1216 2320 1268 2372
rect 6368 2320 6420 2372
rect 6920 2252 6972 2304
rect 14188 2252 14240 2304
rect 23940 2388 23992 2440
rect 27528 2388 27580 2440
rect 28632 2388 28684 2440
rect 30748 2388 30800 2440
rect 33140 2431 33192 2440
rect 33140 2397 33149 2431
rect 33149 2397 33183 2431
rect 33183 2397 33192 2431
rect 33140 2388 33192 2397
rect 34980 2388 35032 2440
rect 18328 2320 18380 2372
rect 26516 2320 26568 2372
rect 38292 2388 38344 2440
rect 42800 2388 42852 2440
rect 49148 2499 49200 2508
rect 49148 2465 49157 2499
rect 49157 2465 49191 2499
rect 49191 2465 49200 2499
rect 49148 2456 49200 2465
rect 48504 2320 48556 2372
rect 37096 2295 37148 2304
rect 37096 2261 37105 2295
rect 37105 2261 37139 2295
rect 37139 2261 37148 2295
rect 37096 2252 37148 2261
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
rect 8760 1708 8812 1760
rect 9588 1708 9640 1760
<< metal2 >>
rect 1582 26200 1638 27000
rect 2226 26200 2282 27000
rect 2870 26200 2926 27000
rect 3514 26200 3570 27000
rect 4158 26200 4214 27000
rect 4802 26330 4858 27000
rect 4802 26302 5120 26330
rect 4802 26200 4858 26302
rect 1596 22438 1624 26200
rect 1768 24608 1820 24614
rect 1768 24550 1820 24556
rect 1780 24410 1808 24550
rect 1768 24404 1820 24410
rect 1768 24346 1820 24352
rect 2136 24200 2188 24206
rect 2136 24142 2188 24148
rect 1768 23112 1820 23118
rect 1768 23054 1820 23060
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1308 22092 1360 22098
rect 1308 22034 1360 22040
rect 1320 20777 1348 22034
rect 1780 21865 1808 23054
rect 1952 22500 2004 22506
rect 1952 22442 2004 22448
rect 1766 21856 1822 21865
rect 1766 21791 1822 21800
rect 1306 20768 1362 20777
rect 1306 20703 1362 20712
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1216 17740 1268 17746
rect 1216 17682 1268 17688
rect 1228 17105 1256 17682
rect 1780 17338 1808 19314
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 1860 17196 1912 17202
rect 1860 17138 1912 17144
rect 1308 17128 1360 17134
rect 1214 17096 1270 17105
rect 1308 17070 1360 17076
rect 1214 17031 1270 17040
rect 1320 16697 1348 17070
rect 1306 16688 1362 16697
rect 1306 16623 1362 16632
rect 1308 16516 1360 16522
rect 1308 16458 1360 16464
rect 1320 16289 1348 16458
rect 1306 16280 1362 16289
rect 1306 16215 1362 16224
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 1320 15881 1348 15982
rect 1306 15872 1362 15881
rect 1306 15807 1362 15816
rect 1308 15564 1360 15570
rect 1308 15506 1360 15512
rect 1320 15473 1348 15506
rect 1306 15464 1362 15473
rect 1306 15399 1362 15408
rect 1780 15337 1808 16050
rect 1766 15328 1822 15337
rect 1766 15263 1822 15272
rect 1306 15056 1362 15065
rect 1306 14991 1362 15000
rect 1320 14958 1348 14991
rect 1308 14952 1360 14958
rect 1308 14894 1360 14900
rect 1306 14648 1362 14657
rect 1306 14583 1362 14592
rect 1320 14482 1348 14583
rect 1308 14476 1360 14482
rect 1308 14418 1360 14424
rect 1768 14272 1820 14278
rect 938 14240 994 14249
rect 1768 14214 1820 14220
rect 938 14175 994 14184
rect 952 13870 980 14175
rect 1780 13938 1808 14214
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 940 13864 992 13870
rect 940 13806 992 13812
rect 1766 13288 1822 13297
rect 1766 13223 1822 13232
rect 1306 13016 1362 13025
rect 1306 12951 1362 12960
rect 1320 12850 1348 12951
rect 1308 12844 1360 12850
rect 1308 12786 1360 12792
rect 1306 12200 1362 12209
rect 1306 12135 1362 12144
rect 1320 11762 1348 12135
rect 1780 11898 1808 13223
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 1872 11762 1900 17138
rect 1964 14550 1992 22442
rect 2044 19304 2096 19310
rect 2044 19246 2096 19252
rect 2056 18329 2084 19246
rect 2042 18320 2098 18329
rect 2042 18255 2098 18264
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 2056 17513 2084 18158
rect 2042 17504 2098 17513
rect 2042 17439 2098 17448
rect 2044 16992 2096 16998
rect 2044 16934 2096 16940
rect 1952 14544 2004 14550
rect 1952 14486 2004 14492
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1308 11756 1360 11762
rect 1308 11698 1360 11704
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1306 10976 1362 10985
rect 1596 10962 1624 11086
rect 1964 11014 1992 14350
rect 2056 12850 2084 16934
rect 2148 13462 2176 24142
rect 2240 22234 2268 26200
rect 2778 24440 2834 24449
rect 2320 24404 2372 24410
rect 2778 24375 2834 24384
rect 2320 24346 2372 24352
rect 2332 23866 2360 24346
rect 2412 24200 2464 24206
rect 2412 24142 2464 24148
rect 2320 23860 2372 23866
rect 2320 23802 2372 23808
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 2320 19236 2372 19242
rect 2320 19178 2372 19184
rect 2228 14544 2280 14550
rect 2228 14486 2280 14492
rect 2136 13456 2188 13462
rect 2136 13398 2188 13404
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1362 10934 1624 10962
rect 1952 11008 2004 11014
rect 1952 10950 2004 10956
rect 1306 10911 1362 10920
rect 1216 10668 1268 10674
rect 1216 10610 1268 10616
rect 1228 10577 1256 10610
rect 1308 10600 1360 10606
rect 1214 10568 1270 10577
rect 1308 10542 1360 10548
rect 1214 10503 1270 10512
rect 1320 10169 1348 10542
rect 1596 10266 1624 10934
rect 1766 10568 1822 10577
rect 1766 10503 1768 10512
rect 1820 10503 1822 10512
rect 1768 10474 1820 10480
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1306 10160 1362 10169
rect 1306 10095 1362 10104
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1596 9761 1624 9998
rect 1582 9752 1638 9761
rect 1582 9687 1638 9696
rect 1216 9580 1268 9586
rect 1216 9522 1268 9528
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 1228 9353 1256 9522
rect 1766 9480 1822 9489
rect 1766 9415 1768 9424
rect 1820 9415 1822 9424
rect 1768 9386 1820 9392
rect 1214 9344 1270 9353
rect 1214 9279 1270 9288
rect 1308 8968 1360 8974
rect 1306 8936 1308 8945
rect 1360 8936 1362 8945
rect 1216 8900 1268 8906
rect 1306 8871 1362 8880
rect 1766 8936 1822 8945
rect 1766 8871 1822 8880
rect 1216 8842 1268 8848
rect 1228 8566 1256 8842
rect 1320 8634 1348 8871
rect 1780 8838 1808 8871
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1308 8628 1360 8634
rect 1308 8570 1360 8576
rect 1216 8560 1268 8566
rect 1214 8528 1216 8537
rect 1268 8528 1270 8537
rect 1214 8463 1270 8472
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1596 8129 1624 8366
rect 1582 8120 1638 8129
rect 2148 8090 2176 9522
rect 2240 9042 2268 14486
rect 2332 12442 2360 19178
rect 2424 16574 2452 24142
rect 2792 23526 2820 24375
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 2884 23186 2912 26200
rect 3422 25664 3478 25673
rect 3422 25599 3478 25608
rect 3436 24886 3464 25599
rect 3424 24880 3476 24886
rect 3424 24822 3476 24828
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 3528 24274 3556 26200
rect 4066 25256 4122 25265
rect 4066 25191 4068 25200
rect 4120 25191 4122 25200
rect 4068 25162 4120 25168
rect 3698 24848 3754 24857
rect 3698 24783 3700 24792
rect 3752 24783 3754 24792
rect 3700 24754 3752 24760
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3608 24132 3660 24138
rect 3608 24074 3660 24080
rect 3330 24032 3386 24041
rect 3330 23967 3386 23976
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 3238 23216 3294 23225
rect 2872 23180 2924 23186
rect 3238 23151 3294 23160
rect 2872 23122 2924 23128
rect 3252 23050 3280 23151
rect 2780 23044 2832 23050
rect 2780 22986 2832 22992
rect 3240 23044 3292 23050
rect 3240 22986 3292 22992
rect 2792 22250 2820 22986
rect 2872 22568 2924 22574
rect 2872 22510 2924 22516
rect 2700 22222 2820 22250
rect 2700 21593 2728 22222
rect 2686 21584 2742 21593
rect 2596 21548 2648 21554
rect 2686 21519 2742 21528
rect 2596 21490 2648 21496
rect 2424 16546 2544 16574
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2424 9722 2452 10542
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2516 9382 2544 16546
rect 2608 11898 2636 21490
rect 2778 21176 2834 21185
rect 2884 21162 2912 22510
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3240 22092 3292 22098
rect 3240 22034 3292 22040
rect 3148 22024 3200 22030
rect 3252 22001 3280 22034
rect 3148 21966 3200 21972
rect 3238 21992 3294 22001
rect 3160 21350 3188 21966
rect 3238 21927 3294 21936
rect 3344 21570 3372 23967
rect 3620 23866 3648 24074
rect 3700 24064 3752 24070
rect 3700 24006 3752 24012
rect 4068 24064 4120 24070
rect 4068 24006 4120 24012
rect 3608 23860 3660 23866
rect 3608 23802 3660 23808
rect 3712 23712 3740 24006
rect 3620 23684 3740 23712
rect 3884 23724 3936 23730
rect 3424 23248 3476 23254
rect 3422 23216 3424 23225
rect 3476 23216 3478 23225
rect 3422 23151 3478 23160
rect 3516 22636 3568 22642
rect 3516 22578 3568 22584
rect 3424 21888 3476 21894
rect 3422 21856 3424 21865
rect 3476 21856 3478 21865
rect 3422 21791 3478 21800
rect 3344 21542 3464 21570
rect 3332 21480 3384 21486
rect 3332 21422 3384 21428
rect 3148 21344 3200 21350
rect 3148 21286 3200 21292
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2834 21134 2912 21162
rect 2778 21111 2834 21120
rect 2872 20868 2924 20874
rect 2872 20810 2924 20816
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2688 20324 2740 20330
rect 2688 20266 2740 20272
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2700 11286 2728 20266
rect 2792 19145 2820 20334
rect 2884 19938 2912 20810
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 3344 19961 3372 21422
rect 3330 19952 3386 19961
rect 2884 19910 3004 19938
rect 2872 19780 2924 19786
rect 2872 19722 2924 19728
rect 2778 19136 2834 19145
rect 2778 19071 2834 19080
rect 2884 18737 2912 19722
rect 2976 19553 3004 19910
rect 3330 19887 3386 19896
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 2962 19544 3018 19553
rect 2962 19479 3018 19488
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2870 18728 2926 18737
rect 2780 18692 2832 18698
rect 2870 18663 2926 18672
rect 2780 18634 2832 18640
rect 2792 17921 2820 18634
rect 2872 18624 2924 18630
rect 2872 18566 2924 18572
rect 2778 17912 2834 17921
rect 2884 17882 2912 18566
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 2778 17847 2834 17856
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 2780 17196 2832 17202
rect 2780 17138 2832 17144
rect 2792 13938 2820 17138
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2884 13938 2912 16730
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 3344 14940 3372 19790
rect 3436 18834 3464 21542
rect 3528 20602 3556 22578
rect 3620 21706 3648 23684
rect 3936 23684 4016 23712
rect 3884 23666 3936 23672
rect 3698 23624 3754 23633
rect 3698 23559 3700 23568
rect 3752 23559 3754 23568
rect 3700 23530 3752 23536
rect 3698 22808 3754 22817
rect 3698 22743 3754 22752
rect 3712 22166 3740 22743
rect 3700 22160 3752 22166
rect 3700 22102 3752 22108
rect 3988 21876 4016 23684
rect 3804 21848 4016 21876
rect 3620 21678 3740 21706
rect 3516 20596 3568 20602
rect 3516 20538 3568 20544
rect 3608 20460 3660 20466
rect 3608 20402 3660 20408
rect 3514 20224 3570 20233
rect 3514 20159 3570 20168
rect 3528 20058 3556 20159
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3516 18896 3568 18902
rect 3516 18838 3568 18844
rect 3424 18828 3476 18834
rect 3424 18770 3476 18776
rect 3424 18692 3476 18698
rect 3424 18634 3476 18640
rect 3436 18601 3464 18634
rect 3422 18592 3478 18601
rect 3422 18527 3478 18536
rect 3528 18426 3556 18838
rect 3620 18426 3648 20402
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 3608 18284 3660 18290
rect 3608 18226 3660 18232
rect 3620 18193 3648 18226
rect 3606 18184 3662 18193
rect 3606 18119 3662 18128
rect 3424 17672 3476 17678
rect 3422 17640 3424 17649
rect 3476 17640 3478 17649
rect 3422 17575 3478 17584
rect 3608 16992 3660 16998
rect 3608 16934 3660 16940
rect 3620 16454 3648 16934
rect 3608 16448 3660 16454
rect 3608 16390 3660 16396
rect 3606 16144 3662 16153
rect 3606 16079 3608 16088
rect 3660 16079 3662 16088
rect 3608 16050 3660 16056
rect 3620 15586 3648 16050
rect 3528 15558 3648 15586
rect 3424 15428 3476 15434
rect 3424 15370 3476 15376
rect 3436 15094 3464 15370
rect 3424 15088 3476 15094
rect 3424 15030 3476 15036
rect 3344 14912 3464 14940
rect 3436 14770 3464 14912
rect 3344 14742 3464 14770
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2778 13832 2834 13841
rect 2778 13767 2834 13776
rect 2792 13394 2820 13767
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2870 13424 2926 13433
rect 2780 13388 2832 13394
rect 2870 13359 2926 13368
rect 2780 13330 2832 13336
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2792 12442 2820 12718
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2884 11830 2912 13359
rect 3056 12912 3108 12918
rect 3054 12880 3056 12889
rect 3108 12880 3110 12889
rect 3054 12815 3110 12824
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2872 11824 2924 11830
rect 2872 11766 2924 11772
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2688 11280 2740 11286
rect 2688 11222 2740 11228
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2792 9450 2820 11018
rect 2884 10810 2912 11630
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 3344 11354 3372 14742
rect 3528 14618 3556 15558
rect 3608 15496 3660 15502
rect 3608 15438 3660 15444
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3620 14074 3648 15438
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 3422 13696 3478 13705
rect 3422 13631 3478 13640
rect 3436 13530 3464 13631
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3422 12336 3478 12345
rect 3422 12271 3424 12280
rect 3476 12271 3478 12280
rect 3424 12242 3476 12248
rect 3620 11898 3648 13874
rect 3712 12238 3740 21678
rect 3700 12232 3752 12238
rect 3700 12174 3752 12180
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3422 11248 3478 11257
rect 3422 11183 3478 11192
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 3332 10736 3384 10742
rect 3332 10678 3384 10684
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2870 9752 2926 9761
rect 2870 9687 2926 9696
rect 2780 9444 2832 9450
rect 2780 9386 2832 9392
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2884 8514 2912 9687
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2792 8486 2912 8514
rect 3148 8492 3200 8498
rect 2792 8362 2820 8486
rect 3148 8434 3200 8440
rect 2872 8424 2924 8430
rect 3160 8378 3188 8434
rect 2924 8372 3188 8378
rect 2872 8366 3188 8372
rect 2780 8356 2832 8362
rect 2884 8350 3188 8366
rect 3344 8362 3372 10678
rect 3436 8974 3464 11183
rect 3620 9722 3648 11834
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 3712 11354 3740 11698
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3804 10674 3832 21848
rect 3976 21344 4028 21350
rect 3976 21286 4028 21292
rect 3884 20392 3936 20398
rect 3882 20360 3884 20369
rect 3936 20360 3938 20369
rect 3882 20295 3938 20304
rect 3884 18760 3936 18766
rect 3884 18702 3936 18708
rect 3896 18154 3924 18702
rect 3884 18148 3936 18154
rect 3884 18090 3936 18096
rect 3882 16960 3938 16969
rect 3882 16895 3938 16904
rect 3896 16590 3924 16895
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3988 16182 4016 21286
rect 3976 16176 4028 16182
rect 3976 16118 4028 16124
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 3896 15706 3924 15982
rect 4080 15706 4108 24006
rect 4172 23798 4200 26200
rect 4344 25696 4396 25702
rect 4344 25638 4396 25644
rect 4252 24200 4304 24206
rect 4252 24142 4304 24148
rect 4160 23792 4212 23798
rect 4160 23734 4212 23740
rect 4160 23656 4212 23662
rect 4160 23598 4212 23604
rect 4172 22778 4200 23598
rect 4264 23497 4292 24142
rect 4250 23488 4306 23497
rect 4250 23423 4306 23432
rect 4356 23338 4384 25638
rect 4712 24948 4764 24954
rect 4712 24890 4764 24896
rect 4264 23310 4384 23338
rect 4618 23352 4674 23361
rect 4264 23118 4292 23310
rect 4618 23287 4674 23296
rect 4436 23180 4488 23186
rect 4436 23122 4488 23128
rect 4252 23112 4304 23118
rect 4250 23080 4252 23089
rect 4344 23112 4396 23118
rect 4304 23080 4306 23089
rect 4344 23054 4396 23060
rect 4250 23015 4306 23024
rect 4160 22772 4212 22778
rect 4160 22714 4212 22720
rect 4356 22624 4384 23054
rect 4264 22596 4384 22624
rect 4158 22128 4214 22137
rect 4158 22063 4214 22072
rect 4172 21010 4200 22063
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 4158 20904 4214 20913
rect 4158 20839 4214 20848
rect 4172 17746 4200 20839
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 3884 15700 3936 15706
rect 3884 15642 3936 15648
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 3976 14544 4028 14550
rect 3974 14512 3976 14521
rect 4028 14512 4030 14521
rect 3974 14447 4030 14456
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 3974 13288 4030 13297
rect 3974 13223 3976 13232
rect 4028 13223 4030 13232
rect 3976 13194 4028 13200
rect 3882 13016 3938 13025
rect 3882 12951 3884 12960
rect 3936 12951 3938 12960
rect 3884 12922 3936 12928
rect 3974 12744 4030 12753
rect 3974 12679 4030 12688
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3896 11558 3924 12174
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3896 11393 3924 11494
rect 3882 11384 3938 11393
rect 3882 11319 3938 11328
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3712 10577 3740 10610
rect 3698 10568 3754 10577
rect 3698 10503 3754 10512
rect 3712 10266 3740 10503
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 3988 9586 4016 12679
rect 4080 12238 4108 13874
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 4080 11830 4108 12038
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 4158 11792 4214 11801
rect 4080 10810 4108 11766
rect 4158 11727 4214 11736
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 4172 9586 4200 11727
rect 4264 10130 4292 22596
rect 4448 22094 4476 23122
rect 4528 22432 4580 22438
rect 4528 22374 4580 22380
rect 4356 22066 4476 22094
rect 4356 21622 4384 22066
rect 4344 21616 4396 21622
rect 4344 21558 4396 21564
rect 4436 21616 4488 21622
rect 4436 21558 4488 21564
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4356 11898 4384 17138
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4356 11150 4384 11494
rect 4448 11354 4476 21558
rect 4540 19446 4568 22374
rect 4528 19440 4580 19446
rect 4528 19382 4580 19388
rect 4632 19242 4660 23287
rect 4724 20942 4752 24890
rect 4804 23724 4856 23730
rect 4804 23666 4856 23672
rect 4816 23633 4844 23666
rect 4802 23624 4858 23633
rect 4802 23559 4858 23568
rect 4804 23248 4856 23254
rect 4804 23190 4856 23196
rect 4712 20936 4764 20942
rect 4712 20878 4764 20884
rect 4620 19236 4672 19242
rect 4620 19178 4672 19184
rect 4710 17912 4766 17921
rect 4710 17847 4766 17856
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4632 17338 4660 17614
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4528 13456 4580 13462
rect 4528 13398 4580 13404
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4540 10810 4568 13398
rect 4632 12918 4660 15438
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4724 12730 4752 17847
rect 4816 17270 4844 23190
rect 5092 22574 5120 26302
rect 5446 26200 5502 27000
rect 6090 26200 6146 27000
rect 6734 26200 6790 27000
rect 6826 26208 6882 26217
rect 5460 23662 5488 26200
rect 5998 24712 6054 24721
rect 5998 24647 6054 24656
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5632 23588 5684 23594
rect 5632 23530 5684 23536
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 4988 22500 5040 22506
rect 4988 22442 5040 22448
rect 4896 22228 4948 22234
rect 4896 22170 4948 22176
rect 4908 19922 4936 22170
rect 5000 20534 5028 22442
rect 5540 21888 5592 21894
rect 5540 21830 5592 21836
rect 5172 20936 5224 20942
rect 5172 20878 5224 20884
rect 4988 20528 5040 20534
rect 4988 20470 5040 20476
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 4896 19780 4948 19786
rect 4896 19722 4948 19728
rect 4804 17264 4856 17270
rect 4804 17206 4856 17212
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4816 15609 4844 15846
rect 4802 15600 4858 15609
rect 4802 15535 4858 15544
rect 4908 14498 4936 19722
rect 5080 19236 5132 19242
rect 5080 19178 5132 19184
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 4816 14470 4936 14498
rect 4816 14346 4844 14470
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 4804 14340 4856 14346
rect 4804 14282 4856 14288
rect 4908 14074 4936 14350
rect 4896 14068 4948 14074
rect 4896 14010 4948 14016
rect 5000 12986 5028 18702
rect 5092 13326 5120 19178
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 4632 12702 4752 12730
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4632 12238 4660 12702
rect 4710 12608 4766 12617
rect 4710 12543 4766 12552
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4632 11626 4660 12038
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 4632 11257 4660 11562
rect 4618 11248 4674 11257
rect 4618 11183 4674 11192
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3528 8401 3556 9522
rect 3620 9178 3648 9522
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 4356 8838 4384 10542
rect 4724 9654 4752 12543
rect 4816 11898 4844 12718
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 5184 11354 5212 20878
rect 5448 19712 5500 19718
rect 5448 19654 5500 19660
rect 5354 19408 5410 19417
rect 5354 19343 5410 19352
rect 5368 16726 5396 19343
rect 5460 18970 5488 19654
rect 5552 18970 5580 21830
rect 5644 21486 5672 23530
rect 5816 22024 5868 22030
rect 5814 21992 5816 22001
rect 5868 21992 5870 22001
rect 5814 21927 5870 21936
rect 6012 21690 6040 24647
rect 6104 23186 6132 26200
rect 6550 25120 6606 25129
rect 6550 25055 6606 25064
rect 6276 24812 6328 24818
rect 6276 24754 6328 24760
rect 6184 23520 6236 23526
rect 6184 23462 6236 23468
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 6092 22024 6144 22030
rect 6092 21966 6144 21972
rect 6000 21684 6052 21690
rect 6000 21626 6052 21632
rect 5908 21548 5960 21554
rect 5908 21490 5960 21496
rect 5632 21480 5684 21486
rect 5632 21422 5684 21428
rect 5632 21344 5684 21350
rect 5632 21286 5684 21292
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5540 18692 5592 18698
rect 5540 18634 5592 18640
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5356 16720 5408 16726
rect 5356 16662 5408 16668
rect 5460 16590 5488 17138
rect 5264 16584 5316 16590
rect 5262 16552 5264 16561
rect 5448 16584 5500 16590
rect 5316 16552 5318 16561
rect 5448 16526 5500 16532
rect 5262 16487 5318 16496
rect 5552 16436 5580 18634
rect 5460 16408 5580 16436
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5276 14550 5304 16050
rect 5354 15736 5410 15745
rect 5354 15671 5356 15680
rect 5408 15671 5410 15680
rect 5356 15642 5408 15648
rect 5356 15428 5408 15434
rect 5356 15370 5408 15376
rect 5264 14544 5316 14550
rect 5264 14486 5316 14492
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5276 11665 5304 11698
rect 5262 11656 5318 11665
rect 5262 11591 5264 11600
rect 5316 11591 5318 11600
rect 5264 11562 5316 11568
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5264 11008 5316 11014
rect 5368 10985 5396 15370
rect 5460 13852 5488 16408
rect 5460 13824 5580 13852
rect 5446 13696 5502 13705
rect 5446 13631 5502 13640
rect 5460 11898 5488 13631
rect 5552 12850 5580 13824
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5644 12730 5672 21286
rect 5722 21040 5778 21049
rect 5722 20975 5778 20984
rect 5736 19786 5764 20975
rect 5724 19780 5776 19786
rect 5724 19722 5776 19728
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 5736 18698 5764 19246
rect 5724 18692 5776 18698
rect 5724 18634 5776 18640
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5828 18329 5856 18566
rect 5814 18320 5870 18329
rect 5814 18255 5870 18264
rect 5920 18086 5948 21490
rect 6000 18284 6052 18290
rect 6000 18226 6052 18232
rect 5724 18080 5776 18086
rect 5724 18022 5776 18028
rect 5908 18080 5960 18086
rect 5908 18022 5960 18028
rect 5736 17678 5764 18022
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 5908 16448 5960 16454
rect 5908 16390 5960 16396
rect 5816 16040 5868 16046
rect 5816 15982 5868 15988
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 5736 14618 5764 15438
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5828 12866 5856 15982
rect 5920 14006 5948 16390
rect 6012 16250 6040 18226
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 6012 14657 6040 14758
rect 5998 14648 6054 14657
rect 5998 14583 6054 14592
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 6012 14074 6040 14350
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 5908 14000 5960 14006
rect 5908 13942 5960 13948
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 6012 12986 6040 13806
rect 6104 13274 6132 21966
rect 6196 19922 6224 23462
rect 6288 20534 6316 24754
rect 6460 23860 6512 23866
rect 6460 23802 6512 23808
rect 6368 22704 6420 22710
rect 6368 22646 6420 22652
rect 6380 22234 6408 22646
rect 6368 22228 6420 22234
rect 6368 22170 6420 22176
rect 6366 22128 6422 22137
rect 6366 22063 6422 22072
rect 6380 21078 6408 22063
rect 6368 21072 6420 21078
rect 6368 21014 6420 21020
rect 6276 20528 6328 20534
rect 6276 20470 6328 20476
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 6276 19780 6328 19786
rect 6276 19722 6328 19728
rect 6184 18692 6236 18698
rect 6184 18634 6236 18640
rect 6196 18465 6224 18634
rect 6182 18456 6238 18465
rect 6182 18391 6238 18400
rect 6182 18184 6238 18193
rect 6182 18119 6238 18128
rect 6196 14958 6224 18119
rect 6184 14952 6236 14958
rect 6184 14894 6236 14900
rect 6104 13246 6224 13274
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 5828 12838 6040 12866
rect 5644 12702 5948 12730
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5722 11792 5778 11801
rect 5722 11727 5778 11736
rect 5540 11620 5592 11626
rect 5540 11562 5592 11568
rect 5552 11286 5580 11562
rect 5736 11354 5764 11727
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5264 10950 5316 10956
rect 5354 10976 5410 10985
rect 5276 10742 5304 10950
rect 5354 10911 5410 10920
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5170 10296 5226 10305
rect 5170 10231 5172 10240
rect 5224 10231 5226 10240
rect 5172 10202 5224 10208
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5368 8838 5396 9522
rect 5552 9382 5580 9998
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5644 8634 5672 9930
rect 5736 9654 5764 10406
rect 5828 10198 5856 12582
rect 5920 10266 5948 12702
rect 6012 10606 6040 12838
rect 6104 11830 6132 13126
rect 6196 12646 6224 13246
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6182 12472 6238 12481
rect 6182 12407 6238 12416
rect 6092 11824 6144 11830
rect 6092 11766 6144 11772
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 6012 9926 6040 10406
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6012 9353 6040 9522
rect 5998 9344 6054 9353
rect 5998 9279 6054 9288
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 6012 8566 6040 9279
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 3514 8392 3570 8401
rect 3332 8356 3384 8362
rect 2780 8298 2832 8304
rect 3514 8327 3570 8336
rect 3332 8298 3384 8304
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 1582 8055 1638 8064
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 1308 7880 1360 7886
rect 1308 7822 1360 7828
rect 1320 7721 1348 7822
rect 1306 7712 1362 7721
rect 1306 7647 1362 7656
rect 6104 7478 6132 11630
rect 6196 10674 6224 12407
rect 6288 11354 6316 19722
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 6380 16697 6408 17274
rect 6366 16688 6422 16697
rect 6366 16623 6422 16632
rect 6368 16516 6420 16522
rect 6368 16458 6420 16464
rect 6380 16250 6408 16458
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6472 16114 6500 23802
rect 6564 23730 6592 25055
rect 6748 24342 6776 26200
rect 7378 26200 7434 27000
rect 8022 26330 8078 27000
rect 7852 26302 8078 26330
rect 6826 26143 6882 26152
rect 6736 24336 6788 24342
rect 6736 24278 6788 24284
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6736 23044 6788 23050
rect 6736 22986 6788 22992
rect 6644 22568 6696 22574
rect 6644 22510 6696 22516
rect 6552 19168 6604 19174
rect 6550 19136 6552 19145
rect 6604 19136 6606 19145
rect 6550 19071 6606 19080
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 6564 18358 6592 18702
rect 6552 18352 6604 18358
rect 6552 18294 6604 18300
rect 6656 17882 6684 22510
rect 6748 21010 6776 22986
rect 6840 22710 6868 26143
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 6828 22704 6880 22710
rect 6826 22672 6828 22681
rect 6880 22672 6882 22681
rect 6826 22607 6882 22616
rect 6828 22160 6880 22166
rect 6826 22128 6828 22137
rect 6880 22128 6882 22137
rect 6826 22063 6882 22072
rect 6736 21004 6788 21010
rect 6736 20946 6788 20952
rect 6736 20868 6788 20874
rect 6736 20810 6788 20816
rect 6644 17876 6696 17882
rect 6644 17818 6696 17824
rect 6748 17762 6776 20810
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 6656 17734 6776 17762
rect 6656 17082 6684 17734
rect 6840 17678 6868 19314
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6564 17054 6684 17082
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6458 15872 6514 15881
rect 6458 15807 6514 15816
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6380 13977 6408 14010
rect 6366 13968 6422 13977
rect 6366 13903 6422 13912
rect 6366 13832 6422 13841
rect 6366 13767 6422 13776
rect 6380 12986 6408 13767
rect 6472 13376 6500 15807
rect 6564 13734 6592 17054
rect 6748 16017 6776 17138
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6734 16008 6790 16017
rect 6734 15943 6790 15952
rect 6840 15502 6868 16390
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6656 14090 6684 15302
rect 6736 15088 6788 15094
rect 6736 15030 6788 15036
rect 6748 14550 6776 15030
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 6656 14062 6776 14090
rect 6840 14074 6868 14962
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6472 13348 6592 13376
rect 6460 13252 6512 13258
rect 6460 13194 6512 13200
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 6472 12866 6500 13194
rect 6380 12838 6500 12866
rect 6380 12442 6408 12838
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6196 9518 6224 10610
rect 6380 9994 6408 12242
rect 6472 11150 6500 12718
rect 6564 12481 6592 13348
rect 6550 12472 6606 12481
rect 6550 12407 6606 12416
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6656 10033 6684 13874
rect 6748 12782 6776 14062
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 12986 6868 13670
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6734 12200 6790 12209
rect 6734 12135 6790 12144
rect 6748 11762 6776 12135
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6932 11014 6960 23598
rect 7010 23488 7066 23497
rect 7010 23423 7066 23432
rect 7024 22710 7052 23423
rect 7288 22772 7340 22778
rect 7288 22714 7340 22720
rect 7012 22704 7064 22710
rect 7012 22646 7064 22652
rect 7300 22386 7328 22714
rect 7392 22574 7420 26200
rect 7654 24848 7710 24857
rect 7654 24783 7710 24792
rect 7472 23112 7524 23118
rect 7472 23054 7524 23060
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 7380 22432 7432 22438
rect 7300 22380 7380 22386
rect 7300 22374 7432 22380
rect 7300 22358 7420 22374
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 7012 19440 7064 19446
rect 7012 19382 7064 19388
rect 7024 18970 7052 19382
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 7010 18864 7066 18873
rect 7116 18834 7144 19110
rect 7010 18799 7066 18808
rect 7104 18828 7156 18834
rect 7024 18290 7052 18799
rect 7104 18770 7156 18776
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 7024 17241 7052 18226
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 7010 17232 7066 17241
rect 7010 17167 7066 17176
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 7024 15162 7052 17070
rect 7116 16182 7144 18158
rect 7208 16726 7236 19790
rect 7196 16720 7248 16726
rect 7196 16662 7248 16668
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7104 16176 7156 16182
rect 7104 16118 7156 16124
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 7104 14884 7156 14890
rect 7104 14826 7156 14832
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 7024 13841 7052 14418
rect 7010 13832 7066 13841
rect 7010 13767 7066 13776
rect 7116 12850 7144 14826
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6932 10674 6960 10950
rect 7116 10742 7144 12582
rect 7208 12306 7236 16390
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6642 10024 6698 10033
rect 6368 9988 6420 9994
rect 6642 9959 6698 9968
rect 6368 9930 6420 9936
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 1308 7404 1360 7410
rect 1308 7346 1360 7352
rect 1320 7313 1348 7346
rect 1306 7304 1362 7313
rect 1306 7239 1362 7248
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1780 7002 1808 7142
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1214 6896 1270 6905
rect 1214 6831 1270 6840
rect 1228 6798 1256 6831
rect 1216 6792 1268 6798
rect 1216 6734 1268 6740
rect 1228 6458 1256 6734
rect 1308 6724 1360 6730
rect 1308 6666 1360 6672
rect 1320 6497 1348 6666
rect 1768 6656 1820 6662
rect 1768 6598 1820 6604
rect 1306 6488 1362 6497
rect 1216 6452 1268 6458
rect 1306 6423 1362 6432
rect 1216 6394 1268 6400
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 1320 6089 1348 6258
rect 1306 6080 1362 6089
rect 1306 6015 1362 6024
rect 1780 5914 1808 6598
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 1308 5704 1360 5710
rect 1306 5672 1308 5681
rect 2780 5704 2832 5710
rect 1360 5672 1362 5681
rect 2780 5646 2832 5652
rect 1306 5607 1362 5616
rect 2792 5273 2820 5646
rect 2778 5264 2834 5273
rect 2778 5199 2834 5208
rect 1308 5160 1360 5166
rect 1308 5102 1360 5108
rect 1320 4865 1348 5102
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 1306 4856 1362 4865
rect 2950 4859 3258 4868
rect 1306 4791 1308 4800
rect 1360 4791 1362 4800
rect 1308 4762 1360 4768
rect 1308 4548 1360 4554
rect 1308 4490 1360 4496
rect 1320 4457 1348 4490
rect 1306 4448 1362 4457
rect 1306 4383 1362 4392
rect 1308 4140 1360 4146
rect 1308 4082 1360 4088
rect 1216 4072 1268 4078
rect 1320 4049 1348 4082
rect 2412 4072 2464 4078
rect 1216 4014 1268 4020
rect 1306 4040 1362 4049
rect 1228 3641 1256 4014
rect 2148 4020 2412 4026
rect 2148 4014 2464 4020
rect 2148 4010 2452 4014
rect 1306 3975 1362 3984
rect 2136 4004 2452 4010
rect 2188 3998 2452 4004
rect 2136 3946 2188 3952
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 3332 3664 3384 3670
rect 1214 3632 1270 3641
rect 3332 3606 3384 3612
rect 1214 3567 1270 3576
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1032 3460 1084 3466
rect 1032 3402 1084 3408
rect 1044 1442 1072 3402
rect 1320 3233 1348 3470
rect 1306 3224 1362 3233
rect 1306 3159 1308 3168
rect 1360 3159 1362 3168
rect 1308 3130 1360 3136
rect 1308 3052 1360 3058
rect 1308 2994 1360 3000
rect 1320 2825 1348 2994
rect 2320 2848 2372 2854
rect 1306 2816 1362 2825
rect 2320 2790 2372 2796
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 1306 2751 1362 2760
rect 2332 2446 2360 2790
rect 2792 2514 2820 2790
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 1308 2440 1360 2446
rect 1306 2408 1308 2417
rect 2320 2440 2372 2446
rect 1360 2408 1362 2417
rect 1216 2372 1268 2378
rect 2320 2382 2372 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 1306 2343 1362 2352
rect 1216 2314 1268 2320
rect 1228 2009 1256 2314
rect 1214 2000 1270 2009
rect 1214 1935 1270 1944
rect 3252 1601 3280 2382
rect 3238 1592 3294 1601
rect 3238 1527 3294 1536
rect 1044 1414 1164 1442
rect 1136 800 1164 1414
rect 3344 1034 3372 3606
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 3252 1006 3372 1034
rect 3252 800 3280 1006
rect 5368 800 5396 3334
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6380 2378 6408 2586
rect 6368 2372 6420 2378
rect 6368 2314 6420 2320
rect 6932 2310 6960 9454
rect 7208 9450 7236 11698
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7300 9042 7328 19858
rect 7392 18408 7420 22358
rect 7484 18737 7512 23054
rect 7564 22772 7616 22778
rect 7564 22714 7616 22720
rect 7576 21842 7604 22714
rect 7668 22030 7696 24783
rect 7852 23186 7880 26302
rect 8022 26200 8078 26302
rect 8666 26200 8722 27000
rect 9310 26330 9366 27000
rect 9140 26302 9366 26330
rect 8680 24274 8708 26200
rect 8852 25220 8904 25226
rect 8852 25162 8904 25168
rect 8668 24268 8720 24274
rect 8668 24210 8720 24216
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8760 23792 8812 23798
rect 8760 23734 8812 23740
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 8300 23112 8352 23118
rect 8300 23054 8352 23060
rect 7748 22976 7800 22982
rect 7748 22918 7800 22924
rect 7760 22545 7788 22918
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7746 22536 7802 22545
rect 7746 22471 7802 22480
rect 7656 22024 7708 22030
rect 7656 21966 7708 21972
rect 7656 21888 7708 21894
rect 7576 21836 7656 21842
rect 7576 21830 7708 21836
rect 7576 21814 7696 21830
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7470 18728 7526 18737
rect 7470 18663 7526 18672
rect 7392 18380 7512 18408
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7392 17338 7420 18226
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7378 17232 7434 17241
rect 7378 17167 7434 17176
rect 7392 15706 7420 17167
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7380 15564 7432 15570
rect 7380 15506 7432 15512
rect 7392 11558 7420 15506
rect 7484 13530 7512 18380
rect 7576 14890 7604 21354
rect 7668 20806 7696 21814
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 7668 19718 7696 20742
rect 7748 20324 7800 20330
rect 7748 20266 7800 20272
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7668 19174 7696 19654
rect 7760 19378 7788 20266
rect 7852 19922 7880 22578
rect 8024 22568 8076 22574
rect 8024 22510 8076 22516
rect 8036 22438 8064 22510
rect 8024 22432 8076 22438
rect 8024 22374 8076 22380
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 7932 21616 7984 21622
rect 7932 21558 7984 21564
rect 7944 20942 7972 21558
rect 7932 20936 7984 20942
rect 7932 20878 7984 20884
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8312 19961 8340 23054
rect 8392 20528 8444 20534
rect 8390 20496 8392 20505
rect 8444 20496 8446 20505
rect 8772 20466 8800 23734
rect 8864 21486 8892 25162
rect 8944 24268 8996 24274
rect 8944 24210 8996 24216
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 8852 21344 8904 21350
rect 8852 21286 8904 21292
rect 8390 20431 8446 20440
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 8772 20369 8800 20402
rect 8758 20360 8814 20369
rect 8758 20295 8814 20304
rect 8864 20210 8892 21286
rect 8956 20534 8984 24210
rect 9036 24200 9088 24206
rect 9036 24142 9088 24148
rect 9048 21554 9076 24142
rect 9140 23798 9168 26302
rect 9310 26200 9366 26302
rect 9954 26330 10010 27000
rect 10598 26330 10654 27000
rect 9954 26302 10272 26330
rect 9954 26200 10010 26302
rect 9864 24880 9916 24886
rect 9864 24822 9916 24828
rect 9312 24064 9364 24070
rect 9312 24006 9364 24012
rect 9404 24064 9456 24070
rect 9404 24006 9456 24012
rect 9128 23792 9180 23798
rect 9128 23734 9180 23740
rect 9220 23724 9272 23730
rect 9220 23666 9272 23672
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 8944 20528 8996 20534
rect 8944 20470 8996 20476
rect 8772 20182 8892 20210
rect 8298 19952 8354 19961
rect 7840 19916 7892 19922
rect 8298 19887 8354 19896
rect 7840 19858 7892 19864
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8206 19408 8262 19417
rect 7748 19372 7800 19378
rect 8206 19343 8208 19352
rect 7748 19314 7800 19320
rect 8260 19343 8262 19352
rect 8208 19314 8260 19320
rect 7748 19236 7800 19242
rect 7748 19178 7800 19184
rect 7840 19236 7892 19242
rect 7840 19178 7892 19184
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7760 18970 7788 19178
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7656 18896 7708 18902
rect 7656 18838 7708 18844
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7576 14278 7604 14418
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7564 13728 7616 13734
rect 7564 13670 7616 13676
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7576 12306 7604 13670
rect 7668 12442 7696 18838
rect 7852 18766 7880 19178
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 8024 19168 8076 19174
rect 8024 19110 8076 19116
rect 7840 18760 7892 18766
rect 7840 18702 7892 18708
rect 7748 18692 7800 18698
rect 7748 18634 7800 18640
rect 7760 17066 7788 18634
rect 7944 18612 7972 19110
rect 8036 18970 8064 19110
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 7852 18584 7972 18612
rect 7852 18154 7880 18584
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8312 18306 8340 19887
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8588 19378 8616 19654
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8484 18692 8536 18698
rect 8484 18634 8536 18640
rect 8312 18278 8432 18306
rect 8496 18290 8524 18634
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 7840 18148 7892 18154
rect 7840 18090 7892 18096
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8116 17264 8168 17270
rect 8114 17232 8116 17241
rect 8168 17232 8170 17241
rect 8114 17167 8170 17176
rect 7748 17060 7800 17066
rect 7748 17002 7800 17008
rect 8312 16794 8340 18090
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8116 16652 8168 16658
rect 7852 16612 8116 16640
rect 7852 16250 7880 16612
rect 8116 16594 8168 16600
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7840 16244 7892 16250
rect 8312 16232 8340 16730
rect 7840 16186 7892 16192
rect 8220 16204 8340 16232
rect 7760 16130 7788 16186
rect 7760 16102 7880 16130
rect 7748 15972 7800 15978
rect 7748 15914 7800 15920
rect 7760 15162 7788 15914
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7852 15094 7880 16102
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 7932 15972 7984 15978
rect 7932 15914 7984 15920
rect 7944 15706 7972 15914
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 8128 15570 8156 16050
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8220 15450 8248 16204
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8312 15570 8340 15846
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8220 15422 8340 15450
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7840 15088 7892 15094
rect 7840 15030 7892 15036
rect 8022 15056 8078 15065
rect 7932 15020 7984 15026
rect 8022 14991 8024 15000
rect 7932 14962 7984 14968
rect 8076 14991 8078 15000
rect 8024 14962 8076 14968
rect 7748 14884 7800 14890
rect 7748 14826 7800 14832
rect 7840 14884 7892 14890
rect 7840 14826 7892 14832
rect 7760 12646 7788 14826
rect 7852 13870 7880 14826
rect 7944 14618 7972 14962
rect 8312 14822 8340 15422
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 8312 14278 8340 14758
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7656 12436 7708 12442
rect 7852 12434 7880 13262
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 7656 12378 7708 12384
rect 7760 12406 7880 12434
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7484 11098 7512 12242
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7392 11082 7512 11098
rect 7380 11076 7512 11082
rect 7432 11070 7512 11076
rect 7380 11018 7432 11024
rect 7378 10296 7434 10305
rect 7378 10231 7380 10240
rect 7432 10231 7434 10240
rect 7380 10202 7432 10208
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7484 7750 7512 11070
rect 7576 8634 7604 12038
rect 7760 11830 7788 12406
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 7852 11694 7880 12174
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 8036 10062 8064 10474
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 8312 9722 8340 10610
rect 8404 10198 8432 18278
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8496 15638 8524 17070
rect 8588 16114 8616 18566
rect 8668 16176 8720 16182
rect 8668 16118 8720 16124
rect 8576 16108 8628 16114
rect 8576 16050 8628 16056
rect 8484 15632 8536 15638
rect 8680 15609 8708 16118
rect 8484 15574 8536 15580
rect 8666 15600 8722 15609
rect 8666 15535 8722 15544
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8496 13462 8524 14962
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8484 13456 8536 13462
rect 8484 13398 8536 13404
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8496 10062 8524 13126
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8404 9897 8432 9998
rect 8390 9888 8446 9897
rect 8390 9823 8446 9832
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 7654 9616 7710 9625
rect 7654 9551 7710 9560
rect 7668 8974 7696 9551
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 7760 9042 7788 9318
rect 8036 9110 8064 9318
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 8404 8090 8432 8842
rect 8496 8809 8524 9114
rect 8588 9042 8616 12038
rect 8680 10266 8708 14554
rect 8772 14414 8800 20182
rect 9048 19394 9076 21490
rect 9128 19712 9180 19718
rect 9126 19680 9128 19689
rect 9180 19680 9182 19689
rect 9126 19615 9182 19624
rect 8956 19366 9076 19394
rect 8956 18850 8984 19366
rect 9034 19272 9090 19281
rect 9232 19258 9260 23666
rect 9324 22778 9352 24006
rect 9416 23769 9444 24006
rect 9402 23760 9458 23769
rect 9402 23695 9458 23704
rect 9680 22976 9732 22982
rect 9680 22918 9732 22924
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 9312 20800 9364 20806
rect 9312 20742 9364 20748
rect 9034 19207 9090 19216
rect 9140 19230 9260 19258
rect 9048 18970 9076 19207
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 8956 18822 9076 18850
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8852 18352 8904 18358
rect 8956 18306 8984 18566
rect 8904 18300 8984 18306
rect 8852 18294 8984 18300
rect 8864 18278 8984 18294
rect 8864 18222 8892 18278
rect 8852 18216 8904 18222
rect 8852 18158 8904 18164
rect 8956 17542 8984 18278
rect 8944 17536 8996 17542
rect 8944 17478 8996 17484
rect 8956 16794 8984 17478
rect 8944 16788 8996 16794
rect 8944 16730 8996 16736
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 8864 15910 8892 16186
rect 8956 16017 8984 16594
rect 9048 16454 9076 18822
rect 9140 17513 9168 19230
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9232 18902 9260 19110
rect 9220 18896 9272 18902
rect 9220 18838 9272 18844
rect 9218 17640 9274 17649
rect 9218 17575 9220 17584
rect 9272 17575 9274 17584
rect 9220 17546 9272 17552
rect 9126 17504 9182 17513
rect 9126 17439 9182 17448
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 9140 16776 9168 16934
rect 9140 16748 9260 16776
rect 9232 16590 9260 16748
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 9036 16040 9088 16046
rect 8942 16008 8998 16017
rect 9036 15982 9088 15988
rect 8942 15943 8998 15952
rect 8956 15910 8984 15943
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8760 13456 8812 13462
rect 8864 13433 8892 15846
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 8760 13398 8812 13404
rect 8850 13424 8906 13433
rect 8772 10690 8800 13398
rect 8850 13359 8906 13368
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 8864 12986 8892 13262
rect 8852 12980 8904 12986
rect 8852 12922 8904 12928
rect 8852 12164 8904 12170
rect 8852 12106 8904 12112
rect 8864 10810 8892 12106
rect 8956 11354 8984 14350
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 8772 10662 8892 10690
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8864 9058 8892 10662
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8772 9030 8892 9058
rect 8576 8832 8628 8838
rect 8482 8800 8538 8809
rect 8576 8774 8628 8780
rect 8482 8735 8538 8744
rect 8588 8430 8616 8774
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 7472 7744 7524 7750
rect 8588 7721 8616 7822
rect 7472 7686 7524 7692
rect 8574 7712 8630 7721
rect 7950 7644 8258 7653
rect 8574 7647 8630 7656
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 8772 6730 8800 9030
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7470 4040 7526 4049
rect 7470 3975 7526 3984
rect 8300 4004 8352 4010
rect 7484 3398 7512 3975
rect 8300 3946 8352 3952
rect 8312 3641 8340 3946
rect 8298 3632 8354 3641
rect 8298 3567 8354 3576
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 7472 2916 7524 2922
rect 7472 2858 7524 2864
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 7484 800 7512 2858
rect 8772 2446 8800 3334
rect 8864 2854 8892 8842
rect 8956 5234 8984 11154
rect 9048 10674 9076 15982
rect 9140 15094 9168 16526
rect 9220 16448 9272 16454
rect 9220 16390 9272 16396
rect 9232 15638 9260 16390
rect 9324 16266 9352 20742
rect 9416 20466 9444 21830
rect 9508 21146 9536 21830
rect 9496 21140 9548 21146
rect 9496 21082 9548 21088
rect 9692 20942 9720 22918
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9784 22409 9812 22578
rect 9770 22400 9826 22409
rect 9770 22335 9826 22344
rect 9772 22094 9824 22098
rect 9876 22094 9904 24822
rect 10140 24336 10192 24342
rect 10140 24278 10192 24284
rect 9956 22228 10008 22234
rect 9956 22170 10008 22176
rect 9772 22092 9904 22094
rect 9824 22066 9904 22092
rect 9772 22034 9824 22040
rect 9770 21448 9826 21457
rect 9770 21383 9826 21392
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9784 20806 9812 21383
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9404 20460 9456 20466
rect 9404 20402 9456 20408
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 9416 17626 9444 18022
rect 9508 17882 9536 18702
rect 9600 18630 9628 19110
rect 9692 18873 9720 20538
rect 9968 20534 9996 22170
rect 10152 21865 10180 24278
rect 10244 22574 10272 26302
rect 10598 26302 10732 26330
rect 10598 26200 10654 26302
rect 10508 24404 10560 24410
rect 10508 24346 10560 24352
rect 10520 23118 10548 24346
rect 10704 23798 10732 26302
rect 11242 26200 11298 27000
rect 11886 26200 11942 27000
rect 12530 26330 12586 27000
rect 12256 26308 12308 26314
rect 12256 26250 12308 26256
rect 12452 26302 12586 26330
rect 10784 24132 10836 24138
rect 10784 24074 10836 24080
rect 10692 23792 10744 23798
rect 10692 23734 10744 23740
rect 10796 23526 10824 24074
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 11256 23186 11284 26200
rect 11518 25256 11574 25265
rect 11518 25191 11574 25200
rect 11336 24608 11388 24614
rect 11336 24550 11388 24556
rect 11244 23180 11296 23186
rect 11244 23122 11296 23128
rect 10508 23112 10560 23118
rect 10508 23054 10560 23060
rect 11060 22704 11112 22710
rect 11058 22672 11060 22681
rect 11112 22672 11114 22681
rect 11058 22607 11114 22616
rect 10232 22568 10284 22574
rect 10232 22510 10284 22516
rect 10324 22228 10376 22234
rect 10324 22170 10376 22176
rect 10138 21856 10194 21865
rect 10138 21791 10194 21800
rect 10152 21690 10180 21791
rect 10140 21684 10192 21690
rect 10140 21626 10192 21632
rect 10336 21146 10364 22170
rect 11348 21962 11376 24550
rect 11428 24064 11480 24070
rect 11428 24006 11480 24012
rect 11440 23662 11468 24006
rect 11428 23656 11480 23662
rect 11428 23598 11480 23604
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 11348 21729 11376 21898
rect 11334 21720 11390 21729
rect 11334 21655 11390 21664
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 10324 21140 10376 21146
rect 10324 21082 10376 21088
rect 10324 20800 10376 20806
rect 10324 20742 10376 20748
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 9956 20392 10008 20398
rect 9956 20334 10008 20340
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9784 19854 9812 20198
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9862 19816 9918 19825
rect 9862 19751 9918 19760
rect 9678 18864 9734 18873
rect 9678 18799 9734 18808
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 9600 17921 9628 18566
rect 9876 18408 9904 19751
rect 9968 19514 9996 20334
rect 10140 20256 10192 20262
rect 10140 20198 10192 20204
rect 10152 19922 10180 20198
rect 10140 19916 10192 19922
rect 10140 19858 10192 19864
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10048 18828 10100 18834
rect 10048 18770 10100 18776
rect 9784 18380 9904 18408
rect 9586 17912 9642 17921
rect 9496 17876 9548 17882
rect 9586 17847 9642 17856
rect 9496 17818 9548 17824
rect 9784 17746 9812 18380
rect 10060 18358 10088 18770
rect 10048 18352 10100 18358
rect 10048 18294 10100 18300
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9956 17672 10008 17678
rect 9416 17610 9628 17626
rect 9956 17614 10008 17620
rect 9416 17604 9640 17610
rect 9416 17598 9588 17604
rect 9588 17546 9640 17552
rect 9968 17270 9996 17614
rect 9956 17264 10008 17270
rect 9956 17206 10008 17212
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 10060 16998 10088 17070
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 9324 16238 9444 16266
rect 9312 15972 9364 15978
rect 9312 15914 9364 15920
rect 9220 15632 9272 15638
rect 9220 15574 9272 15580
rect 9324 15366 9352 15914
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9128 15088 9180 15094
rect 9128 15030 9180 15036
rect 9126 14784 9182 14793
rect 9126 14719 9182 14728
rect 9140 13462 9168 14719
rect 9416 14618 9444 16238
rect 10060 15881 10088 16730
rect 10046 15872 10102 15881
rect 10046 15807 10102 15816
rect 10046 15600 10102 15609
rect 10046 15535 10048 15544
rect 10100 15535 10102 15544
rect 10048 15506 10100 15512
rect 9494 15464 9550 15473
rect 9494 15399 9496 15408
rect 9548 15399 9550 15408
rect 9496 15370 9548 15376
rect 9508 14958 9536 15370
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 9312 13796 9364 13802
rect 9312 13738 9364 13744
rect 9232 13705 9260 13738
rect 9218 13696 9274 13705
rect 9218 13631 9274 13640
rect 9128 13456 9180 13462
rect 9128 13398 9180 13404
rect 9324 12850 9352 13738
rect 9600 13394 9628 15302
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9692 12866 9720 15098
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9784 12986 9812 14758
rect 9876 13734 9904 14894
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9968 14618 9996 14758
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10048 14408 10100 14414
rect 10048 14350 10100 14356
rect 10060 14074 10088 14350
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9968 13462 9996 13942
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9312 12844 9364 12850
rect 9692 12838 9812 12866
rect 9312 12786 9364 12792
rect 9680 12776 9732 12782
rect 9310 12744 9366 12753
rect 9680 12718 9732 12724
rect 9310 12679 9366 12688
rect 9126 12608 9182 12617
rect 9126 12543 9182 12552
rect 9140 11218 9168 12543
rect 9324 11354 9352 12679
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9126 10296 9182 10305
rect 9126 10231 9128 10240
rect 9180 10231 9182 10240
rect 9128 10202 9180 10208
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9232 7546 9260 9522
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9324 6186 9352 10746
rect 9416 10674 9444 11494
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9402 10432 9458 10441
rect 9402 10367 9458 10376
rect 9416 8498 9444 10367
rect 9600 10266 9628 12582
rect 9692 12374 9720 12718
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9692 8974 9720 9930
rect 9784 9704 9812 12838
rect 9876 12442 9904 13262
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9862 12064 9918 12073
rect 9862 11999 9918 12008
rect 9876 11762 9904 11999
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9876 10305 9904 11222
rect 9968 10674 9996 12582
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10060 11218 10088 12378
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9862 10296 9918 10305
rect 9862 10231 9918 10240
rect 9784 9676 9904 9704
rect 9770 9616 9826 9625
rect 9770 9551 9826 9560
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9784 8090 9812 9551
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9508 7313 9536 7346
rect 9494 7304 9550 7313
rect 9494 7239 9550 7248
rect 9508 7002 9536 7239
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9876 6458 9904 9676
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 9968 9382 9996 9454
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 10152 8566 10180 19450
rect 10232 19440 10284 19446
rect 10232 19382 10284 19388
rect 10244 18222 10272 19382
rect 10336 18902 10364 20742
rect 11072 20618 11100 21286
rect 11532 21146 11560 25191
rect 11796 24744 11848 24750
rect 11796 24686 11848 24692
rect 11612 24336 11664 24342
rect 11612 24278 11664 24284
rect 11624 21350 11652 24278
rect 11702 24168 11758 24177
rect 11702 24103 11704 24112
rect 11756 24103 11758 24112
rect 11704 24074 11756 24080
rect 11808 23730 11836 24686
rect 11796 23724 11848 23730
rect 11796 23666 11848 23672
rect 11704 22568 11756 22574
rect 11704 22510 11756 22516
rect 11716 22166 11744 22510
rect 11900 22166 11928 26200
rect 12072 25560 12124 25566
rect 12072 25502 12124 25508
rect 12084 23730 12112 25502
rect 12164 24132 12216 24138
rect 12164 24074 12216 24080
rect 12072 23724 12124 23730
rect 12072 23666 12124 23672
rect 11978 23624 12034 23633
rect 11978 23559 12034 23568
rect 11704 22160 11756 22166
rect 11704 22102 11756 22108
rect 11888 22160 11940 22166
rect 11888 22102 11940 22108
rect 11704 21616 11756 21622
rect 11704 21558 11756 21564
rect 11716 21350 11744 21558
rect 11612 21344 11664 21350
rect 11612 21286 11664 21292
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 11520 21140 11572 21146
rect 11520 21082 11572 21088
rect 11336 21004 11388 21010
rect 11336 20946 11388 20952
rect 11152 20868 11204 20874
rect 11152 20810 11204 20816
rect 10612 20590 11100 20618
rect 10508 19236 10560 19242
rect 10508 19178 10560 19184
rect 10324 18896 10376 18902
rect 10324 18838 10376 18844
rect 10520 18601 10548 19178
rect 10506 18592 10562 18601
rect 10506 18527 10562 18536
rect 10232 18216 10284 18222
rect 10232 18158 10284 18164
rect 10244 17320 10272 18158
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10244 17292 10364 17320
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10244 12782 10272 17138
rect 10336 14958 10364 17292
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10428 13433 10456 16934
rect 10520 16114 10548 17478
rect 10612 17134 10640 20590
rect 11164 20058 11192 20810
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10704 19156 10732 19314
rect 10980 19292 11008 19926
rect 11348 19446 11376 20946
rect 11612 20868 11664 20874
rect 11612 20810 11664 20816
rect 11520 20460 11572 20466
rect 11520 20402 11572 20408
rect 11532 19990 11560 20402
rect 11428 19984 11480 19990
rect 11428 19926 11480 19932
rect 11520 19984 11572 19990
rect 11520 19926 11572 19932
rect 11440 19446 11468 19926
rect 11336 19440 11388 19446
rect 11336 19382 11388 19388
rect 11428 19440 11480 19446
rect 11428 19382 11480 19388
rect 11060 19304 11112 19310
rect 10980 19264 11060 19292
rect 11060 19246 11112 19252
rect 11060 19168 11112 19174
rect 10704 19128 11060 19156
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10520 14074 10548 14350
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10414 13424 10470 13433
rect 10324 13388 10376 13394
rect 10414 13359 10470 13368
rect 10324 13330 10376 13336
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10230 12336 10286 12345
rect 10336 12306 10364 13330
rect 10612 13190 10640 15846
rect 10600 13184 10652 13190
rect 10506 13152 10562 13161
rect 10600 13126 10652 13132
rect 10506 13087 10562 13096
rect 10416 12640 10468 12646
rect 10416 12582 10468 12588
rect 10230 12271 10286 12280
rect 10324 12300 10376 12306
rect 10244 11898 10272 12271
rect 10324 12242 10376 12248
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10336 11694 10364 12242
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10140 8560 10192 8566
rect 10140 8502 10192 8508
rect 9954 8256 10010 8265
rect 9954 8191 10010 8200
rect 9968 7410 9996 8191
rect 10046 7984 10102 7993
rect 10046 7919 10048 7928
rect 10100 7919 10102 7928
rect 10048 7890 10100 7896
rect 10244 7886 10272 11086
rect 10428 10130 10456 12582
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10520 9586 10548 13087
rect 10600 12164 10652 12170
rect 10600 12106 10652 12112
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10336 9178 10364 9522
rect 10612 9178 10640 12106
rect 10704 10538 10732 19128
rect 11060 19110 11112 19116
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11058 19000 11114 19009
rect 11058 18935 11060 18944
rect 11112 18935 11114 18944
rect 11060 18906 11112 18912
rect 11152 18692 11204 18698
rect 11152 18634 11204 18640
rect 10876 18352 10928 18358
rect 10876 18294 10928 18300
rect 11060 18352 11112 18358
rect 11060 18294 11112 18300
rect 10888 17785 10916 18294
rect 11072 17898 11100 18294
rect 10980 17870 11100 17898
rect 10980 17814 11008 17870
rect 10968 17808 11020 17814
rect 10874 17776 10930 17785
rect 10968 17750 11020 17756
rect 11164 17746 11192 18634
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 10874 17711 10930 17720
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 10876 17604 10928 17610
rect 10876 17546 10928 17552
rect 10888 16538 10916 17546
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 10980 16794 11008 17138
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 10968 16584 11020 16590
rect 10796 16510 10916 16538
rect 10966 16552 10968 16561
rect 11020 16552 11022 16561
rect 10796 16182 10824 16510
rect 11072 16522 11100 16730
rect 10966 16487 11022 16496
rect 11060 16516 11112 16522
rect 11060 16458 11112 16464
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 10876 16448 10928 16454
rect 11164 16402 11192 16458
rect 10876 16390 10928 16396
rect 10784 16176 10836 16182
rect 10784 16118 10836 16124
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10796 14414 10824 15506
rect 10888 15094 10916 16390
rect 11072 16374 11192 16402
rect 10966 16008 11022 16017
rect 11072 15978 11100 16374
rect 10966 15943 11022 15952
rect 11060 15972 11112 15978
rect 10876 15088 10928 15094
rect 10876 15030 10928 15036
rect 10980 14940 11008 15943
rect 11060 15914 11112 15920
rect 10888 14912 11008 14940
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10796 13394 10824 14350
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10782 11792 10838 11801
rect 10782 11727 10838 11736
rect 10796 11626 10824 11727
rect 10784 11620 10836 11626
rect 10784 11562 10836 11568
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10796 10742 10824 11086
rect 10784 10736 10836 10742
rect 10784 10678 10836 10684
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10888 10198 10916 14912
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 11058 14240 11114 14249
rect 11058 14175 11114 14184
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10980 12442 11008 12718
rect 11072 12617 11100 14175
rect 11164 13394 11192 14486
rect 11256 14482 11284 18022
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11242 14104 11298 14113
rect 11242 14039 11298 14048
rect 11256 13938 11284 14039
rect 11244 13932 11296 13938
rect 11244 13874 11296 13880
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11152 12912 11204 12918
rect 11152 12854 11204 12860
rect 11058 12608 11114 12617
rect 11058 12543 11114 12552
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10980 11830 11008 12038
rect 10968 11824 11020 11830
rect 10968 11766 11020 11772
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 10980 10606 11008 11562
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10876 10192 10928 10198
rect 10876 10134 10928 10140
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 10704 7342 10732 9998
rect 11072 9654 11100 11494
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 11164 7954 11192 12854
rect 11242 12472 11298 12481
rect 11242 12407 11298 12416
rect 11256 11121 11284 12407
rect 11348 11558 11376 19110
rect 11624 17898 11652 20810
rect 11992 20754 12020 23559
rect 12176 23361 12204 24074
rect 12162 23352 12218 23361
rect 12162 23287 12218 23296
rect 12268 22574 12296 26250
rect 12452 24274 12480 26302
rect 12530 26200 12586 26302
rect 13174 26330 13230 27000
rect 13174 26302 13400 26330
rect 13174 26200 13230 26302
rect 12716 24948 12768 24954
rect 12716 24890 12768 24896
rect 12440 24268 12492 24274
rect 12440 24210 12492 24216
rect 12532 23520 12584 23526
rect 12532 23462 12584 23468
rect 12256 22568 12308 22574
rect 12256 22510 12308 22516
rect 12544 22166 12572 23462
rect 12622 23352 12678 23361
rect 12728 23338 12756 24890
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12806 23760 12862 23769
rect 12806 23695 12862 23704
rect 12820 23497 12848 23695
rect 12806 23488 12862 23497
rect 12806 23423 12862 23432
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12728 23310 12848 23338
rect 12622 23287 12678 23296
rect 12636 23089 12664 23287
rect 12622 23080 12678 23089
rect 12622 23015 12678 23024
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 12532 22160 12584 22166
rect 12728 22137 12756 22578
rect 12532 22102 12584 22108
rect 12714 22128 12770 22137
rect 12714 22063 12770 22072
rect 12348 21956 12400 21962
rect 12348 21898 12400 21904
rect 12624 21956 12676 21962
rect 12624 21898 12676 21904
rect 12084 21554 12296 21570
rect 12084 21548 12308 21554
rect 12084 21542 12256 21548
rect 12084 21486 12112 21542
rect 12256 21490 12308 21496
rect 12072 21480 12124 21486
rect 12072 21422 12124 21428
rect 12256 21412 12308 21418
rect 12256 21354 12308 21360
rect 12268 20806 12296 21354
rect 11900 20726 12020 20754
rect 12256 20800 12308 20806
rect 12256 20742 12308 20748
rect 11900 20466 11928 20726
rect 11888 20460 11940 20466
rect 11888 20402 11940 20408
rect 11900 20233 11928 20402
rect 11886 20224 11942 20233
rect 11886 20159 11942 20168
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11440 17870 11652 17898
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11440 11268 11468 17870
rect 11518 17776 11574 17785
rect 11518 17711 11574 17720
rect 11532 14634 11560 17711
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11624 15348 11652 16594
rect 11716 15706 11744 19450
rect 11794 18320 11850 18329
rect 11794 18255 11796 18264
rect 11848 18255 11850 18264
rect 11796 18226 11848 18232
rect 11808 17785 11836 18226
rect 11992 18222 12020 19790
rect 12256 19780 12308 19786
rect 12256 19722 12308 19728
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 12072 19236 12124 19242
rect 12072 19178 12124 19184
rect 12084 18601 12112 19178
rect 12176 19174 12204 19314
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 12164 18692 12216 18698
rect 12164 18634 12216 18640
rect 12070 18592 12126 18601
rect 12070 18527 12126 18536
rect 12176 18426 12204 18634
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 11794 17776 11850 17785
rect 11992 17746 12020 18158
rect 12176 18154 12204 18362
rect 12164 18148 12216 18154
rect 12164 18090 12216 18096
rect 11794 17711 11850 17720
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 12070 17368 12126 17377
rect 12070 17303 12072 17312
rect 12124 17303 12126 17312
rect 12072 17274 12124 17280
rect 11794 17096 11850 17105
rect 11794 17031 11796 17040
rect 11848 17031 11850 17040
rect 11796 17002 11848 17008
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11808 15638 11836 16390
rect 11900 16250 11928 16390
rect 11978 16280 12034 16289
rect 11888 16244 11940 16250
rect 11978 16215 12034 16224
rect 11888 16186 11940 16192
rect 11992 16130 12020 16215
rect 11900 16102 12020 16130
rect 11900 15910 11928 16102
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11900 15484 11928 15846
rect 11808 15456 11928 15484
rect 11704 15360 11756 15366
rect 11624 15320 11704 15348
rect 11704 15302 11756 15308
rect 11716 15026 11744 15302
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11532 14606 11652 14634
rect 11624 13025 11652 14606
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11716 13938 11744 14214
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 11610 13016 11666 13025
rect 11610 12951 11666 12960
rect 11612 12708 11664 12714
rect 11612 12650 11664 12656
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11532 11336 11560 12582
rect 11624 12374 11652 12650
rect 11612 12368 11664 12374
rect 11612 12310 11664 12316
rect 11716 11937 11744 13194
rect 11808 12073 11836 15456
rect 11978 15328 12034 15337
rect 11978 15263 12034 15272
rect 11888 14340 11940 14346
rect 11888 14282 11940 14288
rect 11900 13530 11928 14282
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11900 12866 11928 13330
rect 11992 13161 12020 15263
rect 12084 13326 12112 16934
rect 12176 16726 12204 17682
rect 12164 16720 12216 16726
rect 12164 16662 12216 16668
rect 12164 16176 12216 16182
rect 12164 16118 12216 16124
rect 12176 15910 12204 16118
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 12176 15026 12204 15302
rect 12268 15065 12296 19722
rect 12360 17649 12388 21898
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 12544 21146 12572 21490
rect 12636 21350 12664 21898
rect 12820 21690 12848 23310
rect 13372 23186 13400 26302
rect 13818 26200 13874 27000
rect 14462 26200 14518 27000
rect 15106 26200 15162 27000
rect 15750 26330 15806 27000
rect 15750 26302 15884 26330
rect 15750 26200 15806 26302
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 13832 22574 13860 26200
rect 14188 24676 14240 24682
rect 14188 24618 14240 24624
rect 14004 24200 14056 24206
rect 14004 24142 14056 24148
rect 13820 22568 13872 22574
rect 13820 22510 13872 22516
rect 13912 22500 13964 22506
rect 13912 22442 13964 22448
rect 13358 22400 13414 22409
rect 12950 22332 13258 22341
rect 13358 22335 13414 22344
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12716 21684 12768 21690
rect 12716 21626 12768 21632
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 12728 21350 12756 21626
rect 12624 21344 12676 21350
rect 12624 21286 12676 21292
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12532 21140 12584 21146
rect 12532 21082 12584 21088
rect 12990 20904 13046 20913
rect 12990 20839 13046 20848
rect 13004 20806 13032 20839
rect 12992 20800 13044 20806
rect 12992 20742 13044 20748
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13372 19446 13400 22335
rect 13636 21888 13688 21894
rect 13636 21830 13688 21836
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13648 21593 13676 21830
rect 13634 21584 13690 21593
rect 13634 21519 13690 21528
rect 13740 21321 13768 21830
rect 13726 21312 13782 21321
rect 13726 21247 13782 21256
rect 13832 21162 13860 21830
rect 13924 21486 13952 22442
rect 13912 21480 13964 21486
rect 13912 21422 13964 21428
rect 13832 21134 13952 21162
rect 13544 21004 13596 21010
rect 13544 20946 13596 20952
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 13556 20641 13584 20946
rect 13542 20632 13598 20641
rect 13542 20567 13598 20576
rect 13832 20534 13860 20946
rect 13924 20806 13952 21134
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13820 20528 13872 20534
rect 13820 20470 13872 20476
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 13360 19440 13412 19446
rect 13360 19382 13412 19388
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12452 17921 12480 19110
rect 12530 18864 12586 18873
rect 12530 18799 12586 18808
rect 12544 18601 12572 18799
rect 12530 18592 12586 18601
rect 12530 18527 12586 18536
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12530 18184 12586 18193
rect 12530 18119 12532 18128
rect 12584 18119 12586 18128
rect 12532 18090 12584 18096
rect 12438 17912 12494 17921
rect 12438 17847 12494 17856
rect 12532 17672 12584 17678
rect 12346 17640 12402 17649
rect 12636 17660 12664 18362
rect 12584 17632 12664 17660
rect 12728 18170 12756 19246
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12820 18465 12848 18566
rect 12806 18456 12862 18465
rect 12806 18391 12862 18400
rect 13372 18358 13400 19246
rect 13360 18352 13412 18358
rect 13360 18294 13412 18300
rect 12900 18216 12952 18222
rect 12728 18164 12900 18170
rect 12728 18158 12952 18164
rect 12728 18142 12940 18158
rect 12532 17614 12584 17620
rect 12346 17575 12402 17584
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12452 17241 12480 17274
rect 12438 17232 12494 17241
rect 12438 17167 12494 17176
rect 12348 16448 12400 16454
rect 12348 16390 12400 16396
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12360 15688 12388 16390
rect 12452 16250 12480 16390
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12440 15700 12492 15706
rect 12360 15660 12440 15688
rect 12440 15642 12492 15648
rect 12440 15428 12492 15434
rect 12544 15416 12572 17614
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12636 16794 12664 17070
rect 12728 16810 12756 18142
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13464 17814 13492 20334
rect 13636 20256 13688 20262
rect 13636 20198 13688 20204
rect 13648 19990 13676 20198
rect 13636 19984 13688 19990
rect 13636 19926 13688 19932
rect 13728 19916 13780 19922
rect 13728 19858 13780 19864
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13556 19718 13584 19790
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13648 19145 13676 19654
rect 13740 19242 13768 19858
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 13634 19136 13690 19145
rect 13832 19122 13860 19654
rect 13924 19553 13952 20334
rect 13910 19544 13966 19553
rect 13910 19479 13966 19488
rect 14016 19310 14044 24142
rect 14200 21690 14228 24618
rect 14476 24274 14504 26200
rect 15016 25084 15068 25090
rect 15016 25026 15068 25032
rect 14832 24608 14884 24614
rect 14832 24550 14884 24556
rect 14464 24268 14516 24274
rect 14464 24210 14516 24216
rect 14648 23724 14700 23730
rect 14648 23666 14700 23672
rect 14660 23322 14688 23666
rect 14556 23316 14608 23322
rect 14556 23258 14608 23264
rect 14648 23316 14700 23322
rect 14648 23258 14700 23264
rect 14740 23316 14792 23322
rect 14740 23258 14792 23264
rect 14568 23202 14596 23258
rect 14752 23202 14780 23258
rect 14568 23174 14780 23202
rect 14556 23112 14608 23118
rect 14556 23054 14608 23060
rect 14462 22264 14518 22273
rect 14462 22199 14464 22208
rect 14516 22199 14518 22208
rect 14464 22170 14516 22176
rect 14568 22137 14596 23054
rect 14646 22808 14702 22817
rect 14646 22743 14702 22752
rect 14554 22128 14610 22137
rect 14554 22063 14610 22072
rect 14372 21956 14424 21962
rect 14372 21898 14424 21904
rect 14188 21684 14240 21690
rect 14188 21626 14240 21632
rect 14280 21684 14332 21690
rect 14280 21626 14332 21632
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 14108 20777 14136 20878
rect 14094 20768 14150 20777
rect 14094 20703 14150 20712
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14200 19786 14228 19994
rect 14096 19780 14148 19786
rect 14096 19722 14148 19728
rect 14188 19780 14240 19786
rect 14188 19722 14240 19728
rect 14108 19310 14136 19722
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 13634 19071 13690 19080
rect 13740 19094 13860 19122
rect 13648 18329 13676 19071
rect 13740 18902 13768 19094
rect 14292 18952 14320 21626
rect 14384 21185 14412 21898
rect 14464 21684 14516 21690
rect 14464 21626 14516 21632
rect 14370 21176 14426 21185
rect 14370 21111 14426 21120
rect 14476 21010 14504 21626
rect 14464 21004 14516 21010
rect 14464 20946 14516 20952
rect 14568 20097 14596 22063
rect 14660 22030 14688 22743
rect 14648 22024 14700 22030
rect 14648 21966 14700 21972
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 14752 21457 14780 21490
rect 14738 21448 14794 21457
rect 14738 21383 14794 21392
rect 14648 20868 14700 20874
rect 14648 20810 14700 20816
rect 14554 20088 14610 20097
rect 14554 20023 14610 20032
rect 14554 19952 14610 19961
rect 14554 19887 14610 19896
rect 14568 19854 14596 19887
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14108 18924 14320 18952
rect 13728 18896 13780 18902
rect 13728 18838 13780 18844
rect 13634 18320 13690 18329
rect 13634 18255 13690 18264
rect 13542 17912 13598 17921
rect 13542 17847 13598 17856
rect 13268 17808 13320 17814
rect 13268 17750 13320 17756
rect 13452 17808 13504 17814
rect 13452 17750 13504 17756
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12820 16969 12848 17682
rect 13280 17270 13308 17750
rect 13556 17610 13584 17847
rect 13544 17604 13596 17610
rect 13544 17546 13596 17552
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 12806 16960 12862 16969
rect 12806 16895 12862 16904
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12624 16788 12676 16794
rect 12728 16782 12848 16810
rect 12624 16730 12676 16736
rect 12820 15688 12848 16782
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 12992 16448 13044 16454
rect 12992 16390 13044 16396
rect 13004 16017 13032 16390
rect 13280 16046 13308 16594
rect 13268 16040 13320 16046
rect 12990 16008 13046 16017
rect 13268 15982 13320 15988
rect 12990 15943 13046 15952
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12820 15660 12940 15688
rect 12806 15600 12862 15609
rect 12806 15535 12808 15544
rect 12860 15535 12862 15544
rect 12808 15506 12860 15512
rect 12492 15388 12572 15416
rect 12440 15370 12492 15376
rect 12254 15056 12310 15065
rect 12164 15020 12216 15026
rect 12254 14991 12310 15000
rect 12164 14962 12216 14968
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12176 13190 12204 13670
rect 12164 13184 12216 13190
rect 11978 13152 12034 13161
rect 12164 13126 12216 13132
rect 11978 13087 12034 13096
rect 11900 12838 12204 12866
rect 12176 12782 12204 12838
rect 11888 12776 11940 12782
rect 12164 12776 12216 12782
rect 11940 12736 12020 12764
rect 11888 12718 11940 12724
rect 11992 12442 12020 12736
rect 12164 12718 12216 12724
rect 12072 12708 12124 12714
rect 12072 12650 12124 12656
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11900 12102 11928 12378
rect 12084 12374 12112 12650
rect 12072 12368 12124 12374
rect 12072 12310 12124 12316
rect 11888 12096 11940 12102
rect 11794 12064 11850 12073
rect 11888 12038 11940 12044
rect 11794 11999 11850 12008
rect 11702 11928 11758 11937
rect 11702 11863 11758 11872
rect 11794 11384 11850 11393
rect 11532 11308 11744 11336
rect 11794 11319 11850 11328
rect 11348 11240 11468 11268
rect 11242 11112 11298 11121
rect 11242 11047 11298 11056
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11256 9654 11284 10406
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11348 7970 11376 11240
rect 11518 11112 11574 11121
rect 11518 11047 11574 11056
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11440 8090 11468 10610
rect 11532 8430 11560 11047
rect 11610 10840 11666 10849
rect 11716 10810 11744 11308
rect 11808 11121 11836 11319
rect 11794 11112 11850 11121
rect 11794 11047 11850 11056
rect 11610 10775 11612 10784
rect 11664 10775 11666 10784
rect 11704 10804 11756 10810
rect 11612 10746 11664 10752
rect 11704 10746 11756 10752
rect 11900 10441 11928 12038
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 11886 10432 11942 10441
rect 11886 10367 11942 10376
rect 11610 10160 11666 10169
rect 11610 10095 11666 10104
rect 11624 8838 11652 10095
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11716 8906 11744 9318
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11256 7942 11376 7970
rect 11256 7546 11284 7942
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11348 7585 11376 7822
rect 11334 7576 11390 7585
rect 11244 7540 11296 7546
rect 11334 7511 11336 7520
rect 11244 7482 11296 7488
rect 11388 7511 11390 7520
rect 11336 7482 11388 7488
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 11334 6896 11390 6905
rect 11334 6831 11390 6840
rect 11348 6798 11376 6831
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9600 3194 9628 3470
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 9692 2446 9720 3878
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9784 2650 9812 2926
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9876 2514 9904 4082
rect 11624 3738 11652 8366
rect 11808 6730 11836 9862
rect 11992 9518 12020 11766
rect 12084 10198 12112 11766
rect 12176 10674 12204 12718
rect 12268 12594 12296 14894
rect 12452 14482 12480 15370
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12348 13728 12400 13734
rect 12346 13696 12348 13705
rect 12400 13696 12402 13705
rect 12346 13631 12402 13640
rect 12452 13530 12480 13942
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12360 12782 12388 13126
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12452 12617 12480 13330
rect 12438 12608 12494 12617
rect 12268 12566 12388 12594
rect 12360 12288 12388 12566
rect 12438 12543 12494 12552
rect 12544 12322 12572 14962
rect 12624 14816 12676 14822
rect 12728 14793 12756 15302
rect 12912 15162 12940 15660
rect 13372 15570 13400 17478
rect 13556 16697 13584 17546
rect 13910 17368 13966 17377
rect 13820 17332 13872 17338
rect 13910 17303 13966 17312
rect 13820 17274 13872 17280
rect 13832 16794 13860 17274
rect 13924 17270 13952 17303
rect 13912 17264 13964 17270
rect 13912 17206 13964 17212
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 13542 16688 13598 16697
rect 13542 16623 13598 16632
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13556 16454 13584 16526
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13464 15706 13492 16186
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 13004 15337 13032 15506
rect 12990 15328 13046 15337
rect 12990 15263 13046 15272
rect 13556 15178 13584 16050
rect 13648 15745 13676 16730
rect 13832 16658 13860 16730
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13820 16516 13872 16522
rect 13820 16458 13872 16464
rect 13728 16040 13780 16046
rect 13832 16017 13860 16458
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13728 15982 13780 15988
rect 13818 16008 13874 16017
rect 13634 15736 13690 15745
rect 13634 15671 13690 15680
rect 13636 15360 13688 15366
rect 13634 15328 13636 15337
rect 13688 15328 13690 15337
rect 13634 15263 13690 15272
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 13268 15156 13320 15162
rect 13556 15150 13676 15178
rect 13268 15098 13320 15104
rect 13280 14958 13308 15098
rect 13542 15056 13598 15065
rect 13542 14991 13544 15000
rect 13596 14991 13598 15000
rect 13544 14962 13596 14968
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 12808 14884 12860 14890
rect 12808 14826 12860 14832
rect 12624 14758 12676 14764
rect 12714 14784 12770 14793
rect 12636 12481 12664 14758
rect 12714 14719 12770 14728
rect 12820 13870 12848 14826
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13450 14648 13506 14657
rect 13450 14583 13506 14592
rect 13360 14408 13412 14414
rect 13464 14385 13492 14583
rect 13360 14350 13412 14356
rect 13450 14376 13506 14385
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12728 13530 12756 13670
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12622 12472 12678 12481
rect 12622 12407 12678 12416
rect 12544 12294 12664 12322
rect 12268 12260 12388 12288
rect 12268 11830 12296 12260
rect 12348 12164 12400 12170
rect 12348 12106 12400 12112
rect 12360 11937 12388 12106
rect 12346 11928 12402 11937
rect 12346 11863 12402 11872
rect 12256 11824 12308 11830
rect 12256 11766 12308 11772
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 12268 10962 12296 11154
rect 12360 11082 12388 11863
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 12452 11014 12480 11494
rect 12440 11008 12492 11014
rect 12268 10934 12388 10962
rect 12440 10950 12492 10956
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12072 10192 12124 10198
rect 12072 10134 12124 10140
rect 12176 10062 12204 10406
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12070 9616 12126 9625
rect 12070 9551 12126 9560
rect 12164 9580 12216 9586
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 11992 7886 12020 8298
rect 12084 7954 12112 9551
rect 12164 9522 12216 9528
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11978 7440 12034 7449
rect 11978 7375 11980 7384
rect 12032 7375 12034 7384
rect 11980 7346 12032 7352
rect 11796 6724 11848 6730
rect 11796 6666 11848 6672
rect 12176 5370 12204 9522
rect 12268 9178 12296 10610
rect 12360 10130 12388 10934
rect 12532 10600 12584 10606
rect 12452 10560 12532 10588
rect 12452 10441 12480 10560
rect 12532 10542 12584 10548
rect 12438 10432 12494 10441
rect 12438 10367 12494 10376
rect 12530 10296 12586 10305
rect 12530 10231 12586 10240
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12544 9761 12572 10231
rect 12530 9752 12586 9761
rect 12530 9687 12586 9696
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 12544 7546 12572 9687
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12346 6760 12402 6769
rect 12346 6695 12402 6704
rect 12360 6662 12388 6695
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12636 6390 12664 12294
rect 12728 11218 12756 13126
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12820 11150 12848 13670
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13084 13456 13136 13462
rect 13084 13398 13136 13404
rect 13174 13424 13230 13433
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 13004 12850 13032 13330
rect 13096 12918 13124 13398
rect 13174 13359 13176 13368
rect 13228 13359 13230 13368
rect 13176 13330 13228 13336
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13188 12764 13216 13126
rect 13266 12880 13322 12889
rect 13372 12866 13400 14350
rect 13450 14311 13506 14320
rect 13450 14240 13506 14249
rect 13450 14175 13506 14184
rect 13464 13462 13492 14175
rect 13556 13938 13584 14758
rect 13648 14278 13676 15150
rect 13740 14498 13768 15982
rect 13818 15943 13874 15952
rect 13924 15910 13952 16050
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13924 15570 13952 15846
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13832 14618 13860 14894
rect 13924 14618 13952 15506
rect 14004 15088 14056 15094
rect 14004 15030 14056 15036
rect 14016 14618 14044 15030
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 13740 14470 13860 14498
rect 13726 14376 13782 14385
rect 13726 14311 13782 14320
rect 13636 14272 13688 14278
rect 13634 14240 13636 14249
rect 13688 14240 13690 14249
rect 13634 14175 13690 14184
rect 13740 14074 13768 14311
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13832 13954 13860 14470
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13740 13926 13860 13954
rect 13544 13796 13596 13802
rect 13544 13738 13596 13744
rect 13452 13456 13504 13462
rect 13452 13398 13504 13404
rect 13464 12986 13492 13398
rect 13556 13394 13584 13738
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13322 12838 13400 12866
rect 13450 12880 13506 12889
rect 13266 12815 13322 12824
rect 13450 12815 13452 12824
rect 13504 12815 13506 12824
rect 13452 12786 13504 12792
rect 13188 12736 13400 12764
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13084 12368 13136 12374
rect 13084 12310 13136 12316
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 13004 12170 13032 12242
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 13096 11558 13124 12310
rect 13372 11694 13400 12736
rect 13452 12640 13504 12646
rect 13556 12617 13584 13330
rect 13740 12782 13768 13926
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13452 12582 13504 12588
rect 13542 12608 13598 12617
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12714 10840 12770 10849
rect 13372 10826 13400 11494
rect 12714 10775 12716 10784
rect 12768 10775 12770 10784
rect 12820 10798 13400 10826
rect 12716 10746 12768 10752
rect 12820 10690 12848 10798
rect 12728 10662 12848 10690
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 12728 8430 12756 10662
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12820 10266 12848 10542
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 13268 10056 13320 10062
rect 13372 10044 13400 10678
rect 13464 10130 13492 12582
rect 13542 12543 13598 12552
rect 13544 12300 13596 12306
rect 13648 12288 13676 12650
rect 13596 12260 13676 12288
rect 13544 12242 13596 12248
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13320 10016 13400 10044
rect 13268 9998 13320 10004
rect 13176 9988 13228 9994
rect 13176 9930 13228 9936
rect 13188 9722 13216 9930
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13280 9586 13308 9998
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13268 9444 13320 9450
rect 13372 9432 13400 9862
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13556 9674 13584 12242
rect 13634 12064 13690 12073
rect 13634 11999 13690 12008
rect 13648 10130 13676 11999
rect 13740 11830 13768 12718
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13320 9404 13400 9432
rect 13268 9386 13320 9392
rect 13372 9353 13400 9404
rect 13358 9344 13414 9353
rect 12950 9276 13258 9285
rect 13358 9279 13414 9288
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 13464 9042 13492 9658
rect 13556 9646 13676 9674
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13280 8786 13308 8910
rect 13452 8832 13504 8838
rect 13280 8780 13452 8786
rect 13280 8774 13504 8780
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 13188 8362 13216 8774
rect 13280 8758 13492 8774
rect 13556 8634 13584 9454
rect 13648 9042 13676 9646
rect 13740 9178 13768 11154
rect 13832 10169 13860 12922
rect 13924 12170 13952 14214
rect 14016 12374 14044 14282
rect 14108 13705 14136 18924
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14188 18692 14240 18698
rect 14188 18634 14240 18640
rect 14200 18358 14228 18634
rect 14188 18352 14240 18358
rect 14188 18294 14240 18300
rect 14292 18086 14320 18770
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 14292 17678 14320 18022
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14292 17377 14320 17614
rect 14278 17368 14334 17377
rect 14476 17338 14504 19314
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14278 17303 14334 17312
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14370 16144 14426 16153
rect 14370 16079 14426 16088
rect 14384 15881 14412 16079
rect 14370 15872 14426 15881
rect 14370 15807 14426 15816
rect 14186 15056 14242 15065
rect 14186 14991 14242 15000
rect 14094 13696 14150 13705
rect 14094 13631 14150 13640
rect 14094 13560 14150 13569
rect 14094 13495 14150 13504
rect 14108 13190 14136 13495
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 14004 12164 14056 12170
rect 14004 12106 14056 12112
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13924 11529 13952 11834
rect 13910 11520 13966 11529
rect 13910 11455 13966 11464
rect 14016 11354 14044 12106
rect 14200 11626 14228 14991
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14292 13326 14320 14894
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14292 12850 14320 13262
rect 14384 13258 14412 15807
rect 14476 14074 14504 16390
rect 14568 16182 14596 18634
rect 14660 18426 14688 20810
rect 14844 19446 14872 24550
rect 15028 23730 15056 25026
rect 15120 23798 15148 26200
rect 15200 25016 15252 25022
rect 15200 24958 15252 24964
rect 15212 24206 15240 24958
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 15108 23792 15160 23798
rect 15108 23734 15160 23740
rect 15016 23724 15068 23730
rect 15016 23666 15068 23672
rect 15752 23180 15804 23186
rect 15752 23122 15804 23128
rect 15290 22808 15346 22817
rect 15290 22743 15346 22752
rect 15108 22636 15160 22642
rect 15108 22578 15160 22584
rect 15016 22092 15068 22098
rect 15120 22094 15148 22578
rect 15304 22234 15332 22743
rect 15292 22228 15344 22234
rect 15292 22170 15344 22176
rect 15120 22066 15240 22094
rect 15016 22034 15068 22040
rect 14924 21888 14976 21894
rect 14924 21830 14976 21836
rect 14936 21486 14964 21830
rect 15028 21690 15056 22034
rect 15016 21684 15068 21690
rect 15016 21626 15068 21632
rect 15108 21684 15160 21690
rect 15108 21626 15160 21632
rect 14924 21480 14976 21486
rect 14924 21422 14976 21428
rect 15014 21040 15070 21049
rect 15014 20975 15070 20984
rect 15028 20874 15056 20975
rect 15016 20868 15068 20874
rect 15016 20810 15068 20816
rect 15016 20460 15068 20466
rect 15016 20402 15068 20408
rect 14832 19440 14884 19446
rect 14832 19382 14884 19388
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 14832 19304 14884 19310
rect 14832 19246 14884 19252
rect 14844 18698 14872 19246
rect 14832 18692 14884 18698
rect 14832 18634 14884 18640
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14648 18148 14700 18154
rect 14648 18090 14700 18096
rect 14660 16590 14688 18090
rect 14832 18080 14884 18086
rect 14830 18048 14832 18057
rect 14884 18048 14886 18057
rect 14830 17983 14886 17992
rect 14936 17882 14964 19314
rect 15028 19310 15056 20402
rect 15016 19304 15068 19310
rect 15016 19246 15068 19252
rect 15120 19122 15148 21626
rect 15212 21049 15240 22066
rect 15384 21956 15436 21962
rect 15384 21898 15436 21904
rect 15396 21486 15424 21898
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15384 21480 15436 21486
rect 15384 21422 15436 21428
rect 15198 21040 15254 21049
rect 15198 20975 15254 20984
rect 15382 20632 15438 20641
rect 15382 20567 15438 20576
rect 15396 20330 15424 20567
rect 15384 20324 15436 20330
rect 15384 20266 15436 20272
rect 15200 19848 15252 19854
rect 15198 19816 15200 19825
rect 15252 19816 15254 19825
rect 15198 19751 15254 19760
rect 15580 19514 15608 21490
rect 15764 21350 15792 23122
rect 15856 22710 15884 26302
rect 16394 26200 16450 27000
rect 17038 26200 17094 27000
rect 17682 26200 17738 27000
rect 18326 26200 18382 27000
rect 18970 26200 19026 27000
rect 19614 26200 19670 27000
rect 20258 26200 20314 27000
rect 20902 26330 20958 27000
rect 20902 26302 21312 26330
rect 20902 26200 20958 26302
rect 16302 23760 16358 23769
rect 16302 23695 16358 23704
rect 16316 23066 16344 23695
rect 16408 23186 16436 26200
rect 16946 24304 17002 24313
rect 16946 24239 17002 24248
rect 16960 24206 16988 24239
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 16764 24064 16816 24070
rect 16764 24006 16816 24012
rect 16776 23594 16804 24006
rect 16854 23760 16910 23769
rect 16854 23695 16856 23704
rect 16908 23695 16910 23704
rect 16856 23666 16908 23672
rect 16672 23588 16724 23594
rect 16672 23530 16724 23536
rect 16764 23588 16816 23594
rect 16764 23530 16816 23536
rect 16578 23216 16634 23225
rect 16396 23180 16448 23186
rect 16578 23151 16634 23160
rect 16396 23122 16448 23128
rect 16592 23118 16620 23151
rect 16580 23112 16632 23118
rect 16316 23038 16436 23066
rect 16580 23054 16632 23060
rect 15844 22704 15896 22710
rect 15844 22646 15896 22652
rect 16028 22500 16080 22506
rect 16028 22442 16080 22448
rect 16040 22234 16068 22442
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 16028 22228 16080 22234
rect 16028 22170 16080 22176
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 15672 20777 15700 21286
rect 15658 20768 15714 20777
rect 15658 20703 15714 20712
rect 15764 20534 15792 21286
rect 15856 20942 15884 21490
rect 16028 21004 16080 21010
rect 16028 20946 16080 20952
rect 15844 20936 15896 20942
rect 15844 20878 15896 20884
rect 15752 20528 15804 20534
rect 15752 20470 15804 20476
rect 15856 20466 15884 20878
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 16040 19825 16068 20946
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 16118 20496 16174 20505
rect 16118 20431 16120 20440
rect 16172 20431 16174 20440
rect 16120 20402 16172 20408
rect 16026 19816 16082 19825
rect 16026 19751 16082 19760
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15028 19094 15148 19122
rect 15028 18873 15056 19094
rect 15106 19000 15162 19009
rect 15106 18935 15108 18944
rect 15160 18935 15162 18944
rect 15108 18906 15160 18912
rect 15014 18864 15070 18873
rect 15014 18799 15070 18808
rect 15016 18692 15068 18698
rect 15016 18634 15068 18640
rect 14740 17876 14792 17882
rect 14740 17818 14792 17824
rect 14924 17876 14976 17882
rect 14924 17818 14976 17824
rect 14752 17542 14780 17818
rect 15028 17610 15056 18634
rect 15016 17604 15068 17610
rect 15016 17546 15068 17552
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 14738 16824 14794 16833
rect 14738 16759 14794 16768
rect 14752 16590 14780 16759
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 15028 16454 15056 17138
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 15120 16697 15148 16934
rect 15106 16688 15162 16697
rect 15106 16623 15162 16632
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 14556 16176 14608 16182
rect 14556 16118 14608 16124
rect 14738 16144 14794 16153
rect 14738 16079 14740 16088
rect 14792 16079 14794 16088
rect 14740 16050 14792 16056
rect 14740 15904 14792 15910
rect 14740 15846 14792 15852
rect 14752 15570 14780 15846
rect 14740 15564 14792 15570
rect 14740 15506 14792 15512
rect 14844 15178 14872 16186
rect 15120 16046 15148 16526
rect 15212 16425 15240 19246
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 15198 16416 15254 16425
rect 15198 16351 15254 16360
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15304 15706 15332 18158
rect 15396 16250 15424 19314
rect 15488 17338 15516 19450
rect 16224 19394 16252 20742
rect 16316 20534 16344 22374
rect 16304 20528 16356 20534
rect 16304 20470 16356 20476
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16316 19718 16344 19858
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 16132 19366 16252 19394
rect 16040 19281 16068 19314
rect 16132 19310 16160 19366
rect 16120 19304 16172 19310
rect 16026 19272 16082 19281
rect 16120 19246 16172 19252
rect 16026 19207 16082 19216
rect 16040 18737 16068 19207
rect 16210 19136 16266 19145
rect 16210 19071 16266 19080
rect 16026 18728 16082 18737
rect 16026 18663 16082 18672
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 15658 18456 15714 18465
rect 15658 18391 15714 18400
rect 15568 18284 15620 18290
rect 15568 18226 15620 18232
rect 15580 18057 15608 18226
rect 15566 18048 15622 18057
rect 15566 17983 15622 17992
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 14752 15162 14872 15178
rect 14740 15156 14872 15162
rect 14792 15150 14872 15156
rect 14740 15098 14792 15104
rect 14830 15056 14886 15065
rect 14830 14991 14886 15000
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14568 14074 14596 14554
rect 14660 14482 14688 14554
rect 14844 14482 14872 14991
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14832 14476 14884 14482
rect 14832 14418 14884 14424
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14372 13252 14424 13258
rect 14372 13194 14424 13200
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14292 12238 14320 12786
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14476 12073 14504 13670
rect 14660 12442 14688 14214
rect 14844 13376 14872 14418
rect 14936 14226 14964 15506
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 15014 14240 15070 14249
rect 14936 14198 15014 14226
rect 15014 14175 15070 14184
rect 15028 13870 15056 14175
rect 15212 13938 15240 15302
rect 15488 14362 15516 17138
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15580 16017 15608 16186
rect 15566 16008 15622 16017
rect 15566 15943 15622 15952
rect 15672 14906 15700 18391
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15856 17490 15884 18158
rect 15936 17536 15988 17542
rect 15856 17484 15936 17490
rect 15856 17478 15988 17484
rect 15856 17462 15976 17478
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15764 16658 15792 17070
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15752 15632 15804 15638
rect 15752 15574 15804 15580
rect 15764 15366 15792 15574
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15856 15201 15884 17462
rect 16132 17134 16160 18566
rect 16224 18222 16252 19071
rect 16302 18456 16358 18465
rect 16302 18391 16358 18400
rect 16316 18290 16344 18391
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 16408 18086 16436 23038
rect 16684 22094 16712 23530
rect 16960 23497 16988 24142
rect 17052 23798 17080 26200
rect 17316 25288 17368 25294
rect 17316 25230 17368 25236
rect 17132 24200 17184 24206
rect 17132 24142 17184 24148
rect 17040 23792 17092 23798
rect 17040 23734 17092 23740
rect 16946 23488 17002 23497
rect 16946 23423 17002 23432
rect 17144 23361 17172 24142
rect 17328 23730 17356 25230
rect 17316 23724 17368 23730
rect 17236 23684 17316 23712
rect 17130 23352 17186 23361
rect 17236 23322 17264 23684
rect 17316 23666 17368 23672
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17130 23287 17186 23296
rect 17224 23316 17276 23322
rect 17224 23258 17276 23264
rect 17040 23248 17092 23254
rect 17040 23190 17092 23196
rect 16764 23180 16816 23186
rect 16764 23122 16816 23128
rect 16776 22982 16804 23122
rect 16764 22976 16816 22982
rect 16764 22918 16816 22924
rect 16592 22066 16712 22094
rect 16486 21720 16542 21729
rect 16486 21655 16542 21664
rect 16500 20233 16528 21655
rect 16592 20346 16620 22066
rect 16776 22030 16804 22918
rect 16856 22568 16908 22574
rect 16856 22510 16908 22516
rect 16868 22166 16896 22510
rect 16856 22160 16908 22166
rect 16856 22102 16908 22108
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16764 22024 16816 22030
rect 16764 21966 16816 21972
rect 16684 21554 16712 21966
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 16762 21448 16818 21457
rect 16762 21383 16818 21392
rect 16776 20874 16804 21383
rect 16764 20868 16816 20874
rect 16764 20810 16816 20816
rect 16672 20800 16724 20806
rect 16672 20742 16724 20748
rect 16684 20448 16712 20742
rect 16868 20466 16896 22102
rect 17052 22094 17080 23190
rect 17132 23112 17184 23118
rect 17132 23054 17184 23060
rect 17144 22778 17172 23054
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17408 22160 17460 22166
rect 17408 22102 17460 22108
rect 17052 22066 17172 22094
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 16960 21457 16988 21490
rect 16946 21448 17002 21457
rect 16946 21383 17002 21392
rect 16960 21146 16988 21383
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 16948 20800 17000 20806
rect 16946 20768 16948 20777
rect 17000 20768 17002 20777
rect 16946 20703 17002 20712
rect 16856 20460 16908 20466
rect 16684 20420 16804 20448
rect 16592 20318 16712 20346
rect 16486 20224 16542 20233
rect 16486 20159 16542 20168
rect 16488 19780 16540 19786
rect 16488 19722 16540 19728
rect 16500 18698 16528 19722
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 16488 18692 16540 18698
rect 16488 18634 16540 18640
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16028 17128 16080 17134
rect 16026 17096 16028 17105
rect 16120 17128 16172 17134
rect 16080 17096 16082 17105
rect 16120 17070 16172 17076
rect 16304 17128 16356 17134
rect 16304 17070 16356 17076
rect 16026 17031 16082 17040
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 16040 16425 16068 16730
rect 16132 16726 16160 17070
rect 16212 17060 16264 17066
rect 16212 17002 16264 17008
rect 16224 16726 16252 17002
rect 16120 16720 16172 16726
rect 16120 16662 16172 16668
rect 16212 16720 16264 16726
rect 16212 16662 16264 16668
rect 16026 16416 16082 16425
rect 16026 16351 16082 16360
rect 16026 16280 16082 16289
rect 15948 16224 16026 16232
rect 15948 16204 16028 16224
rect 15948 16017 15976 16204
rect 16080 16215 16082 16224
rect 16028 16186 16080 16192
rect 16316 16046 16344 17070
rect 16396 16516 16448 16522
rect 16396 16458 16448 16464
rect 16408 16250 16436 16458
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16120 16040 16172 16046
rect 15934 16008 15990 16017
rect 16120 15982 16172 15988
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 15934 15943 15990 15952
rect 16132 15722 16160 15982
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16040 15694 16160 15722
rect 16210 15736 16266 15745
rect 16040 15570 16068 15694
rect 16210 15671 16266 15680
rect 16120 15632 16172 15638
rect 16120 15574 16172 15580
rect 16028 15564 16080 15570
rect 15948 15524 16028 15552
rect 15842 15192 15898 15201
rect 15842 15127 15898 15136
rect 15844 14952 15896 14958
rect 15672 14878 15792 14906
rect 15844 14894 15896 14900
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15396 14334 15516 14362
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14844 13348 14964 13376
rect 14832 13252 14884 13258
rect 14832 13194 14884 13200
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14462 12064 14518 12073
rect 14462 11999 14518 12008
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14370 11792 14426 11801
rect 14280 11756 14332 11762
rect 14370 11727 14426 11736
rect 14280 11698 14332 11704
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 13924 10266 13952 11018
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13818 10160 13874 10169
rect 13818 10095 13874 10104
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12716 7472 12768 7478
rect 12716 7414 12768 7420
rect 12728 7002 12756 7414
rect 12820 7410 12848 8230
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12624 6384 12676 6390
rect 12624 6326 12676 6332
rect 13648 6254 13676 8842
rect 13726 8528 13782 8537
rect 13726 8463 13782 8472
rect 13740 8430 13768 8463
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13726 6896 13782 6905
rect 13726 6831 13728 6840
rect 13780 6831 13782 6840
rect 13728 6802 13780 6808
rect 12348 6248 12400 6254
rect 12346 6216 12348 6225
rect 13636 6248 13688 6254
rect 12400 6216 12402 6225
rect 13636 6190 13688 6196
rect 12346 6151 12402 6160
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 13832 5574 13860 9862
rect 13924 9636 13952 10202
rect 14004 9648 14056 9654
rect 13924 9608 14004 9636
rect 14004 9590 14056 9596
rect 14200 8634 14228 11018
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 14188 8628 14240 8634
rect 14188 8570 14240 8576
rect 14016 5846 14044 8570
rect 14094 7848 14150 7857
rect 14094 7783 14150 7792
rect 14108 7546 14136 7783
rect 14188 7744 14240 7750
rect 14292 7732 14320 11698
rect 14384 8634 14412 11727
rect 14476 11354 14504 11834
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14476 9994 14504 10542
rect 14464 9988 14516 9994
rect 14464 9930 14516 9936
rect 14568 9625 14596 12242
rect 14646 12064 14702 12073
rect 14646 11999 14702 12008
rect 14660 11218 14688 11999
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14554 9616 14610 9625
rect 14554 9551 14610 9560
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14568 8498 14596 9318
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14240 7704 14320 7732
rect 14188 7686 14240 7692
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14108 6662 14136 7482
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 10060 2650 10088 3470
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10520 3058 10548 3334
rect 10704 3126 10732 3334
rect 11164 3194 11192 3470
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 12360 3058 12388 3334
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 10244 2446 10272 2790
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 8772 1766 8800 2382
rect 8760 1760 8812 1766
rect 8760 1702 8812 1708
rect 9588 1760 9640 1766
rect 9588 1702 9640 1708
rect 9600 800 9628 1702
rect 11716 800 11744 2450
rect 12452 2446 12480 3334
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 13832 800 13860 2450
rect 14200 2310 14228 7686
rect 14278 6760 14334 6769
rect 14278 6695 14334 6704
rect 14292 6662 14320 6695
rect 14660 6662 14688 10950
rect 14752 8090 14780 12378
rect 14844 11354 14872 13194
rect 14936 12356 14964 13348
rect 15304 13274 15332 14282
rect 15396 13462 15424 14334
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15488 14074 15516 14214
rect 15672 14074 15700 14758
rect 15764 14278 15792 14878
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 15476 14068 15528 14074
rect 15660 14068 15712 14074
rect 15476 14010 15528 14016
rect 15580 14028 15660 14056
rect 15580 13569 15608 14028
rect 15660 14010 15712 14016
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15566 13560 15622 13569
rect 15488 13518 15566 13546
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 15120 13246 15332 13274
rect 15120 12986 15148 13246
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 14936 12328 15056 12356
rect 15028 11914 15056 12328
rect 15212 12209 15240 13126
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15198 12200 15254 12209
rect 15198 12135 15254 12144
rect 15028 11886 15240 11914
rect 14922 11792 14978 11801
rect 14922 11727 14924 11736
rect 14976 11727 14978 11736
rect 14924 11698 14976 11704
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 15028 11529 15056 11630
rect 15014 11520 15070 11529
rect 15014 11455 15070 11464
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 15212 11286 15240 11886
rect 15304 11830 15332 12242
rect 15292 11824 15344 11830
rect 15292 11766 15344 11772
rect 14924 11280 14976 11286
rect 14924 11222 14976 11228
rect 15200 11280 15252 11286
rect 15200 11222 15252 11228
rect 14832 9988 14884 9994
rect 14832 9930 14884 9936
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14844 7342 14872 9930
rect 14936 9042 14964 11222
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 15028 8922 15056 9522
rect 15120 8974 15148 10610
rect 15212 10606 15240 11222
rect 15304 10742 15332 11766
rect 15488 11336 15516 13518
rect 15566 13495 15622 13504
rect 15566 13424 15622 13433
rect 15566 13359 15622 13368
rect 15580 11694 15608 13359
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15396 11308 15516 11336
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 14936 8894 15056 8922
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15212 8906 15240 10406
rect 15304 10266 15332 10678
rect 15396 10441 15424 11308
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15382 10432 15438 10441
rect 15382 10367 15438 10376
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15304 9994 15332 10202
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15488 9586 15516 11154
rect 15580 10810 15608 11630
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15304 9178 15332 9318
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15200 8900 15252 8906
rect 14936 8838 14964 8894
rect 15200 8842 15252 8848
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14568 6322 14596 6598
rect 14924 6384 14976 6390
rect 14924 6326 14976 6332
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14936 6118 14964 6326
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 15028 5302 15056 8774
rect 15198 8664 15254 8673
rect 15198 8599 15254 8608
rect 15212 8022 15240 8599
rect 15200 8016 15252 8022
rect 15106 7984 15162 7993
rect 15200 7958 15252 7964
rect 15106 7919 15162 7928
rect 15120 7002 15148 7919
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15212 7546 15240 7822
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 15304 6798 15332 9114
rect 15396 8974 15424 9318
rect 15488 9178 15516 9522
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15580 9042 15608 10134
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15580 8634 15608 8978
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15672 8514 15700 13874
rect 15764 11812 15792 13942
rect 15856 12986 15884 14894
rect 15948 14074 15976 15524
rect 16028 15506 16080 15512
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 16040 14618 16068 14962
rect 16132 14958 16160 15574
rect 16224 15094 16252 15671
rect 16212 15088 16264 15094
rect 16212 15030 16264 15036
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 16040 14498 16068 14554
rect 16040 14470 16160 14498
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15856 12238 15884 12718
rect 16040 12714 16068 13466
rect 16132 12850 16160 14470
rect 16224 14414 16252 15030
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 16040 11898 16068 12650
rect 16118 12472 16174 12481
rect 16118 12407 16174 12416
rect 16132 12374 16160 12407
rect 16120 12368 16172 12374
rect 16120 12310 16172 12316
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 15764 11784 15976 11812
rect 15842 11520 15898 11529
rect 15842 11455 15898 11464
rect 15856 11121 15884 11455
rect 15842 11112 15898 11121
rect 15842 11047 15898 11056
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15764 9722 15792 10950
rect 15842 10568 15898 10577
rect 15842 10503 15898 10512
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15856 9602 15884 10503
rect 15580 8486 15700 8514
rect 15764 9574 15884 9602
rect 15580 8430 15608 8486
rect 15568 8424 15620 8430
rect 15568 8366 15620 8372
rect 15764 7478 15792 9574
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15752 7472 15804 7478
rect 15752 7414 15804 7420
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15580 6866 15608 7346
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15856 5778 15884 8434
rect 15948 6322 15976 11784
rect 16224 11694 16252 14010
rect 16316 14006 16344 15846
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16408 15162 16436 15438
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 16408 14793 16436 14962
rect 16394 14784 16450 14793
rect 16394 14719 16450 14728
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16304 14000 16356 14006
rect 16304 13942 16356 13948
rect 16304 12164 16356 12170
rect 16304 12106 16356 12112
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 16118 11112 16174 11121
rect 16118 11047 16120 11056
rect 16172 11047 16174 11056
rect 16120 11018 16172 11024
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16026 9752 16082 9761
rect 16026 9687 16082 9696
rect 16040 9110 16068 9687
rect 16028 9104 16080 9110
rect 16028 9046 16080 9052
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15016 5296 15068 5302
rect 15016 5238 15068 5244
rect 16132 2774 16160 9998
rect 16224 9722 16252 10202
rect 16316 10130 16344 12106
rect 16408 11150 16436 14010
rect 16500 13258 16528 18634
rect 16592 16590 16620 19314
rect 16684 18970 16712 20318
rect 16776 19417 16804 20420
rect 16856 20402 16908 20408
rect 16868 19922 16896 20402
rect 16856 19916 16908 19922
rect 16856 19858 16908 19864
rect 16762 19408 16818 19417
rect 16818 19352 16896 19360
rect 16762 19343 16896 19352
rect 16776 19332 16896 19343
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 16592 15065 16620 15914
rect 16684 15366 16712 17478
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16578 15056 16634 15065
rect 16578 14991 16634 15000
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16580 13728 16632 13734
rect 16684 13716 16712 14962
rect 16776 14482 16804 16526
rect 16868 16454 16896 19332
rect 17144 19145 17172 22066
rect 17316 22024 17368 22030
rect 17316 21966 17368 21972
rect 17224 21956 17276 21962
rect 17224 21898 17276 21904
rect 17236 21622 17264 21898
rect 17224 21616 17276 21622
rect 17224 21558 17276 21564
rect 17328 21486 17356 21966
rect 17316 21480 17368 21486
rect 17316 21422 17368 21428
rect 17224 21344 17276 21350
rect 17224 21286 17276 21292
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 17236 21146 17264 21286
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 17328 20942 17356 21286
rect 17420 21010 17448 22102
rect 17512 22030 17540 23462
rect 17590 22128 17646 22137
rect 17696 22098 17724 26200
rect 18340 24138 18368 26200
rect 18328 24132 18380 24138
rect 18328 24074 18380 24080
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18788 23860 18840 23866
rect 18788 23802 18840 23808
rect 18418 23352 18474 23361
rect 17868 23316 17920 23322
rect 18418 23287 18474 23296
rect 18694 23352 18750 23361
rect 18694 23287 18750 23296
rect 17868 23258 17920 23264
rect 17880 22710 17908 23258
rect 18328 22976 18380 22982
rect 18328 22918 18380 22924
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17868 22704 17920 22710
rect 17868 22646 17920 22652
rect 18142 22672 18198 22681
rect 17590 22063 17646 22072
rect 17684 22092 17736 22098
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17500 21888 17552 21894
rect 17498 21856 17500 21865
rect 17552 21856 17554 21865
rect 17498 21791 17554 21800
rect 17408 21004 17460 21010
rect 17408 20946 17460 20952
rect 17316 20936 17368 20942
rect 17512 20890 17540 21791
rect 17604 21418 17632 22063
rect 17684 22034 17736 22040
rect 17880 22030 17908 22646
rect 18142 22607 18198 22616
rect 18156 22574 18184 22607
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 18144 21616 18196 21622
rect 18142 21584 18144 21593
rect 18196 21584 18198 21593
rect 18142 21519 18198 21528
rect 17684 21480 17736 21486
rect 17684 21422 17736 21428
rect 17868 21480 17920 21486
rect 17868 21422 17920 21428
rect 18236 21480 18288 21486
rect 18340 21468 18368 22918
rect 18432 22681 18460 23287
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 18418 22672 18474 22681
rect 18524 22642 18552 23054
rect 18418 22607 18474 22616
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18288 21440 18368 21468
rect 18524 21604 18552 22578
rect 18604 22432 18656 22438
rect 18604 22374 18656 22380
rect 18616 22234 18644 22374
rect 18604 22228 18656 22234
rect 18604 22170 18656 22176
rect 18604 21616 18656 21622
rect 18524 21576 18604 21604
rect 18236 21422 18288 21428
rect 17592 21412 17644 21418
rect 17592 21354 17644 21360
rect 17696 21298 17724 21422
rect 17316 20878 17368 20884
rect 17420 20862 17540 20890
rect 17604 21270 17724 21298
rect 17130 19136 17186 19145
rect 17130 19071 17186 19080
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 16868 16182 16896 16390
rect 16856 16176 16908 16182
rect 16856 16118 16908 16124
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 16868 14618 16896 15506
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16764 14340 16816 14346
rect 16764 14282 16816 14288
rect 16632 13688 16712 13716
rect 16580 13670 16632 13676
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 16500 12238 16528 13194
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16486 11112 16542 11121
rect 16486 11047 16542 11056
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 16224 9042 16252 9454
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 16224 8401 16252 8978
rect 16210 8392 16266 8401
rect 16210 8327 16266 8336
rect 16316 7886 16344 10066
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16408 8634 16436 9522
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16500 8514 16528 11047
rect 16592 10606 16620 13670
rect 16776 12986 16804 14282
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16868 12306 16896 14350
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16592 10266 16620 10542
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16408 8486 16528 8514
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16224 3534 16252 4014
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16316 3194 16344 7822
rect 16408 6934 16436 8486
rect 16488 8356 16540 8362
rect 16684 8344 16712 11494
rect 16776 9586 16804 11494
rect 16856 11280 16908 11286
rect 16960 11257 16988 18566
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17328 18193 17356 18362
rect 17314 18184 17370 18193
rect 17314 18119 17370 18128
rect 17222 17776 17278 17785
rect 17040 17740 17092 17746
rect 17222 17711 17278 17720
rect 17040 17682 17092 17688
rect 17052 17270 17080 17682
rect 17132 17604 17184 17610
rect 17132 17546 17184 17552
rect 17040 17264 17092 17270
rect 17040 17206 17092 17212
rect 17144 17184 17172 17546
rect 17236 17513 17264 17711
rect 17316 17536 17368 17542
rect 17222 17504 17278 17513
rect 17316 17478 17368 17484
rect 17222 17439 17278 17448
rect 17144 17156 17264 17184
rect 17236 15994 17264 17156
rect 17328 16697 17356 17478
rect 17314 16688 17370 16697
rect 17314 16623 17370 16632
rect 17420 16574 17448 20862
rect 17604 20262 17632 21270
rect 17592 20256 17644 20262
rect 17592 20198 17644 20204
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 17512 18222 17540 18634
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 17512 17377 17540 18158
rect 17498 17368 17554 17377
rect 17498 17303 17554 17312
rect 17512 17270 17540 17303
rect 17500 17264 17552 17270
rect 17500 17206 17552 17212
rect 17604 17082 17632 20198
rect 17880 20058 17908 21422
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18524 20466 18552 21576
rect 18604 21558 18656 21564
rect 18708 21010 18736 23287
rect 18800 21486 18828 23802
rect 18984 23798 19012 26200
rect 19628 25378 19656 26200
rect 19708 25968 19760 25974
rect 19708 25910 19760 25916
rect 19352 25350 19656 25378
rect 19352 24290 19380 25350
rect 19432 24404 19484 24410
rect 19432 24346 19484 24352
rect 19260 24274 19380 24290
rect 19248 24268 19380 24274
rect 19300 24262 19380 24268
rect 19248 24210 19300 24216
rect 19248 24132 19300 24138
rect 19248 24074 19300 24080
rect 18972 23792 19024 23798
rect 18972 23734 19024 23740
rect 19260 23662 19288 24074
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 19062 22944 19118 22953
rect 19062 22879 19118 22888
rect 18970 22808 19026 22817
rect 18970 22743 19026 22752
rect 18878 22536 18934 22545
rect 18984 22522 19012 22743
rect 18934 22494 19012 22522
rect 18878 22471 18934 22480
rect 18892 22438 18920 22471
rect 18880 22432 18932 22438
rect 19076 22409 19104 22879
rect 19260 22778 19288 23598
rect 19248 22772 19300 22778
rect 19248 22714 19300 22720
rect 19260 22642 19288 22714
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 18880 22374 18932 22380
rect 19062 22400 19118 22409
rect 19062 22335 19118 22344
rect 19444 22030 19472 24346
rect 19720 24177 19748 25910
rect 19892 24880 19944 24886
rect 19892 24822 19944 24828
rect 20074 24848 20130 24857
rect 19706 24168 19762 24177
rect 19706 24103 19708 24112
rect 19760 24103 19762 24112
rect 19708 24074 19760 24080
rect 19524 23588 19576 23594
rect 19524 23530 19576 23536
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19352 21729 19380 21830
rect 19338 21720 19394 21729
rect 19338 21655 19394 21664
rect 18788 21480 18840 21486
rect 18788 21422 18840 21428
rect 18800 21010 18828 21422
rect 19156 21412 19208 21418
rect 19156 21354 19208 21360
rect 18696 21004 18748 21010
rect 18696 20946 18748 20952
rect 18788 21004 18840 21010
rect 18788 20946 18840 20952
rect 19168 20913 19196 21354
rect 19154 20904 19210 20913
rect 19154 20839 19210 20848
rect 19248 20868 19300 20874
rect 19248 20810 19300 20816
rect 19064 20800 19116 20806
rect 19064 20742 19116 20748
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 18524 20330 18552 20402
rect 18512 20324 18564 20330
rect 18512 20266 18564 20272
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17880 19378 17908 19994
rect 18420 19848 18472 19854
rect 18524 19836 18552 20266
rect 18880 20256 18932 20262
rect 18602 20224 18658 20233
rect 18880 20198 18932 20204
rect 18602 20159 18658 20168
rect 18472 19808 18552 19836
rect 18420 19790 18472 19796
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18524 19446 18552 19808
rect 18616 19689 18644 20159
rect 18786 20088 18842 20097
rect 18786 20023 18842 20032
rect 18602 19680 18658 19689
rect 18602 19615 18658 19624
rect 18512 19440 18564 19446
rect 18512 19382 18564 19388
rect 17868 19372 17920 19378
rect 18616 19334 18644 19615
rect 17868 19314 17920 19320
rect 18432 19306 18644 19334
rect 17774 19272 17830 19281
rect 17774 19207 17830 19216
rect 17960 19236 18012 19242
rect 17788 18601 17816 19207
rect 17960 19178 18012 19184
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17774 18592 17830 18601
rect 17774 18527 17830 18536
rect 17880 18290 17908 19110
rect 17972 18834 18000 19178
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17958 18320 18014 18329
rect 17868 18284 17920 18290
rect 17958 18255 18014 18264
rect 17868 18226 17920 18232
rect 17972 18086 18000 18255
rect 17960 18080 18012 18086
rect 17774 18048 17830 18057
rect 17960 18022 18012 18028
rect 17774 17983 17830 17992
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17144 15966 17264 15994
rect 17328 16546 17448 16574
rect 17512 17054 17632 17082
rect 17144 15745 17172 15966
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17130 15736 17186 15745
rect 17130 15671 17186 15680
rect 17236 15366 17264 15846
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 17052 14929 17080 14962
rect 17038 14920 17094 14929
rect 17038 14855 17094 14864
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 17052 13870 17080 14350
rect 17144 13938 17172 15302
rect 17222 14920 17278 14929
rect 17222 14855 17278 14864
rect 17236 13977 17264 14855
rect 17222 13968 17278 13977
rect 17132 13932 17184 13938
rect 17222 13903 17278 13912
rect 17132 13874 17184 13880
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 17328 13682 17356 16546
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17420 15570 17448 15982
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 17144 13654 17356 13682
rect 17144 12434 17172 13654
rect 17144 12406 17356 12434
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 16856 11222 16908 11228
rect 16946 11248 17002 11257
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16684 8316 16804 8344
rect 16488 8298 16540 8304
rect 16396 6928 16448 6934
rect 16396 6870 16448 6876
rect 16500 6390 16528 8298
rect 16670 8256 16726 8265
rect 16670 8191 16726 8200
rect 16580 7812 16632 7818
rect 16580 7754 16632 7760
rect 16592 6458 16620 7754
rect 16684 7546 16712 8191
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16776 7342 16804 8316
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16670 7168 16726 7177
rect 16670 7103 16726 7112
rect 16684 6769 16712 7103
rect 16868 6866 16896 11222
rect 16946 11183 17002 11192
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16960 10266 16988 10950
rect 16948 10260 17000 10266
rect 16948 10202 17000 10208
rect 16948 9716 17000 9722
rect 16948 9658 17000 9664
rect 16960 8906 16988 9658
rect 16948 8900 17000 8906
rect 16948 8842 17000 8848
rect 16960 8378 16988 8842
rect 17052 8537 17080 12310
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17144 9722 17172 10406
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17038 8528 17094 8537
rect 17038 8463 17094 8472
rect 16960 8350 17080 8378
rect 17052 7818 17080 8350
rect 17040 7812 17092 7818
rect 17040 7754 17092 7760
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 16670 6760 16726 6769
rect 16670 6695 16726 6704
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16488 6384 16540 6390
rect 16488 6326 16540 6332
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16040 2746 16160 2774
rect 16040 2582 16068 2746
rect 16028 2576 16080 2582
rect 16028 2518 16080 2524
rect 16408 2446 16436 3334
rect 17052 3194 17080 7754
rect 17144 6866 17172 9454
rect 17236 8809 17264 11494
rect 17328 11200 17356 12406
rect 17420 12102 17448 15302
rect 17512 12850 17540 17054
rect 17590 16552 17646 16561
rect 17590 16487 17646 16496
rect 17604 15910 17632 16487
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17590 15328 17646 15337
rect 17590 15263 17646 15272
rect 17604 14362 17632 15263
rect 17696 14618 17724 17478
rect 17788 16794 17816 17983
rect 18340 17898 18368 18566
rect 17880 17870 18368 17898
rect 17880 16794 17908 17870
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 17972 17649 18000 17682
rect 17958 17640 18014 17649
rect 17958 17575 18014 17584
rect 18326 17640 18382 17649
rect 18326 17575 18328 17584
rect 18380 17575 18382 17584
rect 18328 17546 18380 17552
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17972 16998 18000 17206
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 17972 16794 18000 16934
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 17788 16182 17816 16730
rect 18064 16726 18092 16934
rect 18052 16720 18104 16726
rect 17958 16688 18014 16697
rect 18432 16708 18460 19306
rect 18602 19136 18658 19145
rect 18602 19071 18658 19080
rect 18510 17912 18566 17921
rect 18510 17847 18566 17856
rect 18524 17513 18552 17847
rect 18510 17504 18566 17513
rect 18510 17439 18566 17448
rect 18616 17354 18644 19071
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18524 17326 18644 17354
rect 18524 17066 18552 17326
rect 18708 17202 18736 18362
rect 18800 17921 18828 20023
rect 18892 18834 18920 20198
rect 18880 18828 18932 18834
rect 18880 18770 18932 18776
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18786 17912 18842 17921
rect 18786 17847 18842 17856
rect 18788 17604 18840 17610
rect 18788 17546 18840 17552
rect 18696 17196 18748 17202
rect 18616 17156 18696 17184
rect 18512 17060 18564 17066
rect 18512 17002 18564 17008
rect 18432 16680 18552 16708
rect 18052 16662 18104 16668
rect 17958 16623 17960 16632
rect 18012 16623 18014 16632
rect 17960 16594 18012 16600
rect 17868 16516 17920 16522
rect 17868 16458 17920 16464
rect 17776 16176 17828 16182
rect 17776 16118 17828 16124
rect 17880 15978 17908 16458
rect 18236 16448 18288 16454
rect 18288 16408 18368 16436
rect 18236 16390 18288 16396
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17960 16176 18012 16182
rect 18340 16153 18368 16408
rect 17960 16118 18012 16124
rect 18326 16144 18382 16153
rect 17868 15972 17920 15978
rect 17868 15914 17920 15920
rect 17972 15910 18000 16118
rect 18524 16096 18552 16680
rect 18616 16454 18644 17156
rect 18696 17138 18748 17144
rect 18696 17060 18748 17066
rect 18696 17002 18748 17008
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18708 16114 18736 17002
rect 18326 16079 18382 16088
rect 18432 16068 18552 16096
rect 18604 16108 18656 16114
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17866 15736 17922 15745
rect 17866 15671 17922 15680
rect 17776 15088 17828 15094
rect 17776 15030 17828 15036
rect 17684 14612 17736 14618
rect 17684 14554 17736 14560
rect 17604 14346 17724 14362
rect 17604 14340 17736 14346
rect 17604 14334 17684 14340
rect 17684 14282 17736 14288
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17512 11762 17540 12038
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17328 11172 17540 11200
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 17328 10810 17356 11018
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17222 8800 17278 8809
rect 17222 8735 17278 8744
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17328 5778 17356 10610
rect 17512 10554 17540 11172
rect 17604 10713 17632 14214
rect 17684 12844 17736 12850
rect 17684 12786 17736 12792
rect 17696 12646 17724 12786
rect 17684 12640 17736 12646
rect 17684 12582 17736 12588
rect 17788 11558 17816 15030
rect 17880 14550 17908 15671
rect 18432 15502 18460 16068
rect 18604 16050 18656 16056
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18512 15972 18564 15978
rect 18512 15914 18564 15920
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18420 15360 18472 15366
rect 18420 15302 18472 15308
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 17868 14544 17920 14550
rect 17868 14486 17920 14492
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 18340 14006 18368 15098
rect 18432 14793 18460 15302
rect 18524 15201 18552 15914
rect 18510 15192 18566 15201
rect 18510 15127 18566 15136
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18418 14784 18474 14793
rect 18418 14719 18474 14728
rect 18420 14272 18472 14278
rect 18524 14260 18552 14962
rect 18472 14232 18552 14260
rect 18420 14214 18472 14220
rect 18524 14113 18552 14232
rect 18510 14104 18566 14113
rect 18510 14039 18566 14048
rect 18328 14000 18380 14006
rect 18328 13942 18380 13948
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 17868 13796 17920 13802
rect 17868 13738 17920 13744
rect 17880 13530 17908 13738
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17774 10976 17830 10985
rect 17590 10704 17646 10713
rect 17590 10639 17646 10648
rect 17512 10526 17632 10554
rect 17498 10432 17554 10441
rect 17498 10367 17554 10376
rect 17408 10260 17460 10266
rect 17408 10202 17460 10208
rect 17420 10169 17448 10202
rect 17406 10160 17462 10169
rect 17512 10130 17540 10367
rect 17406 10095 17462 10104
rect 17500 10124 17552 10130
rect 17420 8294 17448 10095
rect 17500 10066 17552 10072
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 7478 17448 8230
rect 17512 7478 17540 9658
rect 17604 8650 17632 10526
rect 17696 9353 17724 10950
rect 17774 10911 17830 10920
rect 17788 10810 17816 10911
rect 17776 10804 17828 10810
rect 17776 10746 17828 10752
rect 17774 10704 17830 10713
rect 17774 10639 17776 10648
rect 17828 10639 17830 10648
rect 17776 10610 17828 10616
rect 17880 10606 17908 13466
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18340 12170 18368 13466
rect 18420 12300 18472 12306
rect 18524 12288 18552 13874
rect 18616 12442 18644 16050
rect 18800 16046 18828 17546
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 18696 15632 18748 15638
rect 18696 15574 18748 15580
rect 18708 15473 18736 15574
rect 18694 15464 18750 15473
rect 18694 15399 18750 15408
rect 18696 15020 18748 15026
rect 18696 14962 18748 14968
rect 18708 14822 18736 14962
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18708 13394 18736 14486
rect 18800 14482 18828 15846
rect 18892 15162 18920 18634
rect 18972 18624 19024 18630
rect 18972 18566 19024 18572
rect 18984 16794 19012 18566
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 18970 16688 19026 16697
rect 18970 16623 18972 16632
rect 19024 16623 19026 16632
rect 18972 16594 19024 16600
rect 18970 16552 19026 16561
rect 18970 16487 19026 16496
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18878 15056 18934 15065
rect 18878 14991 18934 15000
rect 18892 14550 18920 14991
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 18788 14476 18840 14482
rect 18788 14418 18840 14424
rect 18984 14362 19012 16487
rect 19076 15994 19104 20742
rect 19260 19990 19288 20810
rect 19432 20800 19484 20806
rect 19430 20768 19432 20777
rect 19484 20768 19486 20777
rect 19430 20703 19486 20712
rect 19338 20360 19394 20369
rect 19338 20295 19340 20304
rect 19392 20295 19394 20304
rect 19340 20266 19392 20272
rect 19248 19984 19300 19990
rect 19248 19926 19300 19932
rect 19536 19854 19564 23530
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19628 22166 19656 22714
rect 19616 22160 19668 22166
rect 19616 22102 19668 22108
rect 19616 21888 19668 21894
rect 19616 21830 19668 21836
rect 19628 21690 19656 21830
rect 19616 21684 19668 21690
rect 19616 21626 19668 21632
rect 19800 21412 19852 21418
rect 19800 21354 19852 21360
rect 19812 21146 19840 21354
rect 19800 21140 19852 21146
rect 19800 21082 19852 21088
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19260 19417 19288 19450
rect 19246 19408 19302 19417
rect 19246 19343 19302 19352
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 19432 19236 19484 19242
rect 19432 19178 19484 19184
rect 19246 18320 19302 18329
rect 19156 18284 19208 18290
rect 19444 18290 19472 19178
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 19246 18255 19302 18264
rect 19432 18284 19484 18290
rect 19156 18226 19208 18232
rect 19168 18086 19196 18226
rect 19156 18080 19208 18086
rect 19260 18057 19288 18255
rect 19432 18226 19484 18232
rect 19536 18057 19564 18634
rect 19156 18022 19208 18028
rect 19246 18048 19302 18057
rect 19168 17610 19196 18022
rect 19246 17983 19302 17992
rect 19522 18048 19578 18057
rect 19522 17983 19578 17992
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19430 17776 19486 17785
rect 19248 17740 19300 17746
rect 19430 17711 19486 17720
rect 19248 17682 19300 17688
rect 19156 17604 19208 17610
rect 19156 17546 19208 17552
rect 19260 17202 19288 17682
rect 19444 17678 19472 17711
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19628 17270 19656 17818
rect 19616 17264 19668 17270
rect 19616 17206 19668 17212
rect 19248 17196 19300 17202
rect 19248 17138 19300 17144
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 19168 16726 19196 16934
rect 19156 16720 19208 16726
rect 19156 16662 19208 16668
rect 19156 16108 19208 16114
rect 19260 16096 19288 17138
rect 19720 16946 19748 19314
rect 19904 17728 19932 24822
rect 20074 24783 20130 24792
rect 19984 24132 20036 24138
rect 19984 24074 20036 24080
rect 19996 23798 20024 24074
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 19996 22982 20024 23734
rect 19984 22976 20036 22982
rect 19984 22918 20036 22924
rect 19996 22710 20024 22918
rect 19984 22704 20036 22710
rect 19984 22646 20036 22652
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 19996 21321 20024 21830
rect 19982 21312 20038 21321
rect 19982 21247 20038 21256
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 19996 21010 20024 21082
rect 20088 21010 20116 24783
rect 20272 23322 20300 26200
rect 21180 26036 21232 26042
rect 21180 25978 21232 25984
rect 20352 25628 20404 25634
rect 20352 25570 20404 25576
rect 20260 23316 20312 23322
rect 20260 23258 20312 23264
rect 20364 21894 20392 25570
rect 21192 24342 21220 25978
rect 21180 24336 21232 24342
rect 21100 24296 21180 24324
rect 21100 23361 21128 24296
rect 21180 24278 21232 24284
rect 21284 24274 21312 26302
rect 21546 26200 21602 27000
rect 22190 26200 22246 27000
rect 22834 26200 22890 27000
rect 23478 26330 23534 27000
rect 23478 26302 24072 26330
rect 23478 26200 23534 26302
rect 21364 24608 21416 24614
rect 21364 24550 21416 24556
rect 21272 24268 21324 24274
rect 21272 24210 21324 24216
rect 21272 24064 21324 24070
rect 21272 24006 21324 24012
rect 21180 23656 21232 23662
rect 21180 23598 21232 23604
rect 21086 23352 21142 23361
rect 21086 23287 21142 23296
rect 21192 23186 21220 23598
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 21086 23080 21142 23089
rect 20812 23044 20864 23050
rect 21086 23015 21088 23024
rect 20812 22986 20864 22992
rect 21140 23015 21142 23024
rect 21088 22986 21140 22992
rect 20824 22710 20852 22986
rect 20812 22704 20864 22710
rect 20812 22646 20864 22652
rect 20904 22568 20956 22574
rect 20904 22510 20956 22516
rect 20352 21888 20404 21894
rect 20352 21830 20404 21836
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 20166 21720 20222 21729
rect 20166 21655 20222 21664
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 20076 21004 20128 21010
rect 20076 20946 20128 20952
rect 20180 20346 20208 21655
rect 20352 21616 20404 21622
rect 20352 21558 20404 21564
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 20272 20641 20300 20742
rect 20258 20632 20314 20641
rect 20258 20567 20314 20576
rect 20088 20318 20208 20346
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 19996 19825 20024 19858
rect 19982 19816 20038 19825
rect 19982 19751 20038 19760
rect 19982 19544 20038 19553
rect 19982 19479 20038 19488
rect 19996 18834 20024 19479
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 20088 17762 20116 20318
rect 20166 20224 20222 20233
rect 20166 20159 20222 20168
rect 20180 19922 20208 20159
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 20180 19281 20208 19858
rect 20166 19272 20222 19281
rect 20166 19207 20222 19216
rect 20166 19136 20222 19145
rect 20166 19071 20222 19080
rect 20180 18970 20208 19071
rect 20168 18964 20220 18970
rect 20168 18906 20220 18912
rect 20272 18873 20300 20567
rect 20258 18864 20314 18873
rect 20258 18799 20314 18808
rect 20364 18766 20392 21558
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20444 19712 20496 19718
rect 20444 19654 20496 19660
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20258 18592 20314 18601
rect 20258 18527 20314 18536
rect 20088 17734 20208 17762
rect 19812 17700 19932 17728
rect 19812 17654 19840 17700
rect 19800 17648 19852 17654
rect 19800 17590 19852 17596
rect 19800 17536 19852 17542
rect 19800 17478 19852 17484
rect 19812 17377 19840 17478
rect 19798 17368 19854 17377
rect 19798 17303 19854 17312
rect 19536 16918 19748 16946
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19208 16068 19288 16096
rect 19156 16050 19208 16056
rect 19076 15966 19196 15994
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 18800 14334 19012 14362
rect 18800 13530 18828 14334
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 18788 13524 18840 13530
rect 18788 13466 18840 13472
rect 18892 13394 18920 14214
rect 19076 14074 19104 14758
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 18696 13388 18748 13394
rect 18880 13388 18932 13394
rect 18748 13348 18828 13376
rect 18696 13330 18748 13336
rect 18696 13252 18748 13258
rect 18696 13194 18748 13200
rect 18708 12918 18736 13194
rect 18696 12912 18748 12918
rect 18696 12854 18748 12860
rect 18604 12436 18656 12442
rect 18604 12378 18656 12384
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 18524 12260 18644 12288
rect 18420 12242 18472 12248
rect 18328 12164 18380 12170
rect 18328 12106 18380 12112
rect 18432 12050 18460 12242
rect 18512 12164 18564 12170
rect 18512 12106 18564 12112
rect 18340 12022 18460 12050
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 17960 11552 18012 11558
rect 17960 11494 18012 11500
rect 17972 11150 18000 11494
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 18248 11082 18276 11766
rect 18236 11076 18288 11082
rect 18236 11018 18288 11024
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 17788 9722 17816 9998
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17776 9376 17828 9382
rect 17682 9344 17738 9353
rect 17776 9318 17828 9324
rect 17682 9279 17738 9288
rect 17696 9178 17724 9279
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17604 8622 17724 8650
rect 17590 8528 17646 8537
rect 17590 8463 17646 8472
rect 17604 8430 17632 8463
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17408 7472 17460 7478
rect 17408 7414 17460 7420
rect 17500 7472 17552 7478
rect 17500 7414 17552 7420
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17604 6458 17632 7346
rect 17696 7274 17724 8622
rect 17788 8294 17816 9318
rect 17776 8288 17828 8294
rect 17776 8230 17828 8236
rect 17776 8016 17828 8022
rect 17776 7958 17828 7964
rect 17684 7268 17736 7274
rect 17684 7210 17736 7216
rect 17788 6848 17816 7958
rect 17880 7342 17908 10542
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 17972 9994 18000 10406
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 17960 9988 18012 9994
rect 17960 9930 18012 9936
rect 18064 9926 18092 10202
rect 18142 10024 18198 10033
rect 18142 9959 18198 9968
rect 18156 9926 18184 9959
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 18144 9716 18196 9722
rect 18196 9664 18276 9674
rect 18144 9658 18276 9664
rect 18156 9646 18276 9658
rect 18248 9382 18276 9646
rect 18340 9602 18368 12022
rect 18524 11354 18552 12106
rect 18616 11354 18644 12260
rect 18708 12102 18736 12310
rect 18800 12306 18828 13348
rect 18880 13330 18932 13336
rect 18880 13252 18932 13258
rect 18880 13194 18932 13200
rect 18892 12986 18920 13194
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18788 12300 18840 12306
rect 18788 12242 18840 12248
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 18420 11280 18472 11286
rect 18420 11222 18472 11228
rect 18602 11248 18658 11257
rect 18432 9722 18460 11222
rect 18512 11212 18564 11218
rect 18602 11183 18604 11192
rect 18512 11154 18564 11160
rect 18656 11183 18658 11192
rect 18604 11154 18656 11160
rect 18524 10985 18552 11154
rect 18708 11098 18736 12038
rect 18800 11529 18828 12038
rect 18786 11520 18842 11529
rect 18786 11455 18842 11464
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18616 11070 18736 11098
rect 18510 10976 18566 10985
rect 18510 10911 18566 10920
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18524 10538 18552 10746
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18616 10266 18644 11070
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18512 10124 18564 10130
rect 18708 10112 18736 10542
rect 18512 10066 18564 10072
rect 18616 10084 18736 10112
rect 18524 9722 18552 10066
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18512 9716 18564 9722
rect 18512 9658 18564 9664
rect 18340 9574 18552 9602
rect 18524 9518 18552 9574
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 18512 9512 18564 9518
rect 18512 9454 18564 9460
rect 18328 9444 18380 9450
rect 18328 9386 18380 9392
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18050 8528 18106 8537
rect 18050 8463 18052 8472
rect 18104 8463 18106 8472
rect 18052 8434 18104 8440
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17972 8090 18000 8366
rect 18156 8265 18184 8570
rect 18248 8362 18276 8570
rect 18340 8566 18368 9386
rect 18432 8673 18460 9454
rect 18524 8974 18552 9454
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18616 8906 18644 10084
rect 18800 9654 18828 11290
rect 18788 9648 18840 9654
rect 18788 9590 18840 9596
rect 18696 9104 18748 9110
rect 18694 9072 18696 9081
rect 18748 9072 18750 9081
rect 18694 9007 18750 9016
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18604 8900 18656 8906
rect 18604 8842 18656 8848
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18418 8664 18474 8673
rect 18418 8599 18474 8608
rect 18328 8560 18380 8566
rect 18328 8502 18380 8508
rect 18418 8392 18474 8401
rect 18236 8356 18288 8362
rect 18418 8327 18474 8336
rect 18236 8298 18288 8304
rect 18432 8294 18460 8327
rect 18420 8288 18472 8294
rect 18142 8256 18198 8265
rect 18420 8230 18472 8236
rect 18142 8191 18198 8200
rect 18432 8090 18460 8230
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17868 6860 17920 6866
rect 17788 6820 17868 6848
rect 17868 6802 17920 6808
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 17696 5302 17724 6734
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 17684 5296 17736 5302
rect 17130 5264 17186 5273
rect 17684 5238 17736 5244
rect 17130 5199 17186 5208
rect 17144 5166 17172 5199
rect 17132 5160 17184 5166
rect 17132 5102 17184 5108
rect 17788 4146 17816 6122
rect 17880 5710 17908 6802
rect 18340 6662 18368 7346
rect 18432 7002 18460 8026
rect 18524 7342 18552 8774
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18524 6798 18552 7142
rect 18512 6792 18564 6798
rect 18512 6734 18564 6740
rect 18328 6656 18380 6662
rect 18616 6610 18644 8842
rect 18708 7818 18736 8910
rect 18800 8634 18828 9590
rect 18892 8809 18920 12582
rect 19076 12170 19104 12718
rect 19064 12164 19116 12170
rect 19064 12106 19116 12112
rect 19064 11620 19116 11626
rect 19064 11562 19116 11568
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 18984 10985 19012 11086
rect 18970 10976 19026 10985
rect 18970 10911 19026 10920
rect 18972 10668 19024 10674
rect 18972 10610 19024 10616
rect 18878 8800 18934 8809
rect 18878 8735 18934 8744
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18878 8528 18934 8537
rect 18878 8463 18934 8472
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18892 6798 18920 8463
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18788 6724 18840 6730
rect 18788 6666 18840 6672
rect 18328 6598 18380 6604
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 18340 3641 18368 6598
rect 18524 6582 18644 6610
rect 18524 6322 18552 6582
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18420 5568 18472 5574
rect 18420 5510 18472 5516
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18432 5234 18460 5510
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 18524 3942 18552 5510
rect 18800 4622 18828 6666
rect 18880 6316 18932 6322
rect 18880 6258 18932 6264
rect 18892 5914 18920 6258
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18984 5778 19012 10610
rect 19076 6730 19104 11562
rect 19168 10577 19196 15966
rect 19248 14544 19300 14550
rect 19248 14486 19300 14492
rect 19260 13977 19288 14486
rect 19246 13968 19302 13977
rect 19246 13903 19302 13912
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 19260 12918 19288 13670
rect 19444 13190 19472 16390
rect 19536 15706 19564 16918
rect 19812 16810 19840 17303
rect 19628 16782 19840 16810
rect 19628 15910 19656 16782
rect 19708 16652 19760 16658
rect 19708 16594 19760 16600
rect 19720 16538 19748 16594
rect 19720 16510 19932 16538
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19628 15162 19656 15302
rect 19616 15156 19668 15162
rect 19616 15098 19668 15104
rect 19524 15088 19576 15094
rect 19524 15030 19576 15036
rect 19536 14958 19564 15030
rect 19524 14952 19576 14958
rect 19522 14920 19524 14929
rect 19576 14920 19578 14929
rect 19522 14855 19578 14864
rect 19628 14657 19656 15098
rect 19720 14890 19748 16510
rect 19904 16454 19932 16510
rect 19800 16448 19852 16454
rect 19800 16390 19852 16396
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 19812 15162 19840 16390
rect 19890 16144 19946 16153
rect 19890 16079 19946 16088
rect 19904 15881 19932 16079
rect 19890 15872 19946 15881
rect 19890 15807 19946 15816
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19800 15156 19852 15162
rect 19800 15098 19852 15104
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19708 14884 19760 14890
rect 19708 14826 19760 14832
rect 19614 14648 19670 14657
rect 19614 14583 19670 14592
rect 19708 14612 19760 14618
rect 19708 14554 19760 14560
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19536 13870 19564 14214
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19536 13530 19564 13806
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19616 13320 19668 13326
rect 19616 13262 19668 13268
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19248 12912 19300 12918
rect 19248 12854 19300 12860
rect 19444 12850 19472 12922
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19338 12744 19394 12753
rect 19338 12679 19340 12688
rect 19392 12679 19394 12688
rect 19340 12650 19392 12656
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19260 11694 19288 12038
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19246 11112 19302 11121
rect 19246 11047 19302 11056
rect 19260 11014 19288 11047
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19352 10810 19380 11494
rect 19444 11354 19472 12786
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 10985 19472 11086
rect 19430 10976 19486 10985
rect 19430 10911 19486 10920
rect 19430 10840 19486 10849
rect 19340 10804 19392 10810
rect 19430 10775 19432 10784
rect 19340 10746 19392 10752
rect 19484 10775 19486 10784
rect 19432 10746 19484 10752
rect 19154 10568 19210 10577
rect 19154 10503 19210 10512
rect 19156 10464 19208 10470
rect 19156 10406 19208 10412
rect 19168 10033 19196 10406
rect 19154 10024 19210 10033
rect 19154 9959 19210 9968
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19156 9920 19208 9926
rect 19156 9862 19208 9868
rect 19168 6866 19196 9862
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19260 9042 19288 9454
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 19260 8430 19288 8978
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 19260 8090 19288 8366
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 19156 6860 19208 6866
rect 19156 6802 19208 6808
rect 19064 6724 19116 6730
rect 19064 6666 19116 6672
rect 19352 6458 19380 9930
rect 19430 9208 19486 9217
rect 19430 9143 19432 9152
rect 19484 9143 19486 9152
rect 19432 9114 19484 9120
rect 19536 7750 19564 12786
rect 19628 11558 19656 13262
rect 19616 11552 19668 11558
rect 19616 11494 19668 11500
rect 19720 11150 19748 14554
rect 19812 13258 19840 14962
rect 19904 14958 19932 15642
rect 20180 15026 20208 17734
rect 20272 15366 20300 18527
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20364 16658 20392 16934
rect 20352 16652 20404 16658
rect 20352 16594 20404 16600
rect 20456 15706 20484 19654
rect 20548 16266 20576 21422
rect 20824 20942 20852 21830
rect 20812 20936 20864 20942
rect 20626 20904 20682 20913
rect 20812 20878 20864 20884
rect 20626 20839 20682 20848
rect 20640 20806 20668 20839
rect 20628 20800 20680 20806
rect 20628 20742 20680 20748
rect 20812 20800 20864 20806
rect 20812 20742 20864 20748
rect 20640 18601 20668 20742
rect 20824 20602 20852 20742
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20732 19922 20760 20538
rect 20720 19916 20772 19922
rect 20720 19858 20772 19864
rect 20626 18592 20682 18601
rect 20626 18527 20682 18536
rect 20732 17592 20760 19858
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 20824 19174 20852 19654
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20916 18714 20944 22510
rect 21088 22160 21140 22166
rect 21088 22102 21140 22108
rect 21100 22012 21128 22102
rect 21192 22094 21220 23122
rect 21284 22574 21312 24006
rect 21376 23866 21404 24550
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 21364 23520 21416 23526
rect 21560 23497 21588 26200
rect 21732 25764 21784 25770
rect 21732 25706 21784 25712
rect 21638 24848 21694 24857
rect 21638 24783 21694 24792
rect 21364 23462 21416 23468
rect 21546 23488 21602 23497
rect 21376 22574 21404 23462
rect 21546 23423 21602 23432
rect 21272 22568 21324 22574
rect 21272 22510 21324 22516
rect 21364 22568 21416 22574
rect 21364 22510 21416 22516
rect 21284 22234 21312 22510
rect 21364 22432 21416 22438
rect 21364 22374 21416 22380
rect 21272 22228 21324 22234
rect 21272 22170 21324 22176
rect 21192 22066 21312 22094
rect 21008 21984 21128 22012
rect 21008 20233 21036 21984
rect 21088 21548 21140 21554
rect 21088 21490 21140 21496
rect 21100 21078 21128 21490
rect 21284 21486 21312 22066
rect 21272 21480 21324 21486
rect 21272 21422 21324 21428
rect 21088 21072 21140 21078
rect 21088 21014 21140 21020
rect 21088 20936 21140 20942
rect 21284 20924 21312 21422
rect 21140 20896 21312 20924
rect 21088 20878 21140 20884
rect 21100 20330 21128 20878
rect 21088 20324 21140 20330
rect 21088 20266 21140 20272
rect 20994 20224 21050 20233
rect 20994 20159 21050 20168
rect 21100 20058 21128 20266
rect 21272 20256 21324 20262
rect 21270 20224 21272 20233
rect 21324 20224 21326 20233
rect 21270 20159 21326 20168
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 21180 20052 21232 20058
rect 21180 19994 21232 20000
rect 20996 19780 21048 19786
rect 20996 19722 21048 19728
rect 21008 18970 21036 19722
rect 21100 19378 21128 19994
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 21192 18766 21220 19994
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21180 18760 21232 18766
rect 20916 18686 21128 18714
rect 21180 18702 21232 18708
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20916 17882 20944 18022
rect 20904 17876 20956 17882
rect 20904 17818 20956 17824
rect 20812 17604 20864 17610
rect 20732 17564 20812 17592
rect 20812 17546 20864 17552
rect 20720 17060 20772 17066
rect 20720 17002 20772 17008
rect 20732 16658 20760 17002
rect 20824 16658 20852 17546
rect 21008 17202 21036 18226
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 20904 17060 20956 17066
rect 20904 17002 20956 17008
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20812 16652 20864 16658
rect 20812 16594 20864 16600
rect 20732 16538 20760 16594
rect 20732 16510 20852 16538
rect 20548 16238 20668 16266
rect 20640 15978 20668 16238
rect 20720 16176 20772 16182
rect 20720 16118 20772 16124
rect 20824 16130 20852 16510
rect 20916 16250 20944 17002
rect 21008 16794 21036 17138
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 20628 15972 20680 15978
rect 20628 15914 20680 15920
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20732 15570 20760 16118
rect 20824 16102 20944 16130
rect 21008 16114 21036 16730
rect 21100 16114 21128 18686
rect 21284 17785 21312 19450
rect 21376 19446 21404 22374
rect 21454 22264 21510 22273
rect 21454 22199 21510 22208
rect 21468 21010 21496 22199
rect 21652 22094 21680 24783
rect 21560 22066 21680 22094
rect 21456 21004 21508 21010
rect 21456 20946 21508 20952
rect 21454 20088 21510 20097
rect 21454 20023 21510 20032
rect 21364 19440 21416 19446
rect 21364 19382 21416 19388
rect 21376 18766 21404 19382
rect 21468 19378 21496 20023
rect 21456 19372 21508 19378
rect 21456 19314 21508 19320
rect 21456 19168 21508 19174
rect 21456 19110 21508 19116
rect 21364 18760 21416 18766
rect 21364 18702 21416 18708
rect 21468 18086 21496 19110
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21270 17776 21326 17785
rect 21270 17711 21326 17720
rect 21272 17604 21324 17610
rect 21272 17546 21324 17552
rect 21284 17134 21312 17546
rect 21364 17536 21416 17542
rect 21364 17478 21416 17484
rect 21376 17377 21404 17478
rect 21362 17368 21418 17377
rect 21362 17303 21418 17312
rect 21272 17128 21324 17134
rect 21272 17070 21324 17076
rect 21362 16280 21418 16289
rect 21180 16244 21232 16250
rect 21362 16215 21418 16224
rect 21180 16186 21232 16192
rect 20916 16046 20944 16102
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 20904 16040 20956 16046
rect 20904 15982 20956 15988
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20824 15094 20852 15506
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19800 13252 19852 13258
rect 19800 13194 19852 13200
rect 19904 12434 19932 14894
rect 20536 14408 20588 14414
rect 20536 14350 20588 14356
rect 19984 14272 20036 14278
rect 20548 14249 20576 14350
rect 19984 14214 20036 14220
rect 20534 14240 20590 14249
rect 19996 13530 20024 14214
rect 20534 14175 20590 14184
rect 20074 13968 20130 13977
rect 20074 13903 20130 13912
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 20088 13394 20116 13903
rect 20350 13696 20406 13705
rect 20350 13631 20406 13640
rect 20168 13456 20220 13462
rect 20220 13404 20300 13410
rect 20168 13398 20300 13404
rect 20076 13388 20128 13394
rect 20180 13382 20300 13398
rect 20076 13330 20128 13336
rect 20088 12434 20116 13330
rect 20272 13190 20300 13382
rect 20168 13184 20220 13190
rect 20168 13126 20220 13132
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20180 12442 20208 13126
rect 19812 12406 19932 12434
rect 19996 12406 20116 12434
rect 20168 12436 20220 12442
rect 19708 11144 19760 11150
rect 19708 11086 19760 11092
rect 19616 10736 19668 10742
rect 19616 10678 19668 10684
rect 19628 7886 19656 10678
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19720 10130 19748 10542
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 19708 9648 19760 9654
rect 19708 9590 19760 9596
rect 19720 9382 19748 9590
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19720 8344 19748 8910
rect 19812 8650 19840 12406
rect 19996 12170 20024 12406
rect 20168 12378 20220 12384
rect 20272 12306 20300 13126
rect 20364 12986 20392 13631
rect 20352 12980 20404 12986
rect 20352 12922 20404 12928
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 20456 12442 20484 12650
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 20260 12300 20312 12306
rect 20260 12242 20312 12248
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 20166 12200 20222 12209
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19904 11354 19932 11494
rect 20088 11354 20116 12174
rect 20166 12135 20222 12144
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 20180 11121 20208 12135
rect 20272 12102 20300 12242
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 20442 11928 20498 11937
rect 20442 11863 20498 11872
rect 20456 11626 20484 11863
rect 20444 11620 20496 11626
rect 20444 11562 20496 11568
rect 20166 11112 20222 11121
rect 20166 11047 20222 11056
rect 20350 10976 20406 10985
rect 20350 10911 20406 10920
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19812 8634 19932 8650
rect 19812 8628 19944 8634
rect 19812 8622 19892 8628
rect 19892 8570 19944 8576
rect 19720 8316 19840 8344
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 19524 7744 19576 7750
rect 19524 7686 19576 7692
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 19720 6458 19748 7346
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19708 6452 19760 6458
rect 19708 6394 19760 6400
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19708 6112 19760 6118
rect 19708 6054 19760 6060
rect 18972 5772 19024 5778
rect 18972 5714 19024 5720
rect 19248 5092 19300 5098
rect 19248 5034 19300 5040
rect 19156 4684 19208 4690
rect 19156 4626 19208 4632
rect 18788 4616 18840 4622
rect 18788 4558 18840 4564
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 19168 3670 19196 4626
rect 19156 3664 19208 3670
rect 18326 3632 18382 3641
rect 19156 3606 19208 3612
rect 18326 3567 18382 3576
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 19260 3482 19288 5034
rect 19524 3528 19576 3534
rect 19260 3476 19524 3482
rect 19260 3470 19576 3476
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 16488 2984 16540 2990
rect 16488 2926 16540 2932
rect 16396 2440 16448 2446
rect 16396 2382 16448 2388
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 15948 870 16068 898
rect 15948 800 15976 870
rect 1122 0 1178 800
rect 3238 0 3294 800
rect 5354 0 5410 800
rect 7470 0 7526 800
rect 9586 0 9642 800
rect 11702 0 11758 800
rect 13818 0 13874 800
rect 15934 0 15990 800
rect 16040 762 16068 870
rect 16500 762 16528 2926
rect 17604 2854 17632 3470
rect 18880 3460 18932 3466
rect 19260 3454 19564 3470
rect 18880 3402 18932 3408
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 18892 3058 18920 3402
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19536 3126 19564 3334
rect 19524 3120 19576 3126
rect 19524 3062 19576 3068
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 19628 2990 19656 6054
rect 19720 4554 19748 6054
rect 19708 4548 19760 4554
rect 19708 4490 19760 4496
rect 19812 3194 19840 8316
rect 19996 7546 20024 10542
rect 20364 10130 20392 10911
rect 20548 10690 20576 12718
rect 20640 11354 20668 14962
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20732 12170 20760 14894
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20824 14074 20852 14350
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20824 13394 20852 14010
rect 20916 13954 20944 15982
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 21008 15706 21036 15846
rect 20996 15700 21048 15706
rect 20996 15642 21048 15648
rect 21086 14376 21142 14385
rect 21086 14311 21088 14320
rect 21140 14311 21142 14320
rect 21088 14282 21140 14288
rect 21192 14226 21220 16186
rect 21376 15910 21404 16215
rect 21364 15904 21416 15910
rect 21364 15846 21416 15852
rect 21468 15570 21496 18022
rect 21560 15745 21588 22066
rect 21640 21888 21692 21894
rect 21640 21830 21692 21836
rect 21652 21690 21680 21830
rect 21640 21684 21692 21690
rect 21640 21626 21692 21632
rect 21640 21412 21692 21418
rect 21640 21354 21692 21360
rect 21652 20890 21680 21354
rect 21744 21298 21772 25706
rect 22098 24304 22154 24313
rect 22098 24239 22154 24248
rect 22112 24206 22140 24239
rect 22100 24200 22152 24206
rect 22100 24142 22152 24148
rect 22204 22658 22232 26200
rect 22558 25256 22614 25265
rect 22558 25191 22614 25200
rect 22282 24712 22338 24721
rect 22282 24647 22338 24656
rect 22112 22630 22232 22658
rect 22112 22624 22140 22630
rect 21928 22596 22140 22624
rect 21824 21956 21876 21962
rect 21824 21898 21876 21904
rect 21836 21434 21864 21898
rect 21928 21554 21956 22596
rect 22192 22568 22244 22574
rect 22192 22510 22244 22516
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22008 21888 22060 21894
rect 22112 21865 22140 21966
rect 22008 21830 22060 21836
rect 22098 21856 22154 21865
rect 22020 21622 22048 21830
rect 22098 21791 22154 21800
rect 22008 21616 22060 21622
rect 22008 21558 22060 21564
rect 21916 21548 21968 21554
rect 21916 21490 21968 21496
rect 22204 21468 22232 22510
rect 22296 21622 22324 24647
rect 22468 23656 22520 23662
rect 22468 23598 22520 23604
rect 22480 23322 22508 23598
rect 22468 23316 22520 23322
rect 22468 23258 22520 23264
rect 22572 23202 22600 25191
rect 22652 23588 22704 23594
rect 22652 23530 22704 23536
rect 22664 23322 22692 23530
rect 22652 23316 22704 23322
rect 22652 23258 22704 23264
rect 22376 23180 22428 23186
rect 22572 23174 22692 23202
rect 22376 23122 22428 23128
rect 22388 22438 22416 23122
rect 22376 22432 22428 22438
rect 22376 22374 22428 22380
rect 22388 21622 22416 22374
rect 22560 22092 22612 22098
rect 22560 22034 22612 22040
rect 22468 21956 22520 21962
rect 22468 21898 22520 21904
rect 22480 21865 22508 21898
rect 22466 21856 22522 21865
rect 22466 21791 22522 21800
rect 22284 21616 22336 21622
rect 22284 21558 22336 21564
rect 22376 21616 22428 21622
rect 22376 21558 22428 21564
rect 22284 21480 22336 21486
rect 22204 21440 22284 21468
rect 21836 21406 22048 21434
rect 22284 21422 22336 21428
rect 21744 21270 21864 21298
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 21744 21010 21772 21082
rect 21732 21004 21784 21010
rect 21732 20946 21784 20952
rect 21652 20862 21772 20890
rect 21640 19916 21692 19922
rect 21640 19858 21692 19864
rect 21652 16833 21680 19858
rect 21744 19446 21772 20862
rect 21732 19440 21784 19446
rect 21732 19382 21784 19388
rect 21730 19272 21786 19281
rect 21730 19207 21732 19216
rect 21784 19207 21786 19216
rect 21732 19178 21784 19184
rect 21732 18896 21784 18902
rect 21732 18838 21784 18844
rect 21638 16824 21694 16833
rect 21744 16794 21772 18838
rect 21638 16759 21694 16768
rect 21732 16788 21784 16794
rect 21732 16730 21784 16736
rect 21640 16108 21692 16114
rect 21640 16050 21692 16056
rect 21652 15910 21680 16050
rect 21640 15904 21692 15910
rect 21692 15852 21772 15858
rect 21640 15846 21772 15852
rect 21652 15830 21772 15846
rect 21546 15736 21602 15745
rect 21546 15671 21602 15680
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 21100 14198 21220 14226
rect 20916 13926 21036 13954
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20904 13252 20956 13258
rect 20904 13194 20956 13200
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20720 12164 20772 12170
rect 20720 12106 20772 12112
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20732 11014 20760 11698
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20732 10742 20760 10950
rect 20720 10736 20772 10742
rect 20548 10662 20668 10690
rect 20720 10678 20772 10684
rect 20640 10606 20668 10662
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20076 9920 20128 9926
rect 20076 9862 20128 9868
rect 20088 9518 20116 9862
rect 20166 9616 20222 9625
rect 20166 9551 20222 9560
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 20180 8537 20208 9551
rect 20166 8528 20222 8537
rect 20166 8463 20222 8472
rect 20260 7744 20312 7750
rect 20260 7686 20312 7692
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 20272 6798 20300 7686
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 20180 4826 20208 5646
rect 20364 5234 20392 10066
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 20456 8430 20484 9658
rect 20536 8900 20588 8906
rect 20536 8842 20588 8848
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20352 5228 20404 5234
rect 20352 5170 20404 5176
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20456 4622 20484 8366
rect 20548 5778 20576 8842
rect 20536 5772 20588 5778
rect 20536 5714 20588 5720
rect 20640 5710 20668 10542
rect 20732 9994 20760 10678
rect 20720 9988 20772 9994
rect 20720 9930 20772 9936
rect 20732 9586 20760 9930
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20732 8906 20760 9522
rect 20824 9178 20852 12582
rect 20812 9172 20864 9178
rect 20812 9114 20864 9120
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20732 8566 20760 8842
rect 20916 8634 20944 13194
rect 21008 12594 21036 13926
rect 21100 12714 21128 14198
rect 21180 13252 21232 13258
rect 21180 13194 21232 13200
rect 21088 12708 21140 12714
rect 21088 12650 21140 12656
rect 21008 12566 21128 12594
rect 20996 12164 21048 12170
rect 20996 12106 21048 12112
rect 21008 11626 21036 12106
rect 21100 11898 21128 12566
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 21100 11762 21128 11834
rect 21088 11756 21140 11762
rect 21088 11698 21140 11704
rect 20996 11620 21048 11626
rect 20996 11562 21048 11568
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 20718 8392 20774 8401
rect 20718 8327 20774 8336
rect 20812 8356 20864 8362
rect 20732 7313 20760 8327
rect 20812 8298 20864 8304
rect 20718 7304 20774 7313
rect 20718 7239 20774 7248
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20824 5234 20852 8298
rect 20902 7712 20958 7721
rect 20902 7647 20958 7656
rect 20916 6254 20944 7647
rect 20996 6316 21048 6322
rect 20996 6258 21048 6264
rect 20904 6248 20956 6254
rect 20904 6190 20956 6196
rect 21008 5914 21036 6258
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 21100 4826 21128 11698
rect 21192 8022 21220 13194
rect 21284 13190 21312 15370
rect 21468 15162 21496 15506
rect 21640 15428 21692 15434
rect 21640 15370 21692 15376
rect 21456 15156 21508 15162
rect 21456 15098 21508 15104
rect 21548 15020 21600 15026
rect 21548 14962 21600 14968
rect 21456 14476 21508 14482
rect 21456 14418 21508 14424
rect 21468 14074 21496 14418
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21364 13728 21416 13734
rect 21560 13705 21588 14962
rect 21364 13670 21416 13676
rect 21546 13696 21602 13705
rect 21376 13274 21404 13670
rect 21546 13631 21602 13640
rect 21652 13530 21680 15370
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21652 13394 21680 13466
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21640 13388 21692 13394
rect 21640 13330 21692 13336
rect 21376 13246 21496 13274
rect 21272 13184 21324 13190
rect 21272 13126 21324 13132
rect 21364 13184 21416 13190
rect 21364 13126 21416 13132
rect 21376 12782 21404 13126
rect 21364 12776 21416 12782
rect 21364 12718 21416 12724
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21284 9994 21312 11630
rect 21376 11218 21404 11630
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 21376 10849 21404 11154
rect 21362 10840 21418 10849
rect 21362 10775 21418 10784
rect 21364 10464 21416 10470
rect 21364 10406 21416 10412
rect 21272 9988 21324 9994
rect 21272 9930 21324 9936
rect 21376 9722 21404 10406
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21468 8090 21496 13246
rect 21560 13025 21588 13330
rect 21546 13016 21602 13025
rect 21546 12951 21602 12960
rect 21560 12434 21588 12951
rect 21560 12406 21680 12434
rect 21652 12170 21680 12406
rect 21640 12164 21692 12170
rect 21640 12106 21692 12112
rect 21652 11694 21680 12106
rect 21640 11688 21692 11694
rect 21744 11665 21772 15830
rect 21836 15638 21864 21270
rect 22020 21146 22048 21406
rect 22100 21344 22152 21350
rect 22388 21332 22416 21558
rect 22100 21286 22152 21292
rect 22204 21304 22416 21332
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 22112 20602 22140 21286
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 22008 19372 22060 19378
rect 22204 19334 22232 21304
rect 22466 20632 22522 20641
rect 22466 20567 22522 20576
rect 22480 20398 22508 20567
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 22284 19440 22336 19446
rect 22284 19382 22336 19388
rect 22008 19314 22060 19320
rect 21916 19304 21968 19310
rect 21916 19246 21968 19252
rect 21928 17542 21956 19246
rect 22020 19174 22048 19314
rect 22112 19306 22232 19334
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 22008 18284 22060 18290
rect 22112 18272 22140 19306
rect 22296 19292 22324 19382
rect 22480 19310 22508 20198
rect 22572 20097 22600 22034
rect 22664 21486 22692 23174
rect 22744 23044 22796 23050
rect 22744 22986 22796 22992
rect 22756 22137 22784 22986
rect 22848 22817 22876 26200
rect 23388 24744 23440 24750
rect 23388 24686 23440 24692
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23202 24032 23258 24041
rect 23202 23967 23258 23976
rect 23216 23730 23244 23967
rect 23204 23724 23256 23730
rect 23204 23666 23256 23672
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22928 23112 22980 23118
rect 22928 23054 22980 23060
rect 22834 22808 22890 22817
rect 22834 22743 22890 22752
rect 22940 22760 22968 23054
rect 23020 22772 23072 22778
rect 22940 22732 23020 22760
rect 22940 22692 22968 22732
rect 23020 22714 23072 22720
rect 22848 22664 22968 22692
rect 22848 22216 22876 22664
rect 23296 22636 23348 22642
rect 23296 22578 23348 22584
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23308 22234 23336 22578
rect 23400 22574 23428 24686
rect 23664 24608 23716 24614
rect 23664 24550 23716 24556
rect 23572 23520 23624 23526
rect 23572 23462 23624 23468
rect 23584 22953 23612 23462
rect 23570 22944 23626 22953
rect 23570 22879 23626 22888
rect 23676 22794 23704 24550
rect 23848 24064 23900 24070
rect 23848 24006 23900 24012
rect 23860 23866 23888 24006
rect 23848 23860 23900 23866
rect 23848 23802 23900 23808
rect 23846 23352 23902 23361
rect 23846 23287 23902 23296
rect 23584 22766 23704 22794
rect 23388 22568 23440 22574
rect 23388 22510 23440 22516
rect 23480 22500 23532 22506
rect 23480 22442 23532 22448
rect 23492 22409 23520 22442
rect 23478 22400 23534 22409
rect 23478 22335 23534 22344
rect 23296 22228 23348 22234
rect 22848 22188 22968 22216
rect 22742 22128 22798 22137
rect 22798 22072 22876 22094
rect 22742 22066 22876 22072
rect 22742 22063 22798 22066
rect 22652 21480 22704 21486
rect 22652 21422 22704 21428
rect 22744 21344 22796 21350
rect 22744 21286 22796 21292
rect 22652 20936 22704 20942
rect 22650 20904 22652 20913
rect 22704 20904 22706 20913
rect 22756 20874 22784 21286
rect 22650 20839 22706 20848
rect 22744 20868 22796 20874
rect 22744 20810 22796 20816
rect 22848 20641 22876 22066
rect 22940 21350 22968 22188
rect 23296 22170 23348 22176
rect 23388 22092 23440 22098
rect 23388 22034 23440 22040
rect 23400 21418 23428 22034
rect 23388 21412 23440 21418
rect 23388 21354 23440 21360
rect 22928 21344 22980 21350
rect 22928 21286 22980 21292
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23296 20868 23348 20874
rect 23296 20810 23348 20816
rect 22928 20800 22980 20806
rect 22928 20742 22980 20748
rect 22650 20632 22706 20641
rect 22834 20632 22890 20641
rect 22706 20590 22784 20618
rect 22650 20567 22706 20576
rect 22652 20460 22704 20466
rect 22652 20402 22704 20408
rect 22558 20088 22614 20097
rect 22558 20023 22614 20032
rect 22572 19990 22600 20023
rect 22560 19984 22612 19990
rect 22560 19926 22612 19932
rect 22560 19848 22612 19854
rect 22560 19790 22612 19796
rect 22468 19304 22520 19310
rect 22296 19264 22416 19292
rect 22284 19168 22336 19174
rect 22284 19110 22336 19116
rect 22190 19000 22246 19009
rect 22296 18970 22324 19110
rect 22190 18935 22246 18944
rect 22284 18964 22336 18970
rect 22204 18426 22232 18935
rect 22284 18906 22336 18912
rect 22296 18630 22324 18906
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 22192 18420 22244 18426
rect 22192 18362 22244 18368
rect 22296 18290 22324 18566
rect 22060 18244 22140 18272
rect 22284 18284 22336 18290
rect 22008 18226 22060 18232
rect 22284 18226 22336 18232
rect 22388 18170 22416 19264
rect 22468 19246 22520 19252
rect 22112 18142 22416 18170
rect 22008 17740 22060 17746
rect 22008 17682 22060 17688
rect 21916 17536 21968 17542
rect 21916 17478 21968 17484
rect 22020 17066 22048 17682
rect 22008 17060 22060 17066
rect 22008 17002 22060 17008
rect 21916 16788 21968 16794
rect 21916 16730 21968 16736
rect 21824 15632 21876 15638
rect 21824 15574 21876 15580
rect 21836 15162 21864 15574
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21928 14521 21956 16730
rect 22008 15156 22060 15162
rect 22008 15098 22060 15104
rect 22020 15026 22048 15098
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 22112 14521 22140 18142
rect 22376 17128 22428 17134
rect 22376 17070 22428 17076
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 22204 15502 22232 16934
rect 22388 16590 22416 17070
rect 22572 16697 22600 19790
rect 22664 17814 22692 20402
rect 22756 19854 22784 20590
rect 22940 20602 22968 20742
rect 22834 20567 22890 20576
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 22836 20528 22888 20534
rect 22836 20470 22888 20476
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 22848 19786 22876 20470
rect 22928 20392 22980 20398
rect 22926 20360 22928 20369
rect 22980 20360 22982 20369
rect 22926 20295 22982 20304
rect 23308 20262 23336 20810
rect 23388 20800 23440 20806
rect 23388 20742 23440 20748
rect 23296 20256 23348 20262
rect 23296 20198 23348 20204
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23296 20052 23348 20058
rect 23296 19994 23348 20000
rect 22836 19780 22888 19786
rect 23308 19768 23336 19994
rect 22888 19740 23336 19768
rect 22836 19722 22888 19728
rect 23400 19334 23428 20742
rect 23584 20534 23612 22766
rect 23664 22432 23716 22438
rect 23664 22374 23716 22380
rect 23676 22273 23704 22374
rect 23662 22264 23718 22273
rect 23860 22234 23888 23287
rect 23940 23180 23992 23186
rect 23940 23122 23992 23128
rect 23952 22273 23980 23122
rect 23938 22264 23994 22273
rect 23662 22199 23718 22208
rect 23848 22228 23900 22234
rect 23938 22199 23994 22208
rect 23848 22170 23900 22176
rect 23860 22098 23888 22170
rect 23940 22160 23992 22166
rect 23940 22102 23992 22108
rect 23756 22092 23808 22098
rect 23756 22034 23808 22040
rect 23848 22092 23900 22098
rect 23848 22034 23900 22040
rect 23768 22001 23796 22034
rect 23754 21992 23810 22001
rect 23754 21927 23810 21936
rect 23768 21554 23796 21927
rect 23756 21548 23808 21554
rect 23756 21490 23808 21496
rect 23664 21412 23716 21418
rect 23664 21354 23716 21360
rect 23676 21128 23704 21354
rect 23676 21100 23796 21128
rect 23572 20528 23624 20534
rect 23572 20470 23624 20476
rect 23480 20256 23532 20262
rect 23480 20198 23532 20204
rect 23492 19553 23520 20198
rect 23768 19922 23796 21100
rect 23848 21004 23900 21010
rect 23848 20946 23900 20952
rect 23860 20874 23888 20946
rect 23848 20868 23900 20874
rect 23848 20810 23900 20816
rect 23846 20768 23902 20777
rect 23846 20703 23902 20712
rect 23756 19916 23808 19922
rect 23756 19858 23808 19864
rect 23572 19848 23624 19854
rect 23572 19790 23624 19796
rect 23478 19544 23534 19553
rect 23478 19479 23534 19488
rect 23478 19408 23534 19417
rect 23478 19343 23480 19352
rect 23308 19306 23428 19334
rect 23532 19343 23534 19352
rect 23480 19314 23532 19320
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22756 18630 22784 18702
rect 22836 18692 22888 18698
rect 22836 18634 22888 18640
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22652 17808 22704 17814
rect 22652 17750 22704 17756
rect 22558 16688 22614 16697
rect 22558 16623 22614 16632
rect 22376 16584 22428 16590
rect 22376 16526 22428 16532
rect 22466 16280 22522 16289
rect 22466 16215 22522 16224
rect 22480 16046 22508 16215
rect 22468 16040 22520 16046
rect 22468 15982 22520 15988
rect 22374 15736 22430 15745
rect 22374 15671 22430 15680
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 22192 14884 22244 14890
rect 22192 14826 22244 14832
rect 21914 14512 21970 14521
rect 21824 14476 21876 14482
rect 21914 14447 21970 14456
rect 22098 14512 22154 14521
rect 22098 14447 22154 14456
rect 21824 14418 21876 14424
rect 21836 14249 21864 14418
rect 22204 14414 22232 14826
rect 22192 14408 22244 14414
rect 22112 14368 22192 14396
rect 21822 14240 21878 14249
rect 21822 14175 21878 14184
rect 21836 11762 21864 14175
rect 22008 14068 22060 14074
rect 22008 14010 22060 14016
rect 22020 13841 22048 14010
rect 22112 13938 22140 14368
rect 22192 14350 22244 14356
rect 22192 14000 22244 14006
rect 22192 13942 22244 13948
rect 22100 13932 22152 13938
rect 22100 13874 22152 13880
rect 22006 13832 22062 13841
rect 22006 13767 22062 13776
rect 22100 13796 22152 13802
rect 22100 13738 22152 13744
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 21824 11756 21876 11762
rect 21824 11698 21876 11704
rect 21640 11630 21692 11636
rect 21730 11656 21786 11665
rect 21652 11150 21680 11630
rect 21730 11591 21786 11600
rect 21640 11144 21692 11150
rect 21640 11086 21692 11092
rect 21546 10840 21602 10849
rect 21652 10810 21680 11086
rect 21824 11076 21876 11082
rect 21824 11018 21876 11024
rect 21916 11076 21968 11082
rect 21916 11018 21968 11024
rect 21546 10775 21602 10784
rect 21640 10804 21692 10810
rect 21560 9654 21588 10775
rect 21640 10746 21692 10752
rect 21836 10742 21864 11018
rect 21824 10736 21876 10742
rect 21824 10678 21876 10684
rect 21548 9648 21600 9654
rect 21548 9590 21600 9596
rect 21824 9444 21876 9450
rect 21824 9386 21876 9392
rect 21836 9042 21864 9386
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21836 8430 21864 8978
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 21730 8120 21786 8129
rect 21456 8084 21508 8090
rect 21730 8055 21786 8064
rect 21456 8026 21508 8032
rect 21180 8016 21232 8022
rect 21180 7958 21232 7964
rect 21744 7886 21772 8055
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21836 7206 21864 8366
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21824 7200 21876 7206
rect 21824 7142 21876 7148
rect 21468 6730 21496 7142
rect 21456 6724 21508 6730
rect 21456 6666 21508 6672
rect 21640 5704 21692 5710
rect 21640 5646 21692 5652
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 21088 4820 21140 4826
rect 21088 4762 21140 4768
rect 20732 4690 20760 4762
rect 20904 4752 20956 4758
rect 20904 4694 20956 4700
rect 20720 4684 20772 4690
rect 20720 4626 20772 4632
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 20088 3738 20116 4082
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 19800 3188 19852 3194
rect 19800 3130 19852 3136
rect 19616 2984 19668 2990
rect 19616 2926 19668 2932
rect 17592 2848 17644 2854
rect 17592 2790 17644 2796
rect 18328 2372 18380 2378
rect 18328 2314 18380 2320
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 16040 734 16528 762
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18340 762 18368 2314
rect 20180 800 20208 4014
rect 20720 4004 20772 4010
rect 20720 3946 20772 3952
rect 20732 3670 20760 3946
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 20916 2514 20944 4694
rect 21272 4548 21324 4554
rect 21272 4490 21324 4496
rect 21284 4282 21312 4490
rect 21272 4276 21324 4282
rect 21272 4218 21324 4224
rect 21652 3670 21680 5646
rect 21836 4690 21864 7142
rect 21928 6458 21956 11018
rect 22020 10130 22048 12786
rect 22112 10198 22140 13738
rect 22204 13138 22232 13942
rect 22296 13240 22324 15574
rect 22388 13734 22416 15671
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22560 15360 22612 15366
rect 22560 15302 22612 15308
rect 22468 14952 22520 14958
rect 22468 14894 22520 14900
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 22296 13212 22416 13240
rect 22204 13110 22324 13138
rect 22192 12912 22244 12918
rect 22192 12854 22244 12860
rect 22204 12646 22232 12854
rect 22192 12640 22244 12646
rect 22192 12582 22244 12588
rect 22296 12238 22324 13110
rect 22388 12714 22416 13212
rect 22376 12708 22428 12714
rect 22376 12650 22428 12656
rect 22480 12434 22508 14894
rect 22572 14278 22600 15302
rect 22560 14272 22612 14278
rect 22560 14214 22612 14220
rect 22664 13938 22692 15438
rect 22756 14006 22784 18566
rect 22848 18222 22876 18634
rect 22836 18216 22888 18222
rect 22836 18158 22888 18164
rect 22848 17678 22876 18158
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22836 17672 22888 17678
rect 22836 17614 22888 17620
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 22848 16658 22876 17614
rect 23124 17202 23152 17614
rect 23112 17196 23164 17202
rect 23112 17138 23164 17144
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22836 16652 22888 16658
rect 22836 16594 22888 16600
rect 23308 16561 23336 19306
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23492 18970 23520 19110
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 23492 18426 23520 18566
rect 23480 18420 23532 18426
rect 23480 18362 23532 18368
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23388 16584 23440 16590
rect 23294 16552 23350 16561
rect 23388 16526 23440 16532
rect 23294 16487 23350 16496
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23308 16250 23336 16390
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 22836 16040 22888 16046
rect 22836 15982 22888 15988
rect 22848 15337 22876 15982
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23308 15502 23336 15846
rect 23296 15496 23348 15502
rect 23296 15438 23348 15444
rect 22834 15328 22890 15337
rect 22834 15263 22890 15272
rect 23110 15328 23166 15337
rect 23110 15263 23166 15272
rect 22836 15088 22888 15094
rect 22836 15030 22888 15036
rect 22848 14074 22876 15030
rect 23124 14958 23152 15263
rect 23202 15056 23258 15065
rect 23202 14991 23258 15000
rect 23112 14952 23164 14958
rect 23112 14894 23164 14900
rect 23216 14822 23244 14991
rect 23204 14816 23256 14822
rect 23400 14804 23428 16526
rect 23492 15366 23520 17478
rect 23584 15978 23612 19790
rect 23860 19310 23888 20703
rect 23952 19961 23980 22102
rect 23938 19952 23994 19961
rect 23938 19887 23994 19896
rect 23952 19310 23980 19887
rect 23848 19304 23900 19310
rect 23848 19246 23900 19252
rect 23940 19304 23992 19310
rect 23940 19246 23992 19252
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23676 17610 23704 18906
rect 23940 18828 23992 18834
rect 23940 18770 23992 18776
rect 23756 18624 23808 18630
rect 23756 18566 23808 18572
rect 23768 17610 23796 18566
rect 23846 17640 23902 17649
rect 23664 17604 23716 17610
rect 23664 17546 23716 17552
rect 23756 17604 23808 17610
rect 23846 17575 23902 17584
rect 23756 17546 23808 17552
rect 23768 16794 23796 17546
rect 23860 17542 23888 17575
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 23952 17320 23980 18770
rect 23860 17292 23980 17320
rect 23756 16788 23808 16794
rect 23756 16730 23808 16736
rect 23860 16522 23888 17292
rect 24044 17048 24072 26302
rect 24122 26200 24178 27000
rect 24216 26376 24268 26382
rect 24766 26330 24822 27000
rect 24216 26318 24268 26324
rect 24136 23497 24164 26200
rect 24228 23769 24256 26318
rect 24688 26302 24822 26330
rect 24308 25832 24360 25838
rect 24308 25774 24360 25780
rect 24214 23760 24270 23769
rect 24214 23695 24216 23704
rect 24268 23695 24270 23704
rect 24216 23666 24268 23672
rect 24122 23488 24178 23497
rect 24122 23423 24178 23432
rect 24124 23248 24176 23254
rect 24124 23190 24176 23196
rect 24136 22114 24164 23190
rect 24320 22658 24348 25774
rect 24584 24880 24636 24886
rect 24584 24822 24636 24828
rect 24400 24336 24452 24342
rect 24400 24278 24452 24284
rect 24228 22630 24348 22658
rect 24412 22642 24440 24278
rect 24492 24064 24544 24070
rect 24492 24006 24544 24012
rect 24504 23254 24532 24006
rect 24492 23248 24544 23254
rect 24492 23190 24544 23196
rect 24400 22636 24452 22642
rect 24228 22234 24256 22630
rect 24400 22578 24452 22584
rect 24308 22568 24360 22574
rect 24308 22510 24360 22516
rect 24216 22228 24268 22234
rect 24216 22170 24268 22176
rect 24136 22086 24256 22114
rect 24124 21888 24176 21894
rect 24124 21830 24176 21836
rect 24136 21729 24164 21830
rect 24122 21720 24178 21729
rect 24122 21655 24178 21664
rect 24124 21548 24176 21554
rect 24124 21490 24176 21496
rect 24136 20482 24164 21490
rect 24228 20874 24256 22086
rect 24320 21554 24348 22510
rect 24596 22386 24624 24822
rect 24412 22358 24624 22386
rect 24308 21548 24360 21554
rect 24308 21490 24360 21496
rect 24306 21448 24362 21457
rect 24306 21383 24308 21392
rect 24360 21383 24362 21392
rect 24308 21354 24360 21360
rect 24216 20868 24268 20874
rect 24216 20810 24268 20816
rect 24308 20800 24360 20806
rect 24308 20742 24360 20748
rect 24136 20454 24256 20482
rect 24124 20392 24176 20398
rect 24124 20334 24176 20340
rect 24136 19446 24164 20334
rect 24124 19440 24176 19446
rect 24124 19382 24176 19388
rect 24228 17882 24256 20454
rect 24320 19990 24348 20742
rect 24308 19984 24360 19990
rect 24308 19926 24360 19932
rect 24308 19712 24360 19718
rect 24308 19654 24360 19660
rect 24320 19446 24348 19654
rect 24308 19440 24360 19446
rect 24308 19382 24360 19388
rect 24308 18624 24360 18630
rect 24308 18566 24360 18572
rect 24216 17876 24268 17882
rect 24216 17818 24268 17824
rect 24320 17626 24348 18566
rect 24228 17598 24348 17626
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 24136 17270 24164 17478
rect 24124 17264 24176 17270
rect 24228 17241 24256 17598
rect 24412 17490 24440 22358
rect 24584 22228 24636 22234
rect 24584 22170 24636 22176
rect 24492 21888 24544 21894
rect 24492 21830 24544 21836
rect 24504 21010 24532 21830
rect 24492 21004 24544 21010
rect 24492 20946 24544 20952
rect 24596 20942 24624 22170
rect 24584 20936 24636 20942
rect 24584 20878 24636 20884
rect 24490 20632 24546 20641
rect 24490 20567 24546 20576
rect 24504 20330 24532 20567
rect 24492 20324 24544 20330
rect 24492 20266 24544 20272
rect 24504 18034 24532 20266
rect 24582 19816 24638 19825
rect 24582 19751 24584 19760
rect 24636 19751 24638 19760
rect 24584 19722 24636 19728
rect 24584 19304 24636 19310
rect 24584 19246 24636 19252
rect 24596 18222 24624 19246
rect 24584 18216 24636 18222
rect 24584 18158 24636 18164
rect 24504 18006 24624 18034
rect 24320 17462 24440 17490
rect 24124 17206 24176 17212
rect 24214 17232 24270 17241
rect 23952 17020 24072 17048
rect 23848 16516 23900 16522
rect 23848 16458 23900 16464
rect 23664 16448 23716 16454
rect 23664 16390 23716 16396
rect 23572 15972 23624 15978
rect 23572 15914 23624 15920
rect 23572 15564 23624 15570
rect 23572 15506 23624 15512
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23584 15026 23612 15506
rect 23572 15020 23624 15026
rect 23572 14962 23624 14968
rect 23480 14816 23532 14822
rect 23400 14776 23480 14804
rect 23204 14758 23256 14764
rect 23480 14758 23532 14764
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22926 14512 22982 14521
rect 22926 14447 22982 14456
rect 22836 14068 22888 14074
rect 22836 14010 22888 14016
rect 22744 14000 22796 14006
rect 22744 13942 22796 13948
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 22940 13818 22968 14447
rect 23386 14376 23442 14385
rect 23386 14311 23442 14320
rect 22652 13796 22704 13802
rect 22652 13738 22704 13744
rect 22756 13790 22968 13818
rect 22388 12406 22508 12434
rect 22284 12232 22336 12238
rect 22284 12174 22336 12180
rect 22284 11824 22336 11830
rect 22284 11766 22336 11772
rect 22296 11558 22324 11766
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 22100 10192 22152 10198
rect 22100 10134 22152 10140
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 22020 9994 22140 10010
rect 22008 9988 22140 9994
rect 22060 9982 22140 9988
rect 22008 9930 22060 9936
rect 22112 9654 22140 9982
rect 22192 9920 22244 9926
rect 22190 9888 22192 9897
rect 22244 9888 22246 9897
rect 22190 9823 22246 9832
rect 22100 9648 22152 9654
rect 22100 9590 22152 9596
rect 22296 9602 22324 11494
rect 22388 11082 22416 12406
rect 22664 12186 22692 13738
rect 22756 13025 22784 13790
rect 22836 13728 22888 13734
rect 22836 13670 22888 13676
rect 22742 13016 22798 13025
rect 22742 12951 22798 12960
rect 22744 12776 22796 12782
rect 22744 12718 22796 12724
rect 22480 12158 22692 12186
rect 22480 11558 22508 12158
rect 22560 12096 22612 12102
rect 22560 12038 22612 12044
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22376 11076 22428 11082
rect 22376 11018 22428 11024
rect 22192 9580 22244 9586
rect 22296 9574 22416 9602
rect 22192 9522 22244 9528
rect 22008 9444 22060 9450
rect 22008 9386 22060 9392
rect 22020 8294 22048 9386
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 22008 8288 22060 8294
rect 22008 8230 22060 8236
rect 22008 7812 22060 7818
rect 22008 7754 22060 7760
rect 22020 6866 22048 7754
rect 22008 6860 22060 6866
rect 22008 6802 22060 6808
rect 21916 6452 21968 6458
rect 21916 6394 21968 6400
rect 22008 5024 22060 5030
rect 22008 4966 22060 4972
rect 21824 4684 21876 4690
rect 21824 4626 21876 4632
rect 22020 4146 22048 4966
rect 22112 4486 22140 9318
rect 22204 8090 22232 9522
rect 22284 9512 22336 9518
rect 22284 9454 22336 9460
rect 22296 9178 22324 9454
rect 22388 9382 22416 9574
rect 22376 9376 22428 9382
rect 22376 9318 22428 9324
rect 22374 9208 22430 9217
rect 22284 9172 22336 9178
rect 22374 9143 22430 9152
rect 22284 9114 22336 9120
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 22204 7478 22232 8026
rect 22192 7472 22244 7478
rect 22192 7414 22244 7420
rect 22296 5710 22324 9114
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22388 5574 22416 9143
rect 22480 6798 22508 11494
rect 22572 7954 22600 12038
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 22664 10130 22692 11154
rect 22756 10606 22784 12718
rect 22848 11098 22876 13670
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23020 13388 23072 13394
rect 23020 13330 23072 13336
rect 23032 13297 23060 13330
rect 23018 13288 23074 13297
rect 23018 13223 23074 13232
rect 23032 12918 23060 13223
rect 23296 13184 23348 13190
rect 23296 13126 23348 13132
rect 23020 12912 23072 12918
rect 23020 12854 23072 12860
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 23308 12102 23336 13126
rect 23296 12096 23348 12102
rect 23296 12038 23348 12044
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23400 11286 23428 14311
rect 23492 13734 23520 14758
rect 23676 14074 23704 16390
rect 23848 16108 23900 16114
rect 23848 16050 23900 16056
rect 23860 15366 23888 16050
rect 23756 15360 23808 15366
rect 23756 15302 23808 15308
rect 23848 15360 23900 15366
rect 23848 15302 23900 15308
rect 23768 15162 23796 15302
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 23756 14952 23808 14958
rect 23756 14894 23808 14900
rect 23664 14068 23716 14074
rect 23664 14010 23716 14016
rect 23480 13728 23532 13734
rect 23480 13670 23532 13676
rect 23492 13326 23520 13670
rect 23480 13320 23532 13326
rect 23480 13262 23532 13268
rect 23664 13184 23716 13190
rect 23478 13152 23534 13161
rect 23664 13126 23716 13132
rect 23478 13087 23534 13096
rect 23492 12918 23520 13087
rect 23480 12912 23532 12918
rect 23480 12854 23532 12860
rect 23572 12844 23624 12850
rect 23572 12786 23624 12792
rect 23584 12434 23612 12786
rect 23492 12406 23612 12434
rect 23492 12306 23520 12406
rect 23480 12300 23532 12306
rect 23480 12242 23532 12248
rect 23492 11506 23520 12242
rect 23676 11626 23704 13126
rect 23768 12714 23796 14894
rect 23860 13977 23888 15302
rect 23846 13968 23902 13977
rect 23846 13903 23902 13912
rect 23756 12708 23808 12714
rect 23756 12650 23808 12656
rect 23756 11824 23808 11830
rect 23756 11766 23808 11772
rect 23664 11620 23716 11626
rect 23664 11562 23716 11568
rect 23492 11478 23704 11506
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 22848 11070 22968 11098
rect 22744 10600 22796 10606
rect 22940 10577 22968 11070
rect 23386 10704 23442 10713
rect 23386 10639 23442 10648
rect 23480 10668 23532 10674
rect 23296 10600 23348 10606
rect 22744 10542 22796 10548
rect 22926 10568 22982 10577
rect 23296 10542 23348 10548
rect 22926 10503 22982 10512
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22652 10124 22704 10130
rect 22704 10084 22784 10112
rect 22652 10066 22704 10072
rect 22652 9988 22704 9994
rect 22652 9930 22704 9936
rect 22664 9382 22692 9930
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22560 7948 22612 7954
rect 22560 7890 22612 7896
rect 22664 7410 22692 9318
rect 22756 9024 22784 10084
rect 23308 10062 23336 10542
rect 23400 10169 23428 10639
rect 23480 10610 23532 10616
rect 23386 10160 23442 10169
rect 23386 10095 23388 10104
rect 23440 10095 23442 10104
rect 23388 10066 23440 10072
rect 23296 10056 23348 10062
rect 23296 9998 23348 10004
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22940 9489 22968 9862
rect 23400 9722 23428 10066
rect 23388 9716 23440 9722
rect 23388 9658 23440 9664
rect 23386 9616 23442 9625
rect 23296 9580 23348 9586
rect 23492 9586 23520 10610
rect 23572 10532 23624 10538
rect 23572 10474 23624 10480
rect 23584 10130 23612 10474
rect 23676 10470 23704 11478
rect 23664 10464 23716 10470
rect 23664 10406 23716 10412
rect 23768 10266 23796 11766
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 23572 10124 23624 10130
rect 23572 10066 23624 10072
rect 23860 9602 23888 13903
rect 23952 12442 23980 17020
rect 24030 16960 24086 16969
rect 24030 16895 24086 16904
rect 24044 15178 24072 16895
rect 24136 16590 24164 17206
rect 24214 17167 24270 17176
rect 24320 16794 24348 17462
rect 24492 17060 24544 17066
rect 24492 17002 24544 17008
rect 24308 16788 24360 16794
rect 24308 16730 24360 16736
rect 24124 16584 24176 16590
rect 24124 16526 24176 16532
rect 24320 16250 24348 16730
rect 24504 16454 24532 17002
rect 24492 16448 24544 16454
rect 24492 16390 24544 16396
rect 24308 16244 24360 16250
rect 24228 16204 24308 16232
rect 24124 15700 24176 15706
rect 24124 15642 24176 15648
rect 24136 15366 24164 15642
rect 24124 15360 24176 15366
rect 24124 15302 24176 15308
rect 24044 15150 24164 15178
rect 24032 15020 24084 15026
rect 24032 14962 24084 14968
rect 23940 12436 23992 12442
rect 23940 12378 23992 12384
rect 23952 12238 23980 12378
rect 23940 12232 23992 12238
rect 23940 12174 23992 12180
rect 23938 11928 23994 11937
rect 23938 11863 23994 11872
rect 23952 11830 23980 11863
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 23386 9551 23442 9560
rect 23480 9580 23532 9586
rect 23296 9522 23348 9528
rect 22926 9480 22982 9489
rect 22926 9415 22982 9424
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22756 8996 22876 9024
rect 22848 7410 22876 8996
rect 22928 8900 22980 8906
rect 22928 8842 22980 8848
rect 22940 8634 22968 8842
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23308 7750 23336 9522
rect 23400 8945 23428 9551
rect 23480 9522 23532 9528
rect 23676 9574 23888 9602
rect 23492 9042 23520 9522
rect 23480 9036 23532 9042
rect 23480 8978 23532 8984
rect 23386 8936 23442 8945
rect 23386 8871 23442 8880
rect 23492 8514 23520 8978
rect 23492 8498 23612 8514
rect 23492 8492 23624 8498
rect 23492 8486 23572 8492
rect 23572 8434 23624 8440
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 22928 7744 22980 7750
rect 22928 7686 22980 7692
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22836 7404 22888 7410
rect 22836 7346 22888 7352
rect 22940 7342 22968 7686
rect 22928 7336 22980 7342
rect 22928 7278 22980 7284
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 23400 6798 23428 7142
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 23492 5914 23520 8230
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 23676 5794 23704 9574
rect 23756 9512 23808 9518
rect 23756 9454 23808 9460
rect 23768 8090 23796 9454
rect 23952 9194 23980 11630
rect 24044 10810 24072 14962
rect 24136 13802 24164 15150
rect 24124 13796 24176 13802
rect 24124 13738 24176 13744
rect 24228 12434 24256 16204
rect 24308 16186 24360 16192
rect 24400 16040 24452 16046
rect 24596 16028 24624 18006
rect 24452 16000 24624 16028
rect 24400 15982 24452 15988
rect 24412 15570 24440 15982
rect 24492 15904 24544 15910
rect 24492 15846 24544 15852
rect 24400 15564 24452 15570
rect 24400 15506 24452 15512
rect 24400 15428 24452 15434
rect 24400 15370 24452 15376
rect 24308 14544 24360 14550
rect 24308 14486 24360 14492
rect 24320 13433 24348 14486
rect 24306 13424 24362 13433
rect 24306 13359 24362 13368
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 24136 12406 24256 12434
rect 24032 10804 24084 10810
rect 24032 10746 24084 10752
rect 24032 10464 24084 10470
rect 24032 10406 24084 10412
rect 24044 10010 24072 10406
rect 24136 10169 24164 12406
rect 24216 12164 24268 12170
rect 24216 12106 24268 12112
rect 24228 10674 24256 12106
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 24228 10266 24256 10610
rect 24320 10470 24348 13126
rect 24412 12986 24440 15370
rect 24504 14414 24532 15846
rect 24688 15434 24716 26302
rect 24766 26200 24822 26302
rect 25410 26200 25466 27000
rect 25502 26616 25558 26625
rect 25502 26551 25558 26560
rect 25424 26092 25452 26200
rect 25516 26092 25544 26551
rect 25778 26344 25834 26353
rect 26054 26330 26110 27000
rect 26698 26330 26754 27000
rect 25834 26302 26110 26330
rect 26344 26314 26754 26330
rect 25778 26279 25834 26288
rect 26054 26200 26110 26302
rect 26332 26308 26754 26314
rect 26384 26302 26754 26308
rect 26332 26250 26384 26256
rect 26698 26200 26754 26302
rect 27342 26200 27398 27000
rect 27986 26330 28042 27000
rect 27632 26302 28042 26330
rect 25424 26064 25544 26092
rect 26884 25900 26936 25906
rect 26884 25842 26936 25848
rect 25136 25492 25188 25498
rect 25136 25434 25188 25440
rect 24860 24676 24912 24682
rect 24860 24618 24912 24624
rect 24872 24206 24900 24618
rect 24860 24200 24912 24206
rect 24860 24142 24912 24148
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 25044 23860 25096 23866
rect 25044 23802 25096 23808
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 24768 23112 24820 23118
rect 24768 23054 24820 23060
rect 24780 22574 24808 23054
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24768 21888 24820 21894
rect 24766 21856 24768 21865
rect 24820 21856 24822 21865
rect 24766 21791 24822 21800
rect 24768 20868 24820 20874
rect 24768 20810 24820 20816
rect 24780 20534 24808 20810
rect 24872 20602 24900 23598
rect 24964 21962 24992 23802
rect 25056 22710 25084 23802
rect 25148 22710 25176 25434
rect 25964 24608 26016 24614
rect 25964 24550 26016 24556
rect 25412 24268 25464 24274
rect 25412 24210 25464 24216
rect 25228 24064 25280 24070
rect 25228 24006 25280 24012
rect 25044 22704 25096 22710
rect 25044 22646 25096 22652
rect 25136 22704 25188 22710
rect 25136 22646 25188 22652
rect 25134 22400 25190 22409
rect 25134 22335 25190 22344
rect 25148 22030 25176 22335
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 24952 21956 25004 21962
rect 24952 21898 25004 21904
rect 25136 21480 25188 21486
rect 25136 21422 25188 21428
rect 25148 20942 25176 21422
rect 25136 20936 25188 20942
rect 25136 20878 25188 20884
rect 25136 20800 25188 20806
rect 25136 20742 25188 20748
rect 24860 20596 24912 20602
rect 24860 20538 24912 20544
rect 24768 20528 24820 20534
rect 24768 20470 24820 20476
rect 24780 20058 24808 20470
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24780 18358 24808 19994
rect 24872 19922 24900 20538
rect 25148 19938 25176 20742
rect 24860 19916 24912 19922
rect 24860 19858 24912 19864
rect 25056 19910 25176 19938
rect 25240 19922 25268 24006
rect 25320 23044 25372 23050
rect 25320 22986 25372 22992
rect 25332 21010 25360 22986
rect 25320 21004 25372 21010
rect 25320 20946 25372 20952
rect 25320 20800 25372 20806
rect 25320 20742 25372 20748
rect 25228 19916 25280 19922
rect 24860 19712 24912 19718
rect 24860 19654 24912 19660
rect 24872 19378 24900 19654
rect 25056 19514 25084 19910
rect 25228 19858 25280 19864
rect 25136 19780 25188 19786
rect 25136 19722 25188 19728
rect 25044 19508 25096 19514
rect 25044 19450 25096 19456
rect 24860 19372 24912 19378
rect 24860 19314 24912 19320
rect 25148 19310 25176 19722
rect 25136 19304 25188 19310
rect 25136 19246 25188 19252
rect 25228 19236 25280 19242
rect 25228 19178 25280 19184
rect 24858 19000 24914 19009
rect 24858 18935 24914 18944
rect 24872 18902 24900 18935
rect 24860 18896 24912 18902
rect 24860 18838 24912 18844
rect 24768 18352 24820 18358
rect 24768 18294 24820 18300
rect 25136 18284 25188 18290
rect 25136 18226 25188 18232
rect 25044 18148 25096 18154
rect 25044 18090 25096 18096
rect 24952 18080 25004 18086
rect 24950 18048 24952 18057
rect 25004 18048 25006 18057
rect 24950 17983 25006 17992
rect 24768 17604 24820 17610
rect 24768 17546 24820 17552
rect 24780 16658 24808 17546
rect 24860 17332 24912 17338
rect 24860 17274 24912 17280
rect 24768 16652 24820 16658
rect 24768 16594 24820 16600
rect 24766 16552 24822 16561
rect 24766 16487 24822 16496
rect 24780 16153 24808 16487
rect 24872 16250 24900 17274
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 24766 16144 24822 16153
rect 24766 16079 24768 16088
rect 24820 16079 24822 16088
rect 24768 16050 24820 16056
rect 24780 15706 24808 16050
rect 24768 15700 24820 15706
rect 24768 15642 24820 15648
rect 24676 15428 24728 15434
rect 24676 15370 24728 15376
rect 24872 15042 24900 16186
rect 25056 16046 25084 18090
rect 25044 16040 25096 16046
rect 25044 15982 25096 15988
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 24688 15014 24900 15042
rect 24688 14958 24716 15014
rect 24676 14952 24728 14958
rect 24860 14952 24912 14958
rect 24676 14894 24728 14900
rect 24780 14912 24860 14940
rect 24780 14550 24808 14912
rect 24860 14894 24912 14900
rect 24768 14544 24820 14550
rect 24964 14521 24992 15438
rect 25056 15366 25084 15982
rect 25044 15360 25096 15366
rect 25044 15302 25096 15308
rect 25148 14618 25176 18226
rect 25240 17513 25268 19178
rect 25332 18834 25360 20742
rect 25320 18828 25372 18834
rect 25320 18770 25372 18776
rect 25226 17504 25282 17513
rect 25226 17439 25282 17448
rect 25240 15434 25268 17439
rect 25424 17338 25452 24210
rect 25976 24206 26004 24550
rect 25964 24200 26016 24206
rect 25964 24142 26016 24148
rect 26424 23792 26476 23798
rect 26424 23734 26476 23740
rect 25686 23624 25742 23633
rect 25686 23559 25742 23568
rect 25502 21992 25558 22001
rect 25502 21927 25504 21936
rect 25556 21927 25558 21936
rect 25504 21898 25556 21904
rect 25596 21004 25648 21010
rect 25596 20946 25648 20952
rect 25504 20256 25556 20262
rect 25504 20198 25556 20204
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 25320 16108 25372 16114
rect 25320 16050 25372 16056
rect 25228 15428 25280 15434
rect 25228 15370 25280 15376
rect 25136 14612 25188 14618
rect 25136 14554 25188 14560
rect 24768 14486 24820 14492
rect 24950 14512 25006 14521
rect 24584 14476 24636 14482
rect 24950 14447 25006 14456
rect 24584 14418 24636 14424
rect 24492 14408 24544 14414
rect 24492 14350 24544 14356
rect 24492 14000 24544 14006
rect 24492 13942 24544 13948
rect 24504 13394 24532 13942
rect 24596 13530 24624 14418
rect 25228 14340 25280 14346
rect 25228 14282 25280 14288
rect 24676 13932 24728 13938
rect 24676 13874 24728 13880
rect 24584 13524 24636 13530
rect 24584 13466 24636 13472
rect 24492 13388 24544 13394
rect 24492 13330 24544 13336
rect 24400 12980 24452 12986
rect 24400 12922 24452 12928
rect 24596 12322 24624 13466
rect 24688 13138 24716 13874
rect 24952 13728 25004 13734
rect 24952 13670 25004 13676
rect 24964 13258 24992 13670
rect 24768 13252 24820 13258
rect 24952 13252 25004 13258
rect 24820 13212 24900 13240
rect 24768 13194 24820 13200
rect 24688 13110 24808 13138
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24400 12300 24452 12306
rect 24400 12242 24452 12248
rect 24504 12294 24624 12322
rect 24412 11762 24440 12242
rect 24400 11756 24452 11762
rect 24400 11698 24452 11704
rect 24400 10736 24452 10742
rect 24400 10678 24452 10684
rect 24308 10464 24360 10470
rect 24308 10406 24360 10412
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 24122 10160 24178 10169
rect 24122 10095 24178 10104
rect 24044 9982 24164 10010
rect 24412 9994 24440 10678
rect 23952 9166 24072 9194
rect 23848 8560 23900 8566
rect 23848 8502 23900 8508
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 23860 8022 23888 8502
rect 23848 8016 23900 8022
rect 23848 7958 23900 7964
rect 24044 6866 24072 9166
rect 24032 6860 24084 6866
rect 24032 6802 24084 6808
rect 23676 5766 23796 5794
rect 23572 5704 23624 5710
rect 23572 5646 23624 5652
rect 23664 5704 23716 5710
rect 23664 5646 23716 5652
rect 22376 5568 22428 5574
rect 22376 5510 22428 5516
rect 22928 5568 22980 5574
rect 22928 5510 22980 5516
rect 22940 5234 22968 5510
rect 23584 5370 23612 5646
rect 23572 5364 23624 5370
rect 23572 5306 23624 5312
rect 22192 5228 22244 5234
rect 22192 5170 22244 5176
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 23572 5228 23624 5234
rect 23572 5170 23624 5176
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 22112 4282 22140 4422
rect 22100 4276 22152 4282
rect 22100 4218 22152 4224
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 21640 3664 21692 3670
rect 21640 3606 21692 3612
rect 22204 3210 22232 5170
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 23296 4684 23348 4690
rect 23296 4626 23348 4632
rect 22836 4548 22888 4554
rect 22836 4490 22888 4496
rect 22744 4480 22796 4486
rect 22744 4422 22796 4428
rect 22756 3942 22784 4422
rect 22744 3936 22796 3942
rect 22744 3878 22796 3884
rect 22112 3182 22232 3210
rect 22848 3194 22876 4490
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 23308 3602 23336 4626
rect 23584 3942 23612 5170
rect 23676 4078 23704 5646
rect 23664 4072 23716 4078
rect 23768 4049 23796 5766
rect 23848 5636 23900 5642
rect 23848 5578 23900 5584
rect 23664 4014 23716 4020
rect 23754 4040 23810 4049
rect 23754 3975 23810 3984
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23572 3936 23624 3942
rect 23572 3878 23624 3884
rect 23296 3596 23348 3602
rect 23296 3538 23348 3544
rect 23308 3194 23336 3538
rect 23400 3534 23428 3878
rect 23388 3528 23440 3534
rect 23388 3470 23440 3476
rect 23584 3398 23612 3878
rect 23572 3392 23624 3398
rect 23572 3334 23624 3340
rect 22652 3188 22704 3194
rect 22112 3126 22140 3182
rect 22652 3130 22704 3136
rect 22836 3188 22888 3194
rect 22836 3130 22888 3136
rect 23296 3188 23348 3194
rect 23296 3130 23348 3136
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 22468 3120 22520 3126
rect 22468 3062 22520 3068
rect 22284 2916 22336 2922
rect 22284 2858 22336 2864
rect 20904 2508 20956 2514
rect 20904 2450 20956 2456
rect 22296 800 22324 2858
rect 22480 2582 22508 3062
rect 22468 2576 22520 2582
rect 22468 2518 22520 2524
rect 22664 2514 22692 3130
rect 23860 3126 23888 5578
rect 24032 4616 24084 4622
rect 24032 4558 24084 4564
rect 23940 4140 23992 4146
rect 23940 4082 23992 4088
rect 23952 3194 23980 4082
rect 24044 3534 24072 4558
rect 24136 3738 24164 9982
rect 24400 9988 24452 9994
rect 24400 9930 24452 9936
rect 24412 9654 24440 9930
rect 24400 9648 24452 9654
rect 24400 9590 24452 9596
rect 24308 9512 24360 9518
rect 24308 9454 24360 9460
rect 24216 8832 24268 8838
rect 24216 8774 24268 8780
rect 24228 6458 24256 8774
rect 24320 8537 24348 9454
rect 24412 8634 24440 9590
rect 24504 8974 24532 12294
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24596 11218 24624 12174
rect 24584 11212 24636 11218
rect 24584 11154 24636 11160
rect 24688 11098 24716 12922
rect 24596 11070 24716 11098
rect 24492 8968 24544 8974
rect 24492 8910 24544 8916
rect 24492 8832 24544 8838
rect 24492 8774 24544 8780
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 24306 8528 24362 8537
rect 24504 8498 24532 8774
rect 24596 8537 24624 11070
rect 24676 10464 24728 10470
rect 24676 10406 24728 10412
rect 24582 8528 24638 8537
rect 24306 8463 24362 8472
rect 24400 8492 24452 8498
rect 24400 8434 24452 8440
rect 24492 8492 24544 8498
rect 24582 8463 24638 8472
rect 24492 8434 24544 8440
rect 24412 8090 24440 8434
rect 24400 8084 24452 8090
rect 24400 8026 24452 8032
rect 24688 7410 24716 10406
rect 24780 10198 24808 13110
rect 24872 12102 24900 13212
rect 24952 13194 25004 13200
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24768 10192 24820 10198
rect 24768 10134 24820 10140
rect 24872 9874 24900 12038
rect 25240 11898 25268 14282
rect 25332 13297 25360 16050
rect 25424 15162 25452 17138
rect 25516 17134 25544 20198
rect 25608 20058 25636 20946
rect 25700 20754 25728 23559
rect 26056 23316 26108 23322
rect 26056 23258 26108 23264
rect 25872 21956 25924 21962
rect 25872 21898 25924 21904
rect 25884 21622 25912 21898
rect 25964 21888 26016 21894
rect 25964 21830 26016 21836
rect 25872 21616 25924 21622
rect 25792 21576 25872 21604
rect 25792 20874 25820 21576
rect 25872 21558 25924 21564
rect 25976 21078 26004 21830
rect 25964 21072 26016 21078
rect 25964 21014 26016 21020
rect 25780 20868 25832 20874
rect 25780 20810 25832 20816
rect 25700 20726 25820 20754
rect 25688 20324 25740 20330
rect 25688 20266 25740 20272
rect 25596 20052 25648 20058
rect 25596 19994 25648 20000
rect 25700 19938 25728 20266
rect 25608 19910 25728 19938
rect 25608 19378 25636 19910
rect 25596 19372 25648 19378
rect 25596 19314 25648 19320
rect 25608 19281 25636 19314
rect 25594 19272 25650 19281
rect 25594 19207 25650 19216
rect 25792 18426 25820 20726
rect 25962 20224 26018 20233
rect 25962 20159 26018 20168
rect 25872 19508 25924 19514
rect 25872 19450 25924 19456
rect 25884 18630 25912 19450
rect 25976 19242 26004 20159
rect 25964 19236 26016 19242
rect 25964 19178 26016 19184
rect 25964 18828 26016 18834
rect 25964 18770 26016 18776
rect 25872 18624 25924 18630
rect 25872 18566 25924 18572
rect 25976 18442 26004 18770
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 25884 18414 26004 18442
rect 25504 17128 25556 17134
rect 25504 17070 25556 17076
rect 25596 17128 25648 17134
rect 25596 17070 25648 17076
rect 25502 16008 25558 16017
rect 25502 15943 25558 15952
rect 25412 15156 25464 15162
rect 25412 15098 25464 15104
rect 25516 14657 25544 15943
rect 25608 15502 25636 17070
rect 25778 16824 25834 16833
rect 25778 16759 25834 16768
rect 25792 16114 25820 16759
rect 25884 16250 25912 18414
rect 25964 18080 26016 18086
rect 25964 18022 26016 18028
rect 25976 16969 26004 18022
rect 25962 16960 26018 16969
rect 25962 16895 26018 16904
rect 25964 16652 26016 16658
rect 25964 16594 26016 16600
rect 25872 16244 25924 16250
rect 25872 16186 25924 16192
rect 25780 16108 25832 16114
rect 25780 16050 25832 16056
rect 25872 16040 25924 16046
rect 25872 15982 25924 15988
rect 25780 15972 25832 15978
rect 25780 15914 25832 15920
rect 25686 15736 25742 15745
rect 25686 15671 25742 15680
rect 25596 15496 25648 15502
rect 25596 15438 25648 15444
rect 25502 14648 25558 14657
rect 25502 14583 25558 14592
rect 25596 14408 25648 14414
rect 25596 14350 25648 14356
rect 25318 13288 25374 13297
rect 25318 13223 25374 13232
rect 25412 12844 25464 12850
rect 25412 12786 25464 12792
rect 25320 12708 25372 12714
rect 25320 12650 25372 12656
rect 25332 12322 25360 12650
rect 25424 12434 25452 12786
rect 25424 12406 25544 12434
rect 25332 12294 25452 12322
rect 25320 12164 25372 12170
rect 25320 12106 25372 12112
rect 25228 11892 25280 11898
rect 25228 11834 25280 11840
rect 25044 11688 25096 11694
rect 25044 11630 25096 11636
rect 24952 11552 25004 11558
rect 24952 11494 25004 11500
rect 24964 11354 24992 11494
rect 24952 11348 25004 11354
rect 24952 11290 25004 11296
rect 24952 11008 25004 11014
rect 24952 10950 25004 10956
rect 24964 10062 24992 10950
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24872 9846 24992 9874
rect 24964 8786 24992 9846
rect 25056 8974 25084 11630
rect 25332 11506 25360 12106
rect 25424 11694 25452 12294
rect 25412 11688 25464 11694
rect 25412 11630 25464 11636
rect 25516 11506 25544 12406
rect 25608 11762 25636 14350
rect 25700 13190 25728 15671
rect 25792 14414 25820 15914
rect 25884 15609 25912 15982
rect 25870 15600 25926 15609
rect 25870 15535 25926 15544
rect 25872 15088 25924 15094
rect 25872 15030 25924 15036
rect 25780 14408 25832 14414
rect 25780 14350 25832 14356
rect 25792 14278 25820 14350
rect 25780 14272 25832 14278
rect 25780 14214 25832 14220
rect 25688 13184 25740 13190
rect 25688 13126 25740 13132
rect 25688 12640 25740 12646
rect 25740 12588 25820 12594
rect 25688 12582 25820 12588
rect 25700 12566 25820 12582
rect 25792 11898 25820 12566
rect 25884 11898 25912 15030
rect 25976 14414 26004 16594
rect 25964 14408 26016 14414
rect 25964 14350 26016 14356
rect 25976 14074 26004 14350
rect 25964 14068 26016 14074
rect 25964 14010 26016 14016
rect 25976 13462 26004 14010
rect 25964 13456 26016 13462
rect 25964 13398 26016 13404
rect 26068 12434 26096 23258
rect 26436 22710 26464 23734
rect 26792 23520 26844 23526
rect 26792 23462 26844 23468
rect 26700 23248 26752 23254
rect 26700 23190 26752 23196
rect 26516 22976 26568 22982
rect 26516 22918 26568 22924
rect 26424 22704 26476 22710
rect 26424 22646 26476 22652
rect 26332 22500 26384 22506
rect 26332 22442 26384 22448
rect 26344 21894 26372 22442
rect 26528 22098 26556 22918
rect 26712 22166 26740 23190
rect 26804 22273 26832 23462
rect 26896 22386 26924 25842
rect 27252 25424 27304 25430
rect 27252 25366 27304 25372
rect 27068 25016 27120 25022
rect 27068 24958 27120 24964
rect 27080 22506 27108 24958
rect 27160 23520 27212 23526
rect 27160 23462 27212 23468
rect 27172 22982 27200 23462
rect 27264 23186 27292 25366
rect 27356 23497 27384 26200
rect 27528 24404 27580 24410
rect 27528 24346 27580 24352
rect 27436 24200 27488 24206
rect 27436 24142 27488 24148
rect 27342 23488 27398 23497
rect 27342 23423 27398 23432
rect 27252 23180 27304 23186
rect 27252 23122 27304 23128
rect 27344 23044 27396 23050
rect 27344 22986 27396 22992
rect 27160 22976 27212 22982
rect 27160 22918 27212 22924
rect 27356 22710 27384 22986
rect 27344 22704 27396 22710
rect 27344 22646 27396 22652
rect 27068 22500 27120 22506
rect 27068 22442 27120 22448
rect 26896 22358 27292 22386
rect 26790 22264 26846 22273
rect 26790 22199 26846 22208
rect 27158 22264 27214 22273
rect 27158 22199 27214 22208
rect 26700 22160 26752 22166
rect 26700 22102 26752 22108
rect 26516 22092 26568 22098
rect 26516 22034 26568 22040
rect 26332 21888 26384 21894
rect 26332 21830 26384 21836
rect 26148 21616 26200 21622
rect 26148 21558 26200 21564
rect 26160 18222 26188 21558
rect 26344 21486 26372 21830
rect 26332 21480 26384 21486
rect 26332 21422 26384 21428
rect 26424 21412 26476 21418
rect 26424 21354 26476 21360
rect 26332 21344 26384 21350
rect 26332 21286 26384 21292
rect 26240 20800 26292 20806
rect 26240 20742 26292 20748
rect 26252 20602 26280 20742
rect 26240 20596 26292 20602
rect 26240 20538 26292 20544
rect 26344 20398 26372 21286
rect 26436 21010 26464 21354
rect 26424 21004 26476 21010
rect 26424 20946 26476 20952
rect 26240 20392 26292 20398
rect 26240 20334 26292 20340
rect 26332 20392 26384 20398
rect 26528 20369 26556 22034
rect 27172 22030 27200 22199
rect 27160 22024 27212 22030
rect 27160 21966 27212 21972
rect 26884 21480 26936 21486
rect 26606 21448 26662 21457
rect 26884 21422 26936 21428
rect 26606 21383 26662 21392
rect 26620 21350 26648 21383
rect 26608 21344 26660 21350
rect 26660 21304 26740 21332
rect 26608 21286 26660 21292
rect 26332 20334 26384 20340
rect 26514 20360 26570 20369
rect 26252 19990 26280 20334
rect 26344 20233 26372 20334
rect 26514 20295 26570 20304
rect 26330 20224 26386 20233
rect 26330 20159 26386 20168
rect 26240 19984 26292 19990
rect 26240 19926 26292 19932
rect 26332 19848 26384 19854
rect 26332 19790 26384 19796
rect 26240 19372 26292 19378
rect 26240 19314 26292 19320
rect 26148 18216 26200 18222
rect 26148 18158 26200 18164
rect 26252 17746 26280 19314
rect 26344 18714 26372 19790
rect 26516 19168 26568 19174
rect 26516 19110 26568 19116
rect 26528 18834 26556 19110
rect 26516 18828 26568 18834
rect 26516 18770 26568 18776
rect 26514 18728 26570 18737
rect 26344 18686 26464 18714
rect 26332 18624 26384 18630
rect 26332 18566 26384 18572
rect 26240 17740 26292 17746
rect 26240 17682 26292 17688
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 26240 17196 26292 17202
rect 26240 17138 26292 17144
rect 26160 16454 26188 17138
rect 26148 16448 26200 16454
rect 26148 16390 26200 16396
rect 26252 15706 26280 17138
rect 26240 15700 26292 15706
rect 26240 15642 26292 15648
rect 26344 15570 26372 18566
rect 26436 18358 26464 18686
rect 26514 18663 26570 18672
rect 26424 18352 26476 18358
rect 26424 18294 26476 18300
rect 26436 17610 26464 18294
rect 26424 17604 26476 17610
rect 26424 17546 26476 17552
rect 26436 17270 26464 17546
rect 26424 17264 26476 17270
rect 26424 17206 26476 17212
rect 26332 15564 26384 15570
rect 26332 15506 26384 15512
rect 26148 15496 26200 15502
rect 26148 15438 26200 15444
rect 26160 12986 26188 15438
rect 26528 15337 26556 18663
rect 26608 18420 26660 18426
rect 26608 18362 26660 18368
rect 26620 18154 26648 18362
rect 26608 18148 26660 18154
rect 26608 18090 26660 18096
rect 26606 18048 26662 18057
rect 26606 17983 26662 17992
rect 26620 17134 26648 17983
rect 26712 17218 26740 21304
rect 26792 20460 26844 20466
rect 26792 20402 26844 20408
rect 26804 17592 26832 20402
rect 26896 19961 26924 21422
rect 27264 21298 27292 22358
rect 27356 22234 27384 22646
rect 27344 22228 27396 22234
rect 27344 22170 27396 22176
rect 27344 21616 27396 21622
rect 27344 21558 27396 21564
rect 27080 21270 27292 21298
rect 27080 20806 27108 21270
rect 27356 21010 27384 21558
rect 27344 21004 27396 21010
rect 27344 20946 27396 20952
rect 26976 20800 27028 20806
rect 26976 20742 27028 20748
rect 27068 20800 27120 20806
rect 27068 20742 27120 20748
rect 27160 20800 27212 20806
rect 27160 20742 27212 20748
rect 26988 19990 27016 20742
rect 27080 20330 27108 20742
rect 27068 20324 27120 20330
rect 27068 20266 27120 20272
rect 26976 19984 27028 19990
rect 26882 19952 26938 19961
rect 27172 19938 27200 20742
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 27356 20233 27384 20402
rect 27342 20224 27398 20233
rect 27342 20159 27398 20168
rect 26976 19926 27028 19932
rect 26882 19887 26938 19896
rect 26884 19236 26936 19242
rect 26884 19178 26936 19184
rect 26896 18465 26924 19178
rect 26882 18456 26938 18465
rect 26882 18391 26938 18400
rect 26988 17882 27016 19926
rect 27080 19910 27200 19938
rect 27080 18902 27108 19910
rect 27160 19848 27212 19854
rect 27160 19790 27212 19796
rect 27068 18896 27120 18902
rect 27068 18838 27120 18844
rect 27066 18456 27122 18465
rect 27066 18391 27068 18400
rect 27120 18391 27122 18400
rect 27068 18362 27120 18368
rect 27172 18290 27200 19790
rect 27356 19689 27384 20159
rect 27448 19922 27476 24142
rect 27540 24041 27568 24346
rect 27526 24032 27582 24041
rect 27526 23967 27582 23976
rect 27528 23792 27580 23798
rect 27528 23734 27580 23740
rect 27436 19916 27488 19922
rect 27436 19858 27488 19864
rect 27342 19680 27398 19689
rect 27342 19615 27398 19624
rect 27252 19304 27304 19310
rect 27252 19246 27304 19252
rect 27264 18426 27292 19246
rect 27436 19236 27488 19242
rect 27436 19178 27488 19184
rect 27344 18828 27396 18834
rect 27344 18770 27396 18776
rect 27356 18465 27384 18770
rect 27448 18766 27476 19178
rect 27436 18760 27488 18766
rect 27436 18702 27488 18708
rect 27342 18456 27398 18465
rect 27252 18420 27304 18426
rect 27342 18391 27398 18400
rect 27252 18362 27304 18368
rect 27068 18284 27120 18290
rect 27068 18226 27120 18232
rect 27160 18284 27212 18290
rect 27212 18244 27292 18272
rect 27160 18226 27212 18232
rect 27080 18034 27108 18226
rect 27080 18006 27200 18034
rect 27066 17912 27122 17921
rect 26976 17876 27028 17882
rect 27066 17847 27122 17856
rect 26976 17818 27028 17824
rect 26804 17564 27016 17592
rect 26790 17368 26846 17377
rect 26988 17354 27016 17564
rect 27080 17542 27108 17847
rect 27068 17536 27120 17542
rect 27068 17478 27120 17484
rect 26988 17326 27108 17354
rect 26790 17303 26792 17312
rect 26844 17303 26846 17312
rect 26792 17274 26844 17280
rect 26712 17190 27016 17218
rect 26608 17128 26660 17134
rect 26700 17128 26752 17134
rect 26608 17070 26660 17076
rect 26698 17096 26700 17105
rect 26752 17096 26754 17105
rect 26698 17031 26754 17040
rect 26712 16794 26740 17031
rect 26608 16788 26660 16794
rect 26608 16730 26660 16736
rect 26700 16788 26752 16794
rect 26700 16730 26752 16736
rect 26620 15706 26648 16730
rect 26700 16448 26752 16454
rect 26700 16390 26752 16396
rect 26712 16250 26740 16390
rect 26700 16244 26752 16250
rect 26700 16186 26752 16192
rect 26884 16176 26936 16182
rect 26698 16144 26754 16153
rect 26884 16118 26936 16124
rect 26698 16079 26700 16088
rect 26752 16079 26754 16088
rect 26700 16050 26752 16056
rect 26792 15904 26844 15910
rect 26792 15846 26844 15852
rect 26608 15700 26660 15706
rect 26608 15642 26660 15648
rect 26514 15328 26570 15337
rect 26514 15263 26570 15272
rect 26606 15056 26662 15065
rect 26606 14991 26662 15000
rect 26620 14958 26648 14991
rect 26240 14952 26292 14958
rect 26240 14894 26292 14900
rect 26424 14952 26476 14958
rect 26424 14894 26476 14900
rect 26608 14952 26660 14958
rect 26608 14894 26660 14900
rect 26252 14793 26280 14894
rect 26238 14784 26294 14793
rect 26238 14719 26294 14728
rect 26148 12980 26200 12986
rect 26148 12922 26200 12928
rect 26240 12776 26292 12782
rect 26240 12718 26292 12724
rect 26332 12776 26384 12782
rect 26332 12718 26384 12724
rect 26068 12406 26188 12434
rect 25780 11892 25832 11898
rect 25780 11834 25832 11840
rect 25872 11892 25924 11898
rect 25872 11834 25924 11840
rect 26056 11824 26108 11830
rect 26056 11766 26108 11772
rect 25596 11756 25648 11762
rect 25596 11698 25648 11704
rect 26068 11665 26096 11766
rect 26054 11656 26110 11665
rect 26054 11591 26110 11600
rect 25332 11478 25544 11506
rect 25228 11348 25280 11354
rect 25228 11290 25280 11296
rect 25136 11076 25188 11082
rect 25136 11018 25188 11024
rect 25148 9178 25176 11018
rect 25240 10130 25268 11290
rect 25332 11064 25360 11478
rect 25412 11076 25464 11082
rect 25332 11036 25412 11064
rect 25412 11018 25464 11024
rect 25228 10124 25280 10130
rect 25228 10066 25280 10072
rect 25136 9172 25188 9178
rect 25136 9114 25188 9120
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 24964 8758 25084 8786
rect 24766 8664 24822 8673
rect 24766 8599 24768 8608
rect 24820 8599 24822 8608
rect 24768 8570 24820 8576
rect 25056 7886 25084 8758
rect 24952 7880 25004 7886
rect 24952 7822 25004 7828
rect 25044 7880 25096 7886
rect 25044 7822 25096 7828
rect 24676 7404 24728 7410
rect 24676 7346 24728 7352
rect 24676 7200 24728 7206
rect 24676 7142 24728 7148
rect 24216 6452 24268 6458
rect 24216 6394 24268 6400
rect 24688 6322 24716 7142
rect 24964 6458 24992 7822
rect 25240 7410 25268 10066
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 25228 7200 25280 7206
rect 25228 7142 25280 7148
rect 25240 6798 25268 7142
rect 25228 6792 25280 6798
rect 25228 6734 25280 6740
rect 24952 6452 25004 6458
rect 24952 6394 25004 6400
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 25332 6118 25360 9998
rect 25424 9994 25452 11018
rect 25872 10600 25924 10606
rect 25872 10542 25924 10548
rect 26056 10600 26108 10606
rect 26056 10542 26108 10548
rect 25412 9988 25464 9994
rect 25412 9930 25464 9936
rect 25884 6866 25912 10542
rect 26068 10282 26096 10542
rect 25976 10266 26096 10282
rect 25964 10260 26096 10266
rect 26016 10254 26096 10260
rect 25964 10202 26016 10208
rect 25962 10160 26018 10169
rect 25962 10095 25964 10104
rect 26016 10095 26018 10104
rect 25964 10066 26016 10072
rect 25962 9888 26018 9897
rect 25962 9823 26018 9832
rect 25976 9586 26004 9823
rect 25964 9580 26016 9586
rect 25964 9522 26016 9528
rect 25976 9110 26004 9522
rect 25964 9104 26016 9110
rect 25964 9046 26016 9052
rect 25964 8832 26016 8838
rect 25964 8774 26016 8780
rect 25976 8498 26004 8774
rect 25964 8492 26016 8498
rect 25964 8434 26016 8440
rect 25872 6860 25924 6866
rect 25872 6802 25924 6808
rect 25320 6112 25372 6118
rect 25320 6054 25372 6060
rect 24676 5228 24728 5234
rect 24676 5170 24728 5176
rect 24308 5160 24360 5166
rect 24308 5102 24360 5108
rect 24320 4078 24348 5102
rect 24688 4826 24716 5170
rect 24768 5024 24820 5030
rect 24768 4966 24820 4972
rect 24860 5024 24912 5030
rect 24860 4966 24912 4972
rect 24676 4820 24728 4826
rect 24676 4762 24728 4768
rect 24780 4690 24808 4966
rect 24768 4684 24820 4690
rect 24768 4626 24820 4632
rect 24584 4276 24636 4282
rect 24584 4218 24636 4224
rect 24308 4072 24360 4078
rect 24308 4014 24360 4020
rect 24124 3732 24176 3738
rect 24124 3674 24176 3680
rect 24492 3664 24544 3670
rect 24492 3606 24544 3612
rect 24032 3528 24084 3534
rect 24032 3470 24084 3476
rect 24400 3460 24452 3466
rect 24400 3402 24452 3408
rect 23940 3188 23992 3194
rect 23940 3130 23992 3136
rect 23572 3120 23624 3126
rect 23572 3062 23624 3068
rect 23848 3120 23900 3126
rect 23848 3062 23900 3068
rect 23584 2938 23612 3062
rect 23848 2984 23900 2990
rect 23584 2932 23848 2938
rect 23584 2926 23900 2932
rect 23584 2910 23888 2926
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 22652 2508 22704 2514
rect 22652 2450 22704 2456
rect 23952 2446 23980 3130
rect 23940 2440 23992 2446
rect 23940 2382 23992 2388
rect 24412 800 24440 3402
rect 24504 3194 24532 3606
rect 24596 3466 24624 4218
rect 24872 3602 24900 4966
rect 25228 4616 25280 4622
rect 25228 4558 25280 4564
rect 25240 4282 25268 4558
rect 25228 4276 25280 4282
rect 25228 4218 25280 4224
rect 24952 4072 25004 4078
rect 24950 4040 24952 4049
rect 25004 4040 25006 4049
rect 24950 3975 25006 3984
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 24584 3460 24636 3466
rect 24584 3402 24636 3408
rect 24492 3188 24544 3194
rect 24492 3130 24544 3136
rect 24596 2774 24624 3402
rect 26068 2990 26096 10254
rect 26160 5302 26188 12406
rect 26252 10810 26280 12718
rect 26344 11354 26372 12718
rect 26436 11626 26464 14894
rect 26516 14272 26568 14278
rect 26516 14214 26568 14220
rect 26528 14074 26556 14214
rect 26516 14068 26568 14074
rect 26516 14010 26568 14016
rect 26804 13394 26832 15846
rect 26792 13388 26844 13394
rect 26792 13330 26844 13336
rect 26516 12844 26568 12850
rect 26516 12786 26568 12792
rect 26424 11620 26476 11626
rect 26424 11562 26476 11568
rect 26332 11348 26384 11354
rect 26332 11290 26384 11296
rect 26240 10804 26292 10810
rect 26240 10746 26292 10752
rect 26436 10713 26464 11562
rect 26528 10810 26556 12786
rect 26896 12714 26924 16118
rect 26988 15201 27016 17190
rect 27080 15609 27108 17326
rect 27172 17105 27200 18006
rect 27264 17814 27292 18244
rect 27540 18222 27568 23734
rect 27632 23254 27660 26302
rect 27986 26200 28042 26302
rect 28630 26200 28686 27000
rect 29274 26200 29330 27000
rect 29366 26208 29422 26217
rect 28356 26104 28408 26110
rect 28356 26046 28408 26052
rect 28264 25152 28316 25158
rect 28264 25094 28316 25100
rect 28276 24206 28304 25094
rect 28264 24200 28316 24206
rect 28264 24142 28316 24148
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 27896 23860 27948 23866
rect 28368 23848 28396 26046
rect 28448 24268 28500 24274
rect 28448 24210 28500 24216
rect 27896 23802 27948 23808
rect 28276 23820 28396 23848
rect 27804 23724 27856 23730
rect 27804 23666 27856 23672
rect 27712 23656 27764 23662
rect 27712 23598 27764 23604
rect 27620 23248 27672 23254
rect 27620 23190 27672 23196
rect 27620 22976 27672 22982
rect 27620 22918 27672 22924
rect 27632 22778 27660 22918
rect 27620 22772 27672 22778
rect 27620 22714 27672 22720
rect 27620 22636 27672 22642
rect 27620 22578 27672 22584
rect 27632 22030 27660 22578
rect 27620 22024 27672 22030
rect 27620 21966 27672 21972
rect 27620 21412 27672 21418
rect 27620 21354 27672 21360
rect 27632 20210 27660 21354
rect 27724 20482 27752 23598
rect 27816 22642 27844 23666
rect 27908 23186 27936 23802
rect 28276 23236 28304 23820
rect 28356 23656 28408 23662
rect 28356 23598 28408 23604
rect 28368 23361 28396 23598
rect 28354 23352 28410 23361
rect 28354 23287 28410 23296
rect 28276 23208 28396 23236
rect 27896 23180 27948 23186
rect 27896 23122 27948 23128
rect 28080 23112 28132 23118
rect 28078 23080 28080 23089
rect 28132 23080 28134 23089
rect 28078 23015 28134 23024
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 27804 22636 27856 22642
rect 27804 22578 27856 22584
rect 28368 22574 28396 23208
rect 28460 23186 28488 24210
rect 28538 24032 28594 24041
rect 28538 23967 28594 23976
rect 28448 23180 28500 23186
rect 28448 23122 28500 23128
rect 28356 22568 28408 22574
rect 28356 22510 28408 22516
rect 28460 22438 28488 23122
rect 28552 23118 28580 23967
rect 28644 23497 28672 26200
rect 28724 24268 28776 24274
rect 28724 24210 28776 24216
rect 28630 23488 28686 23497
rect 28630 23423 28686 23432
rect 28736 23361 28764 24210
rect 29184 24200 29236 24206
rect 29182 24168 29184 24177
rect 29236 24168 29238 24177
rect 29182 24103 29238 24112
rect 29000 24064 29052 24070
rect 29000 24006 29052 24012
rect 28722 23352 28778 23361
rect 28722 23287 28778 23296
rect 28816 23248 28868 23254
rect 28816 23190 28868 23196
rect 28540 23112 28592 23118
rect 28540 23054 28592 23060
rect 28632 23112 28684 23118
rect 28632 23054 28684 23060
rect 28722 23080 28778 23089
rect 28538 22808 28594 22817
rect 28538 22743 28594 22752
rect 28448 22432 28500 22438
rect 28552 22409 28580 22743
rect 28644 22710 28672 23054
rect 28722 23015 28778 23024
rect 28632 22704 28684 22710
rect 28632 22646 28684 22652
rect 28448 22374 28500 22380
rect 28538 22400 28594 22409
rect 28538 22335 28594 22344
rect 28538 22264 28594 22273
rect 28538 22199 28540 22208
rect 28592 22199 28594 22208
rect 28540 22170 28592 22176
rect 28448 22024 28500 22030
rect 28448 21966 28500 21972
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 27804 21480 27856 21486
rect 27804 21422 27856 21428
rect 27816 21146 27844 21422
rect 28172 21344 28224 21350
rect 28172 21286 28224 21292
rect 28356 21344 28408 21350
rect 28356 21286 28408 21292
rect 28184 21146 28212 21286
rect 27804 21140 27856 21146
rect 27804 21082 27856 21088
rect 28172 21140 28224 21146
rect 28172 21082 28224 21088
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 28368 20602 28396 21286
rect 28356 20596 28408 20602
rect 28356 20538 28408 20544
rect 27724 20454 27844 20482
rect 27816 20398 27844 20454
rect 27804 20392 27856 20398
rect 27804 20334 27856 20340
rect 28356 20324 28408 20330
rect 28356 20266 28408 20272
rect 27632 20182 27844 20210
rect 27618 19816 27674 19825
rect 27618 19751 27674 19760
rect 27712 19780 27764 19786
rect 27528 18216 27580 18222
rect 27342 18184 27398 18193
rect 27528 18158 27580 18164
rect 27342 18119 27398 18128
rect 27252 17808 27304 17814
rect 27252 17750 27304 17756
rect 27264 17202 27292 17750
rect 27252 17196 27304 17202
rect 27252 17138 27304 17144
rect 27158 17096 27214 17105
rect 27158 17031 27214 17040
rect 27356 16658 27384 18119
rect 27632 18034 27660 19751
rect 27712 19722 27764 19728
rect 27724 19417 27752 19722
rect 27710 19408 27766 19417
rect 27710 19343 27766 19352
rect 27712 18896 27764 18902
rect 27816 18873 27844 20182
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 28080 19508 28132 19514
rect 28080 19450 28132 19456
rect 27988 19304 28040 19310
rect 27988 19246 28040 19252
rect 27712 18838 27764 18844
rect 27802 18864 27858 18873
rect 27540 18006 27660 18034
rect 27436 17876 27488 17882
rect 27436 17818 27488 17824
rect 27448 17542 27476 17818
rect 27436 17536 27488 17542
rect 27436 17478 27488 17484
rect 27436 17264 27488 17270
rect 27436 17206 27488 17212
rect 27344 16652 27396 16658
rect 27344 16594 27396 16600
rect 27158 16416 27214 16425
rect 27158 16351 27214 16360
rect 27066 15600 27122 15609
rect 27066 15535 27122 15544
rect 26974 15192 27030 15201
rect 26974 15127 27030 15136
rect 26976 15088 27028 15094
rect 26976 15030 27028 15036
rect 26884 12708 26936 12714
rect 26884 12650 26936 12656
rect 26606 12200 26662 12209
rect 26606 12135 26662 12144
rect 26516 10804 26568 10810
rect 26516 10746 26568 10752
rect 26422 10704 26478 10713
rect 26422 10639 26478 10648
rect 26620 9518 26648 12135
rect 26792 11212 26844 11218
rect 26792 11154 26844 11160
rect 26804 10130 26832 11154
rect 26988 10606 27016 15030
rect 27080 12442 27108 15535
rect 27172 14958 27200 16351
rect 27356 16250 27384 16594
rect 27344 16244 27396 16250
rect 27344 16186 27396 16192
rect 27344 16108 27396 16114
rect 27344 16050 27396 16056
rect 27252 15972 27304 15978
rect 27252 15914 27304 15920
rect 27264 15162 27292 15914
rect 27356 15910 27384 16050
rect 27344 15904 27396 15910
rect 27344 15846 27396 15852
rect 27252 15156 27304 15162
rect 27252 15098 27304 15104
rect 27356 15042 27384 15846
rect 27264 15014 27384 15042
rect 27160 14952 27212 14958
rect 27160 14894 27212 14900
rect 27160 13932 27212 13938
rect 27160 13874 27212 13880
rect 27172 13530 27200 13874
rect 27160 13524 27212 13530
rect 27160 13466 27212 13472
rect 27264 12889 27292 15014
rect 27344 14408 27396 14414
rect 27448 14396 27476 17206
rect 27540 16833 27568 18006
rect 27620 17876 27672 17882
rect 27620 17818 27672 17824
rect 27632 17785 27660 17818
rect 27618 17776 27674 17785
rect 27618 17711 27674 17720
rect 27724 17066 27752 18838
rect 27802 18799 27858 18808
rect 28000 18737 28028 19246
rect 27986 18728 28042 18737
rect 27986 18663 28042 18672
rect 28092 18630 28120 19450
rect 28262 19408 28318 19417
rect 28262 19343 28318 19352
rect 28172 19168 28224 19174
rect 28172 19110 28224 19116
rect 28184 18698 28212 19110
rect 28276 19009 28304 19343
rect 28262 19000 28318 19009
rect 28262 18935 28318 18944
rect 28172 18692 28224 18698
rect 28172 18634 28224 18640
rect 28080 18624 28132 18630
rect 28080 18566 28132 18572
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 28080 17876 28132 17882
rect 28080 17818 28132 17824
rect 28092 17746 28120 17818
rect 28080 17740 28132 17746
rect 28080 17682 28132 17688
rect 28368 17678 28396 20266
rect 28460 18057 28488 21966
rect 28552 19854 28580 22170
rect 28644 22166 28672 22646
rect 28632 22160 28684 22166
rect 28632 22102 28684 22108
rect 28632 21344 28684 21350
rect 28632 21286 28684 21292
rect 28644 21078 28672 21286
rect 28632 21072 28684 21078
rect 28632 21014 28684 21020
rect 28736 20942 28764 23015
rect 28828 22234 28856 23190
rect 28908 23044 28960 23050
rect 28908 22986 28960 22992
rect 28816 22228 28868 22234
rect 28816 22170 28868 22176
rect 28814 22128 28870 22137
rect 28814 22063 28870 22072
rect 28828 21554 28856 22063
rect 28920 22001 28948 22986
rect 28906 21992 28962 22001
rect 28906 21927 28962 21936
rect 28908 21888 28960 21894
rect 28908 21830 28960 21836
rect 28816 21548 28868 21554
rect 28816 21490 28868 21496
rect 28920 21418 28948 21830
rect 29012 21622 29040 24006
rect 29090 23216 29146 23225
rect 29090 23151 29092 23160
rect 29144 23151 29146 23160
rect 29092 23122 29144 23128
rect 29196 22778 29224 24103
rect 29288 23322 29316 26200
rect 29918 26200 29974 27000
rect 30562 26330 30618 27000
rect 30562 26302 31064 26330
rect 30562 26200 30618 26302
rect 29366 26143 29422 26152
rect 29276 23316 29328 23322
rect 29276 23258 29328 23264
rect 29184 22772 29236 22778
rect 29184 22714 29236 22720
rect 29092 22568 29144 22574
rect 29092 22510 29144 22516
rect 29104 22273 29132 22510
rect 29090 22264 29146 22273
rect 29090 22199 29146 22208
rect 29092 21956 29144 21962
rect 29092 21898 29144 21904
rect 29000 21616 29052 21622
rect 29000 21558 29052 21564
rect 28908 21412 28960 21418
rect 28908 21354 28960 21360
rect 28816 21140 28868 21146
rect 28816 21082 28868 21088
rect 28828 21049 28856 21082
rect 28814 21040 28870 21049
rect 28814 20975 28870 20984
rect 28724 20936 28776 20942
rect 28724 20878 28776 20884
rect 29012 20806 29040 21558
rect 28908 20800 28960 20806
rect 28908 20742 28960 20748
rect 29000 20800 29052 20806
rect 29000 20742 29052 20748
rect 28920 20602 28948 20742
rect 29104 20618 29132 21898
rect 29380 21570 29408 26143
rect 29460 24200 29512 24206
rect 29460 24142 29512 24148
rect 28724 20596 28776 20602
rect 28724 20538 28776 20544
rect 28908 20596 28960 20602
rect 28908 20538 28960 20544
rect 29012 20590 29132 20618
rect 29196 21542 29408 21570
rect 28632 20460 28684 20466
rect 28632 20402 28684 20408
rect 28540 19848 28592 19854
rect 28540 19790 28592 19796
rect 28540 19304 28592 19310
rect 28540 19246 28592 19252
rect 28446 18048 28502 18057
rect 28446 17983 28502 17992
rect 28356 17672 28408 17678
rect 28356 17614 28408 17620
rect 27896 17604 27948 17610
rect 27816 17564 27896 17592
rect 27712 17060 27764 17066
rect 27712 17002 27764 17008
rect 27710 16960 27766 16969
rect 27710 16895 27766 16904
rect 27526 16824 27582 16833
rect 27526 16759 27582 16768
rect 27540 16726 27568 16759
rect 27528 16720 27580 16726
rect 27528 16662 27580 16668
rect 27620 16516 27672 16522
rect 27620 16458 27672 16464
rect 27632 16046 27660 16458
rect 27724 16454 27752 16895
rect 27712 16448 27764 16454
rect 27712 16390 27764 16396
rect 27620 16040 27672 16046
rect 27620 15982 27672 15988
rect 27724 15910 27752 16390
rect 27712 15904 27764 15910
rect 27712 15846 27764 15852
rect 27528 15632 27580 15638
rect 27526 15600 27528 15609
rect 27580 15600 27582 15609
rect 27526 15535 27582 15544
rect 27620 15564 27672 15570
rect 27620 15506 27672 15512
rect 27712 15564 27764 15570
rect 27712 15506 27764 15512
rect 27528 15428 27580 15434
rect 27528 15370 27580 15376
rect 27540 15337 27568 15370
rect 27526 15328 27582 15337
rect 27526 15263 27582 15272
rect 27526 14920 27582 14929
rect 27526 14855 27582 14864
rect 27396 14368 27476 14396
rect 27344 14350 27396 14356
rect 27356 14006 27384 14350
rect 27344 14000 27396 14006
rect 27344 13942 27396 13948
rect 27436 13252 27488 13258
rect 27436 13194 27488 13200
rect 27250 12880 27306 12889
rect 27250 12815 27306 12824
rect 27068 12436 27120 12442
rect 27068 12378 27120 12384
rect 27068 12096 27120 12102
rect 27252 12096 27304 12102
rect 27068 12038 27120 12044
rect 27250 12064 27252 12073
rect 27304 12064 27306 12073
rect 27080 11558 27108 12038
rect 27250 11999 27306 12008
rect 27264 11830 27292 11999
rect 27252 11824 27304 11830
rect 27252 11766 27304 11772
rect 27344 11620 27396 11626
rect 27344 11562 27396 11568
rect 27068 11552 27120 11558
rect 27068 11494 27120 11500
rect 27160 11552 27212 11558
rect 27160 11494 27212 11500
rect 27252 11552 27304 11558
rect 27252 11494 27304 11500
rect 26976 10600 27028 10606
rect 26976 10542 27028 10548
rect 26792 10124 26844 10130
rect 26792 10066 26844 10072
rect 27080 9674 27108 11494
rect 27172 10742 27200 11494
rect 27264 11218 27292 11494
rect 27252 11212 27304 11218
rect 27252 11154 27304 11160
rect 27160 10736 27212 10742
rect 27160 10678 27212 10684
rect 27356 10033 27384 11562
rect 27342 10024 27398 10033
rect 27342 9959 27398 9968
rect 27080 9646 27200 9674
rect 26608 9512 26660 9518
rect 26608 9454 26660 9460
rect 26620 8498 26648 9454
rect 27068 8968 27120 8974
rect 27068 8910 27120 8916
rect 26608 8492 26660 8498
rect 26608 8434 26660 8440
rect 27080 8090 27108 8910
rect 27068 8084 27120 8090
rect 27068 8026 27120 8032
rect 26976 6656 27028 6662
rect 26976 6598 27028 6604
rect 26988 6390 27016 6598
rect 26976 6384 27028 6390
rect 26976 6326 27028 6332
rect 26148 5296 26200 5302
rect 26148 5238 26200 5244
rect 27172 4486 27200 9646
rect 27252 9512 27304 9518
rect 27252 9454 27304 9460
rect 27264 8906 27292 9454
rect 27252 8900 27304 8906
rect 27252 8842 27304 8848
rect 27448 8022 27476 13194
rect 27436 8016 27488 8022
rect 27436 7958 27488 7964
rect 27540 6118 27568 14855
rect 27632 12782 27660 15506
rect 27724 14618 27752 15506
rect 27816 15094 27844 17564
rect 27896 17546 27948 17552
rect 28552 17542 28580 19246
rect 28644 17898 28672 20402
rect 28736 19514 28764 20538
rect 29012 20482 29040 20590
rect 28920 20454 29040 20482
rect 29090 20496 29146 20505
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 28816 19508 28868 19514
rect 28816 19450 28868 19456
rect 28722 19272 28778 19281
rect 28722 19207 28778 19216
rect 28736 18952 28764 19207
rect 28828 19122 28856 19450
rect 28920 19258 28948 20454
rect 29090 20431 29146 20440
rect 29104 19514 29132 20431
rect 29092 19508 29144 19514
rect 29092 19450 29144 19456
rect 28920 19230 29132 19258
rect 29000 19168 29052 19174
rect 28828 19094 28948 19122
rect 29000 19110 29052 19116
rect 28736 18924 28856 18952
rect 28724 18828 28776 18834
rect 28724 18770 28776 18776
rect 28736 18290 28764 18770
rect 28828 18358 28856 18924
rect 28920 18766 28948 19094
rect 29012 18970 29040 19110
rect 29000 18964 29052 18970
rect 29000 18906 29052 18912
rect 28908 18760 28960 18766
rect 28908 18702 28960 18708
rect 29104 18578 29132 19230
rect 28920 18550 29132 18578
rect 28816 18352 28868 18358
rect 28816 18294 28868 18300
rect 28724 18284 28776 18290
rect 28724 18226 28776 18232
rect 28644 17870 28764 17898
rect 28632 17740 28684 17746
rect 28632 17682 28684 17688
rect 28448 17536 28500 17542
rect 28448 17478 28500 17484
rect 28540 17536 28592 17542
rect 28540 17478 28592 17484
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 27986 17232 28042 17241
rect 27986 17167 28042 17176
rect 28000 16794 28028 17167
rect 28356 16992 28408 16998
rect 28356 16934 28408 16940
rect 27988 16788 28040 16794
rect 27988 16730 28040 16736
rect 27894 16688 27950 16697
rect 28000 16658 28028 16730
rect 27894 16623 27950 16632
rect 27988 16652 28040 16658
rect 27908 16590 27936 16623
rect 27988 16594 28040 16600
rect 27896 16584 27948 16590
rect 27896 16526 27948 16532
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 28368 16114 28396 16934
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 27894 15736 27950 15745
rect 27894 15671 27950 15680
rect 27908 15434 27936 15671
rect 28356 15564 28408 15570
rect 28356 15506 28408 15512
rect 27896 15428 27948 15434
rect 27896 15370 27948 15376
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 27988 15156 28040 15162
rect 27988 15098 28040 15104
rect 27804 15088 27856 15094
rect 27804 15030 27856 15036
rect 27894 15056 27950 15065
rect 27894 14991 27950 15000
rect 27908 14958 27936 14991
rect 27896 14952 27948 14958
rect 28000 14929 28028 15098
rect 28264 15020 28316 15026
rect 28264 14962 28316 14968
rect 28276 14929 28304 14962
rect 27896 14894 27948 14900
rect 27986 14920 28042 14929
rect 27908 14618 27936 14894
rect 27986 14855 28042 14864
rect 28262 14920 28318 14929
rect 28262 14855 28318 14864
rect 27712 14612 27764 14618
rect 27712 14554 27764 14560
rect 27896 14612 27948 14618
rect 27896 14554 27948 14560
rect 28000 14532 28028 14855
rect 28262 14648 28318 14657
rect 28262 14583 28264 14592
rect 28316 14583 28318 14592
rect 28264 14554 28316 14560
rect 28080 14544 28132 14550
rect 27710 14512 27766 14521
rect 28000 14504 28080 14532
rect 28080 14486 28132 14492
rect 27710 14447 27766 14456
rect 27724 14278 27752 14447
rect 28276 14278 28304 14554
rect 27712 14272 27764 14278
rect 27712 14214 27764 14220
rect 28264 14272 28316 14278
rect 28264 14214 28316 14220
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 28368 13410 28396 15506
rect 28460 15337 28488 17478
rect 28540 16652 28592 16658
rect 28540 16594 28592 16600
rect 28446 15328 28502 15337
rect 28446 15263 28502 15272
rect 28448 15156 28500 15162
rect 28448 15098 28500 15104
rect 28460 14822 28488 15098
rect 28552 14822 28580 16594
rect 28448 14816 28500 14822
rect 28540 14816 28592 14822
rect 28448 14758 28500 14764
rect 28538 14784 28540 14793
rect 28592 14784 28594 14793
rect 28538 14719 28594 14728
rect 28368 13382 28488 13410
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 28368 12918 28396 13382
rect 28460 13326 28488 13382
rect 28448 13320 28500 13326
rect 28448 13262 28500 13268
rect 28540 13252 28592 13258
rect 28540 13194 28592 13200
rect 28552 12918 28580 13194
rect 28356 12912 28408 12918
rect 28356 12854 28408 12860
rect 28540 12912 28592 12918
rect 28540 12854 28592 12860
rect 27620 12776 27672 12782
rect 27620 12718 27672 12724
rect 28644 12434 28672 17682
rect 28736 16522 28764 17870
rect 28816 17264 28868 17270
rect 28816 17206 28868 17212
rect 28828 16658 28856 17206
rect 28816 16652 28868 16658
rect 28816 16594 28868 16600
rect 28920 16538 28948 18550
rect 29000 17536 29052 17542
rect 29000 17478 29052 17484
rect 28724 16516 28776 16522
rect 28724 16458 28776 16464
rect 28828 16510 28948 16538
rect 28828 15162 28856 16510
rect 28908 16448 28960 16454
rect 28908 16390 28960 16396
rect 28920 16250 28948 16390
rect 28908 16244 28960 16250
rect 28908 16186 28960 16192
rect 29012 16130 29040 17478
rect 29196 16998 29224 21542
rect 29276 21480 29328 21486
rect 29276 21422 29328 21428
rect 29288 20534 29316 21422
rect 29472 21418 29500 24142
rect 29736 23520 29788 23526
rect 29932 23497 29960 26200
rect 30746 25800 30802 25809
rect 30746 25735 30802 25744
rect 30564 25356 30616 25362
rect 30564 25298 30616 25304
rect 30012 24744 30064 24750
rect 30012 24686 30064 24692
rect 30024 24206 30052 24686
rect 30012 24200 30064 24206
rect 30012 24142 30064 24148
rect 30024 23526 30052 24142
rect 30472 24132 30524 24138
rect 30472 24074 30524 24080
rect 30288 24064 30340 24070
rect 30288 24006 30340 24012
rect 30380 24064 30432 24070
rect 30380 24006 30432 24012
rect 30104 23656 30156 23662
rect 30104 23598 30156 23604
rect 30012 23520 30064 23526
rect 29736 23462 29788 23468
rect 29918 23488 29974 23497
rect 29644 22976 29696 22982
rect 29644 22918 29696 22924
rect 29656 22137 29684 22918
rect 29642 22128 29698 22137
rect 29642 22063 29698 22072
rect 29748 22094 29776 23462
rect 30012 23462 30064 23468
rect 29918 23423 29974 23432
rect 30024 22778 30052 23462
rect 30012 22772 30064 22778
rect 30012 22714 30064 22720
rect 29918 22128 29974 22137
rect 29828 22094 29880 22098
rect 29748 22092 29880 22094
rect 29748 22066 29828 22092
rect 29918 22063 29974 22072
rect 29828 22034 29880 22040
rect 29736 21548 29788 21554
rect 29736 21490 29788 21496
rect 29460 21412 29512 21418
rect 29460 21354 29512 21360
rect 29368 20800 29420 20806
rect 29368 20742 29420 20748
rect 29276 20528 29328 20534
rect 29276 20470 29328 20476
rect 29276 20256 29328 20262
rect 29274 20224 29276 20233
rect 29328 20224 29330 20233
rect 29274 20159 29330 20168
rect 29274 20088 29330 20097
rect 29274 20023 29330 20032
rect 29288 19990 29316 20023
rect 29276 19984 29328 19990
rect 29276 19926 29328 19932
rect 29276 19712 29328 19718
rect 29276 19654 29328 19660
rect 29288 19417 29316 19654
rect 29274 19408 29330 19417
rect 29274 19343 29276 19352
rect 29328 19343 29330 19352
rect 29276 19314 29328 19320
rect 29274 19272 29330 19281
rect 29274 19207 29276 19216
rect 29328 19207 29330 19216
rect 29276 19178 29328 19184
rect 29274 19000 29330 19009
rect 29274 18935 29330 18944
rect 29288 18766 29316 18935
rect 29380 18834 29408 20742
rect 29472 19786 29500 21354
rect 29552 20800 29604 20806
rect 29552 20742 29604 20748
rect 29460 19780 29512 19786
rect 29460 19722 29512 19728
rect 29472 19378 29500 19722
rect 29460 19372 29512 19378
rect 29460 19314 29512 19320
rect 29368 18828 29420 18834
rect 29368 18770 29420 18776
rect 29276 18760 29328 18766
rect 29276 18702 29328 18708
rect 29184 16992 29236 16998
rect 29184 16934 29236 16940
rect 29196 16697 29224 16934
rect 29182 16688 29238 16697
rect 29182 16623 29238 16632
rect 29288 16590 29316 18702
rect 29368 18624 29420 18630
rect 29368 18566 29420 18572
rect 29460 18624 29512 18630
rect 29460 18566 29512 18572
rect 29276 16584 29328 16590
rect 29276 16526 29328 16532
rect 28920 16102 29040 16130
rect 28920 15570 28948 16102
rect 29276 16040 29328 16046
rect 29276 15982 29328 15988
rect 28908 15564 28960 15570
rect 28908 15506 28960 15512
rect 28724 15156 28776 15162
rect 28724 15098 28776 15104
rect 28816 15156 28868 15162
rect 28816 15098 28868 15104
rect 28908 15156 28960 15162
rect 28908 15098 28960 15104
rect 28736 15026 28764 15098
rect 28724 15020 28776 15026
rect 28724 14962 28776 14968
rect 28724 14884 28776 14890
rect 28724 14826 28776 14832
rect 28736 14657 28764 14826
rect 28722 14648 28778 14657
rect 28722 14583 28778 14592
rect 28724 14476 28776 14482
rect 28724 14418 28776 14424
rect 28552 12406 28672 12434
rect 27804 12368 27856 12374
rect 27804 12310 27856 12316
rect 27620 12300 27672 12306
rect 27620 12242 27672 12248
rect 27632 11694 27660 12242
rect 27712 12096 27764 12102
rect 27712 12038 27764 12044
rect 27620 11688 27672 11694
rect 27620 11630 27672 11636
rect 27632 11393 27660 11630
rect 27724 11626 27752 12038
rect 27816 11694 27844 12310
rect 28080 12300 28132 12306
rect 28080 12242 28132 12248
rect 28092 12102 28120 12242
rect 28080 12096 28132 12102
rect 28080 12038 28132 12044
rect 28448 12096 28500 12102
rect 28448 12038 28500 12044
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 28356 11824 28408 11830
rect 28356 11766 28408 11772
rect 27804 11688 27856 11694
rect 27804 11630 27856 11636
rect 27712 11620 27764 11626
rect 27712 11562 27764 11568
rect 27618 11384 27674 11393
rect 27618 11319 27674 11328
rect 27712 11348 27764 11354
rect 27712 11290 27764 11296
rect 27620 9036 27672 9042
rect 27620 8978 27672 8984
rect 27528 6112 27580 6118
rect 27528 6054 27580 6060
rect 26148 4480 26200 4486
rect 26148 4422 26200 4428
rect 27160 4480 27212 4486
rect 27160 4422 27212 4428
rect 26160 4146 26188 4422
rect 27632 4214 27660 8978
rect 27724 7546 27752 11290
rect 27816 10810 27844 11630
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27804 10804 27856 10810
rect 27804 10746 27856 10752
rect 28080 10668 28132 10674
rect 28080 10610 28132 10616
rect 27804 10600 27856 10606
rect 27804 10542 27856 10548
rect 27816 10033 27844 10542
rect 27802 10024 27858 10033
rect 27802 9959 27858 9968
rect 28092 9926 28120 10610
rect 27804 9920 27856 9926
rect 27804 9862 27856 9868
rect 28080 9920 28132 9926
rect 28080 9862 28132 9868
rect 27816 8090 27844 9862
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 27988 8288 28040 8294
rect 27988 8230 28040 8236
rect 27804 8084 27856 8090
rect 27804 8026 27856 8032
rect 28000 7886 28028 8230
rect 28368 8090 28396 11766
rect 28460 10198 28488 12038
rect 28552 10606 28580 12406
rect 28632 11688 28684 11694
rect 28630 11656 28632 11665
rect 28684 11656 28686 11665
rect 28630 11591 28686 11600
rect 28632 11144 28684 11150
rect 28632 11086 28684 11092
rect 28540 10600 28592 10606
rect 28540 10542 28592 10548
rect 28448 10192 28500 10198
rect 28448 10134 28500 10140
rect 28448 9648 28500 9654
rect 28448 9590 28500 9596
rect 28460 8974 28488 9590
rect 28552 9110 28580 10542
rect 28644 9994 28672 11086
rect 28736 10810 28764 14418
rect 28828 13190 28856 15098
rect 28920 15065 28948 15098
rect 29288 15094 29316 15982
rect 29276 15088 29328 15094
rect 28906 15056 28962 15065
rect 28906 14991 28962 15000
rect 29090 15056 29146 15065
rect 29276 15030 29328 15036
rect 29090 14991 29092 15000
rect 29144 14991 29146 15000
rect 29092 14962 29144 14968
rect 29182 14920 29238 14929
rect 29380 14906 29408 18566
rect 29472 17746 29500 18566
rect 29460 17740 29512 17746
rect 29460 17682 29512 17688
rect 29182 14855 29238 14864
rect 29288 14878 29408 14906
rect 29092 14816 29144 14822
rect 29092 14758 29144 14764
rect 28908 14272 28960 14278
rect 29104 14249 29132 14758
rect 28908 14214 28960 14220
rect 29090 14240 29146 14249
rect 28920 13705 28948 14214
rect 29090 14175 29146 14184
rect 28906 13696 28962 13705
rect 28906 13631 28962 13640
rect 28908 13456 28960 13462
rect 28908 13398 28960 13404
rect 28816 13184 28868 13190
rect 28816 13126 28868 13132
rect 28816 12300 28868 12306
rect 28816 12242 28868 12248
rect 28724 10804 28776 10810
rect 28724 10746 28776 10752
rect 28632 9988 28684 9994
rect 28632 9930 28684 9936
rect 28828 9874 28856 12242
rect 28920 10266 28948 13398
rect 29000 13252 29052 13258
rect 29000 13194 29052 13200
rect 29012 12442 29040 13194
rect 29000 12436 29052 12442
rect 29000 12378 29052 12384
rect 28998 12336 29054 12345
rect 28998 12271 29054 12280
rect 29012 11098 29040 12271
rect 29092 12164 29144 12170
rect 29092 12106 29144 12112
rect 29104 11830 29132 12106
rect 29092 11824 29144 11830
rect 29092 11766 29144 11772
rect 29104 11218 29132 11766
rect 29092 11212 29144 11218
rect 29092 11154 29144 11160
rect 29012 11070 29132 11098
rect 29000 11008 29052 11014
rect 29000 10950 29052 10956
rect 28908 10260 28960 10266
rect 28908 10202 28960 10208
rect 28644 9846 28856 9874
rect 28540 9104 28592 9110
rect 28540 9046 28592 9052
rect 28448 8968 28500 8974
rect 28448 8910 28500 8916
rect 28460 8430 28488 8910
rect 28448 8424 28500 8430
rect 28448 8366 28500 8372
rect 28356 8084 28408 8090
rect 28356 8026 28408 8032
rect 27988 7880 28040 7886
rect 27988 7822 28040 7828
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27712 7540 27764 7546
rect 27712 7482 27764 7488
rect 28356 7404 28408 7410
rect 28356 7346 28408 7352
rect 28368 6866 28396 7346
rect 28356 6860 28408 6866
rect 28356 6802 28408 6808
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 27620 4208 27672 4214
rect 27620 4150 27672 4156
rect 26148 4140 26200 4146
rect 26148 4082 26200 4088
rect 27620 4072 27672 4078
rect 27620 4014 27672 4020
rect 27632 3738 27660 4014
rect 27620 3732 27672 3738
rect 27620 3674 27672 3680
rect 27528 3664 27580 3670
rect 27528 3606 27580 3612
rect 26332 3392 26384 3398
rect 26332 3334 26384 3340
rect 26056 2984 26108 2990
rect 26056 2926 26108 2932
rect 24952 2916 25004 2922
rect 24952 2858 25004 2864
rect 24504 2746 24624 2774
rect 24504 2650 24532 2746
rect 24492 2644 24544 2650
rect 24492 2586 24544 2592
rect 24964 2582 24992 2858
rect 26344 2650 26372 3334
rect 27540 3058 27568 3606
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 28460 3058 28488 8366
rect 28552 6798 28580 9046
rect 28540 6792 28592 6798
rect 28540 6734 28592 6740
rect 28644 4622 28672 9846
rect 28724 9376 28776 9382
rect 28724 9318 28776 9324
rect 28816 9376 28868 9382
rect 28816 9318 28868 9324
rect 28736 9042 28764 9318
rect 28828 9110 28856 9318
rect 28816 9104 28868 9110
rect 28816 9046 28868 9052
rect 28920 9042 28948 10202
rect 28724 9036 28776 9042
rect 28724 8978 28776 8984
rect 28908 9036 28960 9042
rect 28908 8978 28960 8984
rect 28920 6322 28948 8978
rect 29012 8634 29040 10950
rect 29000 8628 29052 8634
rect 29000 8570 29052 8576
rect 28908 6316 28960 6322
rect 28908 6258 28960 6264
rect 29104 6254 29132 11070
rect 29196 10674 29224 14855
rect 29288 13274 29316 14878
rect 29368 14816 29420 14822
rect 29366 14784 29368 14793
rect 29420 14784 29422 14793
rect 29366 14719 29422 14728
rect 29368 14408 29420 14414
rect 29368 14350 29420 14356
rect 29380 13938 29408 14350
rect 29368 13932 29420 13938
rect 29368 13874 29420 13880
rect 29380 13394 29408 13874
rect 29368 13388 29420 13394
rect 29368 13330 29420 13336
rect 29288 13246 29408 13274
rect 29472 13258 29500 17682
rect 29564 17626 29592 20742
rect 29644 20460 29696 20466
rect 29644 20402 29696 20408
rect 29656 18630 29684 20402
rect 29748 20058 29776 21490
rect 29840 20942 29868 22034
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 29932 20346 29960 22063
rect 30012 22024 30064 22030
rect 30012 21966 30064 21972
rect 30024 21486 30052 21966
rect 30012 21480 30064 21486
rect 30012 21422 30064 21428
rect 30116 20602 30144 23598
rect 30194 23352 30250 23361
rect 30194 23287 30250 23296
rect 30208 23050 30236 23287
rect 30196 23044 30248 23050
rect 30196 22986 30248 22992
rect 30196 22772 30248 22778
rect 30196 22714 30248 22720
rect 30208 21146 30236 22714
rect 30300 22030 30328 24006
rect 30392 23730 30420 24006
rect 30380 23724 30432 23730
rect 30380 23666 30432 23672
rect 30380 23520 30432 23526
rect 30380 23462 30432 23468
rect 30392 22094 30420 23462
rect 30484 22778 30512 24074
rect 30472 22772 30524 22778
rect 30472 22714 30524 22720
rect 30472 22094 30524 22098
rect 30392 22092 30524 22094
rect 30392 22066 30472 22092
rect 30472 22034 30524 22040
rect 30288 22024 30340 22030
rect 30288 21966 30340 21972
rect 30286 21720 30342 21729
rect 30286 21655 30342 21664
rect 30196 21140 30248 21146
rect 30196 21082 30248 21088
rect 30196 21004 30248 21010
rect 30196 20946 30248 20952
rect 30012 20596 30064 20602
rect 30012 20538 30064 20544
rect 30104 20596 30156 20602
rect 30104 20538 30156 20544
rect 29840 20318 29960 20346
rect 29736 20052 29788 20058
rect 29736 19994 29788 20000
rect 29840 19802 29868 20318
rect 29920 20256 29972 20262
rect 29920 20198 29972 20204
rect 29748 19774 29868 19802
rect 29748 18766 29776 19774
rect 29828 19712 29880 19718
rect 29828 19654 29880 19660
rect 29840 19009 29868 19654
rect 29826 19000 29882 19009
rect 29826 18935 29882 18944
rect 29826 18864 29882 18873
rect 29826 18799 29882 18808
rect 29736 18760 29788 18766
rect 29736 18702 29788 18708
rect 29840 18698 29868 18799
rect 29828 18692 29880 18698
rect 29828 18634 29880 18640
rect 29644 18624 29696 18630
rect 29644 18566 29696 18572
rect 29564 17598 29868 17626
rect 29736 17536 29788 17542
rect 29736 17478 29788 17484
rect 29552 17060 29604 17066
rect 29552 17002 29604 17008
rect 29564 16794 29592 17002
rect 29644 16992 29696 16998
rect 29644 16934 29696 16940
rect 29656 16794 29684 16934
rect 29552 16788 29604 16794
rect 29552 16730 29604 16736
rect 29644 16788 29696 16794
rect 29644 16730 29696 16736
rect 29552 16584 29604 16590
rect 29552 16526 29604 16532
rect 29564 14550 29592 16526
rect 29644 16108 29696 16114
rect 29644 16050 29696 16056
rect 29656 15638 29684 16050
rect 29644 15632 29696 15638
rect 29644 15574 29696 15580
rect 29748 15502 29776 17478
rect 29840 16726 29868 17598
rect 29828 16720 29880 16726
rect 29828 16662 29880 16668
rect 29932 15570 29960 20198
rect 30024 19242 30052 20538
rect 30116 20505 30144 20538
rect 30102 20496 30158 20505
rect 30102 20431 30158 20440
rect 30104 20256 30156 20262
rect 30104 20198 30156 20204
rect 30012 19236 30064 19242
rect 30012 19178 30064 19184
rect 30116 19122 30144 20198
rect 30208 19922 30236 20946
rect 30300 20806 30328 21655
rect 30380 21616 30432 21622
rect 30380 21558 30432 21564
rect 30392 21486 30420 21558
rect 30380 21480 30432 21486
rect 30380 21422 30432 21428
rect 30380 21344 30432 21350
rect 30380 21286 30432 21292
rect 30288 20800 30340 20806
rect 30288 20742 30340 20748
rect 30196 19916 30248 19922
rect 30196 19858 30248 19864
rect 30024 19094 30144 19122
rect 30024 17134 30052 19094
rect 30392 18970 30420 21286
rect 30576 20482 30604 25298
rect 30654 23896 30710 23905
rect 30654 23831 30656 23840
rect 30708 23831 30710 23840
rect 30656 23802 30708 23808
rect 30656 22636 30708 22642
rect 30656 22578 30708 22584
rect 30668 21690 30696 22578
rect 30656 21684 30708 21690
rect 30656 21626 30708 21632
rect 30656 21480 30708 21486
rect 30656 21422 30708 21428
rect 30484 20454 30604 20482
rect 30484 19825 30512 20454
rect 30564 20324 30616 20330
rect 30564 20266 30616 20272
rect 30470 19816 30526 19825
rect 30470 19751 30526 19760
rect 30576 19553 30604 20266
rect 30668 19825 30696 21422
rect 30654 19816 30710 19825
rect 30654 19751 30710 19760
rect 30562 19544 30618 19553
rect 30472 19508 30524 19514
rect 30562 19479 30618 19488
rect 30472 19450 30524 19456
rect 30104 18964 30156 18970
rect 30104 18906 30156 18912
rect 30380 18964 30432 18970
rect 30380 18906 30432 18912
rect 30116 18714 30144 18906
rect 30116 18686 30328 18714
rect 30196 17876 30248 17882
rect 30196 17818 30248 17824
rect 30208 17542 30236 17818
rect 30104 17536 30156 17542
rect 30104 17478 30156 17484
rect 30196 17536 30248 17542
rect 30196 17478 30248 17484
rect 30116 17338 30144 17478
rect 30104 17332 30156 17338
rect 30104 17274 30156 17280
rect 30012 17128 30064 17134
rect 30012 17070 30064 17076
rect 30012 16992 30064 16998
rect 30012 16934 30064 16940
rect 30024 16794 30052 16934
rect 30012 16788 30064 16794
rect 30012 16730 30064 16736
rect 30196 16788 30248 16794
rect 30196 16730 30248 16736
rect 30010 16688 30066 16697
rect 30010 16623 30012 16632
rect 30064 16623 30066 16632
rect 30104 16652 30156 16658
rect 30012 16594 30064 16600
rect 30104 16594 30156 16600
rect 29920 15564 29972 15570
rect 29920 15506 29972 15512
rect 29736 15496 29788 15502
rect 29736 15438 29788 15444
rect 29828 15156 29880 15162
rect 29828 15098 29880 15104
rect 29736 15088 29788 15094
rect 29736 15030 29788 15036
rect 29642 14784 29698 14793
rect 29642 14719 29698 14728
rect 29552 14544 29604 14550
rect 29552 14486 29604 14492
rect 29656 14482 29684 14719
rect 29644 14476 29696 14482
rect 29644 14418 29696 14424
rect 29552 14340 29604 14346
rect 29552 14282 29604 14288
rect 29564 13462 29592 14282
rect 29656 13462 29684 14418
rect 29748 13870 29776 15030
rect 29840 14657 29868 15098
rect 29826 14648 29882 14657
rect 29826 14583 29882 14592
rect 30116 14482 30144 16594
rect 30208 16046 30236 16730
rect 30196 16040 30248 16046
rect 30196 15982 30248 15988
rect 30300 15910 30328 18686
rect 30484 18465 30512 19450
rect 30564 19168 30616 19174
rect 30760 19156 30788 25735
rect 30932 24812 30984 24818
rect 30932 24754 30984 24760
rect 30840 24608 30892 24614
rect 30840 24550 30892 24556
rect 30852 23526 30880 24550
rect 30944 23662 30972 24754
rect 30932 23656 30984 23662
rect 30932 23598 30984 23604
rect 30840 23520 30892 23526
rect 30840 23462 30892 23468
rect 30932 23316 30984 23322
rect 30932 23258 30984 23264
rect 30840 22976 30892 22982
rect 30840 22918 30892 22924
rect 30852 20602 30880 22918
rect 30944 22574 30972 23258
rect 30932 22568 30984 22574
rect 30932 22510 30984 22516
rect 30932 21548 30984 21554
rect 30932 21490 30984 21496
rect 30944 21457 30972 21490
rect 30930 21448 30986 21457
rect 30930 21383 30986 21392
rect 30932 20868 30984 20874
rect 30932 20810 30984 20816
rect 30840 20596 30892 20602
rect 30840 20538 30892 20544
rect 30616 19128 30788 19156
rect 30564 19110 30616 19116
rect 30564 18896 30616 18902
rect 30564 18838 30616 18844
rect 30470 18456 30526 18465
rect 30470 18391 30526 18400
rect 30576 18290 30604 18838
rect 30564 18284 30616 18290
rect 30564 18226 30616 18232
rect 30380 18148 30432 18154
rect 30380 18090 30432 18096
rect 30392 17066 30420 18090
rect 30760 18086 30788 19128
rect 30840 19168 30892 19174
rect 30840 19110 30892 19116
rect 30852 18426 30880 19110
rect 30840 18420 30892 18426
rect 30840 18362 30892 18368
rect 30944 18290 30972 20810
rect 30840 18284 30892 18290
rect 30840 18226 30892 18232
rect 30932 18284 30984 18290
rect 30932 18226 30984 18232
rect 30564 18080 30616 18086
rect 30564 18022 30616 18028
rect 30748 18080 30800 18086
rect 30748 18022 30800 18028
rect 30472 17264 30524 17270
rect 30472 17206 30524 17212
rect 30380 17060 30432 17066
rect 30380 17002 30432 17008
rect 30380 15972 30432 15978
rect 30380 15914 30432 15920
rect 30288 15904 30340 15910
rect 30288 15846 30340 15852
rect 30196 15632 30248 15638
rect 30196 15574 30248 15580
rect 30104 14476 30156 14482
rect 29932 14436 30104 14464
rect 29736 13864 29788 13870
rect 29736 13806 29788 13812
rect 29826 13696 29882 13705
rect 29826 13631 29882 13640
rect 29552 13456 29604 13462
rect 29552 13398 29604 13404
rect 29644 13456 29696 13462
rect 29644 13398 29696 13404
rect 29276 12980 29328 12986
rect 29276 12922 29328 12928
rect 29288 12170 29316 12922
rect 29380 12481 29408 13246
rect 29460 13252 29512 13258
rect 29460 13194 29512 13200
rect 29366 12472 29422 12481
rect 29366 12407 29422 12416
rect 29564 12434 29592 13398
rect 29840 13190 29868 13631
rect 29828 13184 29880 13190
rect 29828 13126 29880 13132
rect 29564 12406 29684 12434
rect 29460 12300 29512 12306
rect 29460 12242 29512 12248
rect 29276 12164 29328 12170
rect 29276 12106 29328 12112
rect 29368 12164 29420 12170
rect 29368 12106 29420 12112
rect 29380 11898 29408 12106
rect 29368 11892 29420 11898
rect 29368 11834 29420 11840
rect 29274 11384 29330 11393
rect 29274 11319 29330 11328
rect 29288 11218 29316 11319
rect 29276 11212 29328 11218
rect 29276 11154 29328 11160
rect 29184 10668 29236 10674
rect 29184 10610 29236 10616
rect 29184 10124 29236 10130
rect 29184 10066 29236 10072
rect 29196 9625 29224 10066
rect 29276 9988 29328 9994
rect 29276 9930 29328 9936
rect 29182 9616 29238 9625
rect 29288 9586 29316 9930
rect 29182 9551 29238 9560
rect 29276 9580 29328 9586
rect 29276 9522 29328 9528
rect 29288 9450 29316 9522
rect 29276 9444 29328 9450
rect 29276 9386 29328 9392
rect 29472 7886 29500 12242
rect 29656 12238 29684 12406
rect 29840 12345 29868 13126
rect 29932 12646 29960 14436
rect 30104 14418 30156 14424
rect 30010 14376 30066 14385
rect 30010 14311 30012 14320
rect 30064 14311 30066 14320
rect 30012 14282 30064 14288
rect 30208 13954 30236 15574
rect 30288 15564 30340 15570
rect 30288 15506 30340 15512
rect 30024 13926 30236 13954
rect 29920 12640 29972 12646
rect 29920 12582 29972 12588
rect 29826 12336 29882 12345
rect 29826 12271 29882 12280
rect 29552 12232 29604 12238
rect 29552 12174 29604 12180
rect 29644 12232 29696 12238
rect 29644 12174 29696 12180
rect 29564 11354 29592 12174
rect 29644 12096 29696 12102
rect 29644 12038 29696 12044
rect 29552 11348 29604 11354
rect 29552 11290 29604 11296
rect 29552 10464 29604 10470
rect 29552 10406 29604 10412
rect 29564 10130 29592 10406
rect 29552 10124 29604 10130
rect 29552 10066 29604 10072
rect 29368 7880 29420 7886
rect 29368 7822 29420 7828
rect 29460 7880 29512 7886
rect 29564 7857 29592 10066
rect 29656 9654 29684 12038
rect 29932 11762 29960 12582
rect 29920 11756 29972 11762
rect 29920 11698 29972 11704
rect 29920 11620 29972 11626
rect 29920 11562 29972 11568
rect 29736 11552 29788 11558
rect 29736 11494 29788 11500
rect 29748 11132 29776 11494
rect 29932 11286 29960 11562
rect 29920 11280 29972 11286
rect 29920 11222 29972 11228
rect 29828 11144 29880 11150
rect 29748 11104 29828 11132
rect 29748 10606 29776 11104
rect 29828 11086 29880 11092
rect 29736 10600 29788 10606
rect 29736 10542 29788 10548
rect 29644 9648 29696 9654
rect 29644 9590 29696 9596
rect 29748 8974 29776 10542
rect 29828 9444 29880 9450
rect 29828 9386 29880 9392
rect 29736 8968 29788 8974
rect 29736 8910 29788 8916
rect 29840 8498 29868 9386
rect 29828 8492 29880 8498
rect 29828 8434 29880 8440
rect 29460 7822 29512 7828
rect 29550 7848 29606 7857
rect 29380 7546 29408 7822
rect 29550 7783 29606 7792
rect 29368 7540 29420 7546
rect 29368 7482 29420 7488
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29288 6458 29316 6734
rect 29276 6452 29328 6458
rect 29276 6394 29328 6400
rect 29092 6248 29144 6254
rect 29092 6190 29144 6196
rect 29564 5846 29592 7783
rect 29552 5840 29604 5846
rect 29552 5782 29604 5788
rect 28632 4616 28684 4622
rect 28632 4558 28684 4564
rect 29092 3392 29144 3398
rect 29092 3334 29144 3340
rect 29104 3126 29132 3334
rect 29840 3126 29868 8434
rect 29932 7410 29960 11222
rect 30024 9722 30052 13926
rect 30196 13864 30248 13870
rect 30300 13818 30328 15506
rect 30392 15502 30420 15914
rect 30380 15496 30432 15502
rect 30380 15438 30432 15444
rect 30380 14952 30432 14958
rect 30380 14894 30432 14900
rect 30392 13841 30420 14894
rect 30248 13812 30328 13818
rect 30196 13806 30328 13812
rect 30208 13790 30328 13806
rect 30378 13832 30434 13841
rect 30104 13524 30156 13530
rect 30104 13466 30156 13472
rect 30012 9716 30064 9722
rect 30012 9658 30064 9664
rect 29920 7404 29972 7410
rect 29920 7346 29972 7352
rect 30116 3466 30144 13466
rect 30208 12306 30236 13790
rect 30378 13767 30434 13776
rect 30392 13462 30420 13767
rect 30484 13705 30512 17206
rect 30576 16114 30604 18022
rect 30656 17876 30708 17882
rect 30656 17818 30708 17824
rect 30668 16522 30696 17818
rect 30760 17202 30788 18022
rect 30748 17196 30800 17202
rect 30748 17138 30800 17144
rect 30748 17060 30800 17066
rect 30748 17002 30800 17008
rect 30656 16516 30708 16522
rect 30656 16458 30708 16464
rect 30656 16244 30708 16250
rect 30656 16186 30708 16192
rect 30564 16108 30616 16114
rect 30564 16050 30616 16056
rect 30564 15904 30616 15910
rect 30564 15846 30616 15852
rect 30576 15638 30604 15846
rect 30564 15632 30616 15638
rect 30564 15574 30616 15580
rect 30564 15496 30616 15502
rect 30564 15438 30616 15444
rect 30470 13696 30526 13705
rect 30470 13631 30526 13640
rect 30380 13456 30432 13462
rect 30380 13398 30432 13404
rect 30288 13184 30340 13190
rect 30288 13126 30340 13132
rect 30300 12442 30328 13126
rect 30472 12980 30524 12986
rect 30472 12922 30524 12928
rect 30484 12782 30512 12922
rect 30472 12776 30524 12782
rect 30472 12718 30524 12724
rect 30288 12436 30340 12442
rect 30288 12378 30340 12384
rect 30576 12374 30604 15438
rect 30668 15026 30696 16186
rect 30656 15020 30708 15026
rect 30656 14962 30708 14968
rect 30656 14816 30708 14822
rect 30656 14758 30708 14764
rect 30668 14482 30696 14758
rect 30656 14476 30708 14482
rect 30656 14418 30708 14424
rect 30760 14362 30788 17002
rect 30852 16250 30880 18226
rect 30932 17536 30984 17542
rect 30932 17478 30984 17484
rect 30840 16244 30892 16250
rect 30840 16186 30892 16192
rect 30840 15904 30892 15910
rect 30840 15846 30892 15852
rect 30852 15502 30880 15846
rect 30840 15496 30892 15502
rect 30840 15438 30892 15444
rect 30840 15360 30892 15366
rect 30840 15302 30892 15308
rect 30852 15201 30880 15302
rect 30838 15192 30894 15201
rect 30838 15127 30894 15136
rect 30840 15020 30892 15026
rect 30840 14962 30892 14968
rect 30668 14334 30788 14362
rect 30564 12368 30616 12374
rect 30564 12310 30616 12316
rect 30196 12300 30248 12306
rect 30196 12242 30248 12248
rect 30380 12232 30432 12238
rect 30576 12209 30604 12310
rect 30380 12174 30432 12180
rect 30562 12200 30618 12209
rect 30196 12164 30248 12170
rect 30248 12124 30328 12152
rect 30196 12106 30248 12112
rect 30194 12064 30250 12073
rect 30194 11999 30250 12008
rect 30208 11898 30236 11999
rect 30196 11892 30248 11898
rect 30196 11834 30248 11840
rect 30196 11688 30248 11694
rect 30300 11676 30328 12124
rect 30248 11648 30328 11676
rect 30196 11630 30248 11636
rect 30208 7449 30236 11630
rect 30392 11506 30420 12174
rect 30562 12135 30618 12144
rect 30300 11478 30420 11506
rect 30300 11150 30328 11478
rect 30668 11370 30696 14334
rect 30748 14272 30800 14278
rect 30748 14214 30800 14220
rect 30760 13938 30788 14214
rect 30748 13932 30800 13938
rect 30748 13874 30800 13880
rect 30852 12764 30880 14962
rect 30760 12736 30880 12764
rect 30760 11898 30788 12736
rect 30840 12640 30892 12646
rect 30840 12582 30892 12588
rect 30748 11892 30800 11898
rect 30748 11834 30800 11840
rect 30392 11342 30696 11370
rect 30288 11144 30340 11150
rect 30288 11086 30340 11092
rect 30392 10130 30420 11342
rect 30470 11112 30526 11121
rect 30470 11047 30526 11056
rect 30748 11076 30800 11082
rect 30380 10124 30432 10130
rect 30380 10066 30432 10072
rect 30392 9897 30420 10066
rect 30378 9888 30434 9897
rect 30378 9823 30434 9832
rect 30484 9586 30512 11047
rect 30748 11018 30800 11024
rect 30656 10600 30708 10606
rect 30656 10542 30708 10548
rect 30562 10432 30618 10441
rect 30562 10367 30618 10376
rect 30576 9761 30604 10367
rect 30668 9926 30696 10542
rect 30656 9920 30708 9926
rect 30656 9862 30708 9868
rect 30562 9752 30618 9761
rect 30562 9687 30618 9696
rect 30472 9580 30524 9586
rect 30472 9522 30524 9528
rect 30564 9512 30616 9518
rect 30564 9454 30616 9460
rect 30288 8424 30340 8430
rect 30288 8366 30340 8372
rect 30194 7440 30250 7449
rect 30194 7375 30250 7384
rect 30300 6662 30328 8366
rect 30380 6792 30432 6798
rect 30380 6734 30432 6740
rect 30288 6656 30340 6662
rect 30288 6598 30340 6604
rect 30392 5914 30420 6734
rect 30472 6656 30524 6662
rect 30472 6598 30524 6604
rect 30484 6322 30512 6598
rect 30576 6458 30604 9454
rect 30760 9194 30788 11018
rect 30852 10656 30880 12582
rect 30944 11558 30972 17478
rect 31036 13938 31064 26302
rect 31206 26200 31262 27000
rect 31850 26330 31906 27000
rect 31850 26302 31984 26330
rect 31850 26200 31906 26302
rect 31116 24064 31168 24070
rect 31116 24006 31168 24012
rect 31128 20466 31156 24006
rect 31220 23497 31248 26200
rect 31760 25084 31812 25090
rect 31760 25026 31812 25032
rect 31300 24608 31352 24614
rect 31300 24550 31352 24556
rect 31206 23488 31262 23497
rect 31206 23423 31262 23432
rect 31312 23338 31340 24550
rect 31392 23860 31444 23866
rect 31392 23802 31444 23808
rect 31220 23310 31340 23338
rect 31220 22094 31248 23310
rect 31220 22066 31340 22094
rect 31208 20868 31260 20874
rect 31208 20810 31260 20816
rect 31116 20460 31168 20466
rect 31116 20402 31168 20408
rect 31116 18692 31168 18698
rect 31116 18634 31168 18640
rect 31024 13932 31076 13938
rect 31024 13874 31076 13880
rect 31024 13252 31076 13258
rect 31024 13194 31076 13200
rect 31036 13161 31064 13194
rect 31022 13152 31078 13161
rect 31022 13087 31078 13096
rect 31128 13002 31156 18634
rect 31220 17270 31248 20810
rect 31312 19922 31340 22066
rect 31404 22080 31432 23802
rect 31772 23798 31800 25026
rect 31852 24404 31904 24410
rect 31852 24346 31904 24352
rect 31760 23792 31812 23798
rect 31760 23734 31812 23740
rect 31576 23724 31628 23730
rect 31576 23666 31628 23672
rect 31588 23497 31616 23666
rect 31574 23488 31630 23497
rect 31574 23423 31630 23432
rect 31482 23352 31538 23361
rect 31482 23287 31538 23296
rect 31496 22234 31524 23287
rect 31760 22976 31812 22982
rect 31760 22918 31812 22924
rect 31574 22672 31630 22681
rect 31574 22607 31576 22616
rect 31628 22607 31630 22616
rect 31576 22578 31628 22584
rect 31668 22568 31720 22574
rect 31772 22556 31800 22918
rect 31864 22642 31892 24346
rect 31852 22636 31904 22642
rect 31852 22578 31904 22584
rect 31720 22528 31800 22556
rect 31668 22510 31720 22516
rect 31576 22500 31628 22506
rect 31576 22442 31628 22448
rect 31484 22228 31536 22234
rect 31484 22170 31536 22176
rect 31404 22052 31524 22080
rect 31392 21956 31444 21962
rect 31392 21898 31444 21904
rect 31404 21865 31432 21898
rect 31390 21856 31446 21865
rect 31390 21791 31446 21800
rect 31496 21486 31524 22052
rect 31588 21690 31616 22442
rect 31666 22400 31722 22409
rect 31666 22335 31722 22344
rect 31576 21684 31628 21690
rect 31576 21626 31628 21632
rect 31576 21548 31628 21554
rect 31576 21490 31628 21496
rect 31392 21480 31444 21486
rect 31392 21422 31444 21428
rect 31484 21480 31536 21486
rect 31484 21422 31536 21428
rect 31404 21078 31432 21422
rect 31392 21072 31444 21078
rect 31392 21014 31444 21020
rect 31392 20800 31444 20806
rect 31390 20768 31392 20777
rect 31444 20768 31446 20777
rect 31390 20703 31446 20712
rect 31300 19916 31352 19922
rect 31300 19858 31352 19864
rect 31496 19446 31524 21422
rect 31588 20874 31616 21490
rect 31576 20868 31628 20874
rect 31576 20810 31628 20816
rect 31680 20806 31708 22335
rect 31772 21962 31800 22528
rect 31956 22386 31984 26302
rect 32494 26200 32550 27000
rect 33138 26330 33194 27000
rect 33138 26302 33364 26330
rect 33138 26200 33194 26302
rect 32034 25392 32090 25401
rect 32034 25327 32090 25336
rect 32048 23361 32076 25327
rect 32220 25084 32272 25090
rect 32220 25026 32272 25032
rect 32128 24404 32180 24410
rect 32128 24346 32180 24352
rect 32034 23352 32090 23361
rect 32034 23287 32090 23296
rect 32140 22710 32168 24346
rect 32128 22704 32180 22710
rect 32128 22646 32180 22652
rect 32126 22536 32182 22545
rect 32126 22471 32182 22480
rect 31864 22358 31984 22386
rect 31864 22137 31892 22358
rect 31850 22128 31906 22137
rect 31850 22063 31906 22072
rect 31760 21956 31812 21962
rect 31760 21898 31812 21904
rect 31760 21684 31812 21690
rect 31760 21626 31812 21632
rect 31852 21684 31904 21690
rect 31852 21626 31904 21632
rect 31668 20800 31720 20806
rect 31668 20742 31720 20748
rect 31576 19780 31628 19786
rect 31576 19722 31628 19728
rect 31484 19440 31536 19446
rect 31484 19382 31536 19388
rect 31300 19372 31352 19378
rect 31300 19314 31352 19320
rect 31392 19372 31444 19378
rect 31392 19314 31444 19320
rect 31208 17264 31260 17270
rect 31208 17206 31260 17212
rect 31208 16992 31260 16998
rect 31208 16934 31260 16940
rect 31036 12974 31156 13002
rect 30932 11552 30984 11558
rect 30932 11494 30984 11500
rect 30852 10628 30972 10656
rect 30944 10266 30972 10628
rect 30932 10260 30984 10266
rect 30932 10202 30984 10208
rect 30840 9920 30892 9926
rect 30840 9862 30892 9868
rect 30668 9166 30788 9194
rect 30668 6730 30696 9166
rect 30748 9036 30800 9042
rect 30748 8978 30800 8984
rect 30656 6724 30708 6730
rect 30656 6666 30708 6672
rect 30564 6452 30616 6458
rect 30564 6394 30616 6400
rect 30472 6316 30524 6322
rect 30472 6258 30524 6264
rect 30760 5914 30788 8978
rect 30852 6458 30880 9862
rect 30944 7886 30972 10202
rect 31036 8809 31064 12974
rect 31116 11552 31168 11558
rect 31116 11494 31168 11500
rect 31128 10713 31156 11494
rect 31114 10704 31170 10713
rect 31114 10639 31170 10648
rect 31116 9920 31168 9926
rect 31116 9862 31168 9868
rect 31220 9874 31248 16934
rect 31312 14006 31340 19314
rect 31404 19281 31432 19314
rect 31390 19272 31446 19281
rect 31390 19207 31446 19216
rect 31588 18766 31616 19722
rect 31666 19136 31722 19145
rect 31666 19071 31722 19080
rect 31576 18760 31628 18766
rect 31576 18702 31628 18708
rect 31588 18426 31616 18702
rect 31576 18420 31628 18426
rect 31576 18362 31628 18368
rect 31392 18216 31444 18222
rect 31392 18158 31444 18164
rect 31404 14958 31432 18158
rect 31680 18086 31708 19071
rect 31772 19009 31800 21626
rect 31758 19000 31814 19009
rect 31758 18935 31814 18944
rect 31864 18873 31892 21626
rect 32036 21616 32088 21622
rect 32036 21558 32088 21564
rect 32048 21146 32076 21558
rect 32036 21140 32088 21146
rect 32036 21082 32088 21088
rect 32140 20806 32168 22471
rect 32232 21876 32260 25026
rect 32312 24064 32364 24070
rect 32312 24006 32364 24012
rect 32324 23769 32352 24006
rect 32310 23760 32366 23769
rect 32310 23695 32366 23704
rect 32404 23724 32456 23730
rect 32404 23666 32456 23672
rect 32312 22500 32364 22506
rect 32312 22442 32364 22448
rect 32324 22273 32352 22442
rect 32310 22264 32366 22273
rect 32310 22199 32366 22208
rect 32310 22128 32366 22137
rect 32416 22098 32444 23666
rect 32508 23497 32536 26200
rect 32770 25528 32826 25537
rect 32770 25463 32826 25472
rect 32678 24848 32734 24857
rect 32678 24783 32734 24792
rect 32692 23798 32720 24783
rect 32680 23792 32732 23798
rect 32680 23734 32732 23740
rect 32784 23610 32812 25463
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 32862 24304 32918 24313
rect 32862 24239 32918 24248
rect 32692 23582 32812 23610
rect 32494 23488 32550 23497
rect 32494 23423 32550 23432
rect 32692 23050 32720 23582
rect 32772 23520 32824 23526
rect 32772 23462 32824 23468
rect 32680 23044 32732 23050
rect 32680 22986 32732 22992
rect 32784 22982 32812 23462
rect 32772 22976 32824 22982
rect 32772 22918 32824 22924
rect 32588 22772 32640 22778
rect 32588 22714 32640 22720
rect 32310 22063 32366 22072
rect 32404 22092 32456 22098
rect 32324 21978 32352 22063
rect 32404 22034 32456 22040
rect 32324 21950 32444 21978
rect 32232 21848 32352 21876
rect 32128 20800 32180 20806
rect 32128 20742 32180 20748
rect 32324 20534 32352 21848
rect 32416 21536 32444 21950
rect 32496 21956 32548 21962
rect 32496 21898 32548 21904
rect 32508 21690 32536 21898
rect 32496 21684 32548 21690
rect 32496 21626 32548 21632
rect 32416 21508 32536 21536
rect 32404 21412 32456 21418
rect 32404 21354 32456 21360
rect 32312 20528 32364 20534
rect 32312 20470 32364 20476
rect 32312 20392 32364 20398
rect 32312 20334 32364 20340
rect 32036 19780 32088 19786
rect 32036 19722 32088 19728
rect 31942 19408 31998 19417
rect 31942 19343 31998 19352
rect 31850 18864 31906 18873
rect 31850 18799 31906 18808
rect 31760 18420 31812 18426
rect 31760 18362 31812 18368
rect 31668 18080 31720 18086
rect 31668 18022 31720 18028
rect 31576 17196 31628 17202
rect 31576 17138 31628 17144
rect 31484 17060 31536 17066
rect 31484 17002 31536 17008
rect 31496 16697 31524 17002
rect 31482 16688 31538 16697
rect 31482 16623 31538 16632
rect 31496 16590 31524 16623
rect 31484 16584 31536 16590
rect 31484 16526 31536 16532
rect 31392 14952 31444 14958
rect 31392 14894 31444 14900
rect 31300 14000 31352 14006
rect 31300 13942 31352 13948
rect 31300 12912 31352 12918
rect 31300 12854 31352 12860
rect 31312 12782 31340 12854
rect 31300 12776 31352 12782
rect 31300 12718 31352 12724
rect 31404 10538 31432 14894
rect 31496 14346 31524 16526
rect 31588 16425 31616 17138
rect 31680 17134 31708 18022
rect 31668 17128 31720 17134
rect 31668 17070 31720 17076
rect 31574 16416 31630 16425
rect 31574 16351 31630 16360
rect 31576 16244 31628 16250
rect 31576 16186 31628 16192
rect 31588 15484 31616 16186
rect 31680 15609 31708 17070
rect 31666 15600 31722 15609
rect 31666 15535 31722 15544
rect 31588 15456 31708 15484
rect 31680 15201 31708 15456
rect 31666 15192 31722 15201
rect 31666 15127 31722 15136
rect 31574 15056 31630 15065
rect 31574 14991 31630 15000
rect 31588 14822 31616 14991
rect 31576 14816 31628 14822
rect 31576 14758 31628 14764
rect 31576 14544 31628 14550
rect 31576 14486 31628 14492
rect 31484 14340 31536 14346
rect 31484 14282 31536 14288
rect 31496 13258 31524 14282
rect 31588 14249 31616 14486
rect 31574 14240 31630 14249
rect 31574 14175 31630 14184
rect 31772 14074 31800 18362
rect 31956 18306 31984 19343
rect 31864 18278 31984 18306
rect 31864 17202 31892 18278
rect 32048 17338 32076 19722
rect 32128 19304 32180 19310
rect 32128 19246 32180 19252
rect 32140 18766 32168 19246
rect 32220 19168 32272 19174
rect 32220 19110 32272 19116
rect 32232 18970 32260 19110
rect 32220 18964 32272 18970
rect 32220 18906 32272 18912
rect 32324 18834 32352 20334
rect 32416 19922 32444 21354
rect 32508 20890 32536 21508
rect 32600 21010 32628 22714
rect 32680 22636 32732 22642
rect 32680 22578 32732 22584
rect 32588 21004 32640 21010
rect 32588 20946 32640 20952
rect 32508 20862 32628 20890
rect 32496 20800 32548 20806
rect 32496 20742 32548 20748
rect 32404 19916 32456 19922
rect 32404 19858 32456 19864
rect 32508 19514 32536 20742
rect 32496 19508 32548 19514
rect 32496 19450 32548 19456
rect 32600 18902 32628 20862
rect 32692 20641 32720 22578
rect 32876 22574 32904 24239
rect 33140 24064 33192 24070
rect 33140 24006 33192 24012
rect 33152 23662 33180 24006
rect 33232 23724 33284 23730
rect 33232 23666 33284 23672
rect 33140 23656 33192 23662
rect 33046 23624 33102 23633
rect 33140 23598 33192 23604
rect 33046 23559 33048 23568
rect 33100 23559 33102 23568
rect 33048 23530 33100 23536
rect 33244 23526 33272 23666
rect 33232 23520 33284 23526
rect 33232 23462 33284 23468
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 33336 23225 33364 26302
rect 33508 26240 33560 26246
rect 33782 26200 33838 27000
rect 34426 26330 34482 27000
rect 33888 26302 34482 26330
rect 33508 26182 33560 26188
rect 33520 24954 33548 26182
rect 33508 24948 33560 24954
rect 33508 24890 33560 24896
rect 33520 24206 33548 24890
rect 33508 24200 33560 24206
rect 33508 24142 33560 24148
rect 33796 23497 33824 26200
rect 33782 23488 33838 23497
rect 33782 23423 33838 23432
rect 33322 23216 33378 23225
rect 33322 23151 33378 23160
rect 33416 23180 33468 23186
rect 33416 23122 33468 23128
rect 33324 22976 33376 22982
rect 33324 22918 33376 22924
rect 32772 22568 32824 22574
rect 32772 22510 32824 22516
rect 32864 22568 32916 22574
rect 32864 22510 32916 22516
rect 32784 22001 32812 22510
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 32864 22092 32916 22098
rect 32864 22034 32916 22040
rect 32770 21992 32826 22001
rect 32770 21927 32826 21936
rect 32876 21593 32904 22034
rect 32956 21616 33008 21622
rect 32862 21584 32918 21593
rect 32784 21542 32862 21570
rect 32678 20632 32734 20641
rect 32678 20567 32734 20576
rect 32784 20058 32812 21542
rect 32956 21558 33008 21564
rect 32862 21519 32918 21528
rect 32968 21468 32996 21558
rect 32876 21440 32996 21468
rect 32772 20052 32824 20058
rect 32772 19994 32824 20000
rect 32678 19952 32734 19961
rect 32678 19887 32734 19896
rect 32588 18896 32640 18902
rect 32588 18838 32640 18844
rect 32312 18828 32364 18834
rect 32312 18770 32364 18776
rect 32128 18760 32180 18766
rect 32128 18702 32180 18708
rect 32220 18692 32272 18698
rect 32220 18634 32272 18640
rect 32232 18290 32260 18634
rect 32220 18284 32272 18290
rect 32220 18226 32272 18232
rect 32128 18216 32180 18222
rect 32128 18158 32180 18164
rect 31944 17332 31996 17338
rect 31944 17274 31996 17280
rect 32036 17332 32088 17338
rect 32036 17274 32088 17280
rect 31852 17196 31904 17202
rect 31852 17138 31904 17144
rect 31852 16992 31904 16998
rect 31852 16934 31904 16940
rect 31864 16250 31892 16934
rect 31956 16697 31984 17274
rect 32140 17218 32168 18158
rect 32232 17921 32260 18226
rect 32218 17912 32274 17921
rect 32218 17847 32274 17856
rect 32324 17746 32352 18770
rect 32404 18692 32456 18698
rect 32404 18634 32456 18640
rect 32312 17740 32364 17746
rect 32312 17682 32364 17688
rect 32048 17190 32168 17218
rect 32324 17202 32352 17682
rect 32312 17196 32364 17202
rect 31942 16688 31998 16697
rect 31942 16623 31998 16632
rect 31944 16584 31996 16590
rect 31944 16526 31996 16532
rect 31956 16250 31984 16526
rect 31852 16244 31904 16250
rect 31852 16186 31904 16192
rect 31944 16244 31996 16250
rect 31944 16186 31996 16192
rect 31944 15904 31996 15910
rect 31944 15846 31996 15852
rect 31956 15570 31984 15846
rect 31944 15564 31996 15570
rect 31944 15506 31996 15512
rect 31942 15328 31998 15337
rect 31942 15263 31998 15272
rect 31956 15178 31984 15263
rect 31864 15150 31984 15178
rect 31760 14068 31812 14074
rect 31760 14010 31812 14016
rect 31668 13864 31720 13870
rect 31668 13806 31720 13812
rect 31484 13252 31536 13258
rect 31484 13194 31536 13200
rect 31496 12170 31524 13194
rect 31484 12164 31536 12170
rect 31484 12106 31536 12112
rect 31680 10810 31708 13806
rect 31760 12912 31812 12918
rect 31760 12854 31812 12860
rect 31772 11082 31800 12854
rect 31864 11694 31892 15150
rect 32048 14940 32076 17190
rect 32312 17138 32364 17144
rect 32128 17128 32180 17134
rect 32128 17070 32180 17076
rect 32140 16980 32168 17070
rect 32140 16952 32352 16980
rect 32220 16244 32272 16250
rect 32220 16186 32272 16192
rect 32128 16040 32180 16046
rect 32128 15982 32180 15988
rect 31956 14912 32076 14940
rect 31852 11688 31904 11694
rect 31852 11630 31904 11636
rect 31956 11540 31984 14912
rect 31864 11512 31984 11540
rect 31760 11076 31812 11082
rect 31760 11018 31812 11024
rect 31668 10804 31720 10810
rect 31668 10746 31720 10752
rect 31772 10690 31800 11018
rect 31484 10668 31536 10674
rect 31588 10662 31800 10690
rect 31588 10656 31616 10662
rect 31536 10628 31616 10656
rect 31484 10610 31536 10616
rect 31392 10532 31444 10538
rect 31392 10474 31444 10480
rect 31392 10124 31444 10130
rect 31392 10066 31444 10072
rect 31300 9920 31352 9926
rect 31220 9868 31300 9874
rect 31220 9862 31352 9868
rect 31022 8800 31078 8809
rect 31022 8735 31078 8744
rect 31128 8022 31156 9862
rect 31220 9846 31340 9862
rect 31206 9752 31262 9761
rect 31404 9738 31432 10066
rect 31206 9687 31262 9696
rect 31312 9710 31432 9738
rect 31116 8016 31168 8022
rect 31116 7958 31168 7964
rect 30932 7880 30984 7886
rect 30932 7822 30984 7828
rect 30932 7744 30984 7750
rect 30932 7686 30984 7692
rect 30944 7410 30972 7686
rect 30932 7404 30984 7410
rect 30932 7346 30984 7352
rect 30840 6452 30892 6458
rect 30840 6394 30892 6400
rect 30380 5908 30432 5914
rect 30380 5850 30432 5856
rect 30748 5908 30800 5914
rect 30748 5850 30800 5856
rect 31220 5794 31248 9687
rect 31312 9110 31340 9710
rect 31392 9580 31444 9586
rect 31392 9522 31444 9528
rect 31300 9104 31352 9110
rect 31300 9046 31352 9052
rect 30760 5766 31248 5794
rect 30104 3460 30156 3466
rect 30104 3402 30156 3408
rect 29092 3120 29144 3126
rect 29092 3062 29144 3068
rect 29828 3120 29880 3126
rect 29828 3062 29880 3068
rect 27528 3052 27580 3058
rect 27528 2994 27580 3000
rect 28448 3052 28500 3058
rect 28448 2994 28500 3000
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 24952 2576 25004 2582
rect 24952 2518 25004 2524
rect 27540 2446 27568 2994
rect 30760 2582 30788 5766
rect 31312 5710 31340 9046
rect 31404 8650 31432 9522
rect 31496 8974 31524 10610
rect 31758 9752 31814 9761
rect 31758 9687 31814 9696
rect 31772 9518 31800 9687
rect 31760 9512 31812 9518
rect 31760 9454 31812 9460
rect 31484 8968 31536 8974
rect 31484 8910 31536 8916
rect 31404 8622 31524 8650
rect 31392 8492 31444 8498
rect 31392 8434 31444 8440
rect 31404 5778 31432 8434
rect 31392 5772 31444 5778
rect 31392 5714 31444 5720
rect 31300 5704 31352 5710
rect 31300 5646 31352 5652
rect 31496 5370 31524 8622
rect 31760 8424 31812 8430
rect 31760 8366 31812 8372
rect 31772 7954 31800 8366
rect 31760 7948 31812 7954
rect 31760 7890 31812 7896
rect 31576 7880 31628 7886
rect 31576 7822 31628 7828
rect 31588 7546 31616 7822
rect 31576 7540 31628 7546
rect 31576 7482 31628 7488
rect 31864 6934 31892 11512
rect 32140 11218 32168 15982
rect 32232 15162 32260 16186
rect 32324 15978 32352 16952
rect 32416 16250 32444 18634
rect 32692 18222 32720 19887
rect 32772 19712 32824 19718
rect 32772 19654 32824 19660
rect 32680 18216 32732 18222
rect 32680 18158 32732 18164
rect 32680 18080 32732 18086
rect 32680 18022 32732 18028
rect 32588 17808 32640 17814
rect 32508 17768 32588 17796
rect 32508 16946 32536 17768
rect 32588 17750 32640 17756
rect 32588 17672 32640 17678
rect 32588 17614 32640 17620
rect 32600 17066 32628 17614
rect 32692 17338 32720 18022
rect 32680 17332 32732 17338
rect 32680 17274 32732 17280
rect 32588 17060 32640 17066
rect 32588 17002 32640 17008
rect 32508 16918 32720 16946
rect 32404 16244 32456 16250
rect 32404 16186 32456 16192
rect 32404 16108 32456 16114
rect 32404 16050 32456 16056
rect 32312 15972 32364 15978
rect 32312 15914 32364 15920
rect 32416 15722 32444 16050
rect 32416 15694 32536 15722
rect 32312 15632 32364 15638
rect 32312 15574 32364 15580
rect 32220 15156 32272 15162
rect 32220 15098 32272 15104
rect 32220 14884 32272 14890
rect 32220 14826 32272 14832
rect 32232 14550 32260 14826
rect 32324 14550 32352 15574
rect 32508 15434 32536 15694
rect 32588 15564 32640 15570
rect 32588 15506 32640 15512
rect 32496 15428 32548 15434
rect 32496 15370 32548 15376
rect 32600 15314 32628 15506
rect 32416 15286 32628 15314
rect 32220 14544 32272 14550
rect 32220 14486 32272 14492
rect 32312 14544 32364 14550
rect 32312 14486 32364 14492
rect 32312 13320 32364 13326
rect 32312 13262 32364 13268
rect 32218 12880 32274 12889
rect 32324 12850 32352 13262
rect 32218 12815 32220 12824
rect 32272 12815 32274 12824
rect 32312 12844 32364 12850
rect 32220 12786 32272 12792
rect 32312 12786 32364 12792
rect 32324 12306 32352 12786
rect 32312 12300 32364 12306
rect 32312 12242 32364 12248
rect 32220 11280 32272 11286
rect 32220 11222 32272 11228
rect 32128 11212 32180 11218
rect 32128 11154 32180 11160
rect 31944 10532 31996 10538
rect 31944 10474 31996 10480
rect 31956 9042 31984 10474
rect 32036 10464 32088 10470
rect 32036 10406 32088 10412
rect 31944 9036 31996 9042
rect 31944 8978 31996 8984
rect 31852 6928 31904 6934
rect 31852 6870 31904 6876
rect 32048 6322 32076 10406
rect 32232 9674 32260 11222
rect 32140 9646 32260 9674
rect 32140 8430 32168 9646
rect 32324 9586 32352 12242
rect 32416 12102 32444 15286
rect 32496 15020 32548 15026
rect 32496 14962 32548 14968
rect 32404 12096 32456 12102
rect 32404 12038 32456 12044
rect 32416 10674 32444 12038
rect 32404 10668 32456 10674
rect 32404 10610 32456 10616
rect 32404 9988 32456 9994
rect 32404 9930 32456 9936
rect 32416 9722 32444 9930
rect 32404 9716 32456 9722
rect 32404 9658 32456 9664
rect 32312 9580 32364 9586
rect 32312 9522 32364 9528
rect 32220 8900 32272 8906
rect 32220 8842 32272 8848
rect 32128 8424 32180 8430
rect 32128 8366 32180 8372
rect 32232 6866 32260 8842
rect 32508 8634 32536 14962
rect 32692 14793 32720 16918
rect 32784 15502 32812 19654
rect 32876 18873 32904 21440
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 33336 21128 33364 22918
rect 33428 22642 33456 23122
rect 33692 22976 33744 22982
rect 33692 22918 33744 22924
rect 33416 22636 33468 22642
rect 33416 22578 33468 22584
rect 33600 22636 33652 22642
rect 33600 22578 33652 22584
rect 33416 21888 33468 21894
rect 33416 21830 33468 21836
rect 33508 21888 33560 21894
rect 33508 21830 33560 21836
rect 33428 21690 33456 21830
rect 33416 21684 33468 21690
rect 33416 21626 33468 21632
rect 33520 21593 33548 21830
rect 33506 21584 33562 21593
rect 33612 21554 33640 22578
rect 33506 21519 33562 21528
rect 33600 21548 33652 21554
rect 33600 21490 33652 21496
rect 33612 21418 33640 21490
rect 33600 21412 33652 21418
rect 33600 21354 33652 21360
rect 33244 21100 33364 21128
rect 33244 20534 33272 21100
rect 33704 21078 33732 22918
rect 33888 22817 33916 26302
rect 34426 26200 34482 26302
rect 35070 26330 35126 27000
rect 35714 26330 35770 27000
rect 36082 26344 36138 26353
rect 35070 26302 35480 26330
rect 35070 26200 35126 26302
rect 34702 25256 34758 25265
rect 34702 25191 34758 25200
rect 34426 24848 34482 24857
rect 33968 24812 34020 24818
rect 34426 24783 34482 24792
rect 33968 24754 34020 24760
rect 33980 24313 34008 24754
rect 34152 24676 34204 24682
rect 34152 24618 34204 24624
rect 34164 24410 34192 24618
rect 34152 24404 34204 24410
rect 34152 24346 34204 24352
rect 33966 24304 34022 24313
rect 33966 24239 34022 24248
rect 33968 24064 34020 24070
rect 33968 24006 34020 24012
rect 34150 24032 34206 24041
rect 33874 22808 33930 22817
rect 33874 22743 33930 22752
rect 33980 21894 34008 24006
rect 34150 23967 34206 23976
rect 34060 23792 34112 23798
rect 34060 23734 34112 23740
rect 34072 23254 34100 23734
rect 34164 23254 34192 23967
rect 34336 23656 34388 23662
rect 34336 23598 34388 23604
rect 34242 23352 34298 23361
rect 34242 23287 34298 23296
rect 34060 23248 34112 23254
rect 34060 23190 34112 23196
rect 34152 23248 34204 23254
rect 34152 23190 34204 23196
rect 34164 22817 34192 23190
rect 34150 22808 34206 22817
rect 34150 22743 34206 22752
rect 34256 22166 34284 23287
rect 34244 22160 34296 22166
rect 34244 22102 34296 22108
rect 33784 21888 33836 21894
rect 33782 21856 33784 21865
rect 33968 21888 34020 21894
rect 33836 21856 33838 21865
rect 33968 21830 34020 21836
rect 34058 21856 34114 21865
rect 33782 21791 33838 21800
rect 33796 21350 33824 21791
rect 33784 21344 33836 21350
rect 33784 21286 33836 21292
rect 33782 21176 33838 21185
rect 33782 21111 33784 21120
rect 33836 21111 33838 21120
rect 33784 21082 33836 21088
rect 33692 21072 33744 21078
rect 33692 21014 33744 21020
rect 33508 21004 33560 21010
rect 33508 20946 33560 20952
rect 33324 20800 33376 20806
rect 33324 20742 33376 20748
rect 33232 20528 33284 20534
rect 33232 20470 33284 20476
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 33230 19952 33286 19961
rect 33140 19916 33192 19922
rect 33230 19887 33286 19896
rect 33140 19858 33192 19864
rect 33152 19786 33180 19858
rect 33140 19780 33192 19786
rect 33140 19722 33192 19728
rect 33244 19718 33272 19887
rect 33232 19712 33284 19718
rect 33232 19654 33284 19660
rect 33336 19514 33364 20742
rect 33520 19802 33548 20946
rect 33690 20904 33746 20913
rect 33690 20839 33746 20848
rect 33428 19774 33548 19802
rect 33598 19816 33654 19825
rect 33048 19508 33100 19514
rect 33048 19450 33100 19456
rect 33324 19508 33376 19514
rect 33324 19450 33376 19456
rect 32954 19408 33010 19417
rect 32954 19343 33010 19352
rect 32968 19310 32996 19343
rect 32956 19304 33008 19310
rect 32956 19246 33008 19252
rect 33060 19224 33088 19450
rect 33060 19196 33364 19224
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 33336 18952 33364 19196
rect 33060 18924 33364 18952
rect 32862 18864 32918 18873
rect 32862 18799 32918 18808
rect 33060 18601 33088 18924
rect 33324 18624 33376 18630
rect 33046 18592 33102 18601
rect 33324 18566 33376 18572
rect 33046 18527 33102 18536
rect 33060 18329 33088 18527
rect 33336 18358 33364 18566
rect 33324 18352 33376 18358
rect 33046 18320 33102 18329
rect 33324 18294 33376 18300
rect 33046 18255 33102 18264
rect 33428 18222 33456 19774
rect 33598 19751 33600 19760
rect 33652 19751 33654 19760
rect 33600 19722 33652 19728
rect 33508 19712 33560 19718
rect 33508 19654 33560 19660
rect 33232 18216 33284 18222
rect 33230 18184 33232 18193
rect 33324 18216 33376 18222
rect 33284 18184 33286 18193
rect 33324 18158 33376 18164
rect 33416 18216 33468 18222
rect 33416 18158 33468 18164
rect 33230 18119 33286 18128
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 32864 17264 32916 17270
rect 32862 17232 32864 17241
rect 32916 17232 32918 17241
rect 33336 17218 33364 18158
rect 33428 17814 33456 18158
rect 33416 17808 33468 17814
rect 33416 17750 33468 17756
rect 33336 17190 33456 17218
rect 32862 17167 32918 17176
rect 33324 17128 33376 17134
rect 33324 17070 33376 17076
rect 32864 16992 32916 16998
rect 32864 16934 32916 16940
rect 32876 16250 32904 16934
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 33336 16794 33364 17070
rect 33324 16788 33376 16794
rect 33324 16730 33376 16736
rect 33336 16658 33364 16730
rect 33428 16658 33456 17190
rect 33324 16652 33376 16658
rect 33324 16594 33376 16600
rect 33416 16652 33468 16658
rect 33416 16594 33468 16600
rect 33414 16552 33470 16561
rect 33414 16487 33470 16496
rect 33324 16448 33376 16454
rect 33324 16390 33376 16396
rect 32864 16244 32916 16250
rect 32864 16186 32916 16192
rect 32876 16153 32904 16186
rect 32862 16144 32918 16153
rect 32862 16079 32918 16088
rect 32862 16008 32918 16017
rect 32862 15943 32918 15952
rect 32772 15496 32824 15502
rect 32772 15438 32824 15444
rect 32876 14822 32904 15943
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 32956 15360 33008 15366
rect 32954 15328 32956 15337
rect 33008 15328 33010 15337
rect 32954 15263 33010 15272
rect 33232 15156 33284 15162
rect 33232 15098 33284 15104
rect 33244 14822 33272 15098
rect 32864 14816 32916 14822
rect 32678 14784 32734 14793
rect 32864 14758 32916 14764
rect 33232 14816 33284 14822
rect 33232 14758 33284 14764
rect 32678 14719 32734 14728
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32770 14648 32826 14657
rect 32950 14651 33258 14660
rect 33336 14618 33364 16390
rect 33428 15570 33456 16487
rect 33520 15910 33548 19654
rect 33598 19272 33654 19281
rect 33598 19207 33654 19216
rect 33612 18834 33640 19207
rect 33600 18828 33652 18834
rect 33600 18770 33652 18776
rect 33598 18728 33654 18737
rect 33598 18663 33654 18672
rect 33612 18358 33640 18663
rect 33600 18352 33652 18358
rect 33600 18294 33652 18300
rect 33612 17746 33640 18294
rect 33600 17740 33652 17746
rect 33600 17682 33652 17688
rect 33704 16794 33732 20839
rect 33796 20806 33824 21082
rect 33784 20800 33836 20806
rect 33784 20742 33836 20748
rect 33980 20505 34008 21830
rect 34058 21791 34114 21800
rect 34072 21622 34100 21791
rect 34060 21616 34112 21622
rect 34060 21558 34112 21564
rect 34060 21140 34112 21146
rect 34060 21082 34112 21088
rect 34072 20942 34100 21082
rect 34060 20936 34112 20942
rect 34060 20878 34112 20884
rect 33966 20496 34022 20505
rect 33888 20454 33966 20482
rect 33784 20052 33836 20058
rect 33784 19994 33836 20000
rect 33796 19786 33824 19994
rect 33784 19780 33836 19786
rect 33784 19722 33836 19728
rect 33782 19272 33838 19281
rect 33782 19207 33784 19216
rect 33836 19207 33838 19216
rect 33784 19178 33836 19184
rect 33888 18952 33916 20454
rect 33966 20431 34022 20440
rect 34072 20398 34100 20878
rect 34256 20534 34284 22102
rect 34348 21894 34376 23598
rect 34440 22438 34468 24783
rect 34716 23712 34744 25191
rect 34980 24268 35032 24274
rect 34980 24210 35032 24216
rect 34716 23684 34836 23712
rect 34704 23588 34756 23594
rect 34704 23530 34756 23536
rect 34612 23180 34664 23186
rect 34612 23122 34664 23128
rect 34520 23044 34572 23050
rect 34520 22986 34572 22992
rect 34532 22953 34560 22986
rect 34518 22944 34574 22953
rect 34518 22879 34574 22888
rect 34624 22545 34652 23122
rect 34610 22536 34666 22545
rect 34610 22471 34666 22480
rect 34428 22432 34480 22438
rect 34428 22374 34480 22380
rect 34428 22160 34480 22166
rect 34428 22102 34480 22108
rect 34336 21888 34388 21894
rect 34336 21830 34388 21836
rect 34440 21729 34468 22102
rect 34716 22094 34744 23530
rect 34624 22066 34744 22094
rect 34624 22030 34652 22066
rect 34612 22024 34664 22030
rect 34612 21966 34664 21972
rect 34702 21992 34758 22001
rect 34702 21927 34758 21936
rect 34426 21720 34482 21729
rect 34426 21655 34482 21664
rect 34440 20913 34468 21655
rect 34426 20904 34482 20913
rect 34426 20839 34482 20848
rect 34428 20800 34480 20806
rect 34428 20742 34480 20748
rect 34244 20528 34296 20534
rect 34164 20488 34244 20516
rect 34060 20392 34112 20398
rect 34060 20334 34112 20340
rect 34060 20256 34112 20262
rect 34060 20198 34112 20204
rect 33968 20052 34020 20058
rect 33968 19994 34020 20000
rect 33796 18924 33916 18952
rect 33692 16788 33744 16794
rect 33692 16730 33744 16736
rect 33600 16448 33652 16454
rect 33600 16390 33652 16396
rect 33692 16448 33744 16454
rect 33692 16390 33744 16396
rect 33508 15904 33560 15910
rect 33508 15846 33560 15852
rect 33416 15564 33468 15570
rect 33416 15506 33468 15512
rect 33416 15020 33468 15026
rect 33416 14962 33468 14968
rect 32770 14583 32826 14592
rect 33324 14612 33376 14618
rect 32784 14482 32812 14583
rect 33324 14554 33376 14560
rect 32588 14476 32640 14482
rect 32588 14418 32640 14424
rect 32772 14476 32824 14482
rect 32772 14418 32824 14424
rect 32600 13530 32628 14418
rect 32680 14340 32732 14346
rect 32680 14282 32732 14288
rect 32692 14006 32720 14282
rect 32772 14068 32824 14074
rect 32772 14010 32824 14016
rect 32680 14000 32732 14006
rect 32680 13942 32732 13948
rect 32588 13524 32640 13530
rect 32588 13466 32640 13472
rect 32680 13456 32732 13462
rect 32680 13398 32732 13404
rect 32692 13190 32720 13398
rect 32784 13258 32812 14010
rect 33140 13932 33192 13938
rect 33192 13892 33364 13920
rect 33140 13874 33192 13880
rect 32864 13796 32916 13802
rect 32864 13738 32916 13744
rect 32876 13433 32904 13738
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 33336 13530 33364 13892
rect 33324 13524 33376 13530
rect 33324 13466 33376 13472
rect 32862 13424 32918 13433
rect 32862 13359 32918 13368
rect 32772 13252 32824 13258
rect 32772 13194 32824 13200
rect 32680 13184 32732 13190
rect 32680 13126 32732 13132
rect 32784 11898 32812 13194
rect 33324 12640 33376 12646
rect 33324 12582 33376 12588
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 32864 12096 32916 12102
rect 32864 12038 32916 12044
rect 32876 11898 32904 12038
rect 32772 11892 32824 11898
rect 32772 11834 32824 11840
rect 32864 11892 32916 11898
rect 32864 11834 32916 11840
rect 32680 11756 32732 11762
rect 32680 11698 32732 11704
rect 32588 11008 32640 11014
rect 32588 10950 32640 10956
rect 32600 9761 32628 10950
rect 32692 10606 32720 11698
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32770 11384 32826 11393
rect 32950 11387 33258 11396
rect 32770 11319 32772 11328
rect 32824 11319 32826 11328
rect 32772 11290 32824 11296
rect 32784 10690 32812 11290
rect 32784 10674 32904 10690
rect 32784 10668 32916 10674
rect 32784 10662 32864 10668
rect 32864 10610 32916 10616
rect 32680 10600 32732 10606
rect 32680 10542 32732 10548
rect 32772 10600 32824 10606
rect 32772 10542 32824 10548
rect 32586 9752 32642 9761
rect 32586 9687 32642 9696
rect 32588 9648 32640 9654
rect 32588 9590 32640 9596
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 32600 7546 32628 9590
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 32588 7540 32640 7546
rect 32588 7482 32640 7488
rect 32220 6860 32272 6866
rect 32220 6802 32272 6808
rect 32312 6792 32364 6798
rect 32312 6734 32364 6740
rect 32324 6458 32352 6734
rect 32312 6452 32364 6458
rect 32312 6394 32364 6400
rect 32036 6316 32088 6322
rect 32036 6258 32088 6264
rect 31484 5364 31536 5370
rect 31484 5306 31536 5312
rect 32692 5302 32720 8434
rect 32784 7410 32812 10542
rect 33336 10470 33364 12582
rect 33428 11150 33456 14962
rect 33508 14952 33560 14958
rect 33508 14894 33560 14900
rect 33520 14074 33548 14894
rect 33508 14068 33560 14074
rect 33508 14010 33560 14016
rect 33508 13388 33560 13394
rect 33508 13330 33560 13336
rect 33520 12238 33548 13330
rect 33508 12232 33560 12238
rect 33508 12174 33560 12180
rect 33520 11694 33548 12174
rect 33508 11688 33560 11694
rect 33508 11630 33560 11636
rect 33416 11144 33468 11150
rect 33416 11086 33468 11092
rect 33520 10538 33548 11630
rect 33508 10532 33560 10538
rect 33508 10474 33560 10480
rect 33324 10464 33376 10470
rect 33324 10406 33376 10412
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 33520 10130 33548 10474
rect 33508 10124 33560 10130
rect 33508 10066 33560 10072
rect 32864 9716 32916 9722
rect 32864 9658 32916 9664
rect 32876 8634 32904 9658
rect 33324 9648 33376 9654
rect 33324 9590 33376 9596
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 33336 8974 33364 9590
rect 33612 9194 33640 16390
rect 33704 16182 33732 16390
rect 33692 16176 33744 16182
rect 33692 16118 33744 16124
rect 33690 15192 33746 15201
rect 33690 15127 33746 15136
rect 33704 15026 33732 15127
rect 33692 15020 33744 15026
rect 33692 14962 33744 14968
rect 33704 14396 33732 14962
rect 33796 14498 33824 18924
rect 33876 18828 33928 18834
rect 33876 18770 33928 18776
rect 33888 17066 33916 18770
rect 33980 18086 34008 19994
rect 34072 19446 34100 20198
rect 34164 19990 34192 20488
rect 34244 20470 34296 20476
rect 34152 19984 34204 19990
rect 34152 19926 34204 19932
rect 34244 19916 34296 19922
rect 34244 19858 34296 19864
rect 34060 19440 34112 19446
rect 34060 19382 34112 19388
rect 34256 19378 34284 19858
rect 34440 19446 34468 20742
rect 34716 20534 34744 21927
rect 34704 20528 34756 20534
rect 34704 20470 34756 20476
rect 34520 19780 34572 19786
rect 34520 19722 34572 19728
rect 34428 19440 34480 19446
rect 34428 19382 34480 19388
rect 34152 19372 34204 19378
rect 34152 19314 34204 19320
rect 34244 19372 34296 19378
rect 34244 19314 34296 19320
rect 34060 19168 34112 19174
rect 34060 19110 34112 19116
rect 34072 18698 34100 19110
rect 34060 18692 34112 18698
rect 34060 18634 34112 18640
rect 34060 18216 34112 18222
rect 34060 18158 34112 18164
rect 33968 18080 34020 18086
rect 33968 18022 34020 18028
rect 34072 17728 34100 18158
rect 34164 17882 34192 19314
rect 34336 19304 34388 19310
rect 34334 19272 34336 19281
rect 34388 19272 34390 19281
rect 34334 19207 34390 19216
rect 34244 18828 34296 18834
rect 34244 18770 34296 18776
rect 34152 17876 34204 17882
rect 34152 17818 34204 17824
rect 34152 17740 34204 17746
rect 34072 17700 34152 17728
rect 34152 17682 34204 17688
rect 34256 17649 34284 18770
rect 34334 18728 34390 18737
rect 34334 18663 34336 18672
rect 34388 18663 34390 18672
rect 34336 18634 34388 18640
rect 34440 18426 34468 19382
rect 34428 18420 34480 18426
rect 34428 18362 34480 18368
rect 34336 18352 34388 18358
rect 34336 18294 34388 18300
rect 34348 17921 34376 18294
rect 34428 18216 34480 18222
rect 34428 18158 34480 18164
rect 34334 17912 34390 17921
rect 34334 17847 34390 17856
rect 34440 17678 34468 18158
rect 34532 17746 34560 19722
rect 34808 19718 34836 23684
rect 34992 23526 35020 24210
rect 35256 24200 35308 24206
rect 35256 24142 35308 24148
rect 35072 23656 35124 23662
rect 35072 23598 35124 23604
rect 34888 23520 34940 23526
rect 34888 23462 34940 23468
rect 34980 23520 35032 23526
rect 34980 23462 35032 23468
rect 34900 23186 34928 23462
rect 34888 23180 34940 23186
rect 34888 23122 34940 23128
rect 34900 21010 34928 23122
rect 34980 22432 35032 22438
rect 34980 22374 35032 22380
rect 34992 22234 35020 22374
rect 34980 22228 35032 22234
rect 34980 22170 35032 22176
rect 34980 22024 35032 22030
rect 34980 21966 35032 21972
rect 34888 21004 34940 21010
rect 34888 20946 34940 20952
rect 34888 20256 34940 20262
rect 34888 20198 34940 20204
rect 34796 19712 34848 19718
rect 34796 19654 34848 19660
rect 34796 19372 34848 19378
rect 34796 19314 34848 19320
rect 34702 19272 34758 19281
rect 34702 19207 34758 19216
rect 34612 18828 34664 18834
rect 34612 18770 34664 18776
rect 34520 17740 34572 17746
rect 34520 17682 34572 17688
rect 34428 17672 34480 17678
rect 34242 17640 34298 17649
rect 34428 17614 34480 17620
rect 34242 17575 34298 17584
rect 34060 17536 34112 17542
rect 34060 17478 34112 17484
rect 33876 17060 33928 17066
rect 33876 17002 33928 17008
rect 34072 16697 34100 17478
rect 34336 16992 34388 16998
rect 34334 16960 34336 16969
rect 34388 16960 34390 16969
rect 34334 16895 34390 16904
rect 34244 16788 34296 16794
rect 34244 16730 34296 16736
rect 34058 16688 34114 16697
rect 34058 16623 34114 16632
rect 33968 16040 34020 16046
rect 33968 15982 34020 15988
rect 33980 14618 34008 15982
rect 34072 15366 34100 16623
rect 34152 16108 34204 16114
rect 34152 16050 34204 16056
rect 34164 15570 34192 16050
rect 34152 15564 34204 15570
rect 34152 15506 34204 15512
rect 34060 15360 34112 15366
rect 34060 15302 34112 15308
rect 33968 14612 34020 14618
rect 33968 14554 34020 14560
rect 33796 14470 33916 14498
rect 33784 14408 33836 14414
rect 33704 14368 33784 14396
rect 33704 13394 33732 14368
rect 33784 14350 33836 14356
rect 33782 13968 33838 13977
rect 33782 13903 33838 13912
rect 33692 13388 33744 13394
rect 33692 13330 33744 13336
rect 33796 12170 33824 13903
rect 33784 12164 33836 12170
rect 33784 12106 33836 12112
rect 33796 12073 33824 12106
rect 33782 12064 33838 12073
rect 33782 11999 33838 12008
rect 33690 11928 33746 11937
rect 33690 11863 33746 11872
rect 33704 11121 33732 11863
rect 33784 11688 33836 11694
rect 33784 11630 33836 11636
rect 33690 11112 33746 11121
rect 33690 11047 33746 11056
rect 33796 10266 33824 11630
rect 33784 10260 33836 10266
rect 33784 10202 33836 10208
rect 33690 9888 33746 9897
rect 33690 9823 33746 9832
rect 33428 9166 33640 9194
rect 33324 8968 33376 8974
rect 33324 8910 33376 8916
rect 32864 8628 32916 8634
rect 32864 8570 32916 8576
rect 32864 8424 32916 8430
rect 33048 8424 33100 8430
rect 32864 8366 32916 8372
rect 33046 8392 33048 8401
rect 33100 8392 33102 8401
rect 32876 7970 32904 8366
rect 33046 8327 33102 8336
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 32876 7942 32996 7970
rect 32968 7886 32996 7942
rect 32956 7880 33008 7886
rect 33324 7880 33376 7886
rect 32956 7822 33008 7828
rect 33322 7848 33324 7857
rect 33376 7848 33378 7857
rect 32864 7812 32916 7818
rect 33322 7783 33378 7792
rect 32864 7754 32916 7760
rect 32772 7404 32824 7410
rect 32772 7346 32824 7352
rect 32876 6390 32904 7754
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 32864 6384 32916 6390
rect 32864 6326 32916 6332
rect 33428 6089 33456 9166
rect 33704 9110 33732 9823
rect 33888 9586 33916 14470
rect 34060 14408 34112 14414
rect 34060 14350 34112 14356
rect 33966 13832 34022 13841
rect 33966 13767 34022 13776
rect 33980 12617 34008 13767
rect 34072 13569 34100 14350
rect 34058 13560 34114 13569
rect 34058 13495 34060 13504
rect 34112 13495 34114 13504
rect 34060 13466 34112 13472
rect 34256 13394 34284 16730
rect 34348 16046 34376 16895
rect 34440 16658 34468 17614
rect 34532 17202 34560 17682
rect 34520 17196 34572 17202
rect 34520 17138 34572 17144
rect 34428 16652 34480 16658
rect 34428 16594 34480 16600
rect 34336 16040 34388 16046
rect 34336 15982 34388 15988
rect 34624 15892 34652 18770
rect 34716 18737 34744 19207
rect 34808 19145 34836 19314
rect 34794 19136 34850 19145
rect 34794 19071 34850 19080
rect 34702 18728 34758 18737
rect 34702 18663 34758 18672
rect 34796 18624 34848 18630
rect 34796 18566 34848 18572
rect 34704 18352 34756 18358
rect 34702 18320 34704 18329
rect 34756 18320 34758 18329
rect 34702 18255 34758 18264
rect 34704 17740 34756 17746
rect 34704 17682 34756 17688
rect 34716 17105 34744 17682
rect 34702 17096 34758 17105
rect 34702 17031 34758 17040
rect 34704 16788 34756 16794
rect 34704 16730 34756 16736
rect 34716 16250 34744 16730
rect 34704 16244 34756 16250
rect 34704 16186 34756 16192
rect 34808 16182 34836 18566
rect 34900 17338 34928 20198
rect 34992 17882 35020 21966
rect 35084 21457 35112 23598
rect 35164 22704 35216 22710
rect 35164 22646 35216 22652
rect 35176 21554 35204 22646
rect 35268 21978 35296 24142
rect 35348 22568 35400 22574
rect 35348 22510 35400 22516
rect 35360 22234 35388 22510
rect 35348 22228 35400 22234
rect 35348 22170 35400 22176
rect 35268 21950 35388 21978
rect 35256 21888 35308 21894
rect 35256 21830 35308 21836
rect 35268 21593 35296 21830
rect 35254 21584 35310 21593
rect 35164 21548 35216 21554
rect 35254 21519 35310 21528
rect 35164 21490 35216 21496
rect 35256 21480 35308 21486
rect 35070 21448 35126 21457
rect 35256 21422 35308 21428
rect 35070 21383 35126 21392
rect 35084 20856 35112 21383
rect 35084 20828 35204 20856
rect 35070 20496 35126 20505
rect 35070 20431 35072 20440
rect 35124 20431 35126 20440
rect 35072 20402 35124 20408
rect 35176 20097 35204 20828
rect 35162 20088 35218 20097
rect 35162 20023 35218 20032
rect 35164 19984 35216 19990
rect 35070 19952 35126 19961
rect 35164 19926 35216 19932
rect 35070 19887 35126 19896
rect 34980 17876 35032 17882
rect 34980 17818 35032 17824
rect 34888 17332 34940 17338
rect 34888 17274 34940 17280
rect 34888 16584 34940 16590
rect 34888 16526 34940 16532
rect 34796 16176 34848 16182
rect 34796 16118 34848 16124
rect 34900 16114 34928 16526
rect 34888 16108 34940 16114
rect 34888 16050 34940 16056
rect 34704 15904 34756 15910
rect 34624 15864 34704 15892
rect 34756 15864 34928 15892
rect 34704 15846 34756 15852
rect 34716 15706 34744 15846
rect 34900 15722 34928 15864
rect 34704 15700 34756 15706
rect 34900 15694 35020 15722
rect 34704 15642 34756 15648
rect 34336 15564 34388 15570
rect 34336 15506 34388 15512
rect 34348 14958 34376 15506
rect 34612 15360 34664 15366
rect 34612 15302 34664 15308
rect 34336 14952 34388 14958
rect 34388 14912 34468 14940
rect 34336 14894 34388 14900
rect 34336 14816 34388 14822
rect 34336 14758 34388 14764
rect 34348 14278 34376 14758
rect 34336 14272 34388 14278
rect 34336 14214 34388 14220
rect 34244 13388 34296 13394
rect 34244 13330 34296 13336
rect 34060 13320 34112 13326
rect 34060 13262 34112 13268
rect 33966 12608 34022 12617
rect 33966 12543 34022 12552
rect 34072 12102 34100 13262
rect 34244 12776 34296 12782
rect 34244 12718 34296 12724
rect 33968 12096 34020 12102
rect 33968 12038 34020 12044
rect 34060 12096 34112 12102
rect 34060 12038 34112 12044
rect 33980 11529 34008 12038
rect 33966 11520 34022 11529
rect 33966 11455 34022 11464
rect 34072 11370 34100 12038
rect 33980 11342 34100 11370
rect 33876 9580 33928 9586
rect 33876 9522 33928 9528
rect 33784 9512 33836 9518
rect 33980 9466 34008 11342
rect 34060 11280 34112 11286
rect 34060 11222 34112 11228
rect 33784 9454 33836 9460
rect 33796 9217 33824 9454
rect 33888 9438 34008 9466
rect 33782 9208 33838 9217
rect 33782 9143 33838 9152
rect 33692 9104 33744 9110
rect 33692 9046 33744 9052
rect 33508 8968 33560 8974
rect 33508 8910 33560 8916
rect 33520 6458 33548 8910
rect 33704 6798 33732 9046
rect 33692 6792 33744 6798
rect 33692 6734 33744 6740
rect 33508 6452 33560 6458
rect 33508 6394 33560 6400
rect 33414 6080 33470 6089
rect 32950 6012 33258 6021
rect 33414 6015 33470 6024
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 32680 5296 32732 5302
rect 32680 5238 32732 5244
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 32864 4276 32916 4282
rect 32864 4218 32916 4224
rect 30840 3936 30892 3942
rect 30840 3878 30892 3884
rect 30852 2650 30880 3878
rect 32876 2650 32904 4218
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 33888 3738 33916 9438
rect 33968 9376 34020 9382
rect 33968 9318 34020 9324
rect 33980 8634 34008 9318
rect 34072 8634 34100 11222
rect 34152 11144 34204 11150
rect 34150 11112 34152 11121
rect 34204 11112 34206 11121
rect 34150 11047 34206 11056
rect 34152 9920 34204 9926
rect 34152 9862 34204 9868
rect 34164 9042 34192 9862
rect 34256 9722 34284 12718
rect 34348 12102 34376 14214
rect 34440 13818 34468 14912
rect 34624 14278 34652 15302
rect 34888 15020 34940 15026
rect 34888 14962 34940 14968
rect 34796 14340 34848 14346
rect 34796 14282 34848 14288
rect 34612 14272 34664 14278
rect 34612 14214 34664 14220
rect 34440 13790 34560 13818
rect 34428 13728 34480 13734
rect 34426 13696 34428 13705
rect 34480 13696 34482 13705
rect 34426 13631 34482 13640
rect 34428 13388 34480 13394
rect 34428 13330 34480 13336
rect 34336 12096 34388 12102
rect 34336 12038 34388 12044
rect 34334 11520 34390 11529
rect 34334 11455 34390 11464
rect 34348 10169 34376 11455
rect 34334 10160 34390 10169
rect 34334 10095 34390 10104
rect 34244 9716 34296 9722
rect 34244 9658 34296 9664
rect 34244 9376 34296 9382
rect 34244 9318 34296 9324
rect 34152 9036 34204 9042
rect 34152 8978 34204 8984
rect 34256 8906 34284 9318
rect 34244 8900 34296 8906
rect 34244 8842 34296 8848
rect 33968 8628 34020 8634
rect 33968 8570 34020 8576
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 34256 8430 34284 8842
rect 34244 8424 34296 8430
rect 34244 8366 34296 8372
rect 34348 6390 34376 10095
rect 34440 9518 34468 13330
rect 34532 13258 34560 13790
rect 34624 13734 34652 14214
rect 34704 13864 34756 13870
rect 34704 13806 34756 13812
rect 34612 13728 34664 13734
rect 34612 13670 34664 13676
rect 34520 13252 34572 13258
rect 34520 13194 34572 13200
rect 34612 12776 34664 12782
rect 34612 12718 34664 12724
rect 34624 12306 34652 12718
rect 34612 12300 34664 12306
rect 34612 12242 34664 12248
rect 34518 12200 34574 12209
rect 34518 12135 34574 12144
rect 34532 11694 34560 12135
rect 34520 11688 34572 11694
rect 34572 11648 34652 11676
rect 34520 11630 34572 11636
rect 34518 10296 34574 10305
rect 34518 10231 34574 10240
rect 34532 10198 34560 10231
rect 34520 10192 34572 10198
rect 34520 10134 34572 10140
rect 34428 9512 34480 9518
rect 34428 9454 34480 9460
rect 34426 7984 34482 7993
rect 34426 7919 34482 7928
rect 34440 7750 34468 7919
rect 34520 7880 34572 7886
rect 34624 7868 34652 11648
rect 34716 9110 34744 13806
rect 34808 9654 34836 14282
rect 34900 13530 34928 14962
rect 34888 13524 34940 13530
rect 34888 13466 34940 13472
rect 34900 13297 34928 13466
rect 34886 13288 34942 13297
rect 34886 13223 34942 13232
rect 34992 13172 35020 15694
rect 34900 13144 35020 13172
rect 34900 11354 34928 13144
rect 35084 13002 35112 19887
rect 35176 19242 35204 19926
rect 35164 19236 35216 19242
rect 35164 19178 35216 19184
rect 35268 19009 35296 21422
rect 35360 21049 35388 21950
rect 35346 21040 35402 21049
rect 35346 20975 35402 20984
rect 35348 20392 35400 20398
rect 35346 20360 35348 20369
rect 35400 20360 35402 20369
rect 35346 20295 35402 20304
rect 35348 20256 35400 20262
rect 35348 20198 35400 20204
rect 35254 19000 35310 19009
rect 35254 18935 35310 18944
rect 35268 18698 35296 18935
rect 35256 18692 35308 18698
rect 35256 18634 35308 18640
rect 35164 16176 35216 16182
rect 35164 16118 35216 16124
rect 35176 13326 35204 16118
rect 35254 16008 35310 16017
rect 35254 15943 35310 15952
rect 35164 13320 35216 13326
rect 35164 13262 35216 13268
rect 35084 12974 35204 13002
rect 35072 12912 35124 12918
rect 35072 12854 35124 12860
rect 34980 12096 35032 12102
rect 34980 12038 35032 12044
rect 34888 11348 34940 11354
rect 34888 11290 34940 11296
rect 34992 11286 35020 12038
rect 35084 11354 35112 12854
rect 35176 11354 35204 12974
rect 35268 12782 35296 15943
rect 35360 15162 35388 20198
rect 35452 19122 35480 26302
rect 35714 26302 35848 26330
rect 35714 26200 35770 26302
rect 35820 26178 35848 26302
rect 36082 26279 36138 26288
rect 36358 26330 36414 27000
rect 36358 26302 36768 26330
rect 35808 26172 35860 26178
rect 35808 26114 35860 26120
rect 35900 25220 35952 25226
rect 35900 25162 35952 25168
rect 35532 24676 35584 24682
rect 35532 24618 35584 24624
rect 35544 24274 35572 24618
rect 35532 24268 35584 24274
rect 35532 24210 35584 24216
rect 35808 24268 35860 24274
rect 35808 24210 35860 24216
rect 35544 22982 35572 24210
rect 35624 24200 35676 24206
rect 35624 24142 35676 24148
rect 35636 23594 35664 24142
rect 35716 24064 35768 24070
rect 35716 24006 35768 24012
rect 35624 23588 35676 23594
rect 35624 23530 35676 23536
rect 35532 22976 35584 22982
rect 35532 22918 35584 22924
rect 35728 22273 35756 24006
rect 35714 22264 35770 22273
rect 35714 22199 35770 22208
rect 35530 22128 35586 22137
rect 35530 22063 35586 22072
rect 35544 21350 35572 22063
rect 35624 21548 35676 21554
rect 35624 21490 35676 21496
rect 35532 21344 35584 21350
rect 35532 21286 35584 21292
rect 35544 19990 35572 21286
rect 35636 20874 35664 21490
rect 35624 20868 35676 20874
rect 35624 20810 35676 20816
rect 35532 19984 35584 19990
rect 35532 19926 35584 19932
rect 35622 19680 35678 19689
rect 35622 19615 35678 19624
rect 35636 19242 35664 19615
rect 35624 19236 35676 19242
rect 35624 19178 35676 19184
rect 35452 19094 35572 19122
rect 35438 18864 35494 18873
rect 35438 18799 35494 18808
rect 35452 18698 35480 18799
rect 35440 18692 35492 18698
rect 35440 18634 35492 18640
rect 35544 18057 35572 19094
rect 35530 18048 35586 18057
rect 35530 17983 35586 17992
rect 35532 17740 35584 17746
rect 35532 17682 35584 17688
rect 35544 17338 35572 17682
rect 35728 17377 35756 22199
rect 35820 21690 35848 24210
rect 35912 21865 35940 25162
rect 35992 22500 36044 22506
rect 35992 22442 36044 22448
rect 35898 21856 35954 21865
rect 35898 21791 35954 21800
rect 35808 21684 35860 21690
rect 35808 21626 35860 21632
rect 35898 20632 35954 20641
rect 35898 20567 35954 20576
rect 35912 20466 35940 20567
rect 35900 20460 35952 20466
rect 35900 20402 35952 20408
rect 35808 20392 35860 20398
rect 36004 20346 36032 22442
rect 36096 22094 36124 26279
rect 36358 26200 36414 26302
rect 36174 25120 36230 25129
rect 36174 25055 36230 25064
rect 36188 22438 36216 25055
rect 36452 24064 36504 24070
rect 36452 24006 36504 24012
rect 36544 24064 36596 24070
rect 36544 24006 36596 24012
rect 36464 23905 36492 24006
rect 36450 23896 36506 23905
rect 36556 23866 36584 24006
rect 36450 23831 36506 23840
rect 36544 23860 36596 23866
rect 36544 23802 36596 23808
rect 36360 23724 36412 23730
rect 36360 23666 36412 23672
rect 36372 23633 36400 23666
rect 36452 23656 36504 23662
rect 36358 23624 36414 23633
rect 36452 23598 36504 23604
rect 36358 23559 36414 23568
rect 36268 23248 36320 23254
rect 36268 23190 36320 23196
rect 36176 22432 36228 22438
rect 36176 22374 36228 22380
rect 36096 22066 36216 22094
rect 36188 21010 36216 22066
rect 36280 21622 36308 23190
rect 36360 22092 36412 22098
rect 36360 22034 36412 22040
rect 36372 21894 36400 22034
rect 36360 21888 36412 21894
rect 36360 21830 36412 21836
rect 36268 21616 36320 21622
rect 36268 21558 36320 21564
rect 36360 21548 36412 21554
rect 36360 21490 36412 21496
rect 36268 21480 36320 21486
rect 36268 21422 36320 21428
rect 36176 21004 36228 21010
rect 36176 20946 36228 20952
rect 36174 20768 36230 20777
rect 36174 20703 36230 20712
rect 36082 20632 36138 20641
rect 36082 20567 36138 20576
rect 35808 20334 35860 20340
rect 35820 18193 35848 20334
rect 35912 20318 36032 20346
rect 35912 19689 35940 20318
rect 35990 19816 36046 19825
rect 35990 19751 36046 19760
rect 35898 19680 35954 19689
rect 35898 19615 35954 19624
rect 35900 19168 35952 19174
rect 35900 19110 35952 19116
rect 35806 18184 35862 18193
rect 35806 18119 35862 18128
rect 35820 17746 35848 18119
rect 35912 17814 35940 19110
rect 36004 18086 36032 19751
rect 36096 19378 36124 20567
rect 36188 19378 36216 20703
rect 36280 19922 36308 21422
rect 36372 21350 36400 21490
rect 36360 21344 36412 21350
rect 36360 21286 36412 21292
rect 36268 19916 36320 19922
rect 36268 19858 36320 19864
rect 36372 19786 36400 21286
rect 36464 20330 36492 23598
rect 36740 23361 36768 26302
rect 37002 26200 37058 27000
rect 37646 26200 37702 27000
rect 38290 26200 38346 27000
rect 38934 26200 38990 27000
rect 39578 26330 39634 27000
rect 39316 26302 39634 26330
rect 36820 24880 36872 24886
rect 36820 24822 36872 24828
rect 36832 24274 36860 24822
rect 36820 24268 36872 24274
rect 36820 24210 36872 24216
rect 36818 23624 36874 23633
rect 36818 23559 36874 23568
rect 36726 23352 36782 23361
rect 36832 23322 36860 23559
rect 36912 23520 36964 23526
rect 37016 23497 37044 26200
rect 37556 24676 37608 24682
rect 37556 24618 37608 24624
rect 37464 24608 37516 24614
rect 37464 24550 37516 24556
rect 37476 24410 37504 24550
rect 37464 24404 37516 24410
rect 37464 24346 37516 24352
rect 37188 23656 37240 23662
rect 37188 23598 37240 23604
rect 37464 23656 37516 23662
rect 37464 23598 37516 23604
rect 36912 23462 36964 23468
rect 37002 23488 37058 23497
rect 36726 23287 36782 23296
rect 36820 23316 36872 23322
rect 36820 23258 36872 23264
rect 36544 23044 36596 23050
rect 36544 22986 36596 22992
rect 36556 22710 36584 22986
rect 36544 22704 36596 22710
rect 36544 22646 36596 22652
rect 36544 22568 36596 22574
rect 36544 22510 36596 22516
rect 36636 22568 36688 22574
rect 36636 22510 36688 22516
rect 36556 21690 36584 22510
rect 36544 21684 36596 21690
rect 36544 21626 36596 21632
rect 36648 21321 36676 22510
rect 36820 22092 36872 22098
rect 36820 22034 36872 22040
rect 36832 21418 36860 22034
rect 36924 21978 36952 23462
rect 37002 23423 37058 23432
rect 37096 22976 37148 22982
rect 37096 22918 37148 22924
rect 37108 22094 37136 22918
rect 37200 22438 37228 23598
rect 37280 23520 37332 23526
rect 37280 23462 37332 23468
rect 37292 22642 37320 23462
rect 37476 23186 37504 23598
rect 37464 23180 37516 23186
rect 37464 23122 37516 23128
rect 37476 22642 37504 23122
rect 37280 22636 37332 22642
rect 37280 22578 37332 22584
rect 37464 22636 37516 22642
rect 37464 22578 37516 22584
rect 37188 22432 37240 22438
rect 37188 22374 37240 22380
rect 37108 22066 37228 22094
rect 36924 21950 37044 21978
rect 36912 21888 36964 21894
rect 36912 21830 36964 21836
rect 36820 21412 36872 21418
rect 36820 21354 36872 21360
rect 36634 21312 36690 21321
rect 36634 21247 36690 21256
rect 36648 20806 36676 21247
rect 36636 20800 36688 20806
rect 36636 20742 36688 20748
rect 36544 20528 36596 20534
rect 36542 20496 36544 20505
rect 36596 20496 36598 20505
rect 36542 20431 36598 20440
rect 36648 20346 36676 20742
rect 36728 20528 36780 20534
rect 36728 20470 36780 20476
rect 36452 20324 36504 20330
rect 36452 20266 36504 20272
rect 36556 20318 36676 20346
rect 36452 19916 36504 19922
rect 36452 19858 36504 19864
rect 36360 19780 36412 19786
rect 36360 19722 36412 19728
rect 36084 19372 36136 19378
rect 36084 19314 36136 19320
rect 36176 19372 36228 19378
rect 36464 19334 36492 19858
rect 36176 19314 36228 19320
rect 36188 19224 36216 19314
rect 36372 19306 36492 19334
rect 36188 19196 36308 19224
rect 36280 18834 36308 19196
rect 36084 18828 36136 18834
rect 36084 18770 36136 18776
rect 36268 18828 36320 18834
rect 36268 18770 36320 18776
rect 36096 18601 36124 18770
rect 36176 18760 36228 18766
rect 36176 18702 36228 18708
rect 36082 18592 36138 18601
rect 36082 18527 36138 18536
rect 36096 18306 36124 18527
rect 36188 18426 36216 18702
rect 36176 18420 36228 18426
rect 36176 18362 36228 18368
rect 36096 18278 36216 18306
rect 36188 18154 36216 18278
rect 36266 18184 36322 18193
rect 36176 18148 36228 18154
rect 36266 18119 36322 18128
rect 36176 18090 36228 18096
rect 35992 18080 36044 18086
rect 35992 18022 36044 18028
rect 36004 17882 36032 18022
rect 35992 17876 36044 17882
rect 35992 17818 36044 17824
rect 35900 17808 35952 17814
rect 35900 17750 35952 17756
rect 35808 17740 35860 17746
rect 35808 17682 35860 17688
rect 35992 17740 36044 17746
rect 35992 17682 36044 17688
rect 35808 17604 35860 17610
rect 35808 17546 35860 17552
rect 35714 17368 35770 17377
rect 35532 17332 35584 17338
rect 35714 17303 35770 17312
rect 35532 17274 35584 17280
rect 35532 17196 35584 17202
rect 35532 17138 35584 17144
rect 35544 16794 35572 17138
rect 35716 17128 35768 17134
rect 35820 17105 35848 17546
rect 35716 17070 35768 17076
rect 35806 17096 35862 17105
rect 35532 16788 35584 16794
rect 35532 16730 35584 16736
rect 35624 15904 35676 15910
rect 35624 15846 35676 15852
rect 35532 15360 35584 15366
rect 35438 15328 35494 15337
rect 35532 15302 35584 15308
rect 35438 15263 35494 15272
rect 35348 15156 35400 15162
rect 35348 15098 35400 15104
rect 35346 14104 35402 14113
rect 35346 14039 35348 14048
rect 35400 14039 35402 14048
rect 35348 14010 35400 14016
rect 35348 13796 35400 13802
rect 35348 13738 35400 13744
rect 35256 12776 35308 12782
rect 35256 12718 35308 12724
rect 35360 12646 35388 13738
rect 35452 13258 35480 15263
rect 35544 15065 35572 15302
rect 35530 15056 35586 15065
rect 35530 14991 35586 15000
rect 35636 14958 35664 15846
rect 35532 14952 35584 14958
rect 35532 14894 35584 14900
rect 35624 14952 35676 14958
rect 35624 14894 35676 14900
rect 35440 13252 35492 13258
rect 35440 13194 35492 13200
rect 35348 12640 35400 12646
rect 35348 12582 35400 12588
rect 35544 12434 35572 14894
rect 35636 14346 35664 14894
rect 35728 14482 35756 17070
rect 35806 17031 35862 17040
rect 35900 16992 35952 16998
rect 35900 16934 35952 16940
rect 35808 16516 35860 16522
rect 35808 16458 35860 16464
rect 35820 16182 35848 16458
rect 35808 16176 35860 16182
rect 35808 16118 35860 16124
rect 35820 15910 35848 16118
rect 35808 15904 35860 15910
rect 35808 15846 35860 15852
rect 35808 15564 35860 15570
rect 35808 15506 35860 15512
rect 35820 14793 35848 15506
rect 35912 15314 35940 16934
rect 36004 16017 36032 17682
rect 36176 17536 36228 17542
rect 36176 17478 36228 17484
rect 35990 16008 36046 16017
rect 35990 15943 36046 15952
rect 35912 15286 36124 15314
rect 35992 15156 36044 15162
rect 35992 15098 36044 15104
rect 35900 14816 35952 14822
rect 35806 14784 35862 14793
rect 35900 14758 35952 14764
rect 35806 14719 35862 14728
rect 35716 14476 35768 14482
rect 35716 14418 35768 14424
rect 35624 14340 35676 14346
rect 35624 14282 35676 14288
rect 35624 13388 35676 13394
rect 35624 13330 35676 13336
rect 35360 12406 35572 12434
rect 35360 12102 35388 12406
rect 35440 12164 35492 12170
rect 35440 12106 35492 12112
rect 35348 12096 35400 12102
rect 35348 12038 35400 12044
rect 35072 11348 35124 11354
rect 35072 11290 35124 11296
rect 35164 11348 35216 11354
rect 35164 11290 35216 11296
rect 34980 11280 35032 11286
rect 34980 11222 35032 11228
rect 35176 11150 35204 11290
rect 35256 11212 35308 11218
rect 35256 11154 35308 11160
rect 35164 11144 35216 11150
rect 35268 11121 35296 11154
rect 35164 11086 35216 11092
rect 35254 11112 35310 11121
rect 35254 11047 35310 11056
rect 35072 10804 35124 10810
rect 35072 10746 35124 10752
rect 34980 9920 35032 9926
rect 34980 9862 35032 9868
rect 34796 9648 34848 9654
rect 34796 9590 34848 9596
rect 34888 9580 34940 9586
rect 34888 9522 34940 9528
rect 34900 9178 34928 9522
rect 34888 9172 34940 9178
rect 34888 9114 34940 9120
rect 34704 9104 34756 9110
rect 34704 9046 34756 9052
rect 34992 8838 35020 9862
rect 35084 9654 35112 10746
rect 35452 10742 35480 12106
rect 35636 11642 35664 13330
rect 35728 12866 35756 14418
rect 35912 13870 35940 14758
rect 36004 14006 36032 15098
rect 35992 14000 36044 14006
rect 35992 13942 36044 13948
rect 35900 13864 35952 13870
rect 35900 13806 35952 13812
rect 36004 12918 36032 13942
rect 36096 13841 36124 15286
rect 36188 13938 36216 17478
rect 36280 14822 36308 18119
rect 36372 16833 36400 19306
rect 36452 19236 36504 19242
rect 36556 19224 36584 20318
rect 36740 19961 36768 20470
rect 36820 20324 36872 20330
rect 36820 20266 36872 20272
rect 36726 19952 36782 19961
rect 36726 19887 36782 19896
rect 36636 19848 36688 19854
rect 36688 19796 36768 19802
rect 36636 19790 36768 19796
rect 36648 19774 36768 19790
rect 36636 19712 36688 19718
rect 36636 19654 36688 19660
rect 36504 19196 36584 19224
rect 36452 19178 36504 19184
rect 36450 19136 36506 19145
rect 36450 19071 36506 19080
rect 36464 18465 36492 19071
rect 36450 18456 36506 18465
rect 36648 18426 36676 19654
rect 36740 18737 36768 19774
rect 36726 18728 36782 18737
rect 36832 18698 36860 20266
rect 36726 18663 36782 18672
rect 36820 18692 36872 18698
rect 36820 18634 36872 18640
rect 36728 18624 36780 18630
rect 36728 18566 36780 18572
rect 36740 18426 36768 18566
rect 36818 18456 36874 18465
rect 36450 18391 36506 18400
rect 36636 18420 36688 18426
rect 36636 18362 36688 18368
rect 36728 18420 36780 18426
rect 36818 18391 36874 18400
rect 36728 18362 36780 18368
rect 36728 18284 36780 18290
rect 36728 18226 36780 18232
rect 36450 17912 36506 17921
rect 36450 17847 36506 17856
rect 36464 17814 36492 17847
rect 36452 17808 36504 17814
rect 36452 17750 36504 17756
rect 36358 16824 36414 16833
rect 36358 16759 36414 16768
rect 36360 15496 36412 15502
rect 36360 15438 36412 15444
rect 36372 14890 36400 15438
rect 36464 15178 36492 17750
rect 36740 17649 36768 18226
rect 36832 18154 36860 18391
rect 36820 18148 36872 18154
rect 36820 18090 36872 18096
rect 36924 17785 36952 21830
rect 37016 21162 37044 21950
rect 37200 21350 37228 22066
rect 37280 21956 37332 21962
rect 37280 21898 37332 21904
rect 37292 21486 37320 21898
rect 37476 21486 37504 22578
rect 37280 21480 37332 21486
rect 37280 21422 37332 21428
rect 37464 21480 37516 21486
rect 37464 21422 37516 21428
rect 37188 21344 37240 21350
rect 37188 21286 37240 21292
rect 37016 21134 37228 21162
rect 37096 20800 37148 20806
rect 37096 20742 37148 20748
rect 37108 20602 37136 20742
rect 37096 20596 37148 20602
rect 37096 20538 37148 20544
rect 37004 20460 37056 20466
rect 37004 20402 37056 20408
rect 37016 19961 37044 20402
rect 37200 20262 37228 21134
rect 37476 21010 37504 21422
rect 37464 21004 37516 21010
rect 37464 20946 37516 20952
rect 37476 20777 37504 20946
rect 37462 20768 37518 20777
rect 37462 20703 37518 20712
rect 37278 20632 37334 20641
rect 37278 20567 37334 20576
rect 37096 20256 37148 20262
rect 37096 20198 37148 20204
rect 37188 20256 37240 20262
rect 37188 20198 37240 20204
rect 37002 19952 37058 19961
rect 37002 19887 37058 19896
rect 37004 19780 37056 19786
rect 37004 19722 37056 19728
rect 36910 17776 36966 17785
rect 36910 17711 36966 17720
rect 36726 17640 36782 17649
rect 36726 17575 36782 17584
rect 36820 17604 36872 17610
rect 36820 17546 36872 17552
rect 36544 17196 36596 17202
rect 36544 17138 36596 17144
rect 36556 16969 36584 17138
rect 36832 17134 36860 17546
rect 36636 17128 36688 17134
rect 36820 17128 36872 17134
rect 36636 17070 36688 17076
rect 36740 17088 36820 17116
rect 36542 16960 36598 16969
rect 36542 16895 36598 16904
rect 36648 16454 36676 17070
rect 36636 16448 36688 16454
rect 36636 16390 36688 16396
rect 36648 16046 36676 16390
rect 36636 16040 36688 16046
rect 36636 15982 36688 15988
rect 36464 15150 36676 15178
rect 36452 15020 36504 15026
rect 36452 14962 36504 14968
rect 36360 14884 36412 14890
rect 36360 14826 36412 14832
rect 36268 14816 36320 14822
rect 36268 14758 36320 14764
rect 36266 13968 36322 13977
rect 36176 13932 36228 13938
rect 36266 13903 36322 13912
rect 36176 13874 36228 13880
rect 36082 13832 36138 13841
rect 36082 13767 36138 13776
rect 36174 13560 36230 13569
rect 36174 13495 36230 13504
rect 36188 13394 36216 13495
rect 36176 13388 36228 13394
rect 36176 13330 36228 13336
rect 36176 13184 36228 13190
rect 36176 13126 36228 13132
rect 35992 12912 36044 12918
rect 35728 12838 35848 12866
rect 35992 12854 36044 12860
rect 35716 12776 35768 12782
rect 35716 12718 35768 12724
rect 35728 12306 35756 12718
rect 35820 12424 35848 12838
rect 36188 12481 36216 13126
rect 36174 12472 36230 12481
rect 35820 12396 35940 12424
rect 36174 12407 36230 12416
rect 35716 12300 35768 12306
rect 35716 12242 35768 12248
rect 35808 12300 35860 12306
rect 35808 12242 35860 12248
rect 35544 11614 35664 11642
rect 35728 11626 35756 12242
rect 35820 12102 35848 12242
rect 35808 12096 35860 12102
rect 35808 12038 35860 12044
rect 35808 11756 35860 11762
rect 35808 11698 35860 11704
rect 35716 11620 35768 11626
rect 35544 10810 35572 11614
rect 35716 11562 35768 11568
rect 35624 11552 35676 11558
rect 35624 11494 35676 11500
rect 35532 10804 35584 10810
rect 35532 10746 35584 10752
rect 35440 10736 35492 10742
rect 35440 10678 35492 10684
rect 35348 10532 35400 10538
rect 35348 10474 35400 10480
rect 35072 9648 35124 9654
rect 35072 9590 35124 9596
rect 35072 9512 35124 9518
rect 35072 9454 35124 9460
rect 35162 9480 35218 9489
rect 34980 8832 35032 8838
rect 34980 8774 35032 8780
rect 35084 8616 35112 9454
rect 35162 9415 35218 9424
rect 35176 9042 35204 9415
rect 35256 9104 35308 9110
rect 35256 9046 35308 9052
rect 35164 9036 35216 9042
rect 35164 8978 35216 8984
rect 34900 8588 35112 8616
rect 34900 8294 34928 8588
rect 34888 8288 34940 8294
rect 34888 8230 34940 8236
rect 34900 7886 34928 8230
rect 34572 7840 34652 7868
rect 34888 7880 34940 7886
rect 34520 7822 34572 7828
rect 34888 7822 34940 7828
rect 34428 7744 34480 7750
rect 34428 7686 34480 7692
rect 34532 7546 34560 7822
rect 34520 7540 34572 7546
rect 34520 7482 34572 7488
rect 34888 7200 34940 7206
rect 34888 7142 34940 7148
rect 34900 6798 34928 7142
rect 34888 6792 34940 6798
rect 34888 6734 34940 6740
rect 34336 6384 34388 6390
rect 34336 6326 34388 6332
rect 35176 5273 35204 8978
rect 35268 8838 35296 9046
rect 35256 8832 35308 8838
rect 35256 8774 35308 8780
rect 35360 8566 35388 10474
rect 35544 9908 35572 10746
rect 35452 9880 35572 9908
rect 35348 8560 35400 8566
rect 35348 8502 35400 8508
rect 35452 8430 35480 9880
rect 35532 9512 35584 9518
rect 35530 9480 35532 9489
rect 35584 9480 35586 9489
rect 35530 9415 35586 9424
rect 35636 9110 35664 11494
rect 35728 11218 35756 11562
rect 35820 11257 35848 11698
rect 35912 11694 35940 12396
rect 35992 12096 36044 12102
rect 36188 12073 36216 12407
rect 35992 12038 36044 12044
rect 36174 12064 36230 12073
rect 36004 11830 36032 12038
rect 36174 11999 36230 12008
rect 35992 11824 36044 11830
rect 35992 11766 36044 11772
rect 35900 11688 35952 11694
rect 36280 11676 36308 13903
rect 36360 13456 36412 13462
rect 36360 13398 36412 13404
rect 35900 11630 35952 11636
rect 36004 11648 36308 11676
rect 36004 11354 36032 11648
rect 35992 11348 36044 11354
rect 35992 11290 36044 11296
rect 35806 11248 35862 11257
rect 35716 11212 35768 11218
rect 35806 11183 35862 11192
rect 36082 11248 36138 11257
rect 36082 11183 36138 11192
rect 35716 11154 35768 11160
rect 35808 11144 35860 11150
rect 35808 11086 35860 11092
rect 35716 9444 35768 9450
rect 35716 9386 35768 9392
rect 35624 9104 35676 9110
rect 35624 9046 35676 9052
rect 35532 9036 35584 9042
rect 35532 8978 35584 8984
rect 35440 8424 35492 8430
rect 35440 8366 35492 8372
rect 35544 7410 35572 8978
rect 35624 8968 35676 8974
rect 35624 8910 35676 8916
rect 35636 7954 35664 8910
rect 35624 7948 35676 7954
rect 35624 7890 35676 7896
rect 35728 7410 35756 9386
rect 35820 8974 35848 11086
rect 35900 9580 35952 9586
rect 35900 9522 35952 9528
rect 35912 9489 35940 9522
rect 35898 9480 35954 9489
rect 35898 9415 35954 9424
rect 35992 9376 36044 9382
rect 35992 9318 36044 9324
rect 35808 8968 35860 8974
rect 35808 8910 35860 8916
rect 35898 8936 35954 8945
rect 35898 8871 35954 8880
rect 35808 8356 35860 8362
rect 35808 8298 35860 8304
rect 35820 7478 35848 8298
rect 35912 8294 35940 8871
rect 35900 8288 35952 8294
rect 35900 8230 35952 8236
rect 35898 8120 35954 8129
rect 36004 8090 36032 9318
rect 36096 9058 36124 11183
rect 36176 11008 36228 11014
rect 36176 10950 36228 10956
rect 36188 10674 36216 10950
rect 36176 10668 36228 10674
rect 36176 10610 36228 10616
rect 36188 9994 36216 10610
rect 36268 10600 36320 10606
rect 36268 10542 36320 10548
rect 36176 9988 36228 9994
rect 36176 9930 36228 9936
rect 36096 9030 36216 9058
rect 36084 8968 36136 8974
rect 36084 8910 36136 8916
rect 35898 8055 35900 8064
rect 35952 8055 35954 8064
rect 35992 8084 36044 8090
rect 35900 8026 35952 8032
rect 35992 8026 36044 8032
rect 35808 7472 35860 7478
rect 35808 7414 35860 7420
rect 35532 7404 35584 7410
rect 35532 7346 35584 7352
rect 35716 7404 35768 7410
rect 35716 7346 35768 7352
rect 35808 7268 35860 7274
rect 35808 7210 35860 7216
rect 35624 6860 35676 6866
rect 35624 6802 35676 6808
rect 35636 6497 35664 6802
rect 35820 6769 35848 7210
rect 35806 6760 35862 6769
rect 36096 6730 36124 8910
rect 36188 7818 36216 9030
rect 36280 8498 36308 10542
rect 36372 9674 36400 13398
rect 36464 12238 36492 14962
rect 36544 12640 36596 12646
rect 36544 12582 36596 12588
rect 36452 12232 36504 12238
rect 36452 12174 36504 12180
rect 36556 12170 36584 12582
rect 36544 12164 36596 12170
rect 36544 12106 36596 12112
rect 36450 12064 36506 12073
rect 36450 11999 36506 12008
rect 36464 10690 36492 11999
rect 36556 11694 36584 12106
rect 36544 11688 36596 11694
rect 36544 11630 36596 11636
rect 36556 11014 36584 11630
rect 36544 11008 36596 11014
rect 36544 10950 36596 10956
rect 36648 10810 36676 15150
rect 36740 12782 36768 17088
rect 36820 17070 36872 17076
rect 36910 16960 36966 16969
rect 36910 16895 36966 16904
rect 36818 16416 36874 16425
rect 36818 16351 36874 16360
rect 36832 16114 36860 16351
rect 36820 16108 36872 16114
rect 36820 16050 36872 16056
rect 36818 16008 36874 16017
rect 36818 15943 36820 15952
rect 36872 15943 36874 15952
rect 36820 15914 36872 15920
rect 36820 15360 36872 15366
rect 36820 15302 36872 15308
rect 36832 14958 36860 15302
rect 36820 14952 36872 14958
rect 36820 14894 36872 14900
rect 36820 14476 36872 14482
rect 36820 14418 36872 14424
rect 36832 14006 36860 14418
rect 36820 14000 36872 14006
rect 36820 13942 36872 13948
rect 36832 13394 36860 13942
rect 36820 13388 36872 13394
rect 36820 13330 36872 13336
rect 36832 12850 36860 13330
rect 36924 12918 36952 16895
rect 37016 16289 37044 19722
rect 37002 16280 37058 16289
rect 37002 16215 37058 16224
rect 37004 15972 37056 15978
rect 37004 15914 37056 15920
rect 37016 15450 37044 15914
rect 37108 15638 37136 20198
rect 37200 19553 37228 20198
rect 37186 19544 37242 19553
rect 37186 19479 37242 19488
rect 37200 17116 37228 19479
rect 37292 18737 37320 20567
rect 37476 20466 37504 20703
rect 37568 20602 37596 24618
rect 37660 23497 37688 26200
rect 38304 26081 38332 26200
rect 38290 26072 38346 26081
rect 38290 26007 38346 26016
rect 37830 24984 37886 24993
rect 37830 24919 37886 24928
rect 37738 23896 37794 23905
rect 37844 23866 37872 24919
rect 38660 24268 38712 24274
rect 38660 24210 38712 24216
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 38382 23896 38438 23905
rect 37738 23831 37794 23840
rect 37832 23860 37884 23866
rect 37752 23746 37780 23831
rect 37832 23802 37884 23808
rect 37924 23860 37976 23866
rect 38382 23831 38438 23840
rect 37924 23802 37976 23808
rect 37936 23746 37964 23802
rect 37752 23718 37964 23746
rect 37646 23488 37702 23497
rect 37646 23423 37702 23432
rect 38396 22982 38424 23831
rect 38566 23352 38622 23361
rect 38566 23287 38622 23296
rect 38384 22976 38436 22982
rect 38384 22918 38436 22924
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 37740 22568 37792 22574
rect 37740 22510 37792 22516
rect 38476 22568 38528 22574
rect 38476 22510 38528 22516
rect 37752 22409 37780 22510
rect 37738 22400 37794 22409
rect 37738 22335 37794 22344
rect 38488 22234 38516 22510
rect 38476 22228 38528 22234
rect 38476 22170 38528 22176
rect 38106 21992 38162 22001
rect 37752 21950 37964 21978
rect 37752 21729 37780 21950
rect 37936 21894 37964 21950
rect 38580 21978 38608 23287
rect 38672 23254 38700 24210
rect 38844 23724 38896 23730
rect 38844 23666 38896 23672
rect 38660 23248 38712 23254
rect 38660 23190 38712 23196
rect 38856 23118 38884 23666
rect 38948 23497 38976 26200
rect 38934 23488 38990 23497
rect 38934 23423 38990 23432
rect 38844 23112 38896 23118
rect 38844 23054 38896 23060
rect 38934 23080 38990 23089
rect 38660 23044 38712 23050
rect 38660 22986 38712 22992
rect 38672 22681 38700 22986
rect 38750 22944 38806 22953
rect 38750 22879 38806 22888
rect 38658 22672 38714 22681
rect 38658 22607 38714 22616
rect 38660 22092 38712 22098
rect 38660 22034 38712 22040
rect 38162 21950 38608 21978
rect 38106 21927 38162 21936
rect 37832 21888 37884 21894
rect 37832 21830 37884 21836
rect 37924 21888 37976 21894
rect 37924 21830 37976 21836
rect 38382 21856 38438 21865
rect 37738 21720 37794 21729
rect 37844 21690 37872 21830
rect 37950 21788 38258 21797
rect 38382 21791 38438 21800
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 37738 21655 37794 21664
rect 37832 21684 37884 21690
rect 37832 21626 37884 21632
rect 37830 21584 37886 21593
rect 37648 21548 37700 21554
rect 37830 21519 37832 21528
rect 37648 21490 37700 21496
rect 37884 21519 37886 21528
rect 37832 21490 37884 21496
rect 37660 21457 37688 21490
rect 37646 21448 37702 21457
rect 37646 21383 37702 21392
rect 37844 21049 37872 21490
rect 37830 21040 37886 21049
rect 37830 20975 37886 20984
rect 38292 20868 38344 20874
rect 38396 20856 38424 21791
rect 38476 21616 38528 21622
rect 38568 21616 38620 21622
rect 38476 21558 38528 21564
rect 38566 21584 38568 21593
rect 38620 21584 38622 21593
rect 38488 21468 38516 21558
rect 38566 21519 38622 21528
rect 38568 21480 38620 21486
rect 38488 21440 38568 21468
rect 38568 21422 38620 21428
rect 38344 20828 38424 20856
rect 38292 20810 38344 20816
rect 38672 20806 38700 22034
rect 38764 21010 38792 22879
rect 38856 22642 38884 23054
rect 38934 23015 38990 23024
rect 38948 22982 38976 23015
rect 38936 22976 38988 22982
rect 38936 22918 38988 22924
rect 39028 22704 39080 22710
rect 39028 22646 39080 22652
rect 38844 22636 38896 22642
rect 38896 22596 38976 22624
rect 38844 22578 38896 22584
rect 38844 22160 38896 22166
rect 38842 22128 38844 22137
rect 38896 22128 38898 22137
rect 38842 22063 38898 22072
rect 38844 21888 38896 21894
rect 38844 21830 38896 21836
rect 38752 21004 38804 21010
rect 38752 20946 38804 20952
rect 38660 20800 38712 20806
rect 38660 20742 38712 20748
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 38474 20632 38530 20641
rect 37556 20596 37608 20602
rect 38474 20567 38530 20576
rect 37556 20538 37608 20544
rect 37464 20460 37516 20466
rect 37464 20402 37516 20408
rect 37832 20460 37884 20466
rect 37832 20402 37884 20408
rect 37648 20256 37700 20262
rect 37648 20198 37700 20204
rect 37740 20256 37792 20262
rect 37740 20198 37792 20204
rect 37372 19780 37424 19786
rect 37372 19722 37424 19728
rect 37384 19378 37412 19722
rect 37660 19417 37688 20198
rect 37752 20058 37780 20198
rect 37740 20052 37792 20058
rect 37740 19994 37792 20000
rect 37646 19408 37702 19417
rect 37359 19372 37412 19378
rect 37411 19320 37412 19372
rect 37359 19314 37412 19320
rect 37464 19372 37516 19378
rect 37844 19378 37872 20402
rect 38382 20224 38438 20233
rect 38382 20159 38438 20168
rect 38292 19780 38344 19786
rect 38292 19722 38344 19728
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 38198 19408 38254 19417
rect 37646 19343 37702 19352
rect 37832 19372 37884 19378
rect 37516 19320 37596 19334
rect 37464 19314 37596 19320
rect 37278 18728 37334 18737
rect 37278 18663 37334 18672
rect 37280 18284 37332 18290
rect 37280 18226 37332 18232
rect 37292 17270 37320 18226
rect 37280 17264 37332 17270
rect 37280 17206 37332 17212
rect 37200 17088 37320 17116
rect 37096 15632 37148 15638
rect 37292 15586 37320 17088
rect 37096 15574 37148 15580
rect 37200 15558 37320 15586
rect 37016 15422 37136 15450
rect 37004 15360 37056 15366
rect 37004 15302 37056 15308
rect 37016 14929 37044 15302
rect 37108 15026 37136 15422
rect 37096 15020 37148 15026
rect 37096 14962 37148 14968
rect 37002 14920 37058 14929
rect 37002 14855 37058 14864
rect 37096 13864 37148 13870
rect 37096 13806 37148 13812
rect 36912 12912 36964 12918
rect 36912 12854 36964 12860
rect 36820 12844 36872 12850
rect 36820 12786 36872 12792
rect 36728 12776 36780 12782
rect 36728 12718 36780 12724
rect 36924 11898 36952 12854
rect 37108 12434 37136 13806
rect 37200 13682 37228 15558
rect 37280 15428 37332 15434
rect 37280 15370 37332 15376
rect 37292 13802 37320 15370
rect 37384 15162 37412 19314
rect 37476 19306 37596 19314
rect 37464 18080 37516 18086
rect 37464 18022 37516 18028
rect 37476 17202 37504 18022
rect 37568 17338 37596 19306
rect 37660 18057 37688 19343
rect 38198 19343 38254 19352
rect 37832 19314 37884 19320
rect 38212 19174 38240 19343
rect 38200 19168 38252 19174
rect 38200 19110 38252 19116
rect 37832 18692 37884 18698
rect 37832 18634 37884 18640
rect 37844 18358 37872 18634
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 37832 18352 37884 18358
rect 37884 18312 38056 18340
rect 37832 18294 37884 18300
rect 37646 18048 37702 18057
rect 37646 17983 37702 17992
rect 37924 17876 37976 17882
rect 37924 17818 37976 17824
rect 37936 17626 37964 17818
rect 38028 17678 38056 18312
rect 38304 18222 38332 19722
rect 38396 19417 38424 20159
rect 38488 19922 38516 20567
rect 38856 20380 38884 21830
rect 38948 20534 38976 22596
rect 39040 22234 39068 22646
rect 39028 22228 39080 22234
rect 39028 22170 39080 22176
rect 39212 22160 39264 22166
rect 39212 22102 39264 22108
rect 39028 21480 39080 21486
rect 39028 21422 39080 21428
rect 39120 21480 39172 21486
rect 39120 21422 39172 21428
rect 39040 21010 39068 21422
rect 39028 21004 39080 21010
rect 39028 20946 39080 20952
rect 39132 20942 39160 21422
rect 39120 20936 39172 20942
rect 39120 20878 39172 20884
rect 38936 20528 38988 20534
rect 38988 20488 39160 20516
rect 38936 20470 38988 20476
rect 38856 20352 39068 20380
rect 38750 20224 38806 20233
rect 38750 20159 38806 20168
rect 38568 20052 38620 20058
rect 38568 19994 38620 20000
rect 38476 19916 38528 19922
rect 38476 19858 38528 19864
rect 38474 19816 38530 19825
rect 38474 19751 38530 19760
rect 38382 19408 38438 19417
rect 38382 19343 38438 19352
rect 38292 18216 38344 18222
rect 38292 18158 38344 18164
rect 38304 17746 38332 18158
rect 38488 17814 38516 19751
rect 38580 18902 38608 19994
rect 38764 19972 38792 20159
rect 38672 19944 38792 19972
rect 38672 19854 38700 19944
rect 38660 19848 38712 19854
rect 38660 19790 38712 19796
rect 38752 19712 38804 19718
rect 38752 19654 38804 19660
rect 38568 18896 38620 18902
rect 38568 18838 38620 18844
rect 38764 18834 38792 19654
rect 38752 18828 38804 18834
rect 38752 18770 38804 18776
rect 38660 18760 38712 18766
rect 38660 18702 38712 18708
rect 38672 18426 38700 18702
rect 38752 18624 38804 18630
rect 38750 18592 38752 18601
rect 38844 18624 38896 18630
rect 38804 18592 38806 18601
rect 38844 18566 38896 18572
rect 38936 18624 38988 18630
rect 38936 18566 38988 18572
rect 38750 18527 38806 18536
rect 38660 18420 38712 18426
rect 38660 18362 38712 18368
rect 38476 17808 38528 17814
rect 38476 17750 38528 17756
rect 38568 17808 38620 17814
rect 38568 17750 38620 17756
rect 38292 17740 38344 17746
rect 38292 17682 38344 17688
rect 38384 17740 38436 17746
rect 38384 17682 38436 17688
rect 37752 17598 37964 17626
rect 38016 17672 38068 17678
rect 38016 17614 38068 17620
rect 37556 17332 37608 17338
rect 37556 17274 37608 17280
rect 37464 17196 37516 17202
rect 37464 17138 37516 17144
rect 37648 17060 37700 17066
rect 37648 17002 37700 17008
rect 37462 16688 37518 16697
rect 37462 16623 37518 16632
rect 37476 15745 37504 16623
rect 37462 15736 37518 15745
rect 37462 15671 37518 15680
rect 37464 15496 37516 15502
rect 37464 15438 37516 15444
rect 37372 15156 37424 15162
rect 37372 15098 37424 15104
rect 37476 15026 37504 15438
rect 37464 15020 37516 15026
rect 37464 14962 37516 14968
rect 37476 14482 37504 14962
rect 37556 14952 37608 14958
rect 37556 14894 37608 14900
rect 37464 14476 37516 14482
rect 37464 14418 37516 14424
rect 37372 14340 37424 14346
rect 37372 14282 37424 14288
rect 37280 13796 37332 13802
rect 37280 13738 37332 13744
rect 37200 13654 37320 13682
rect 37292 13394 37320 13654
rect 37384 13569 37412 14282
rect 37370 13560 37426 13569
rect 37370 13495 37426 13504
rect 37280 13388 37332 13394
rect 37280 13330 37332 13336
rect 37568 13274 37596 14894
rect 37292 13246 37596 13274
rect 37108 12406 37228 12434
rect 37200 12374 37228 12406
rect 37188 12368 37240 12374
rect 37002 12336 37058 12345
rect 37188 12310 37240 12316
rect 37002 12271 37058 12280
rect 36912 11892 36964 11898
rect 36912 11834 36964 11840
rect 36910 11112 36966 11121
rect 36910 11047 36966 11056
rect 36726 10976 36782 10985
rect 36726 10911 36782 10920
rect 36636 10804 36688 10810
rect 36636 10746 36688 10752
rect 36464 10662 36676 10690
rect 36648 10606 36676 10662
rect 36544 10600 36596 10606
rect 36544 10542 36596 10548
rect 36636 10600 36688 10606
rect 36636 10542 36688 10548
rect 36556 10441 36584 10542
rect 36542 10432 36598 10441
rect 36542 10367 36598 10376
rect 36648 10266 36676 10542
rect 36452 10260 36504 10266
rect 36636 10260 36688 10266
rect 36452 10202 36504 10208
rect 36556 10220 36636 10248
rect 36464 10062 36492 10202
rect 36452 10056 36504 10062
rect 36452 9998 36504 10004
rect 36372 9654 36492 9674
rect 36372 9648 36504 9654
rect 36372 9646 36452 9648
rect 36452 9590 36504 9596
rect 36360 9580 36412 9586
rect 36360 9522 36412 9528
rect 36372 8634 36400 9522
rect 36556 9178 36584 10220
rect 36636 10202 36688 10208
rect 36636 9920 36688 9926
rect 36634 9888 36636 9897
rect 36688 9888 36690 9897
rect 36634 9823 36690 9832
rect 36648 9586 36676 9823
rect 36636 9580 36688 9586
rect 36636 9522 36688 9528
rect 36544 9172 36596 9178
rect 36544 9114 36596 9120
rect 36636 9104 36688 9110
rect 36636 9046 36688 9052
rect 36452 8968 36504 8974
rect 36452 8910 36504 8916
rect 36360 8628 36412 8634
rect 36360 8570 36412 8576
rect 36268 8492 36320 8498
rect 36268 8434 36320 8440
rect 36176 7812 36228 7818
rect 36176 7754 36228 7760
rect 35806 6695 35862 6704
rect 36084 6724 36136 6730
rect 36084 6666 36136 6672
rect 35622 6488 35678 6497
rect 35622 6423 35678 6432
rect 35898 5944 35954 5953
rect 35898 5879 35954 5888
rect 35162 5264 35218 5273
rect 35162 5199 35218 5208
rect 35912 5098 35940 5879
rect 36464 5710 36492 8910
rect 36648 8566 36676 9046
rect 36740 8945 36768 10911
rect 36924 10674 36952 11047
rect 37016 10962 37044 12271
rect 37188 11688 37240 11694
rect 37188 11630 37240 11636
rect 37200 11098 37228 11630
rect 37292 11268 37320 13246
rect 37372 12708 37424 12714
rect 37372 12650 37424 12656
rect 37384 11393 37412 12650
rect 37556 12300 37608 12306
rect 37556 12242 37608 12248
rect 37464 12096 37516 12102
rect 37464 12038 37516 12044
rect 37476 11937 37504 12038
rect 37462 11928 37518 11937
rect 37462 11863 37518 11872
rect 37370 11384 37426 11393
rect 37370 11319 37426 11328
rect 37292 11240 37412 11268
rect 37476 11257 37504 11863
rect 37568 11286 37596 12242
rect 37660 11642 37688 17002
rect 37752 16522 37780 17598
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 38200 17332 38252 17338
rect 38200 17274 38252 17280
rect 38212 17082 38240 17274
rect 38304 17202 38332 17682
rect 38292 17196 38344 17202
rect 38292 17138 38344 17144
rect 38120 17054 38240 17082
rect 38120 16794 38148 17054
rect 38200 16992 38252 16998
rect 38200 16934 38252 16940
rect 38108 16788 38160 16794
rect 38108 16730 38160 16736
rect 38212 16726 38240 16934
rect 38200 16720 38252 16726
rect 38200 16662 38252 16668
rect 37740 16516 37792 16522
rect 37740 16458 37792 16464
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 38304 16114 38332 17138
rect 38396 17134 38424 17682
rect 38580 17626 38608 17750
rect 38488 17598 38608 17626
rect 38488 17542 38516 17598
rect 38476 17536 38528 17542
rect 38476 17478 38528 17484
rect 38384 17128 38436 17134
rect 38384 17070 38436 17076
rect 38384 16448 38436 16454
rect 38384 16390 38436 16396
rect 38292 16108 38344 16114
rect 38292 16050 38344 16056
rect 37740 15904 37792 15910
rect 37740 15846 37792 15852
rect 37752 12345 37780 15846
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 37832 15088 37884 15094
rect 37832 15030 37884 15036
rect 38198 15056 38254 15065
rect 37844 14822 37872 15030
rect 38198 14991 38254 15000
rect 37832 14816 37884 14822
rect 37832 14758 37884 14764
rect 38212 14532 38240 14991
rect 38396 14958 38424 16390
rect 38488 16182 38516 17478
rect 38750 17368 38806 17377
rect 38856 17338 38884 18566
rect 38948 18426 38976 18566
rect 38936 18420 38988 18426
rect 38936 18362 38988 18368
rect 39040 17728 39068 20352
rect 39132 19961 39160 20488
rect 39118 19952 39174 19961
rect 39118 19887 39174 19896
rect 39132 19446 39160 19887
rect 39120 19440 39172 19446
rect 39120 19382 39172 19388
rect 39118 18592 39174 18601
rect 39118 18527 39174 18536
rect 39132 18358 39160 18527
rect 39120 18352 39172 18358
rect 39120 18294 39172 18300
rect 38948 17700 39068 17728
rect 38948 17513 38976 17700
rect 39224 17626 39252 22102
rect 39040 17598 39252 17626
rect 38934 17504 38990 17513
rect 38934 17439 38990 17448
rect 38750 17303 38806 17312
rect 38844 17332 38896 17338
rect 38764 16794 38792 17303
rect 38844 17274 38896 17280
rect 38752 16788 38804 16794
rect 38752 16730 38804 16736
rect 38568 16720 38620 16726
rect 38568 16662 38620 16668
rect 38580 16182 38608 16662
rect 38844 16652 38896 16658
rect 38844 16594 38896 16600
rect 38658 16552 38714 16561
rect 38658 16487 38714 16496
rect 38672 16454 38700 16487
rect 38660 16448 38712 16454
rect 38660 16390 38712 16396
rect 38752 16448 38804 16454
rect 38856 16425 38884 16594
rect 38752 16390 38804 16396
rect 38842 16416 38898 16425
rect 38764 16266 38792 16390
rect 38842 16351 38898 16360
rect 38948 16266 38976 17439
rect 39040 17338 39068 17598
rect 39224 17542 39252 17598
rect 39120 17536 39172 17542
rect 39120 17478 39172 17484
rect 39212 17536 39264 17542
rect 39212 17478 39264 17484
rect 39132 17338 39160 17478
rect 39028 17332 39080 17338
rect 39028 17274 39080 17280
rect 39120 17332 39172 17338
rect 39120 17274 39172 17280
rect 39316 17218 39344 26302
rect 39578 26200 39634 26302
rect 40222 26200 40278 27000
rect 40958 26752 41014 26761
rect 40958 26687 41014 26696
rect 39946 24440 40002 24449
rect 39946 24375 40002 24384
rect 39960 24342 39988 24375
rect 39948 24336 40000 24342
rect 39948 24278 40000 24284
rect 39396 24268 39448 24274
rect 39396 24210 39448 24216
rect 39408 24154 39436 24210
rect 39672 24200 39724 24206
rect 39408 24126 39620 24154
rect 39672 24142 39724 24148
rect 39592 23202 39620 24126
rect 39408 23174 39620 23202
rect 39408 22710 39436 23174
rect 39488 23112 39540 23118
rect 39488 23054 39540 23060
rect 39396 22704 39448 22710
rect 39396 22646 39448 22652
rect 39396 22432 39448 22438
rect 39396 22374 39448 22380
rect 39408 22234 39436 22374
rect 39396 22228 39448 22234
rect 39396 22170 39448 22176
rect 39396 21888 39448 21894
rect 39396 21830 39448 21836
rect 39408 20913 39436 21830
rect 39394 20904 39450 20913
rect 39394 20839 39450 20848
rect 39394 20632 39450 20641
rect 39394 20567 39450 20576
rect 39408 20330 39436 20567
rect 39396 20324 39448 20330
rect 39396 20266 39448 20272
rect 39500 18193 39528 23054
rect 39592 22234 39620 23174
rect 39684 22778 39712 24142
rect 39948 23724 40000 23730
rect 39948 23666 40000 23672
rect 39856 23656 39908 23662
rect 39856 23598 39908 23604
rect 39764 23248 39816 23254
rect 39764 23190 39816 23196
rect 39672 22772 39724 22778
rect 39672 22714 39724 22720
rect 39580 22228 39632 22234
rect 39580 22170 39632 22176
rect 39578 21040 39634 21049
rect 39578 20975 39634 20984
rect 39592 19281 39620 20975
rect 39776 20890 39804 23190
rect 39868 22098 39896 23598
rect 39960 22681 39988 23666
rect 40040 23112 40092 23118
rect 40040 23054 40092 23060
rect 39946 22672 40002 22681
rect 39946 22607 40002 22616
rect 40052 22545 40080 23054
rect 40132 22704 40184 22710
rect 40132 22646 40184 22652
rect 40038 22536 40094 22545
rect 40038 22471 40094 22480
rect 39856 22092 39908 22098
rect 39856 22034 39908 22040
rect 40040 21888 40092 21894
rect 40040 21830 40092 21836
rect 40052 21622 40080 21830
rect 40040 21616 40092 21622
rect 40040 21558 40092 21564
rect 39948 21548 40000 21554
rect 39948 21490 40000 21496
rect 39960 21418 39988 21490
rect 39948 21412 40000 21418
rect 39948 21354 40000 21360
rect 40144 21146 40172 22646
rect 40132 21140 40184 21146
rect 40132 21082 40184 21088
rect 39684 20862 39804 20890
rect 39684 20466 39712 20862
rect 39764 20800 39816 20806
rect 39764 20742 39816 20748
rect 39672 20460 39724 20466
rect 39672 20402 39724 20408
rect 39672 19916 39724 19922
rect 39672 19858 39724 19864
rect 39578 19272 39634 19281
rect 39578 19207 39634 19216
rect 39592 18902 39620 19207
rect 39684 18902 39712 19858
rect 39580 18896 39632 18902
rect 39580 18838 39632 18844
rect 39672 18896 39724 18902
rect 39672 18838 39724 18844
rect 39486 18184 39542 18193
rect 39486 18119 39542 18128
rect 39684 17814 39712 18838
rect 39776 18766 39804 20742
rect 40236 20641 40264 26200
rect 40868 25832 40920 25838
rect 40868 25774 40920 25780
rect 40316 25288 40368 25294
rect 40316 25230 40368 25236
rect 40328 23118 40356 25230
rect 40684 24676 40736 24682
rect 40684 24618 40736 24624
rect 40696 24410 40724 24618
rect 40684 24404 40736 24410
rect 40684 24346 40736 24352
rect 40696 24274 40724 24346
rect 40684 24268 40736 24274
rect 40684 24210 40736 24216
rect 40408 24064 40460 24070
rect 40408 24006 40460 24012
rect 40420 23497 40448 24006
rect 40684 23656 40736 23662
rect 40684 23598 40736 23604
rect 40776 23656 40828 23662
rect 40776 23598 40828 23604
rect 40406 23488 40462 23497
rect 40406 23423 40462 23432
rect 40408 23248 40460 23254
rect 40696 23225 40724 23598
rect 40788 23526 40816 23598
rect 40776 23520 40828 23526
rect 40776 23462 40828 23468
rect 40880 23338 40908 25774
rect 40788 23310 40908 23338
rect 40408 23190 40460 23196
rect 40682 23216 40738 23225
rect 40316 23112 40368 23118
rect 40316 23054 40368 23060
rect 40316 22568 40368 22574
rect 40316 22510 40368 22516
rect 40328 22409 40356 22510
rect 40314 22400 40370 22409
rect 40420 22386 40448 23190
rect 40682 23151 40738 23160
rect 40498 23080 40554 23089
rect 40498 23015 40554 23024
rect 40512 22642 40540 23015
rect 40696 22817 40724 23151
rect 40682 22808 40738 22817
rect 40682 22743 40738 22752
rect 40500 22636 40552 22642
rect 40500 22578 40552 22584
rect 40684 22568 40736 22574
rect 40684 22510 40736 22516
rect 40420 22358 40540 22386
rect 40314 22335 40370 22344
rect 40406 22128 40462 22137
rect 40406 22063 40462 22072
rect 40512 22094 40540 22358
rect 40512 22066 40632 22094
rect 40420 21962 40448 22063
rect 40316 21956 40368 21962
rect 40316 21898 40368 21904
rect 40408 21956 40460 21962
rect 40408 21898 40460 21904
rect 40328 21536 40356 21898
rect 40500 21888 40552 21894
rect 40500 21830 40552 21836
rect 40512 21729 40540 21830
rect 40498 21720 40554 21729
rect 40498 21655 40554 21664
rect 40408 21548 40460 21554
rect 40328 21508 40408 21536
rect 40408 21490 40460 21496
rect 40222 20632 40278 20641
rect 40420 20618 40448 21490
rect 40512 20913 40540 21655
rect 40498 20904 40554 20913
rect 40498 20839 40554 20848
rect 40420 20590 40540 20618
rect 40222 20567 40278 20576
rect 40316 20528 40368 20534
rect 40316 20470 40368 20476
rect 40406 20496 40462 20505
rect 40132 20460 40184 20466
rect 40132 20402 40184 20408
rect 40040 20256 40092 20262
rect 39854 20224 39910 20233
rect 39854 20159 39910 20168
rect 40038 20224 40040 20233
rect 40092 20224 40094 20233
rect 40038 20159 40094 20168
rect 39868 20058 39896 20159
rect 39856 20052 39908 20058
rect 39856 19994 39908 20000
rect 39854 19952 39910 19961
rect 39854 19887 39910 19896
rect 39868 19334 39896 19887
rect 40144 19666 40172 20402
rect 40328 20398 40356 20470
rect 40406 20431 40462 20440
rect 40420 20398 40448 20431
rect 40316 20392 40368 20398
rect 40316 20334 40368 20340
rect 40408 20392 40460 20398
rect 40408 20334 40460 20340
rect 40224 20256 40276 20262
rect 40224 20198 40276 20204
rect 40316 20256 40368 20262
rect 40512 20244 40540 20590
rect 40604 20262 40632 22066
rect 40316 20198 40368 20204
rect 40420 20216 40540 20244
rect 40592 20256 40644 20262
rect 40236 19854 40264 20198
rect 40328 19854 40356 20198
rect 40224 19848 40276 19854
rect 40224 19790 40276 19796
rect 40316 19848 40368 19854
rect 40316 19790 40368 19796
rect 40420 19718 40448 20216
rect 40592 20198 40644 20204
rect 40590 19952 40646 19961
rect 40590 19887 40646 19896
rect 40498 19816 40554 19825
rect 40498 19751 40554 19760
rect 40316 19712 40368 19718
rect 40144 19638 40264 19666
rect 40316 19654 40368 19660
rect 40408 19712 40460 19718
rect 40408 19654 40460 19660
rect 40236 19378 40264 19638
rect 40224 19372 40276 19378
rect 39868 19306 39988 19334
rect 40224 19314 40276 19320
rect 40328 19310 40356 19654
rect 40512 19514 40540 19751
rect 40604 19718 40632 19887
rect 40592 19712 40644 19718
rect 40592 19654 40644 19660
rect 40500 19508 40552 19514
rect 40500 19450 40552 19456
rect 40408 19372 40460 19378
rect 40408 19314 40460 19320
rect 39856 18828 39908 18834
rect 39856 18770 39908 18776
rect 39764 18760 39816 18766
rect 39764 18702 39816 18708
rect 39672 17808 39724 17814
rect 39672 17750 39724 17756
rect 39396 17604 39448 17610
rect 39396 17546 39448 17552
rect 38764 16238 38976 16266
rect 39040 17190 39344 17218
rect 38476 16176 38528 16182
rect 38476 16118 38528 16124
rect 38568 16176 38620 16182
rect 38568 16118 38620 16124
rect 38474 15464 38530 15473
rect 38474 15399 38530 15408
rect 38292 14952 38344 14958
rect 38292 14894 38344 14900
rect 38384 14952 38436 14958
rect 38384 14894 38436 14900
rect 38304 14657 38332 14894
rect 38290 14648 38346 14657
rect 38290 14583 38346 14592
rect 38384 14544 38436 14550
rect 38212 14504 38384 14532
rect 38384 14486 38436 14492
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 38488 14074 38516 15399
rect 38764 15337 38792 16238
rect 38842 15872 38898 15881
rect 38842 15807 38898 15816
rect 38856 15502 38884 15807
rect 38844 15496 38896 15502
rect 38844 15438 38896 15444
rect 38750 15328 38806 15337
rect 38750 15263 38806 15272
rect 38752 15088 38804 15094
rect 38856 15076 38884 15438
rect 38934 15192 38990 15201
rect 38934 15127 38990 15136
rect 38804 15048 38884 15076
rect 38752 15030 38804 15036
rect 38856 14414 38884 15048
rect 38948 14414 38976 15127
rect 38844 14408 38896 14414
rect 38844 14350 38896 14356
rect 38936 14408 38988 14414
rect 38936 14350 38988 14356
rect 38936 14272 38988 14278
rect 38936 14214 38988 14220
rect 38476 14068 38528 14074
rect 38476 14010 38528 14016
rect 38292 13864 38344 13870
rect 38290 13832 38292 13841
rect 38344 13832 38346 13841
rect 38016 13796 38068 13802
rect 38016 13738 38068 13744
rect 38200 13796 38252 13802
rect 38290 13767 38346 13776
rect 38200 13738 38252 13744
rect 38028 13546 38056 13738
rect 37936 13518 38056 13546
rect 38212 13530 38240 13738
rect 38292 13728 38344 13734
rect 38292 13670 38344 13676
rect 38568 13728 38620 13734
rect 38948 13705 38976 14214
rect 38568 13670 38620 13676
rect 38934 13696 38990 13705
rect 38200 13524 38252 13530
rect 37936 13240 37964 13518
rect 38200 13466 38252 13472
rect 37844 13212 37964 13240
rect 37844 12986 37872 13212
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 37832 12980 37884 12986
rect 37832 12922 37884 12928
rect 37832 12640 37884 12646
rect 37832 12582 37884 12588
rect 37738 12336 37794 12345
rect 37738 12271 37794 12280
rect 37740 12164 37792 12170
rect 37740 12106 37792 12112
rect 37752 11830 37780 12106
rect 37740 11824 37792 11830
rect 37740 11766 37792 11772
rect 37740 11688 37792 11694
rect 37660 11636 37740 11642
rect 37660 11630 37792 11636
rect 37660 11614 37780 11630
rect 37556 11280 37608 11286
rect 37280 11144 37332 11150
rect 37200 11092 37280 11098
rect 37200 11086 37332 11092
rect 37200 11070 37320 11086
rect 37016 10934 37228 10962
rect 37094 10840 37150 10849
rect 37004 10804 37056 10810
rect 37094 10775 37096 10784
rect 37004 10746 37056 10752
rect 37148 10775 37150 10784
rect 37096 10746 37148 10752
rect 36912 10668 36964 10674
rect 36912 10610 36964 10616
rect 36912 10464 36964 10470
rect 36912 10406 36964 10412
rect 36924 10130 36952 10406
rect 36912 10124 36964 10130
rect 36912 10066 36964 10072
rect 37016 9908 37044 10746
rect 37108 10441 37136 10746
rect 37094 10432 37150 10441
rect 37094 10367 37150 10376
rect 37200 9926 37228 10934
rect 37096 9920 37148 9926
rect 37016 9880 37096 9908
rect 37096 9862 37148 9868
rect 37188 9920 37240 9926
rect 37188 9862 37240 9868
rect 37004 9716 37056 9722
rect 37004 9658 37056 9664
rect 37016 9382 37044 9658
rect 37004 9376 37056 9382
rect 37004 9318 37056 9324
rect 37016 9081 37044 9318
rect 37002 9072 37058 9081
rect 37002 9007 37058 9016
rect 36726 8936 36782 8945
rect 36726 8871 36782 8880
rect 36636 8560 36688 8566
rect 36636 8502 36688 8508
rect 36452 5704 36504 5710
rect 36452 5646 36504 5652
rect 35900 5092 35952 5098
rect 35900 5034 35952 5040
rect 34428 4004 34480 4010
rect 34428 3946 34480 3952
rect 33876 3732 33928 3738
rect 33876 3674 33928 3680
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 34440 2650 34468 3946
rect 36820 3664 36872 3670
rect 36820 3606 36872 3612
rect 30840 2644 30892 2650
rect 30840 2586 30892 2592
rect 32864 2644 32916 2650
rect 32864 2586 32916 2592
rect 34428 2644 34480 2650
rect 34428 2586 34480 2592
rect 30748 2576 30800 2582
rect 30748 2518 30800 2524
rect 36832 2514 36860 3606
rect 37108 3602 37136 9862
rect 37278 9752 37334 9761
rect 37278 9687 37334 9696
rect 37188 9648 37240 9654
rect 37188 9590 37240 9596
rect 37200 9489 37228 9590
rect 37292 9586 37320 9687
rect 37280 9580 37332 9586
rect 37280 9522 37332 9528
rect 37186 9480 37242 9489
rect 37186 9415 37242 9424
rect 37280 9376 37332 9382
rect 37280 9318 37332 9324
rect 37188 9172 37240 9178
rect 37188 9114 37240 9120
rect 37200 8809 37228 9114
rect 37186 8800 37242 8809
rect 37186 8735 37242 8744
rect 37188 7744 37240 7750
rect 37188 7686 37240 7692
rect 37200 6730 37228 7686
rect 37292 7342 37320 9318
rect 37384 9217 37412 11240
rect 37462 11248 37518 11257
rect 37556 11222 37608 11228
rect 37462 11183 37518 11192
rect 37568 10810 37596 11222
rect 37648 11076 37700 11082
rect 37648 11018 37700 11024
rect 37556 10804 37608 10810
rect 37556 10746 37608 10752
rect 37464 10736 37516 10742
rect 37464 10678 37516 10684
rect 37476 9897 37504 10678
rect 37660 10674 37688 11018
rect 37738 10976 37794 10985
rect 37738 10911 37794 10920
rect 37648 10668 37700 10674
rect 37648 10610 37700 10616
rect 37462 9888 37518 9897
rect 37462 9823 37518 9832
rect 37556 9444 37608 9450
rect 37556 9386 37608 9392
rect 37370 9208 37426 9217
rect 37370 9143 37426 9152
rect 37372 9104 37424 9110
rect 37372 9046 37424 9052
rect 37384 7546 37412 9046
rect 37568 8974 37596 9386
rect 37556 8968 37608 8974
rect 37556 8910 37608 8916
rect 37648 8832 37700 8838
rect 37648 8774 37700 8780
rect 37464 8492 37516 8498
rect 37464 8434 37516 8440
rect 37476 8362 37504 8434
rect 37464 8356 37516 8362
rect 37464 8298 37516 8304
rect 37372 7540 37424 7546
rect 37372 7482 37424 7488
rect 37280 7336 37332 7342
rect 37280 7278 37332 7284
rect 37188 6724 37240 6730
rect 37188 6666 37240 6672
rect 37660 5370 37688 8774
rect 37752 7868 37780 10911
rect 37844 10674 37872 12582
rect 38304 12345 38332 13670
rect 38476 13388 38528 13394
rect 38476 13330 38528 13336
rect 38382 12608 38438 12617
rect 38382 12543 38438 12552
rect 38290 12336 38346 12345
rect 38290 12271 38346 12280
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 38292 11144 38344 11150
rect 38292 11086 38344 11092
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 38016 10804 38068 10810
rect 38016 10746 38068 10752
rect 37832 10668 37884 10674
rect 37832 10610 37884 10616
rect 37844 9722 37872 10610
rect 38028 10130 38056 10746
rect 38304 10690 38332 11086
rect 38396 10985 38424 12543
rect 38488 12345 38516 13330
rect 38474 12336 38530 12345
rect 38580 12306 38608 13670
rect 38934 13631 38990 13640
rect 38936 13320 38988 13326
rect 38936 13262 38988 13268
rect 38752 12912 38804 12918
rect 38752 12854 38804 12860
rect 38474 12271 38530 12280
rect 38568 12300 38620 12306
rect 38568 12242 38620 12248
rect 38476 12096 38528 12102
rect 38476 12038 38528 12044
rect 38660 12096 38712 12102
rect 38660 12038 38712 12044
rect 38382 10976 38438 10985
rect 38382 10911 38438 10920
rect 38304 10662 38424 10690
rect 38108 10600 38160 10606
rect 38108 10542 38160 10548
rect 38292 10600 38344 10606
rect 38292 10542 38344 10548
rect 38016 10124 38068 10130
rect 38016 10066 38068 10072
rect 38120 9926 38148 10542
rect 38108 9920 38160 9926
rect 38108 9862 38160 9868
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 37832 9716 37884 9722
rect 37832 9658 37884 9664
rect 37844 9586 37872 9658
rect 37832 9580 37884 9586
rect 37832 9522 37884 9528
rect 37830 9480 37886 9489
rect 37830 9415 37886 9424
rect 37844 8430 37872 9415
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 38304 8634 38332 10542
rect 38396 9110 38424 10662
rect 38488 9450 38516 12038
rect 38568 11348 38620 11354
rect 38568 11290 38620 11296
rect 38580 11150 38608 11290
rect 38568 11144 38620 11150
rect 38568 11086 38620 11092
rect 38580 10674 38608 11086
rect 38568 10668 38620 10674
rect 38568 10610 38620 10616
rect 38568 10532 38620 10538
rect 38568 10474 38620 10480
rect 38580 9586 38608 10474
rect 38672 10266 38700 12038
rect 38764 11744 38792 12854
rect 38844 11756 38896 11762
rect 38764 11716 38844 11744
rect 38844 11698 38896 11704
rect 38856 11082 38884 11698
rect 38844 11076 38896 11082
rect 38844 11018 38896 11024
rect 38660 10260 38712 10266
rect 38660 10202 38712 10208
rect 38660 10056 38712 10062
rect 38660 9998 38712 10004
rect 38672 9722 38700 9998
rect 38948 9908 38976 13262
rect 39040 11014 39068 17190
rect 39304 16652 39356 16658
rect 39304 16594 39356 16600
rect 39120 15496 39172 15502
rect 39120 15438 39172 15444
rect 39132 15366 39160 15438
rect 39316 15366 39344 16594
rect 39408 15502 39436 17546
rect 39488 17536 39540 17542
rect 39488 17478 39540 17484
rect 39500 16658 39528 17478
rect 39488 16652 39540 16658
rect 39488 16594 39540 16600
rect 39488 16516 39540 16522
rect 39488 16458 39540 16464
rect 39500 15638 39528 16458
rect 39672 16448 39724 16454
rect 39776 16425 39804 18702
rect 39868 18193 39896 18770
rect 39960 18698 39988 19306
rect 40132 19304 40184 19310
rect 40038 19272 40094 19281
rect 40132 19246 40184 19252
rect 40316 19304 40368 19310
rect 40316 19246 40368 19252
rect 40038 19207 40094 19216
rect 40052 19174 40080 19207
rect 40040 19168 40092 19174
rect 40040 19110 40092 19116
rect 40040 18760 40092 18766
rect 40040 18702 40092 18708
rect 39948 18692 40000 18698
rect 39948 18634 40000 18640
rect 39960 18290 39988 18634
rect 39948 18284 40000 18290
rect 39948 18226 40000 18232
rect 39854 18184 39910 18193
rect 39854 18119 39910 18128
rect 40052 18086 40080 18702
rect 40144 18465 40172 19246
rect 40224 19168 40276 19174
rect 40224 19110 40276 19116
rect 40130 18456 40186 18465
rect 40130 18391 40186 18400
rect 40132 18352 40184 18358
rect 40132 18294 40184 18300
rect 40144 18086 40172 18294
rect 40040 18080 40092 18086
rect 40040 18022 40092 18028
rect 40132 18080 40184 18086
rect 40132 18022 40184 18028
rect 40052 17746 40080 18022
rect 40236 17954 40264 19110
rect 40316 18692 40368 18698
rect 40316 18634 40368 18640
rect 40328 18290 40356 18634
rect 40316 18284 40368 18290
rect 40316 18226 40368 18232
rect 40314 18184 40370 18193
rect 40314 18119 40316 18128
rect 40368 18119 40370 18128
rect 40316 18090 40368 18096
rect 40144 17926 40264 17954
rect 39856 17740 39908 17746
rect 39856 17682 39908 17688
rect 40040 17740 40092 17746
rect 40040 17682 40092 17688
rect 39672 16390 39724 16396
rect 39762 16416 39818 16425
rect 39684 16114 39712 16390
rect 39762 16351 39818 16360
rect 39672 16108 39724 16114
rect 39672 16050 39724 16056
rect 39684 15881 39712 16050
rect 39868 15910 39896 17682
rect 40040 16448 40092 16454
rect 40040 16390 40092 16396
rect 40052 16250 40080 16390
rect 40144 16289 40172 17926
rect 40420 16810 40448 19314
rect 40500 19304 40552 19310
rect 40500 19246 40552 19252
rect 40512 18193 40540 19246
rect 40592 18624 40644 18630
rect 40592 18566 40644 18572
rect 40604 18426 40632 18566
rect 40592 18420 40644 18426
rect 40592 18362 40644 18368
rect 40592 18284 40644 18290
rect 40592 18226 40644 18232
rect 40498 18184 40554 18193
rect 40498 18119 40554 18128
rect 40604 16969 40632 18226
rect 40590 16960 40646 16969
rect 40590 16895 40646 16904
rect 40328 16782 40448 16810
rect 40498 16824 40554 16833
rect 40224 16652 40276 16658
rect 40224 16594 40276 16600
rect 40130 16280 40186 16289
rect 40040 16244 40092 16250
rect 40130 16215 40186 16224
rect 40040 16186 40092 16192
rect 39856 15904 39908 15910
rect 39670 15872 39726 15881
rect 39856 15846 39908 15852
rect 39670 15807 39726 15816
rect 39488 15632 39540 15638
rect 39488 15574 39540 15580
rect 39396 15496 39448 15502
rect 39396 15438 39448 15444
rect 39120 15360 39172 15366
rect 39120 15302 39172 15308
rect 39304 15360 39356 15366
rect 39304 15302 39356 15308
rect 39316 14890 39344 15302
rect 39304 14884 39356 14890
rect 39304 14826 39356 14832
rect 39132 14606 39436 14634
rect 39132 14346 39160 14606
rect 39408 14550 39436 14606
rect 39212 14544 39264 14550
rect 39304 14544 39356 14550
rect 39212 14486 39264 14492
rect 39302 14512 39304 14521
rect 39396 14544 39448 14550
rect 39356 14512 39358 14521
rect 39224 14346 39252 14486
rect 39396 14486 39448 14492
rect 39302 14447 39358 14456
rect 39120 14340 39172 14346
rect 39120 14282 39172 14288
rect 39212 14340 39264 14346
rect 39212 14282 39264 14288
rect 39224 12434 39252 14282
rect 39304 13184 39356 13190
rect 39304 13126 39356 13132
rect 39316 12889 39344 13126
rect 39302 12880 39358 12889
rect 39302 12815 39358 12824
rect 39224 12406 39344 12434
rect 39212 12300 39264 12306
rect 39212 12242 39264 12248
rect 39224 11898 39252 12242
rect 39212 11892 39264 11898
rect 39212 11834 39264 11840
rect 39118 11384 39174 11393
rect 39118 11319 39120 11328
rect 39172 11319 39174 11328
rect 39120 11290 39172 11296
rect 39028 11008 39080 11014
rect 39028 10950 39080 10956
rect 39026 10024 39082 10033
rect 39026 9959 39082 9968
rect 38764 9880 38976 9908
rect 38660 9716 38712 9722
rect 38660 9658 38712 9664
rect 38568 9580 38620 9586
rect 38568 9522 38620 9528
rect 38476 9444 38528 9450
rect 38476 9386 38528 9392
rect 38660 9444 38712 9450
rect 38660 9386 38712 9392
rect 38568 9172 38620 9178
rect 38568 9114 38620 9120
rect 38384 9104 38436 9110
rect 38384 9046 38436 9052
rect 38476 8832 38528 8838
rect 38476 8774 38528 8780
rect 38292 8628 38344 8634
rect 38292 8570 38344 8576
rect 38384 8628 38436 8634
rect 38384 8570 38436 8576
rect 38016 8560 38068 8566
rect 38016 8502 38068 8508
rect 37832 8424 37884 8430
rect 37832 8366 37884 8372
rect 38028 8362 38056 8502
rect 38016 8356 38068 8362
rect 38016 8298 38068 8304
rect 38396 8294 38424 8570
rect 38488 8344 38516 8774
rect 38580 8548 38608 9114
rect 38672 8945 38700 9386
rect 38658 8936 38714 8945
rect 38658 8871 38714 8880
rect 38764 8809 38792 9880
rect 38842 9616 38898 9625
rect 38842 9551 38898 9560
rect 38936 9580 38988 9586
rect 38856 9178 38884 9551
rect 38936 9522 38988 9528
rect 38948 9489 38976 9522
rect 38934 9480 38990 9489
rect 38934 9415 38990 9424
rect 38936 9376 38988 9382
rect 38936 9318 38988 9324
rect 38844 9172 38896 9178
rect 38844 9114 38896 9120
rect 38948 9110 38976 9318
rect 38936 9104 38988 9110
rect 38936 9046 38988 9052
rect 38948 8906 38976 9046
rect 38936 8900 38988 8906
rect 38936 8842 38988 8848
rect 38750 8800 38806 8809
rect 38750 8735 38806 8744
rect 39040 8634 39068 9959
rect 39120 9648 39172 9654
rect 39120 9590 39172 9596
rect 39132 9489 39160 9590
rect 39118 9480 39174 9489
rect 39118 9415 39174 9424
rect 39316 9058 39344 12406
rect 39500 12288 39528 15574
rect 39578 15192 39634 15201
rect 39578 15127 39634 15136
rect 39592 13977 39620 15127
rect 39578 13968 39634 13977
rect 39578 13903 39634 13912
rect 39684 13530 39712 15807
rect 39764 15360 39816 15366
rect 39764 15302 39816 15308
rect 39776 14822 39804 15302
rect 39948 15020 40000 15026
rect 39948 14962 40000 14968
rect 39764 14816 39816 14822
rect 39764 14758 39816 14764
rect 39856 14816 39908 14822
rect 39856 14758 39908 14764
rect 39868 14550 39896 14758
rect 39856 14544 39908 14550
rect 39762 14512 39818 14521
rect 39856 14486 39908 14492
rect 39762 14447 39764 14456
rect 39816 14447 39818 14456
rect 39764 14418 39816 14424
rect 39856 14340 39908 14346
rect 39960 14328 39988 14962
rect 40236 14793 40264 16594
rect 40328 15201 40356 16782
rect 40498 16759 40554 16768
rect 40512 16658 40540 16759
rect 40500 16652 40552 16658
rect 40500 16594 40552 16600
rect 40408 16108 40460 16114
rect 40408 16050 40460 16056
rect 40314 15192 40370 15201
rect 40314 15127 40370 15136
rect 40222 14784 40278 14793
rect 40222 14719 40278 14728
rect 40224 14544 40276 14550
rect 40224 14486 40276 14492
rect 39908 14300 39988 14328
rect 40130 14376 40186 14385
rect 40130 14311 40132 14320
rect 39856 14282 39908 14288
rect 39960 13938 39988 14300
rect 40184 14311 40186 14320
rect 40132 14282 40184 14288
rect 39764 13932 39816 13938
rect 39764 13874 39816 13880
rect 39856 13932 39908 13938
rect 39856 13874 39908 13880
rect 39948 13932 40000 13938
rect 39948 13874 40000 13880
rect 39672 13524 39724 13530
rect 39672 13466 39724 13472
rect 39684 13326 39712 13466
rect 39672 13320 39724 13326
rect 39672 13262 39724 13268
rect 39580 12776 39632 12782
rect 39580 12718 39632 12724
rect 39592 12646 39620 12718
rect 39580 12640 39632 12646
rect 39578 12608 39580 12617
rect 39632 12608 39634 12617
rect 39578 12543 39634 12552
rect 39408 12260 39528 12288
rect 39408 10130 39436 12260
rect 39684 12238 39712 13262
rect 39672 12232 39724 12238
rect 39672 12174 39724 12180
rect 39488 12096 39540 12102
rect 39488 12038 39540 12044
rect 39672 12096 39724 12102
rect 39672 12038 39724 12044
rect 39500 11257 39528 12038
rect 39684 11370 39712 12038
rect 39776 11558 39804 13874
rect 39868 13530 39896 13874
rect 39856 13524 39908 13530
rect 39856 13466 39908 13472
rect 40040 13320 40092 13326
rect 40040 13262 40092 13268
rect 39948 13184 40000 13190
rect 39948 13126 40000 13132
rect 39960 12850 39988 13126
rect 40052 12918 40080 13262
rect 40040 12912 40092 12918
rect 40040 12854 40092 12860
rect 39948 12844 40000 12850
rect 39948 12786 40000 12792
rect 39856 12232 39908 12238
rect 39856 12174 39908 12180
rect 40132 12232 40184 12238
rect 40132 12174 40184 12180
rect 39868 11830 39896 12174
rect 39856 11824 39908 11830
rect 39856 11766 39908 11772
rect 39764 11552 39816 11558
rect 39764 11494 39816 11500
rect 39592 11342 39712 11370
rect 39868 11354 39896 11766
rect 40144 11370 40172 12174
rect 40236 11762 40264 14486
rect 40316 13252 40368 13258
rect 40316 13194 40368 13200
rect 40328 11898 40356 13194
rect 40420 12434 40448 16050
rect 40590 13968 40646 13977
rect 40590 13903 40646 13912
rect 40500 13864 40552 13870
rect 40500 13806 40552 13812
rect 40512 13433 40540 13806
rect 40604 13734 40632 13903
rect 40592 13728 40644 13734
rect 40592 13670 40644 13676
rect 40498 13424 40554 13433
rect 40498 13359 40554 13368
rect 40590 13288 40646 13297
rect 40590 13223 40646 13232
rect 40604 12986 40632 13223
rect 40592 12980 40644 12986
rect 40592 12922 40644 12928
rect 40420 12406 40540 12434
rect 40512 12073 40540 12406
rect 40498 12064 40554 12073
rect 40498 11999 40554 12008
rect 40316 11892 40368 11898
rect 40316 11834 40368 11840
rect 40224 11756 40276 11762
rect 40224 11698 40276 11704
rect 39856 11348 39908 11354
rect 39486 11248 39542 11257
rect 39486 11183 39542 11192
rect 39396 10124 39448 10130
rect 39396 10066 39448 10072
rect 39120 9036 39172 9042
rect 39120 8978 39172 8984
rect 39224 9030 39344 9058
rect 39028 8628 39080 8634
rect 39028 8570 39080 8576
rect 38936 8560 38988 8566
rect 38580 8520 38654 8548
rect 38626 8514 38654 8520
rect 38856 8520 38936 8548
rect 38626 8486 38700 8514
rect 38672 8412 38700 8486
rect 38856 8412 38884 8520
rect 38936 8502 38988 8508
rect 38672 8384 38884 8412
rect 38936 8356 38988 8362
rect 38488 8316 38936 8344
rect 38936 8298 38988 8304
rect 38304 8266 38424 8294
rect 37832 7880 37884 7886
rect 37752 7840 37832 7868
rect 37752 7342 37780 7840
rect 37832 7822 37884 7828
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 38014 7440 38070 7449
rect 38014 7375 38016 7384
rect 38068 7375 38070 7384
rect 38016 7346 38068 7352
rect 37740 7336 37792 7342
rect 37740 7278 37792 7284
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 38304 5710 38332 8266
rect 39040 7818 39068 8570
rect 39132 8430 39160 8978
rect 39120 8424 39172 8430
rect 39120 8366 39172 8372
rect 39028 7812 39080 7818
rect 39028 7754 39080 7760
rect 39132 7313 39160 8366
rect 39224 8265 39252 9030
rect 39304 8900 39356 8906
rect 39304 8842 39356 8848
rect 39210 8256 39266 8265
rect 39210 8191 39266 8200
rect 39212 7744 39264 7750
rect 39212 7686 39264 7692
rect 39118 7304 39174 7313
rect 39118 7239 39174 7248
rect 38384 6248 38436 6254
rect 38384 6190 38436 6196
rect 38396 5778 38424 6190
rect 38384 5772 38436 5778
rect 38384 5714 38436 5720
rect 38292 5704 38344 5710
rect 38292 5646 38344 5652
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 37648 5364 37700 5370
rect 37648 5306 37700 5312
rect 38106 5264 38162 5273
rect 38106 5199 38108 5208
rect 38160 5199 38162 5208
rect 38108 5170 38160 5176
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 39224 4078 39252 7686
rect 39316 7002 39344 8842
rect 39304 6996 39356 7002
rect 39304 6938 39356 6944
rect 39408 5681 39436 10066
rect 39500 8430 39528 11183
rect 39592 10674 39620 11342
rect 40144 11342 40264 11370
rect 39856 11290 39908 11296
rect 39672 11144 39724 11150
rect 39672 11086 39724 11092
rect 40132 11144 40184 11150
rect 40132 11086 40184 11092
rect 39580 10668 39632 10674
rect 39580 10610 39632 10616
rect 39578 9208 39634 9217
rect 39578 9143 39634 9152
rect 39592 8906 39620 9143
rect 39580 8900 39632 8906
rect 39580 8842 39632 8848
rect 39592 8634 39620 8842
rect 39580 8628 39632 8634
rect 39580 8570 39632 8576
rect 39488 8424 39540 8430
rect 39488 8366 39540 8372
rect 39394 5672 39450 5681
rect 39394 5607 39450 5616
rect 39396 4480 39448 4486
rect 39396 4422 39448 4428
rect 39212 4072 39264 4078
rect 39212 4014 39264 4020
rect 37096 3596 37148 3602
rect 37096 3538 37148 3544
rect 39212 3460 39264 3466
rect 39212 3402 39264 3408
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 38292 2848 38344 2854
rect 38292 2790 38344 2796
rect 36820 2508 36872 2514
rect 36820 2450 36872 2456
rect 38304 2446 38332 2790
rect 27528 2440 27580 2446
rect 27528 2382 27580 2388
rect 28632 2440 28684 2446
rect 28632 2382 28684 2388
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 33140 2440 33192 2446
rect 33140 2382 33192 2388
rect 34980 2440 35032 2446
rect 34980 2382 35032 2388
rect 38292 2440 38344 2446
rect 38292 2382 38344 2388
rect 26516 2372 26568 2378
rect 26516 2314 26568 2320
rect 26528 800 26556 2314
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 28644 800 28672 2382
rect 30760 800 30788 2382
rect 33152 1578 33180 2382
rect 32876 1550 33180 1578
rect 32876 800 32904 1550
rect 34992 800 35020 2382
rect 37096 2304 37148 2310
rect 37096 2246 37148 2252
rect 37108 800 37136 2246
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 39224 800 39252 3402
rect 39408 3058 39436 4422
rect 39684 3670 39712 11086
rect 39856 10600 39908 10606
rect 39856 10542 39908 10548
rect 39868 10441 39896 10542
rect 39854 10432 39910 10441
rect 39854 10367 39910 10376
rect 39868 9994 39896 10367
rect 39856 9988 39908 9994
rect 39856 9930 39908 9936
rect 40144 9722 40172 11086
rect 40132 9716 40184 9722
rect 40132 9658 40184 9664
rect 39856 9648 39908 9654
rect 39856 9590 39908 9596
rect 39764 9580 39816 9586
rect 39764 9522 39816 9528
rect 39776 9178 39804 9522
rect 39868 9489 39896 9590
rect 39948 9512 40000 9518
rect 39854 9480 39910 9489
rect 39948 9454 40000 9460
rect 39854 9415 39910 9424
rect 39856 9376 39908 9382
rect 39856 9318 39908 9324
rect 39764 9172 39816 9178
rect 39764 9114 39816 9120
rect 39868 9110 39896 9318
rect 39856 9104 39908 9110
rect 39856 9046 39908 9052
rect 39960 8294 39988 9454
rect 40040 8560 40092 8566
rect 40038 8528 40040 8537
rect 40092 8528 40094 8537
rect 40038 8463 40094 8472
rect 39948 8288 40000 8294
rect 39948 8230 40000 8236
rect 40236 8129 40264 11342
rect 40408 10464 40460 10470
rect 40408 10406 40460 10412
rect 40420 10198 40448 10406
rect 40408 10192 40460 10198
rect 40408 10134 40460 10140
rect 40316 8900 40368 8906
rect 40316 8842 40368 8848
rect 40222 8120 40278 8129
rect 40222 8055 40278 8064
rect 40224 7880 40276 7886
rect 40130 7848 40186 7857
rect 40224 7822 40276 7828
rect 40130 7783 40132 7792
rect 40184 7783 40186 7792
rect 40132 7754 40184 7760
rect 40144 7478 40172 7754
rect 40132 7472 40184 7478
rect 40132 7414 40184 7420
rect 40132 7336 40184 7342
rect 40132 7278 40184 7284
rect 40038 6352 40094 6361
rect 40038 6287 40040 6296
rect 40092 6287 40094 6296
rect 40040 6258 40092 6264
rect 40144 5234 40172 7278
rect 40132 5228 40184 5234
rect 40132 5170 40184 5176
rect 40236 4690 40264 7822
rect 40328 6662 40356 8842
rect 40316 6656 40368 6662
rect 40316 6598 40368 6604
rect 40408 5160 40460 5166
rect 40408 5102 40460 5108
rect 40224 4684 40276 4690
rect 40224 4626 40276 4632
rect 39672 3664 39724 3670
rect 39672 3606 39724 3612
rect 40420 3534 40448 5102
rect 40512 4010 40540 11999
rect 40592 11756 40644 11762
rect 40592 11698 40644 11704
rect 40604 11354 40632 11698
rect 40592 11348 40644 11354
rect 40592 11290 40644 11296
rect 40696 11257 40724 22510
rect 40788 20466 40816 23310
rect 40972 23254 41000 26687
rect 42154 26330 42210 27000
rect 42154 26302 42472 26330
rect 42154 26200 42210 26302
rect 41880 25492 41932 25498
rect 41880 25434 41932 25440
rect 41420 25152 41472 25158
rect 41420 25094 41472 25100
rect 41328 25016 41380 25022
rect 41328 24958 41380 24964
rect 41144 24064 41196 24070
rect 41144 24006 41196 24012
rect 41052 23724 41104 23730
rect 41052 23666 41104 23672
rect 40960 23248 41012 23254
rect 40960 23190 41012 23196
rect 40960 22976 41012 22982
rect 40960 22918 41012 22924
rect 40972 22001 41000 22918
rect 40958 21992 41014 22001
rect 40868 21956 40920 21962
rect 40958 21927 41014 21936
rect 40868 21898 40920 21904
rect 40776 20460 40828 20466
rect 40776 20402 40828 20408
rect 40776 19984 40828 19990
rect 40776 19926 40828 19932
rect 40788 18222 40816 19926
rect 40776 18216 40828 18222
rect 40776 18158 40828 18164
rect 40776 17604 40828 17610
rect 40776 17546 40828 17552
rect 40788 17270 40816 17546
rect 40776 17264 40828 17270
rect 40776 17206 40828 17212
rect 40788 15881 40816 17206
rect 40774 15872 40830 15881
rect 40774 15807 40830 15816
rect 40880 15162 40908 21898
rect 40972 21729 41000 21927
rect 40958 21720 41014 21729
rect 40958 21655 41014 21664
rect 41064 19904 41092 23666
rect 41156 20942 41184 24006
rect 41236 23588 41288 23594
rect 41236 23530 41288 23536
rect 41248 22574 41276 23530
rect 41236 22568 41288 22574
rect 41234 22536 41236 22545
rect 41288 22536 41290 22545
rect 41234 22471 41290 22480
rect 41234 22400 41290 22409
rect 41234 22335 41290 22344
rect 41248 22137 41276 22335
rect 41234 22128 41290 22137
rect 41234 22063 41290 22072
rect 41236 21888 41288 21894
rect 41236 21830 41288 21836
rect 41248 21690 41276 21830
rect 41236 21684 41288 21690
rect 41236 21626 41288 21632
rect 41236 21412 41288 21418
rect 41236 21354 41288 21360
rect 41248 21146 41276 21354
rect 41236 21140 41288 21146
rect 41236 21082 41288 21088
rect 41144 20936 41196 20942
rect 41144 20878 41196 20884
rect 41234 20904 41290 20913
rect 41234 20839 41290 20848
rect 41142 20496 41198 20505
rect 41142 20431 41144 20440
rect 41196 20431 41198 20440
rect 41144 20402 41196 20408
rect 41064 19876 41184 19904
rect 41156 19666 41184 19876
rect 41064 19638 41184 19666
rect 41248 19666 41276 20839
rect 41340 20233 41368 24958
rect 41432 24274 41460 25094
rect 41420 24268 41472 24274
rect 41420 24210 41472 24216
rect 41432 22001 41460 24210
rect 41696 24132 41748 24138
rect 41696 24074 41748 24080
rect 41604 22432 41656 22438
rect 41604 22374 41656 22380
rect 41512 22024 41564 22030
rect 41418 21992 41474 22001
rect 41512 21966 41564 21972
rect 41418 21927 41474 21936
rect 41524 21486 41552 21966
rect 41616 21729 41644 22374
rect 41708 22030 41736 24074
rect 41892 23866 41920 25434
rect 41972 25084 42024 25090
rect 41972 25026 42024 25032
rect 41880 23860 41932 23866
rect 41880 23802 41932 23808
rect 41880 22500 41932 22506
rect 41880 22442 41932 22448
rect 41892 22273 41920 22442
rect 41878 22264 41934 22273
rect 41878 22199 41934 22208
rect 41696 22024 41748 22030
rect 41696 21966 41748 21972
rect 41880 22024 41932 22030
rect 41880 21966 41932 21972
rect 41602 21720 41658 21729
rect 41602 21655 41658 21664
rect 41604 21616 41656 21622
rect 41604 21558 41656 21564
rect 41512 21480 41564 21486
rect 41512 21422 41564 21428
rect 41420 21072 41472 21078
rect 41420 21014 41472 21020
rect 41432 20942 41460 21014
rect 41420 20936 41472 20942
rect 41420 20878 41472 20884
rect 41512 20800 41564 20806
rect 41512 20742 41564 20748
rect 41418 20360 41474 20369
rect 41418 20295 41474 20304
rect 41326 20224 41382 20233
rect 41326 20159 41382 20168
rect 41432 20074 41460 20295
rect 41340 20046 41460 20074
rect 41340 19786 41368 20046
rect 41328 19780 41380 19786
rect 41328 19722 41380 19728
rect 41248 19638 41460 19666
rect 40960 19508 41012 19514
rect 40960 19450 41012 19456
rect 40972 18086 41000 19450
rect 40960 18080 41012 18086
rect 40960 18022 41012 18028
rect 40958 17368 41014 17377
rect 40958 17303 40960 17312
rect 41012 17303 41014 17312
rect 40960 17274 41012 17280
rect 40960 16992 41012 16998
rect 40960 16934 41012 16940
rect 40972 16658 41000 16934
rect 40960 16652 41012 16658
rect 40960 16594 41012 16600
rect 40960 15904 41012 15910
rect 40960 15846 41012 15852
rect 40868 15156 40920 15162
rect 40868 15098 40920 15104
rect 40776 15088 40828 15094
rect 40776 15030 40828 15036
rect 40866 15056 40922 15065
rect 40682 11248 40738 11257
rect 40682 11183 40738 11192
rect 40684 10464 40736 10470
rect 40684 10406 40736 10412
rect 40696 10062 40724 10406
rect 40684 10056 40736 10062
rect 40684 9998 40736 10004
rect 40592 9580 40644 9586
rect 40592 9522 40644 9528
rect 40604 8022 40632 9522
rect 40592 8016 40644 8022
rect 40592 7958 40644 7964
rect 40788 7478 40816 15030
rect 40866 14991 40922 15000
rect 40880 9042 40908 14991
rect 40972 11121 41000 15846
rect 40958 11112 41014 11121
rect 40958 11047 41014 11056
rect 40960 10668 41012 10674
rect 40960 10610 41012 10616
rect 40972 10305 41000 10610
rect 40958 10296 41014 10305
rect 40958 10231 41014 10240
rect 40868 9036 40920 9042
rect 40868 8978 40920 8984
rect 40868 8424 40920 8430
rect 40868 8366 40920 8372
rect 40880 8022 40908 8366
rect 41064 8022 41092 19638
rect 41144 19440 41196 19446
rect 41142 19408 41144 19417
rect 41328 19440 41380 19446
rect 41196 19408 41198 19417
rect 41142 19343 41198 19352
rect 41264 19388 41328 19394
rect 41264 19382 41380 19388
rect 41264 19366 41368 19382
rect 41264 19334 41292 19366
rect 41248 19306 41292 19334
rect 41248 19242 41276 19306
rect 41328 19304 41380 19310
rect 41432 19292 41460 19638
rect 41380 19264 41460 19292
rect 41328 19246 41380 19252
rect 41236 19236 41288 19242
rect 41236 19178 41288 19184
rect 41248 18680 41276 19178
rect 41248 18652 41460 18680
rect 41236 18352 41288 18358
rect 41236 18294 41288 18300
rect 41144 18080 41196 18086
rect 41248 18057 41276 18294
rect 41432 18222 41460 18652
rect 41524 18306 41552 20742
rect 41616 19145 41644 21558
rect 41708 20913 41736 21966
rect 41788 21956 41840 21962
rect 41788 21898 41840 21904
rect 41694 20904 41750 20913
rect 41694 20839 41750 20848
rect 41800 19334 41828 21898
rect 41892 21146 41920 21966
rect 41880 21140 41932 21146
rect 41880 21082 41932 21088
rect 41878 20768 41934 20777
rect 41878 20703 41934 20712
rect 41892 20602 41920 20703
rect 41984 20602 42012 25026
rect 42246 24032 42302 24041
rect 42246 23967 42302 23976
rect 42260 23866 42288 23967
rect 42248 23860 42300 23866
rect 42248 23802 42300 23808
rect 42444 23497 42472 26302
rect 42798 26200 42854 27000
rect 43442 26200 43498 27000
rect 43812 26376 43864 26382
rect 44086 26330 44142 27000
rect 44730 26330 44786 27000
rect 43864 26324 44142 26330
rect 43812 26318 44142 26324
rect 43824 26302 44142 26318
rect 44086 26200 44142 26302
rect 44652 26302 44786 26330
rect 43352 26104 43404 26110
rect 43352 26046 43404 26052
rect 43534 26072 43590 26081
rect 42524 25220 42576 25226
rect 42524 25162 42576 25168
rect 42430 23488 42486 23497
rect 42430 23423 42486 23432
rect 42340 23316 42392 23322
rect 42340 23258 42392 23264
rect 42064 22976 42116 22982
rect 42064 22918 42116 22924
rect 42076 21978 42104 22918
rect 42352 22522 42380 23258
rect 42430 22672 42486 22681
rect 42430 22607 42432 22616
rect 42484 22607 42486 22616
rect 42432 22578 42484 22584
rect 42352 22494 42472 22522
rect 42246 22264 42302 22273
rect 42246 22199 42302 22208
rect 42260 22098 42288 22199
rect 42248 22092 42300 22098
rect 42248 22034 42300 22040
rect 42076 21950 42380 21978
rect 42156 21888 42208 21894
rect 42156 21830 42208 21836
rect 42168 21418 42196 21830
rect 42246 21720 42302 21729
rect 42246 21655 42302 21664
rect 42156 21412 42208 21418
rect 42156 21354 42208 21360
rect 42064 21344 42116 21350
rect 42260 21298 42288 21655
rect 42064 21286 42116 21292
rect 41880 20596 41932 20602
rect 41880 20538 41932 20544
rect 41972 20596 42024 20602
rect 41972 20538 42024 20544
rect 42076 20466 42104 21286
rect 42168 21270 42288 21298
rect 42064 20460 42116 20466
rect 42064 20402 42116 20408
rect 42064 20052 42116 20058
rect 42064 19994 42116 20000
rect 41880 19848 41932 19854
rect 41880 19790 41932 19796
rect 41892 19514 41920 19790
rect 42076 19786 42104 19994
rect 42064 19780 42116 19786
rect 42064 19722 42116 19728
rect 41880 19508 41932 19514
rect 41880 19450 41932 19456
rect 41708 19306 41828 19334
rect 41708 19258 41736 19306
rect 41972 19304 42024 19310
rect 41970 19272 41972 19281
rect 42024 19272 42026 19281
rect 41708 19230 41828 19258
rect 41696 19168 41748 19174
rect 41602 19136 41658 19145
rect 41696 19110 41748 19116
rect 41602 19071 41658 19080
rect 41604 18828 41656 18834
rect 41604 18770 41656 18776
rect 41616 18630 41644 18770
rect 41708 18630 41736 19110
rect 41604 18624 41656 18630
rect 41604 18566 41656 18572
rect 41696 18624 41748 18630
rect 41696 18566 41748 18572
rect 41524 18278 41736 18306
rect 41420 18216 41472 18222
rect 41512 18216 41564 18222
rect 41420 18158 41472 18164
rect 41510 18184 41512 18193
rect 41604 18216 41656 18222
rect 41564 18184 41566 18193
rect 41604 18158 41656 18164
rect 41510 18119 41566 18128
rect 41144 18022 41196 18028
rect 41234 18048 41290 18057
rect 41156 17270 41184 18022
rect 41234 17983 41290 17992
rect 41512 17808 41564 17814
rect 41512 17750 41564 17756
rect 41144 17264 41196 17270
rect 41144 17206 41196 17212
rect 41236 17196 41288 17202
rect 41236 17138 41288 17144
rect 41144 16108 41196 16114
rect 41144 16050 41196 16056
rect 41156 15337 41184 16050
rect 41142 15328 41198 15337
rect 41142 15263 41198 15272
rect 41248 14793 41276 17138
rect 41524 17134 41552 17750
rect 41512 17128 41564 17134
rect 41340 17088 41512 17116
rect 41340 16794 41368 17088
rect 41512 17070 41564 17076
rect 41420 16992 41472 16998
rect 41420 16934 41472 16940
rect 41328 16788 41380 16794
rect 41328 16730 41380 16736
rect 41326 16552 41382 16561
rect 41326 16487 41382 16496
rect 41340 16250 41368 16487
rect 41328 16244 41380 16250
rect 41328 16186 41380 16192
rect 41328 16040 41380 16046
rect 41328 15982 41380 15988
rect 41340 15638 41368 15982
rect 41432 15910 41460 16934
rect 41420 15904 41472 15910
rect 41420 15846 41472 15852
rect 41328 15632 41380 15638
rect 41328 15574 41380 15580
rect 41234 14784 41290 14793
rect 41234 14719 41290 14728
rect 41340 13977 41368 15574
rect 41512 14408 41564 14414
rect 41512 14350 41564 14356
rect 41524 14074 41552 14350
rect 41512 14068 41564 14074
rect 41512 14010 41564 14016
rect 41326 13968 41382 13977
rect 41326 13903 41382 13912
rect 41234 13696 41290 13705
rect 41234 13631 41290 13640
rect 41144 12844 41196 12850
rect 41144 12786 41196 12792
rect 41156 12646 41184 12786
rect 41144 12640 41196 12646
rect 41144 12582 41196 12588
rect 41156 12238 41184 12582
rect 41248 12434 41276 13631
rect 41420 13252 41472 13258
rect 41420 13194 41472 13200
rect 41248 12406 41368 12434
rect 41144 12232 41196 12238
rect 41144 12174 41196 12180
rect 41144 11144 41196 11150
rect 41144 11086 41196 11092
rect 41156 10266 41184 11086
rect 41144 10260 41196 10266
rect 41144 10202 41196 10208
rect 41236 9512 41288 9518
rect 41236 9454 41288 9460
rect 41248 8566 41276 9454
rect 41236 8560 41288 8566
rect 41236 8502 41288 8508
rect 41340 8378 41368 12406
rect 41432 12374 41460 13194
rect 41420 12368 41472 12374
rect 41420 12310 41472 12316
rect 41420 12232 41472 12238
rect 41420 12174 41472 12180
rect 41432 11898 41460 12174
rect 41420 11892 41472 11898
rect 41420 11834 41472 11840
rect 41512 11756 41564 11762
rect 41512 11698 41564 11704
rect 41418 9616 41474 9625
rect 41418 9551 41420 9560
rect 41472 9551 41474 9560
rect 41420 9522 41472 9528
rect 41248 8362 41368 8378
rect 41248 8356 41380 8362
rect 41248 8350 41328 8356
rect 41248 8022 41276 8350
rect 41328 8298 41380 8304
rect 41420 8288 41472 8294
rect 41340 8236 41420 8242
rect 41340 8230 41472 8236
rect 41524 8242 41552 11698
rect 41616 11082 41644 18158
rect 41708 16289 41736 18278
rect 41694 16280 41750 16289
rect 41694 16215 41750 16224
rect 41694 15872 41750 15881
rect 41694 15807 41750 15816
rect 41708 15434 41736 15807
rect 41696 15428 41748 15434
rect 41696 15370 41748 15376
rect 41708 13870 41736 15370
rect 41696 13864 41748 13870
rect 41696 13806 41748 13812
rect 41696 13320 41748 13326
rect 41696 13262 41748 13268
rect 41708 12986 41736 13262
rect 41696 12980 41748 12986
rect 41696 12922 41748 12928
rect 41696 11620 41748 11626
rect 41696 11562 41748 11568
rect 41604 11076 41656 11082
rect 41604 11018 41656 11024
rect 41602 10976 41658 10985
rect 41602 10911 41658 10920
rect 41616 8378 41644 10911
rect 41708 8650 41736 11562
rect 41800 11506 41828 19230
rect 41970 19207 42026 19216
rect 41972 19168 42024 19174
rect 41878 19136 41934 19145
rect 41972 19110 42024 19116
rect 41878 19071 41934 19080
rect 41892 16522 41920 19071
rect 41984 18465 42012 19110
rect 42062 19000 42118 19009
rect 42168 18986 42196 21270
rect 42248 20528 42300 20534
rect 42248 20470 42300 20476
rect 42260 20058 42288 20470
rect 42248 20052 42300 20058
rect 42248 19994 42300 20000
rect 42248 19168 42300 19174
rect 42246 19136 42248 19145
rect 42300 19136 42302 19145
rect 42246 19071 42302 19080
rect 42352 18986 42380 21950
rect 42118 18958 42196 18986
rect 42260 18958 42380 18986
rect 42062 18935 42118 18944
rect 41970 18456 42026 18465
rect 41970 18391 42026 18400
rect 41970 17912 42026 17921
rect 41970 17847 42026 17856
rect 41984 16658 42012 17847
rect 41972 16652 42024 16658
rect 41972 16594 42024 16600
rect 41880 16516 41932 16522
rect 41880 16458 41932 16464
rect 42076 16046 42104 18935
rect 42260 18766 42288 18958
rect 42156 18760 42208 18766
rect 42156 18702 42208 18708
rect 42248 18760 42300 18766
rect 42248 18702 42300 18708
rect 42338 18728 42394 18737
rect 42168 18465 42196 18702
rect 42260 18601 42288 18702
rect 42338 18663 42394 18672
rect 42246 18592 42302 18601
rect 42246 18527 42302 18536
rect 42154 18456 42210 18465
rect 42154 18391 42210 18400
rect 42168 18358 42196 18391
rect 42156 18352 42208 18358
rect 42156 18294 42208 18300
rect 42154 18184 42210 18193
rect 42154 18119 42210 18128
rect 42168 17649 42196 18119
rect 42352 18086 42380 18663
rect 42340 18080 42392 18086
rect 42340 18022 42392 18028
rect 42248 17672 42300 17678
rect 42154 17640 42210 17649
rect 42352 17649 42380 18022
rect 42248 17614 42300 17620
rect 42338 17640 42394 17649
rect 42154 17575 42210 17584
rect 42168 17202 42196 17575
rect 42156 17196 42208 17202
rect 42156 17138 42208 17144
rect 42260 16794 42288 17614
rect 42338 17575 42394 17584
rect 42248 16788 42300 16794
rect 42248 16730 42300 16736
rect 42248 16448 42300 16454
rect 42248 16390 42300 16396
rect 42064 16040 42116 16046
rect 42064 15982 42116 15988
rect 41880 15904 41932 15910
rect 41880 15846 41932 15852
rect 41892 14090 41920 15846
rect 42260 15502 42288 16390
rect 42340 16040 42392 16046
rect 42340 15982 42392 15988
rect 42248 15496 42300 15502
rect 42248 15438 42300 15444
rect 42154 15328 42210 15337
rect 42154 15263 42210 15272
rect 41972 14816 42024 14822
rect 41972 14758 42024 14764
rect 42064 14816 42116 14822
rect 42064 14758 42116 14764
rect 41984 14278 42012 14758
rect 42076 14618 42104 14758
rect 42064 14612 42116 14618
rect 42064 14554 42116 14560
rect 41972 14272 42024 14278
rect 41972 14214 42024 14220
rect 41892 14062 42012 14090
rect 41880 12776 41932 12782
rect 41880 12718 41932 12724
rect 41892 11898 41920 12718
rect 41880 11892 41932 11898
rect 41880 11834 41932 11840
rect 41800 11478 41920 11506
rect 41788 11348 41840 11354
rect 41788 11290 41840 11296
rect 41800 8809 41828 11290
rect 41892 11286 41920 11478
rect 41880 11280 41932 11286
rect 41880 11222 41932 11228
rect 41984 11218 42012 14062
rect 42062 13288 42118 13297
rect 42062 13223 42118 13232
rect 42076 12322 42104 13223
rect 42168 12442 42196 15263
rect 42156 12436 42208 12442
rect 42156 12378 42208 12384
rect 42076 12294 42288 12322
rect 42062 12200 42118 12209
rect 42062 12135 42118 12144
rect 41972 11212 42024 11218
rect 41972 11154 42024 11160
rect 42076 11150 42104 12135
rect 42156 11756 42208 11762
rect 42156 11698 42208 11704
rect 42064 11144 42116 11150
rect 42064 11086 42116 11092
rect 42076 10810 42104 11086
rect 42064 10804 42116 10810
rect 42064 10746 42116 10752
rect 42168 10606 42196 11698
rect 41880 10600 41932 10606
rect 41880 10542 41932 10548
rect 42156 10600 42208 10606
rect 42156 10542 42208 10548
rect 41786 8800 41842 8809
rect 41786 8735 41842 8744
rect 41708 8622 41828 8650
rect 41616 8350 41736 8378
rect 41340 8214 41460 8230
rect 41524 8214 41644 8242
rect 40868 8016 40920 8022
rect 40868 7958 40920 7964
rect 41052 8016 41104 8022
rect 41052 7958 41104 7964
rect 41236 8016 41288 8022
rect 41236 7958 41288 7964
rect 41064 7886 41092 7958
rect 41052 7880 41104 7886
rect 41248 7857 41276 7958
rect 41052 7822 41104 7828
rect 41234 7848 41290 7857
rect 41340 7834 41368 8214
rect 41510 8120 41566 8129
rect 41510 8055 41566 8064
rect 41340 7806 41460 7834
rect 41234 7783 41290 7792
rect 40776 7472 40828 7478
rect 40776 7414 40828 7420
rect 41432 5273 41460 7806
rect 41524 7750 41552 8055
rect 41512 7744 41564 7750
rect 41512 7686 41564 7692
rect 41524 5642 41552 7686
rect 41616 6089 41644 8214
rect 41708 8022 41736 8350
rect 41696 8016 41748 8022
rect 41696 7958 41748 7964
rect 41800 6934 41828 8622
rect 41788 6928 41840 6934
rect 41788 6870 41840 6876
rect 41892 6118 41920 10542
rect 42064 10124 42116 10130
rect 41984 10084 42064 10112
rect 41984 9926 42012 10084
rect 42064 10066 42116 10072
rect 41972 9920 42024 9926
rect 41972 9862 42024 9868
rect 42064 9920 42116 9926
rect 42064 9862 42116 9868
rect 41972 8968 42024 8974
rect 41972 8910 42024 8916
rect 41984 8838 42012 8910
rect 41972 8832 42024 8838
rect 41972 8774 42024 8780
rect 41984 8022 42012 8774
rect 42076 8362 42104 9862
rect 42154 8664 42210 8673
rect 42154 8599 42210 8608
rect 42168 8498 42196 8599
rect 42156 8492 42208 8498
rect 42156 8434 42208 8440
rect 42064 8356 42116 8362
rect 42064 8298 42116 8304
rect 42168 8022 42196 8434
rect 41972 8016 42024 8022
rect 41972 7958 42024 7964
rect 42156 8016 42208 8022
rect 42156 7958 42208 7964
rect 42260 7410 42288 12294
rect 42352 8634 42380 15982
rect 42444 14822 42472 22494
rect 42536 21690 42564 25162
rect 42800 24744 42852 24750
rect 42800 24686 42852 24692
rect 42812 24410 42840 24686
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 42800 24404 42852 24410
rect 42800 24346 42852 24352
rect 42706 24304 42762 24313
rect 42706 24239 42762 24248
rect 42720 24206 42748 24239
rect 42708 24200 42760 24206
rect 42708 24142 42760 24148
rect 42708 23520 42760 23526
rect 42708 23462 42760 23468
rect 42720 23361 42748 23462
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42706 23352 42762 23361
rect 42950 23355 43258 23364
rect 42706 23287 42762 23296
rect 42616 23180 42668 23186
rect 42616 23122 42668 23128
rect 42524 21684 42576 21690
rect 42524 21626 42576 21632
rect 42524 21548 42576 21554
rect 42524 21490 42576 21496
rect 42536 21418 42564 21490
rect 42524 21412 42576 21418
rect 42524 21354 42576 21360
rect 42628 21060 42656 23122
rect 43258 23080 43314 23089
rect 43258 23015 43260 23024
rect 43312 23015 43314 23024
rect 43260 22986 43312 22992
rect 43272 22710 43300 22986
rect 43260 22704 43312 22710
rect 43260 22646 43312 22652
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 43364 22098 43392 26046
rect 43534 26007 43590 26016
rect 43444 24880 43496 24886
rect 43444 24822 43496 24828
rect 43456 23186 43484 24822
rect 43444 23180 43496 23186
rect 43444 23122 43496 23128
rect 43352 22092 43404 22098
rect 43352 22034 43404 22040
rect 42892 22024 42944 22030
rect 42892 21966 42944 21972
rect 42904 21706 42932 21966
rect 42720 21678 42932 21706
rect 42720 21185 42748 21678
rect 42800 21548 42852 21554
rect 42800 21490 42852 21496
rect 42812 21321 42840 21490
rect 42798 21312 42854 21321
rect 42798 21247 42854 21256
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42706 21176 42762 21185
rect 42950 21179 43258 21188
rect 42706 21111 42762 21120
rect 42628 21032 42748 21060
rect 42524 21004 42576 21010
rect 42524 20946 42576 20952
rect 42536 18873 42564 20946
rect 42616 19508 42668 19514
rect 42616 19450 42668 19456
rect 42628 19378 42656 19450
rect 42616 19372 42668 19378
rect 42616 19314 42668 19320
rect 42616 19236 42668 19242
rect 42616 19178 42668 19184
rect 42522 18864 42578 18873
rect 42628 18834 42656 19178
rect 42522 18799 42578 18808
rect 42616 18828 42668 18834
rect 42536 15910 42564 18799
rect 42616 18770 42668 18776
rect 42616 18624 42668 18630
rect 42616 18566 42668 18572
rect 42628 18290 42656 18566
rect 42720 18358 42748 21032
rect 43456 21026 43484 23122
rect 43364 20998 43484 21026
rect 42984 20800 43036 20806
rect 42984 20742 43036 20748
rect 42996 20466 43024 20742
rect 42984 20460 43036 20466
rect 42984 20402 43036 20408
rect 42800 20256 42852 20262
rect 42800 20198 42852 20204
rect 42812 19718 42840 20198
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 43364 19938 43392 20998
rect 43444 20936 43496 20942
rect 43444 20878 43496 20884
rect 43456 20058 43484 20878
rect 43548 20482 43576 26007
rect 44180 25696 44232 25702
rect 44180 25638 44232 25644
rect 44086 25256 44142 25265
rect 44086 25191 44142 25200
rect 44100 24342 44128 25191
rect 44088 24336 44140 24342
rect 44088 24278 44140 24284
rect 43720 24064 43772 24070
rect 43720 24006 43772 24012
rect 43812 24064 43864 24070
rect 43812 24006 43864 24012
rect 43732 23730 43760 24006
rect 43720 23724 43772 23730
rect 43720 23666 43772 23672
rect 43824 23202 43852 24006
rect 43902 23760 43958 23769
rect 43902 23695 43958 23704
rect 43640 23174 43852 23202
rect 43640 22030 43668 23174
rect 43720 23044 43772 23050
rect 43720 22986 43772 22992
rect 43732 22817 43760 22986
rect 43718 22808 43774 22817
rect 43718 22743 43774 22752
rect 43720 22636 43772 22642
rect 43720 22578 43772 22584
rect 43628 22024 43680 22030
rect 43628 21966 43680 21972
rect 43732 21894 43760 22578
rect 43812 22568 43864 22574
rect 43812 22510 43864 22516
rect 43720 21888 43772 21894
rect 43720 21830 43772 21836
rect 43720 21548 43772 21554
rect 43720 21490 43772 21496
rect 43732 20602 43760 21490
rect 43720 20596 43772 20602
rect 43720 20538 43772 20544
rect 43548 20454 43668 20482
rect 43444 20052 43496 20058
rect 43444 19994 43496 20000
rect 43364 19910 43576 19938
rect 43260 19848 43312 19854
rect 43260 19790 43312 19796
rect 43442 19816 43498 19825
rect 42800 19712 42852 19718
rect 42800 19654 42852 19660
rect 43272 19514 43300 19790
rect 43442 19751 43498 19760
rect 43352 19712 43404 19718
rect 43352 19654 43404 19660
rect 43260 19508 43312 19514
rect 43260 19450 43312 19456
rect 42800 19304 42852 19310
rect 42800 19246 42852 19252
rect 42812 18426 42840 19246
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 42800 18420 42852 18426
rect 42800 18362 42852 18368
rect 42708 18352 42760 18358
rect 42708 18294 42760 18300
rect 42616 18284 42668 18290
rect 42616 18226 42668 18232
rect 42800 18080 42852 18086
rect 42800 18022 42852 18028
rect 42616 17536 42668 17542
rect 42616 17478 42668 17484
rect 42628 17202 42656 17478
rect 42812 17241 42840 18022
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 43364 17921 43392 19654
rect 43456 19514 43484 19751
rect 43444 19508 43496 19514
rect 43444 19450 43496 19456
rect 43350 17912 43406 17921
rect 43350 17847 43406 17856
rect 43352 17536 43404 17542
rect 43352 17478 43404 17484
rect 42890 17368 42946 17377
rect 42890 17303 42946 17312
rect 42798 17232 42854 17241
rect 42616 17196 42668 17202
rect 42798 17167 42854 17176
rect 42616 17138 42668 17144
rect 42904 16980 42932 17303
rect 43260 17128 43312 17134
rect 43258 17096 43260 17105
rect 43312 17096 43314 17105
rect 43258 17031 43314 17040
rect 42812 16952 42932 16980
rect 42812 16833 42840 16952
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42798 16824 42854 16833
rect 42950 16827 43258 16836
rect 42798 16759 42854 16768
rect 43364 16590 43392 17478
rect 43352 16584 43404 16590
rect 43352 16526 43404 16532
rect 42708 16176 42760 16182
rect 42708 16118 42760 16124
rect 42616 16108 42668 16114
rect 42616 16050 42668 16056
rect 42628 16017 42656 16050
rect 42614 16008 42670 16017
rect 42614 15943 42670 15952
rect 42524 15904 42576 15910
rect 42524 15846 42576 15852
rect 42720 15638 42748 16118
rect 42800 15904 42852 15910
rect 42800 15846 42852 15852
rect 42708 15632 42760 15638
rect 42708 15574 42760 15580
rect 42812 15094 42840 15846
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 43444 15428 43496 15434
rect 43444 15370 43496 15376
rect 42800 15088 42852 15094
rect 42800 15030 42852 15036
rect 42432 14816 42484 14822
rect 42432 14758 42484 14764
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42798 14648 42854 14657
rect 42950 14651 43258 14660
rect 42798 14583 42800 14592
rect 42852 14583 42854 14592
rect 42800 14554 42852 14560
rect 43166 14512 43222 14521
rect 43166 14447 43168 14456
rect 43220 14447 43222 14456
rect 43168 14418 43220 14424
rect 43260 14408 43312 14414
rect 43260 14350 43312 14356
rect 42798 14104 42854 14113
rect 43272 14074 43300 14350
rect 42798 14039 42854 14048
rect 43260 14068 43312 14074
rect 42706 13968 42762 13977
rect 42706 13903 42708 13912
rect 42760 13903 42762 13912
rect 42708 13874 42760 13880
rect 42616 13796 42668 13802
rect 42616 13738 42668 13744
rect 42524 13728 42576 13734
rect 42524 13670 42576 13676
rect 42432 12436 42484 12442
rect 42432 12378 42484 12384
rect 42444 11898 42472 12378
rect 42432 11892 42484 11898
rect 42432 11834 42484 11840
rect 42430 11792 42486 11801
rect 42430 11727 42486 11736
rect 42444 11558 42472 11727
rect 42432 11552 42484 11558
rect 42432 11494 42484 11500
rect 42430 10840 42486 10849
rect 42430 10775 42486 10784
rect 42444 9042 42472 10775
rect 42536 9518 42564 13670
rect 42628 12850 42656 13738
rect 42812 13682 42840 14039
rect 43260 14010 43312 14016
rect 43352 14000 43404 14006
rect 43352 13942 43404 13948
rect 42720 13654 42840 13682
rect 42720 13410 42748 13654
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42798 13560 42854 13569
rect 42950 13563 43258 13572
rect 42798 13495 42800 13504
rect 42852 13495 42854 13504
rect 42800 13466 42852 13472
rect 42720 13382 42840 13410
rect 42706 12880 42762 12889
rect 42616 12844 42668 12850
rect 42706 12815 42762 12824
rect 42616 12786 42668 12792
rect 42614 11384 42670 11393
rect 42720 11354 42748 12815
rect 42614 11319 42670 11328
rect 42708 11348 42760 11354
rect 42628 10606 42656 11319
rect 42708 11290 42760 11296
rect 42708 11076 42760 11082
rect 42708 11018 42760 11024
rect 42616 10600 42668 10606
rect 42616 10542 42668 10548
rect 42614 10160 42670 10169
rect 42614 10095 42670 10104
rect 42628 10062 42656 10095
rect 42616 10056 42668 10062
rect 42616 9998 42668 10004
rect 42720 9518 42748 11018
rect 42524 9512 42576 9518
rect 42524 9454 42576 9460
rect 42616 9512 42668 9518
rect 42616 9454 42668 9460
rect 42708 9512 42760 9518
rect 42708 9454 42760 9460
rect 42432 9036 42484 9042
rect 42432 8978 42484 8984
rect 42340 8628 42392 8634
rect 42340 8570 42392 8576
rect 42628 8514 42656 9454
rect 42628 8486 42748 8514
rect 42720 8430 42748 8486
rect 42524 8424 42576 8430
rect 42524 8366 42576 8372
rect 42708 8424 42760 8430
rect 42708 8366 42760 8372
rect 42248 7404 42300 7410
rect 42248 7346 42300 7352
rect 42536 6186 42564 8366
rect 42616 7812 42668 7818
rect 42616 7754 42668 7760
rect 42628 6934 42656 7754
rect 42616 6928 42668 6934
rect 42616 6870 42668 6876
rect 42524 6180 42576 6186
rect 42524 6122 42576 6128
rect 41880 6112 41932 6118
rect 41602 6080 41658 6089
rect 41880 6054 41932 6060
rect 41602 6015 41658 6024
rect 41512 5636 41564 5642
rect 41512 5578 41564 5584
rect 41418 5264 41474 5273
rect 41418 5199 41474 5208
rect 42720 4729 42748 8366
rect 42812 7342 42840 13382
rect 43260 13320 43312 13326
rect 43260 13262 43312 13268
rect 43272 12986 43300 13262
rect 43260 12980 43312 12986
rect 43260 12922 43312 12928
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 43076 12368 43128 12374
rect 43076 12310 43128 12316
rect 42984 12096 43036 12102
rect 42984 12038 43036 12044
rect 42996 11694 43024 12038
rect 42984 11688 43036 11694
rect 42984 11630 43036 11636
rect 43088 11626 43116 12310
rect 43076 11620 43128 11626
rect 43076 11562 43128 11568
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 43258 11248 43314 11257
rect 43258 11183 43314 11192
rect 43272 11082 43300 11183
rect 43364 11150 43392 13942
rect 43456 11354 43484 15370
rect 43548 12424 43576 19910
rect 43640 12617 43668 20454
rect 43718 19408 43774 19417
rect 43718 19343 43774 19352
rect 43732 18834 43760 19343
rect 43720 18828 43772 18834
rect 43720 18770 43772 18776
rect 43720 18624 43772 18630
rect 43720 18566 43772 18572
rect 43732 18290 43760 18566
rect 43720 18284 43772 18290
rect 43720 18226 43772 18232
rect 43824 18193 43852 22510
rect 43916 18766 43944 23695
rect 44192 23322 44220 25638
rect 44456 25560 44508 25566
rect 44456 25502 44508 25508
rect 44364 25424 44416 25430
rect 44364 25366 44416 25372
rect 44270 24984 44326 24993
rect 44270 24919 44326 24928
rect 44180 23316 44232 23322
rect 44180 23258 44232 23264
rect 43996 22976 44048 22982
rect 43996 22918 44048 22924
rect 44008 18986 44036 22918
rect 44086 22808 44142 22817
rect 44086 22743 44142 22752
rect 44100 20262 44128 22743
rect 44180 22500 44232 22506
rect 44180 22442 44232 22448
rect 44192 21962 44220 22442
rect 44180 21956 44232 21962
rect 44180 21898 44232 21904
rect 44284 21078 44312 24919
rect 44376 23730 44404 25366
rect 44364 23724 44416 23730
rect 44364 23666 44416 23672
rect 44468 23118 44496 25502
rect 44546 24712 44602 24721
rect 44546 24647 44602 24656
rect 44560 23730 44588 24647
rect 44548 23724 44600 23730
rect 44548 23666 44600 23672
rect 44456 23112 44508 23118
rect 44454 23080 44456 23089
rect 44508 23080 44510 23089
rect 44454 23015 44510 23024
rect 44456 22500 44508 22506
rect 44456 22442 44508 22448
rect 44468 22098 44496 22442
rect 44456 22092 44508 22098
rect 44456 22034 44508 22040
rect 44548 22092 44600 22098
rect 44548 22034 44600 22040
rect 44560 21978 44588 22034
rect 44468 21950 44588 21978
rect 44468 21622 44496 21950
rect 44548 21888 44600 21894
rect 44548 21830 44600 21836
rect 44456 21616 44508 21622
rect 44456 21558 44508 21564
rect 44272 21072 44324 21078
rect 44272 21014 44324 21020
rect 44180 20800 44232 20806
rect 44180 20742 44232 20748
rect 44088 20256 44140 20262
rect 44088 20198 44140 20204
rect 44192 19854 44220 20742
rect 44364 20392 44416 20398
rect 44362 20360 44364 20369
rect 44416 20360 44418 20369
rect 44362 20295 44418 20304
rect 44272 20256 44324 20262
rect 44560 20244 44588 21830
rect 44652 21457 44680 26302
rect 44730 26200 44786 26302
rect 45374 26200 45430 27000
rect 45650 26344 45706 26353
rect 45650 26279 45706 26288
rect 45192 25900 45244 25906
rect 45192 25842 45244 25848
rect 45006 25528 45062 25537
rect 45006 25463 45062 25472
rect 44732 23724 44784 23730
rect 44784 23684 44956 23712
rect 44732 23666 44784 23672
rect 44824 22976 44876 22982
rect 44824 22918 44876 22924
rect 44836 22409 44864 22918
rect 44822 22400 44878 22409
rect 44822 22335 44878 22344
rect 44824 22228 44876 22234
rect 44824 22170 44876 22176
rect 44732 22024 44784 22030
rect 44732 21966 44784 21972
rect 44638 21448 44694 21457
rect 44638 21383 44694 21392
rect 44652 21185 44680 21383
rect 44638 21176 44694 21185
rect 44638 21111 44694 21120
rect 44744 20806 44772 21966
rect 44836 21554 44864 22170
rect 44824 21548 44876 21554
rect 44824 21490 44876 21496
rect 44732 20800 44784 20806
rect 44732 20742 44784 20748
rect 44272 20198 44324 20204
rect 44376 20216 44588 20244
rect 44284 20058 44312 20198
rect 44272 20052 44324 20058
rect 44272 19994 44324 20000
rect 44180 19848 44232 19854
rect 44180 19790 44232 19796
rect 44088 19440 44140 19446
rect 44088 19382 44140 19388
rect 44100 19310 44128 19382
rect 44088 19304 44140 19310
rect 44088 19246 44140 19252
rect 44008 18970 44220 18986
rect 44008 18964 44232 18970
rect 44008 18958 44180 18964
rect 44180 18906 44232 18912
rect 44284 18873 44312 19994
rect 44376 19553 44404 20216
rect 44456 19780 44508 19786
rect 44456 19722 44508 19728
rect 44362 19544 44418 19553
rect 44362 19479 44418 19488
rect 44270 18864 44326 18873
rect 44270 18799 44326 18808
rect 43904 18760 43956 18766
rect 44376 18714 44404 19479
rect 44468 19310 44496 19722
rect 44456 19304 44508 19310
rect 44456 19246 44508 19252
rect 44744 19145 44772 20742
rect 44928 20641 44956 23684
rect 45020 22506 45048 25463
rect 45204 23866 45232 25842
rect 45192 23860 45244 23866
rect 45192 23802 45244 23808
rect 45190 23624 45246 23633
rect 45190 23559 45246 23568
rect 45100 23180 45152 23186
rect 45100 23122 45152 23128
rect 45112 22642 45140 23122
rect 45204 23118 45232 23559
rect 45388 23497 45416 26200
rect 45560 25968 45612 25974
rect 45560 25910 45612 25916
rect 45468 23792 45520 23798
rect 45468 23734 45520 23740
rect 45374 23488 45430 23497
rect 45374 23423 45430 23432
rect 45192 23112 45244 23118
rect 45192 23054 45244 23060
rect 45100 22636 45152 22642
rect 45100 22578 45152 22584
rect 45008 22500 45060 22506
rect 45008 22442 45060 22448
rect 45284 22500 45336 22506
rect 45284 22442 45336 22448
rect 45192 22432 45244 22438
rect 45192 22374 45244 22380
rect 45204 22030 45232 22374
rect 45192 22024 45244 22030
rect 45192 21966 45244 21972
rect 45006 21856 45062 21865
rect 45006 21791 45062 21800
rect 45020 20942 45048 21791
rect 45192 21412 45244 21418
rect 45192 21354 45244 21360
rect 45008 20936 45060 20942
rect 45008 20878 45060 20884
rect 45100 20936 45152 20942
rect 45100 20878 45152 20884
rect 44914 20632 44970 20641
rect 44914 20567 44970 20576
rect 44916 20392 44968 20398
rect 44916 20334 44968 20340
rect 44730 19136 44786 19145
rect 44730 19071 44786 19080
rect 44928 18986 44956 20334
rect 43904 18702 43956 18708
rect 44284 18686 44404 18714
rect 44652 18958 44956 18986
rect 44284 18630 44312 18686
rect 44272 18624 44324 18630
rect 43902 18592 43958 18601
rect 44272 18566 44324 18572
rect 43902 18527 43958 18536
rect 43810 18184 43866 18193
rect 43810 18119 43866 18128
rect 43720 17196 43772 17202
rect 43720 17138 43772 17144
rect 43732 16794 43760 17138
rect 43720 16788 43772 16794
rect 43720 16730 43772 16736
rect 43810 16280 43866 16289
rect 43810 16215 43866 16224
rect 43824 13462 43852 16215
rect 43916 14006 43944 18527
rect 43996 18148 44048 18154
rect 43996 18090 44048 18096
rect 44008 17746 44036 18090
rect 44178 18048 44234 18057
rect 44178 17983 44234 17992
rect 44086 17776 44142 17785
rect 43996 17740 44048 17746
rect 44086 17711 44142 17720
rect 43996 17682 44048 17688
rect 44100 17134 44128 17711
rect 44088 17128 44140 17134
rect 44088 17070 44140 17076
rect 44088 16992 44140 16998
rect 44088 16934 44140 16940
rect 43996 15360 44048 15366
rect 43996 15302 44048 15308
rect 44008 15026 44036 15302
rect 43996 15020 44048 15026
rect 43996 14962 44048 14968
rect 44100 14906 44128 16934
rect 44192 15450 44220 17983
rect 44284 16998 44312 18566
rect 44362 18320 44418 18329
rect 44362 18255 44364 18264
rect 44416 18255 44418 18264
rect 44548 18284 44600 18290
rect 44364 18226 44416 18232
rect 44548 18226 44600 18232
rect 44456 17876 44508 17882
rect 44456 17818 44508 17824
rect 44468 17746 44496 17818
rect 44456 17740 44508 17746
rect 44456 17682 44508 17688
rect 44272 16992 44324 16998
rect 44272 16934 44324 16940
rect 44560 16726 44588 18226
rect 44548 16720 44600 16726
rect 44548 16662 44600 16668
rect 44272 16652 44324 16658
rect 44272 16594 44324 16600
rect 44284 15570 44312 16594
rect 44364 16584 44416 16590
rect 44364 16526 44416 16532
rect 44456 16584 44508 16590
rect 44456 16526 44508 16532
rect 44376 16250 44404 16526
rect 44364 16244 44416 16250
rect 44364 16186 44416 16192
rect 44468 16130 44496 16526
rect 44546 16416 44602 16425
rect 44546 16351 44602 16360
rect 44560 16250 44588 16351
rect 44548 16244 44600 16250
rect 44548 16186 44600 16192
rect 44376 16102 44496 16130
rect 44376 16046 44404 16102
rect 44364 16040 44416 16046
rect 44364 15982 44416 15988
rect 44272 15564 44324 15570
rect 44272 15506 44324 15512
rect 44192 15422 44312 15450
rect 44008 14878 44128 14906
rect 43904 14000 43956 14006
rect 43904 13942 43956 13948
rect 43812 13456 43864 13462
rect 44008 13433 44036 14878
rect 44180 14816 44232 14822
rect 44086 14784 44142 14793
rect 44180 14758 44232 14764
rect 44086 14719 44142 14728
rect 44100 14550 44128 14719
rect 44088 14544 44140 14550
rect 44088 14486 44140 14492
rect 43812 13398 43864 13404
rect 43994 13424 44050 13433
rect 44192 13394 44220 14758
rect 43994 13359 44050 13368
rect 44180 13388 44232 13394
rect 44180 13330 44232 13336
rect 44284 13274 44312 15422
rect 44376 15094 44404 15982
rect 44652 15586 44680 18958
rect 44824 18828 44876 18834
rect 44824 18770 44876 18776
rect 44732 17604 44784 17610
rect 44732 17546 44784 17552
rect 44744 17066 44772 17546
rect 44732 17060 44784 17066
rect 44732 17002 44784 17008
rect 44730 16824 44786 16833
rect 44836 16794 44864 18770
rect 44916 18420 44968 18426
rect 44916 18362 44968 18368
rect 44730 16759 44786 16768
rect 44824 16788 44876 16794
rect 44560 15558 44680 15586
rect 44456 15360 44508 15366
rect 44456 15302 44508 15308
rect 44364 15088 44416 15094
rect 44364 15030 44416 15036
rect 44364 14408 44416 14414
rect 44364 14350 44416 14356
rect 44376 14074 44404 14350
rect 44364 14068 44416 14074
rect 44364 14010 44416 14016
rect 44100 13246 44312 13274
rect 43720 13184 43772 13190
rect 43720 13126 43772 13132
rect 43732 12850 43760 13126
rect 43720 12844 43772 12850
rect 43720 12786 43772 12792
rect 43626 12608 43682 12617
rect 43626 12543 43682 12552
rect 43548 12396 43760 12424
rect 43534 12200 43590 12209
rect 43534 12135 43590 12144
rect 43444 11348 43496 11354
rect 43444 11290 43496 11296
rect 43442 11248 43498 11257
rect 43442 11183 43498 11192
rect 43456 11150 43484 11183
rect 43352 11144 43404 11150
rect 43352 11086 43404 11092
rect 43444 11144 43496 11150
rect 43444 11086 43496 11092
rect 43260 11076 43312 11082
rect 43260 11018 43312 11024
rect 43456 10810 43484 11086
rect 43444 10804 43496 10810
rect 43444 10746 43496 10752
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 43258 10160 43314 10169
rect 43258 10095 43314 10104
rect 42890 9616 42946 9625
rect 43272 9586 43300 10095
rect 42890 9551 42892 9560
rect 42944 9551 42946 9560
rect 43260 9580 43312 9586
rect 42892 9522 42944 9528
rect 43260 9522 43312 9528
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 43548 9058 43576 12135
rect 43732 12050 43760 12396
rect 43996 12096 44048 12102
rect 43732 12022 43944 12050
rect 43996 12038 44048 12044
rect 43628 10736 43680 10742
rect 43628 10678 43680 10684
rect 43364 9030 43576 9058
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 42890 7984 42946 7993
rect 42890 7919 42946 7928
rect 42904 7886 42932 7919
rect 42892 7880 42944 7886
rect 43364 7834 43392 9030
rect 43536 8968 43588 8974
rect 43534 8936 43536 8945
rect 43588 8936 43590 8945
rect 43534 8871 43590 8880
rect 43442 8800 43498 8809
rect 43442 8735 43498 8744
rect 43456 8430 43484 8735
rect 43444 8424 43496 8430
rect 43444 8366 43496 8372
rect 42892 7822 42944 7828
rect 42996 7806 43392 7834
rect 42800 7336 42852 7342
rect 42800 7278 42852 7284
rect 42996 7206 43024 7806
rect 43168 7744 43220 7750
rect 43168 7686 43220 7692
rect 43352 7744 43404 7750
rect 43352 7686 43404 7692
rect 43180 7206 43208 7686
rect 43364 7478 43392 7686
rect 43352 7472 43404 7478
rect 43352 7414 43404 7420
rect 42984 7200 43036 7206
rect 42984 7142 43036 7148
rect 43168 7200 43220 7206
rect 43168 7142 43220 7148
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 43350 6896 43406 6905
rect 43350 6831 43352 6840
rect 43404 6831 43406 6840
rect 43352 6802 43404 6808
rect 43260 6656 43312 6662
rect 43260 6598 43312 6604
rect 43272 6390 43300 6598
rect 43260 6384 43312 6390
rect 43260 6326 43312 6332
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 43456 5137 43484 8366
rect 43536 7880 43588 7886
rect 43536 7822 43588 7828
rect 43548 7478 43576 7822
rect 43536 7472 43588 7478
rect 43536 7414 43588 7420
rect 43534 7032 43590 7041
rect 43534 6967 43590 6976
rect 43548 6798 43576 6967
rect 43640 6866 43668 10678
rect 43720 10600 43772 10606
rect 43720 10542 43772 10548
rect 43732 10266 43760 10542
rect 43720 10260 43772 10266
rect 43720 10202 43772 10208
rect 43812 10056 43864 10062
rect 43812 9998 43864 10004
rect 43720 9580 43772 9586
rect 43720 9522 43772 9528
rect 43732 9058 43760 9522
rect 43824 9178 43852 9998
rect 43916 9674 43944 12022
rect 44008 10538 44036 12038
rect 44100 10674 44128 13246
rect 44180 12164 44232 12170
rect 44180 12106 44232 12112
rect 44192 11762 44220 12106
rect 44362 11928 44418 11937
rect 44272 11892 44324 11898
rect 44362 11863 44364 11872
rect 44272 11834 44324 11840
rect 44416 11863 44418 11872
rect 44364 11834 44416 11840
rect 44180 11756 44232 11762
rect 44180 11698 44232 11704
rect 44178 11656 44234 11665
rect 44178 11591 44234 11600
rect 44192 11218 44220 11591
rect 44284 11558 44312 11834
rect 44272 11552 44324 11558
rect 44272 11494 44324 11500
rect 44180 11212 44232 11218
rect 44180 11154 44232 11160
rect 44088 10668 44140 10674
rect 44088 10610 44140 10616
rect 43996 10532 44048 10538
rect 43996 10474 44048 10480
rect 44088 10464 44140 10470
rect 44088 10406 44140 10412
rect 43916 9646 44036 9674
rect 43904 9512 43956 9518
rect 43904 9454 43956 9460
rect 43812 9172 43864 9178
rect 43812 9114 43864 9120
rect 43732 9030 43852 9058
rect 43720 8832 43772 8838
rect 43720 8774 43772 8780
rect 43732 7818 43760 8774
rect 43824 8566 43852 9030
rect 43916 8838 43944 9454
rect 43904 8832 43956 8838
rect 43904 8774 43956 8780
rect 44008 8786 44036 9646
rect 44100 8974 44128 10406
rect 44468 10062 44496 15302
rect 44560 14074 44588 15558
rect 44640 15496 44692 15502
rect 44638 15464 44640 15473
rect 44692 15464 44694 15473
rect 44638 15399 44694 15408
rect 44640 15088 44692 15094
rect 44640 15030 44692 15036
rect 44548 14068 44600 14074
rect 44548 14010 44600 14016
rect 44652 13870 44680 15030
rect 44640 13864 44692 13870
rect 44640 13806 44692 13812
rect 44548 13388 44600 13394
rect 44548 13330 44600 13336
rect 44560 11937 44588 13330
rect 44652 12646 44680 13806
rect 44744 12918 44772 16759
rect 44824 16730 44876 16736
rect 44824 16108 44876 16114
rect 44824 16050 44876 16056
rect 44836 15162 44864 16050
rect 44824 15156 44876 15162
rect 44824 15098 44876 15104
rect 44822 13696 44878 13705
rect 44822 13631 44878 13640
rect 44732 12912 44784 12918
rect 44732 12854 44784 12860
rect 44732 12708 44784 12714
rect 44732 12650 44784 12656
rect 44640 12640 44692 12646
rect 44640 12582 44692 12588
rect 44546 11928 44602 11937
rect 44546 11863 44602 11872
rect 44548 11348 44600 11354
rect 44548 11290 44600 11296
rect 44560 11150 44588 11290
rect 44548 11144 44600 11150
rect 44548 11086 44600 11092
rect 44548 11008 44600 11014
rect 44548 10950 44600 10956
rect 44560 10674 44588 10950
rect 44548 10668 44600 10674
rect 44548 10610 44600 10616
rect 44456 10056 44508 10062
rect 44456 9998 44508 10004
rect 44560 9654 44588 10610
rect 44548 9648 44600 9654
rect 44178 9616 44234 9625
rect 44548 9590 44600 9596
rect 44178 9551 44234 9560
rect 44088 8968 44140 8974
rect 44088 8910 44140 8916
rect 43812 8560 43864 8566
rect 43812 8502 43864 8508
rect 43720 7812 43772 7818
rect 43720 7754 43772 7760
rect 43824 6866 43852 8502
rect 43916 8401 43944 8774
rect 44008 8758 44128 8786
rect 43996 8560 44048 8566
rect 43996 8502 44048 8508
rect 43902 8392 43958 8401
rect 43902 8327 43958 8336
rect 44008 8022 44036 8502
rect 43996 8016 44048 8022
rect 43996 7958 44048 7964
rect 44100 7750 44128 8758
rect 44192 8634 44220 9551
rect 44548 9036 44600 9042
rect 44548 8978 44600 8984
rect 44180 8628 44232 8634
rect 44180 8570 44232 8576
rect 44362 8528 44418 8537
rect 44180 8492 44232 8498
rect 44362 8463 44418 8472
rect 44180 8434 44232 8440
rect 44088 7744 44140 7750
rect 44088 7686 44140 7692
rect 44192 7342 44220 8434
rect 44376 7410 44404 8463
rect 44560 7954 44588 8978
rect 44652 8090 44680 12582
rect 44744 11898 44772 12650
rect 44732 11892 44784 11898
rect 44732 11834 44784 11840
rect 44732 11280 44784 11286
rect 44732 11222 44784 11228
rect 44744 11121 44772 11222
rect 44730 11112 44786 11121
rect 44730 11047 44786 11056
rect 44732 10600 44784 10606
rect 44732 10542 44784 10548
rect 44640 8084 44692 8090
rect 44640 8026 44692 8032
rect 44548 7948 44600 7954
rect 44548 7890 44600 7896
rect 44560 7721 44588 7890
rect 44546 7712 44602 7721
rect 44546 7647 44602 7656
rect 44364 7404 44416 7410
rect 44364 7346 44416 7352
rect 44180 7336 44232 7342
rect 44180 7278 44232 7284
rect 44272 7336 44324 7342
rect 44272 7278 44324 7284
rect 43628 6860 43680 6866
rect 43628 6802 43680 6808
rect 43812 6860 43864 6866
rect 43812 6802 43864 6808
rect 43536 6792 43588 6798
rect 43536 6734 43588 6740
rect 43996 6792 44048 6798
rect 43996 6734 44048 6740
rect 44008 6458 44036 6734
rect 44284 6458 44312 7278
rect 44376 6882 44404 7346
rect 44640 7336 44692 7342
rect 44454 7304 44510 7313
rect 44640 7278 44692 7284
rect 44454 7239 44510 7248
rect 44468 7206 44496 7239
rect 44456 7200 44508 7206
rect 44456 7142 44508 7148
rect 44376 6854 44496 6882
rect 44362 6760 44418 6769
rect 44362 6695 44418 6704
rect 44376 6458 44404 6695
rect 44468 6458 44496 6854
rect 43996 6452 44048 6458
rect 43996 6394 44048 6400
rect 44272 6452 44324 6458
rect 44272 6394 44324 6400
rect 44364 6452 44416 6458
rect 44364 6394 44416 6400
rect 44456 6452 44508 6458
rect 44456 6394 44508 6400
rect 44652 5914 44680 7278
rect 44640 5908 44692 5914
rect 44640 5850 44692 5856
rect 43442 5128 43498 5137
rect 43442 5063 43498 5072
rect 44272 5092 44324 5098
rect 44272 5034 44324 5040
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 42706 4720 42762 4729
rect 42706 4655 42762 4664
rect 42800 4548 42852 4554
rect 42800 4490 42852 4496
rect 40500 4004 40552 4010
rect 40500 3946 40552 3952
rect 40408 3528 40460 3534
rect 40408 3470 40460 3476
rect 39396 3052 39448 3058
rect 39396 2994 39448 3000
rect 41328 2508 41380 2514
rect 41328 2450 41380 2456
rect 41340 800 41368 2450
rect 42812 2446 42840 4490
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 43444 3732 43496 3738
rect 43444 3674 43496 3680
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 42800 2440 42852 2446
rect 42800 2382 42852 2388
rect 43456 800 43484 3674
rect 44284 2514 44312 5034
rect 44744 4593 44772 10542
rect 44836 7478 44864 13631
rect 44928 13462 44956 18362
rect 45020 16402 45048 20878
rect 45112 16561 45140 20878
rect 45204 20262 45232 21354
rect 45296 21010 45324 22442
rect 45376 22432 45428 22438
rect 45376 22374 45428 22380
rect 45284 21004 45336 21010
rect 45284 20946 45336 20952
rect 45296 20398 45324 20946
rect 45284 20392 45336 20398
rect 45284 20334 45336 20340
rect 45192 20256 45244 20262
rect 45192 20198 45244 20204
rect 45192 19712 45244 19718
rect 45192 19654 45244 19660
rect 45204 18465 45232 19654
rect 45282 19408 45338 19417
rect 45282 19343 45338 19352
rect 45190 18456 45246 18465
rect 45190 18391 45246 18400
rect 45204 16726 45232 18391
rect 45192 16720 45244 16726
rect 45192 16662 45244 16668
rect 45192 16584 45244 16590
rect 45098 16552 45154 16561
rect 45192 16526 45244 16532
rect 45098 16487 45154 16496
rect 45020 16374 45140 16402
rect 45008 15564 45060 15570
rect 45008 15506 45060 15512
rect 45020 13530 45048 15506
rect 45008 13524 45060 13530
rect 45008 13466 45060 13472
rect 44916 13456 44968 13462
rect 44916 13398 44968 13404
rect 44916 13320 44968 13326
rect 44916 13262 44968 13268
rect 44928 12986 44956 13262
rect 44916 12980 44968 12986
rect 44916 12922 44968 12928
rect 45008 12164 45060 12170
rect 45008 12106 45060 12112
rect 44914 11792 44970 11801
rect 44914 11727 44916 11736
rect 44968 11727 44970 11736
rect 44916 11698 44968 11704
rect 44928 8022 44956 11698
rect 45020 9178 45048 12106
rect 45112 9586 45140 16374
rect 45204 15978 45232 16526
rect 45192 15972 45244 15978
rect 45192 15914 45244 15920
rect 45192 14816 45244 14822
rect 45192 14758 45244 14764
rect 45204 12714 45232 14758
rect 45296 13938 45324 19343
rect 45388 19334 45416 22374
rect 45480 21690 45508 23734
rect 45572 23730 45600 25910
rect 45664 24290 45692 26279
rect 46018 26200 46074 27000
rect 46662 26330 46718 27000
rect 46662 26302 46796 26330
rect 46662 26200 46718 26302
rect 45742 25936 45798 25945
rect 45742 25871 45798 25880
rect 45756 24410 45784 25871
rect 45926 25800 45982 25809
rect 45926 25735 45982 25744
rect 45834 25120 45890 25129
rect 45834 25055 45890 25064
rect 45848 25022 45876 25055
rect 45836 25016 45888 25022
rect 45836 24958 45888 24964
rect 45744 24404 45796 24410
rect 45744 24346 45796 24352
rect 45664 24262 45876 24290
rect 45652 24200 45704 24206
rect 45652 24142 45704 24148
rect 45560 23724 45612 23730
rect 45560 23666 45612 23672
rect 45664 22778 45692 24142
rect 45744 23656 45796 23662
rect 45744 23598 45796 23604
rect 45652 22772 45704 22778
rect 45652 22714 45704 22720
rect 45560 21888 45612 21894
rect 45560 21830 45612 21836
rect 45468 21684 45520 21690
rect 45468 21626 45520 21632
rect 45468 20936 45520 20942
rect 45468 20878 45520 20884
rect 45480 20602 45508 20878
rect 45468 20596 45520 20602
rect 45468 20538 45520 20544
rect 45572 19417 45600 21830
rect 45650 20632 45706 20641
rect 45650 20567 45652 20576
rect 45704 20567 45706 20576
rect 45652 20538 45704 20544
rect 45558 19408 45614 19417
rect 45558 19343 45614 19352
rect 45388 19306 45508 19334
rect 45376 18080 45428 18086
rect 45376 18022 45428 18028
rect 45388 16522 45416 18022
rect 45480 17513 45508 19306
rect 45652 19236 45704 19242
rect 45652 19178 45704 19184
rect 45466 17504 45522 17513
rect 45466 17439 45522 17448
rect 45664 17377 45692 19178
rect 45650 17368 45706 17377
rect 45650 17303 45706 17312
rect 45468 17196 45520 17202
rect 45468 17138 45520 17144
rect 45480 16590 45508 17138
rect 45560 16992 45612 16998
rect 45560 16934 45612 16940
rect 45468 16584 45520 16590
rect 45468 16526 45520 16532
rect 45376 16516 45428 16522
rect 45376 16458 45428 16464
rect 45468 16448 45520 16454
rect 45374 16416 45430 16425
rect 45430 16396 45468 16402
rect 45430 16390 45520 16396
rect 45430 16374 45508 16390
rect 45374 16351 45430 16360
rect 45480 16046 45508 16374
rect 45572 16182 45600 16934
rect 45560 16176 45612 16182
rect 45560 16118 45612 16124
rect 45468 16040 45520 16046
rect 45468 15982 45520 15988
rect 45468 15904 45520 15910
rect 45468 15846 45520 15852
rect 45480 15706 45508 15846
rect 45468 15700 45520 15706
rect 45468 15642 45520 15648
rect 45466 15600 45522 15609
rect 45466 15535 45468 15544
rect 45520 15535 45522 15544
rect 45468 15506 45520 15512
rect 45374 15192 45430 15201
rect 45664 15178 45692 17303
rect 45374 15127 45430 15136
rect 45480 15150 45692 15178
rect 45388 14414 45416 15127
rect 45480 14822 45508 15150
rect 45652 15020 45704 15026
rect 45652 14962 45704 14968
rect 45664 14822 45692 14962
rect 45468 14816 45520 14822
rect 45468 14758 45520 14764
rect 45652 14816 45704 14822
rect 45652 14758 45704 14764
rect 45376 14408 45428 14414
rect 45376 14350 45428 14356
rect 45560 14068 45612 14074
rect 45560 14010 45612 14016
rect 45284 13932 45336 13938
rect 45284 13874 45336 13880
rect 45282 13832 45338 13841
rect 45282 13767 45338 13776
rect 45192 12708 45244 12714
rect 45192 12650 45244 12656
rect 45296 12322 45324 13767
rect 45572 12918 45600 14010
rect 45560 12912 45612 12918
rect 45560 12854 45612 12860
rect 45376 12844 45428 12850
rect 45376 12786 45428 12792
rect 45388 12442 45416 12786
rect 45664 12764 45692 14758
rect 45756 14074 45784 23598
rect 45848 21010 45876 24262
rect 45940 22094 45968 25735
rect 46032 23497 46060 26200
rect 46662 25528 46718 25537
rect 46662 25463 46718 25472
rect 46570 25392 46626 25401
rect 46570 25327 46626 25336
rect 46204 24268 46256 24274
rect 46204 24210 46256 24216
rect 46018 23488 46074 23497
rect 46018 23423 46074 23432
rect 46110 22672 46166 22681
rect 46216 22642 46244 24210
rect 46296 24200 46348 24206
rect 46296 24142 46348 24148
rect 46308 23322 46336 24142
rect 46296 23316 46348 23322
rect 46296 23258 46348 23264
rect 46388 23316 46440 23322
rect 46388 23258 46440 23264
rect 46110 22607 46166 22616
rect 46204 22636 46256 22642
rect 46124 22574 46152 22607
rect 46204 22578 46256 22584
rect 46112 22568 46164 22574
rect 46112 22510 46164 22516
rect 46216 22098 46244 22578
rect 46294 22264 46350 22273
rect 46294 22199 46350 22208
rect 45940 22066 46152 22094
rect 46020 22024 46072 22030
rect 46020 21966 46072 21972
rect 45836 21004 45888 21010
rect 45836 20946 45888 20952
rect 45928 20868 45980 20874
rect 45928 20810 45980 20816
rect 45836 20460 45888 20466
rect 45836 20402 45888 20408
rect 45848 20058 45876 20402
rect 45836 20052 45888 20058
rect 45836 19994 45888 20000
rect 45940 19378 45968 20810
rect 46032 20641 46060 21966
rect 46018 20632 46074 20641
rect 46018 20567 46074 20576
rect 46124 20466 46152 22066
rect 46204 22092 46256 22098
rect 46204 22034 46256 22040
rect 46202 21448 46258 21457
rect 46202 21383 46258 21392
rect 46112 20460 46164 20466
rect 46112 20402 46164 20408
rect 46020 20392 46072 20398
rect 46020 20334 46072 20340
rect 46032 20233 46060 20334
rect 46112 20256 46164 20262
rect 46018 20224 46074 20233
rect 46112 20198 46164 20204
rect 46018 20159 46074 20168
rect 46124 19825 46152 20198
rect 46110 19816 46166 19825
rect 46110 19751 46166 19760
rect 45928 19372 45980 19378
rect 45928 19314 45980 19320
rect 46020 17808 46072 17814
rect 46020 17750 46072 17756
rect 46032 17678 46060 17750
rect 46020 17672 46072 17678
rect 46020 17614 46072 17620
rect 45836 17536 45888 17542
rect 45836 17478 45888 17484
rect 45928 17536 45980 17542
rect 45928 17478 45980 17484
rect 45848 17270 45876 17478
rect 45836 17264 45888 17270
rect 45836 17206 45888 17212
rect 45940 17202 45968 17478
rect 45928 17196 45980 17202
rect 45928 17138 45980 17144
rect 46018 16960 46074 16969
rect 46018 16895 46074 16904
rect 45836 16720 45888 16726
rect 45836 16662 45888 16668
rect 45848 15994 45876 16662
rect 45928 16448 45980 16454
rect 45928 16390 45980 16396
rect 45940 16114 45968 16390
rect 45928 16108 45980 16114
rect 45928 16050 45980 16056
rect 45848 15966 45968 15994
rect 45834 15464 45890 15473
rect 45834 15399 45890 15408
rect 45744 14068 45796 14074
rect 45744 14010 45796 14016
rect 45848 13818 45876 15399
rect 45940 15026 45968 15966
rect 45928 15020 45980 15026
rect 45928 14962 45980 14968
rect 45926 14920 45982 14929
rect 45926 14855 45982 14864
rect 45572 12736 45692 12764
rect 45756 13790 45876 13818
rect 45376 12436 45428 12442
rect 45376 12378 45428 12384
rect 45296 12294 45416 12322
rect 45284 12232 45336 12238
rect 45284 12174 45336 12180
rect 45192 11688 45244 11694
rect 45192 11630 45244 11636
rect 45204 11286 45232 11630
rect 45296 11354 45324 12174
rect 45388 11762 45416 12294
rect 45468 12096 45520 12102
rect 45468 12038 45520 12044
rect 45376 11756 45428 11762
rect 45376 11698 45428 11704
rect 45480 11626 45508 12038
rect 45468 11620 45520 11626
rect 45468 11562 45520 11568
rect 45284 11348 45336 11354
rect 45284 11290 45336 11296
rect 45192 11280 45244 11286
rect 45192 11222 45244 11228
rect 45204 10266 45232 11222
rect 45468 11144 45520 11150
rect 45468 11086 45520 11092
rect 45284 11076 45336 11082
rect 45284 11018 45336 11024
rect 45192 10260 45244 10266
rect 45192 10202 45244 10208
rect 45100 9580 45152 9586
rect 45100 9522 45152 9528
rect 45192 9512 45244 9518
rect 45190 9480 45192 9489
rect 45244 9480 45246 9489
rect 45190 9415 45246 9424
rect 45008 9172 45060 9178
rect 45008 9114 45060 9120
rect 45204 8090 45232 9415
rect 45192 8084 45244 8090
rect 45192 8026 45244 8032
rect 44916 8016 44968 8022
rect 44916 7958 44968 7964
rect 45296 7546 45324 11018
rect 45376 10532 45428 10538
rect 45376 10474 45428 10480
rect 45388 8566 45416 10474
rect 45376 8560 45428 8566
rect 45376 8502 45428 8508
rect 45376 7948 45428 7954
rect 45376 7890 45428 7896
rect 45284 7540 45336 7546
rect 45284 7482 45336 7488
rect 44824 7472 44876 7478
rect 45008 7472 45060 7478
rect 44824 7414 44876 7420
rect 45006 7440 45008 7449
rect 45060 7440 45062 7449
rect 44836 6866 44864 7414
rect 45006 7375 45062 7384
rect 45190 7304 45246 7313
rect 45190 7239 45246 7248
rect 44824 6860 44876 6866
rect 44824 6802 44876 6808
rect 45008 6656 45060 6662
rect 45008 6598 45060 6604
rect 45020 5817 45048 6598
rect 45100 6112 45152 6118
rect 45098 6080 45100 6089
rect 45152 6080 45154 6089
rect 45098 6015 45154 6024
rect 45204 5914 45232 7239
rect 45284 6792 45336 6798
rect 45284 6734 45336 6740
rect 45296 6118 45324 6734
rect 45284 6112 45336 6118
rect 45284 6054 45336 6060
rect 45388 5914 45416 7890
rect 45480 6798 45508 11086
rect 45572 10742 45600 12736
rect 45652 12368 45704 12374
rect 45652 12310 45704 12316
rect 45560 10736 45612 10742
rect 45560 10678 45612 10684
rect 45558 10160 45614 10169
rect 45558 10095 45614 10104
rect 45572 10062 45600 10095
rect 45560 10056 45612 10062
rect 45560 9998 45612 10004
rect 45468 6792 45520 6798
rect 45468 6734 45520 6740
rect 45468 6656 45520 6662
rect 45466 6624 45468 6633
rect 45520 6624 45522 6633
rect 45466 6559 45522 6568
rect 45468 6316 45520 6322
rect 45468 6258 45520 6264
rect 45480 6118 45508 6258
rect 45468 6112 45520 6118
rect 45468 6054 45520 6060
rect 45192 5908 45244 5914
rect 45192 5850 45244 5856
rect 45376 5908 45428 5914
rect 45376 5850 45428 5856
rect 45480 5846 45508 6054
rect 45572 5914 45600 9998
rect 45664 6458 45692 12310
rect 45756 9738 45784 13790
rect 45756 9710 45876 9738
rect 45744 9580 45796 9586
rect 45744 9522 45796 9528
rect 45652 6452 45704 6458
rect 45652 6394 45704 6400
rect 45560 5908 45612 5914
rect 45560 5850 45612 5856
rect 45756 5846 45784 9522
rect 45468 5840 45520 5846
rect 45006 5808 45062 5817
rect 45468 5782 45520 5788
rect 45744 5840 45796 5846
rect 45744 5782 45796 5788
rect 45006 5743 45062 5752
rect 45558 5672 45614 5681
rect 45558 5607 45614 5616
rect 45744 5636 45796 5642
rect 45572 5370 45600 5607
rect 45744 5578 45796 5584
rect 45560 5364 45612 5370
rect 45560 5306 45612 5312
rect 44730 4584 44786 4593
rect 44730 4519 44786 4528
rect 45560 4004 45612 4010
rect 45560 3946 45612 3952
rect 44272 2508 44324 2514
rect 44272 2450 44324 2456
rect 45572 800 45600 3946
rect 45756 3058 45784 5578
rect 45848 5370 45876 9710
rect 45940 9178 45968 14855
rect 45928 9172 45980 9178
rect 45928 9114 45980 9120
rect 45926 8256 45982 8265
rect 45926 8191 45982 8200
rect 45940 7410 45968 8191
rect 45928 7404 45980 7410
rect 45928 7346 45980 7352
rect 45926 6896 45982 6905
rect 46032 6866 46060 16895
rect 46124 11830 46152 19751
rect 46216 12434 46244 21383
rect 46308 19938 46336 22199
rect 46400 20913 46428 23258
rect 46478 22128 46534 22137
rect 46478 22063 46534 22072
rect 46492 22030 46520 22063
rect 46480 22024 46532 22030
rect 46480 21966 46532 21972
rect 46584 21690 46612 25327
rect 46676 24070 46704 25463
rect 46664 24064 46716 24070
rect 46662 24032 46664 24041
rect 46716 24032 46718 24041
rect 46662 23967 46718 23976
rect 46664 23180 46716 23186
rect 46664 23122 46716 23128
rect 46480 21684 46532 21690
rect 46480 21626 46532 21632
rect 46572 21684 46624 21690
rect 46572 21626 46624 21632
rect 46386 20904 46442 20913
rect 46386 20839 46442 20848
rect 46492 20330 46520 21626
rect 46676 21049 46704 23122
rect 46662 21040 46718 21049
rect 46662 20975 46718 20984
rect 46664 20936 46716 20942
rect 46664 20878 46716 20884
rect 46572 20868 46624 20874
rect 46572 20810 46624 20816
rect 46480 20324 46532 20330
rect 46480 20266 46532 20272
rect 46308 19910 46428 19938
rect 46296 19848 46348 19854
rect 46296 19790 46348 19796
rect 46308 18970 46336 19790
rect 46296 18964 46348 18970
rect 46296 18906 46348 18912
rect 46296 18760 46348 18766
rect 46296 18702 46348 18708
rect 46308 18222 46336 18702
rect 46296 18216 46348 18222
rect 46296 18158 46348 18164
rect 46294 17776 46350 17785
rect 46294 17711 46350 17720
rect 46308 16425 46336 17711
rect 46294 16416 46350 16425
rect 46294 16351 46350 16360
rect 46400 13938 46428 19910
rect 46480 18352 46532 18358
rect 46480 18294 46532 18300
rect 46492 17882 46520 18294
rect 46480 17876 46532 17882
rect 46480 17818 46532 17824
rect 46584 17785 46612 20810
rect 46676 18086 46704 20878
rect 46664 18080 46716 18086
rect 46664 18022 46716 18028
rect 46570 17776 46626 17785
rect 46570 17711 46626 17720
rect 46480 17060 46532 17066
rect 46480 17002 46532 17008
rect 46296 13932 46348 13938
rect 46296 13874 46348 13880
rect 46388 13932 46440 13938
rect 46388 13874 46440 13880
rect 46308 12753 46336 13874
rect 46294 12744 46350 12753
rect 46294 12679 46350 12688
rect 46216 12406 46336 12434
rect 46112 11824 46164 11830
rect 46112 11766 46164 11772
rect 46112 11144 46164 11150
rect 46110 11112 46112 11121
rect 46164 11112 46166 11121
rect 46110 11047 46166 11056
rect 46204 10736 46256 10742
rect 46110 10704 46166 10713
rect 46204 10678 46256 10684
rect 46110 10639 46112 10648
rect 46164 10639 46166 10648
rect 46112 10610 46164 10616
rect 46216 10577 46244 10678
rect 46202 10568 46258 10577
rect 46202 10503 46258 10512
rect 46216 10198 46244 10503
rect 46204 10192 46256 10198
rect 46204 10134 46256 10140
rect 46202 7440 46258 7449
rect 46308 7410 46336 12406
rect 46388 12232 46440 12238
rect 46388 12174 46440 12180
rect 46400 8362 46428 12174
rect 46492 9586 46520 17002
rect 46676 16946 46704 18022
rect 46768 17066 46796 26302
rect 47216 26240 47268 26246
rect 47306 26200 47362 27000
rect 47950 26330 48006 27000
rect 47872 26302 48006 26330
rect 47216 26182 47268 26188
rect 47124 26036 47176 26042
rect 47124 25978 47176 25984
rect 46938 24848 46994 24857
rect 46938 24783 46994 24792
rect 46848 24132 46900 24138
rect 46848 24074 46900 24080
rect 46860 23497 46888 24074
rect 46846 23488 46902 23497
rect 46846 23423 46902 23432
rect 46952 23254 46980 24783
rect 47030 24168 47086 24177
rect 47030 24103 47086 24112
rect 47044 23633 47072 24103
rect 47030 23624 47086 23633
rect 47030 23559 47086 23568
rect 47136 23254 47164 25978
rect 47228 24410 47256 26182
rect 47216 24404 47268 24410
rect 47216 24346 47268 24352
rect 47214 23896 47270 23905
rect 47214 23831 47270 23840
rect 47228 23730 47256 23831
rect 47216 23724 47268 23730
rect 47216 23666 47268 23672
rect 47214 23624 47270 23633
rect 47214 23559 47270 23568
rect 46940 23248 46992 23254
rect 46940 23190 46992 23196
rect 47124 23248 47176 23254
rect 47124 23190 47176 23196
rect 47136 23118 47164 23190
rect 46848 23112 46900 23118
rect 46848 23054 46900 23060
rect 47124 23112 47176 23118
rect 47124 23054 47176 23060
rect 46860 22778 46888 23054
rect 47032 23044 47084 23050
rect 47032 22986 47084 22992
rect 47044 22953 47072 22986
rect 47030 22944 47086 22953
rect 47030 22879 47086 22888
rect 46848 22772 46900 22778
rect 46848 22714 46900 22720
rect 46940 22704 46992 22710
rect 46940 22646 46992 22652
rect 46846 21040 46902 21049
rect 46846 20975 46902 20984
rect 46756 17060 46808 17066
rect 46756 17002 46808 17008
rect 46584 16918 46704 16946
rect 46584 16182 46612 16918
rect 46860 16776 46888 20975
rect 46952 20942 46980 22646
rect 47228 22094 47256 23559
rect 47320 23322 47348 26200
rect 47492 26172 47544 26178
rect 47492 26114 47544 26120
rect 47400 23520 47452 23526
rect 47400 23462 47452 23468
rect 47308 23316 47360 23322
rect 47308 23258 47360 23264
rect 47044 22066 47256 22094
rect 47044 21690 47072 22066
rect 47124 21956 47176 21962
rect 47124 21898 47176 21904
rect 47032 21684 47084 21690
rect 47032 21626 47084 21632
rect 46940 20936 46992 20942
rect 46940 20878 46992 20884
rect 46940 20800 46992 20806
rect 46938 20768 46940 20777
rect 46992 20768 46994 20777
rect 46938 20703 46994 20712
rect 47136 20346 47164 21898
rect 47308 21888 47360 21894
rect 47308 21830 47360 21836
rect 47136 20318 47256 20346
rect 47124 20256 47176 20262
rect 47124 20198 47176 20204
rect 47032 19712 47084 19718
rect 46938 19680 46994 19689
rect 47032 19654 47084 19660
rect 46938 19615 46994 19624
rect 46952 19378 46980 19615
rect 46940 19372 46992 19378
rect 46940 19314 46992 19320
rect 46940 19168 46992 19174
rect 46940 19110 46992 19116
rect 46952 18873 46980 19110
rect 46938 18864 46994 18873
rect 46938 18799 46994 18808
rect 46940 18352 46992 18358
rect 46940 18294 46992 18300
rect 46676 16748 46888 16776
rect 46572 16176 46624 16182
rect 46572 16118 46624 16124
rect 46572 15904 46624 15910
rect 46572 15846 46624 15852
rect 46584 15638 46612 15846
rect 46572 15632 46624 15638
rect 46572 15574 46624 15580
rect 46572 12844 46624 12850
rect 46572 12786 46624 12792
rect 46584 11354 46612 12786
rect 46572 11348 46624 11354
rect 46572 11290 46624 11296
rect 46480 9580 46532 9586
rect 46480 9522 46532 9528
rect 46676 9058 46704 16748
rect 46754 16552 46810 16561
rect 46754 16487 46810 16496
rect 46768 12918 46796 16487
rect 46952 16289 46980 18294
rect 47044 18290 47072 19654
rect 47136 18986 47164 20198
rect 47228 19174 47256 20318
rect 47216 19168 47268 19174
rect 47216 19110 47268 19116
rect 47136 18958 47256 18986
rect 47124 18896 47176 18902
rect 47124 18838 47176 18844
rect 47136 18290 47164 18838
rect 47032 18284 47084 18290
rect 47032 18226 47084 18232
rect 47124 18284 47176 18290
rect 47124 18226 47176 18232
rect 47124 18148 47176 18154
rect 47124 18090 47176 18096
rect 47136 18057 47164 18090
rect 47122 18048 47178 18057
rect 47122 17983 47178 17992
rect 47124 17536 47176 17542
rect 47124 17478 47176 17484
rect 47136 17270 47164 17478
rect 47124 17264 47176 17270
rect 47124 17206 47176 17212
rect 47124 17128 47176 17134
rect 47124 17070 47176 17076
rect 47032 16448 47084 16454
rect 47032 16390 47084 16396
rect 46938 16280 46994 16289
rect 46938 16215 46994 16224
rect 47044 16096 47072 16390
rect 46952 16068 47072 16096
rect 46848 15360 46900 15366
rect 46848 15302 46900 15308
rect 46756 12912 46808 12918
rect 46756 12854 46808 12860
rect 46754 12336 46810 12345
rect 46754 12271 46756 12280
rect 46808 12271 46810 12280
rect 46756 12242 46808 12248
rect 46860 12238 46888 15302
rect 46952 13462 46980 16068
rect 47030 16008 47086 16017
rect 47030 15943 47086 15952
rect 47044 15910 47072 15943
rect 47032 15904 47084 15910
rect 47032 15846 47084 15852
rect 47032 14952 47084 14958
rect 47032 14894 47084 14900
rect 47044 14074 47072 14894
rect 47032 14068 47084 14074
rect 47032 14010 47084 14016
rect 46940 13456 46992 13462
rect 46992 13404 47072 13410
rect 46940 13398 47072 13404
rect 46952 13382 47072 13398
rect 46940 13320 46992 13326
rect 46940 13262 46992 13268
rect 46952 12986 46980 13262
rect 47044 12986 47072 13382
rect 46940 12980 46992 12986
rect 46940 12922 46992 12928
rect 47032 12980 47084 12986
rect 47032 12922 47084 12928
rect 46848 12232 46900 12238
rect 46848 12174 46900 12180
rect 47136 12050 47164 17070
rect 47228 16833 47256 18958
rect 47214 16824 47270 16833
rect 47214 16759 47270 16768
rect 47216 16720 47268 16726
rect 47214 16688 47216 16697
rect 47268 16688 47270 16697
rect 47214 16623 47270 16632
rect 47216 16584 47268 16590
rect 47216 16526 47268 16532
rect 47228 12186 47256 16526
rect 47320 14414 47348 21830
rect 47412 21690 47440 23462
rect 47504 22094 47532 26114
rect 47768 24812 47820 24818
rect 47768 24754 47820 24760
rect 47780 23866 47808 24754
rect 47768 23860 47820 23866
rect 47768 23802 47820 23808
rect 47768 23656 47820 23662
rect 47768 23598 47820 23604
rect 47584 23588 47636 23594
rect 47636 23548 47716 23576
rect 47584 23530 47636 23536
rect 47504 22066 47624 22094
rect 47400 21684 47452 21690
rect 47400 21626 47452 21632
rect 47492 21548 47544 21554
rect 47492 21490 47544 21496
rect 47400 21344 47452 21350
rect 47400 21286 47452 21292
rect 47412 20942 47440 21286
rect 47400 20936 47452 20942
rect 47400 20878 47452 20884
rect 47398 20632 47454 20641
rect 47398 20567 47454 20576
rect 47412 18970 47440 20567
rect 47400 18964 47452 18970
rect 47400 18906 47452 18912
rect 47398 18728 47454 18737
rect 47398 18663 47454 18672
rect 47412 16454 47440 18663
rect 47400 16448 47452 16454
rect 47400 16390 47452 16396
rect 47400 16176 47452 16182
rect 47400 16118 47452 16124
rect 47308 14408 47360 14414
rect 47308 14350 47360 14356
rect 47412 14226 47440 16118
rect 47504 14618 47532 21490
rect 47596 18222 47624 22066
rect 47688 21962 47716 23548
rect 47780 22778 47808 23598
rect 47872 23322 47900 26302
rect 47950 26200 48006 26302
rect 48594 26200 48650 27000
rect 49238 26330 49294 27000
rect 49238 26302 49556 26330
rect 49238 26200 49294 26302
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 47860 23316 47912 23322
rect 47860 23258 47912 23264
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 47768 22772 47820 22778
rect 47768 22714 47820 22720
rect 47768 22636 47820 22642
rect 47768 22578 47820 22584
rect 47676 21956 47728 21962
rect 47676 21898 47728 21904
rect 47676 21684 47728 21690
rect 47676 21626 47728 21632
rect 47584 18216 47636 18222
rect 47584 18158 47636 18164
rect 47584 17604 47636 17610
rect 47584 17546 47636 17552
rect 47492 14612 47544 14618
rect 47492 14554 47544 14560
rect 47412 14198 47532 14226
rect 47400 14068 47452 14074
rect 47400 14010 47452 14016
rect 47306 13968 47362 13977
rect 47306 13903 47362 13912
rect 47320 12374 47348 13903
rect 47412 13308 47440 14010
rect 47504 13734 47532 14198
rect 47492 13728 47544 13734
rect 47492 13670 47544 13676
rect 47492 13456 47544 13462
rect 47490 13424 47492 13433
rect 47544 13424 47546 13433
rect 47490 13359 47546 13368
rect 47412 13280 47532 13308
rect 47308 12368 47360 12374
rect 47308 12310 47360 12316
rect 47228 12158 47348 12186
rect 47136 12022 47256 12050
rect 47122 11928 47178 11937
rect 47122 11863 47124 11872
rect 47176 11863 47178 11872
rect 47124 11834 47176 11840
rect 46848 11756 46900 11762
rect 46848 11698 46900 11704
rect 46940 11756 46992 11762
rect 46940 11698 46992 11704
rect 47032 11756 47084 11762
rect 47032 11698 47084 11704
rect 46860 11218 46888 11698
rect 46848 11212 46900 11218
rect 46848 11154 46900 11160
rect 46848 10124 46900 10130
rect 46848 10066 46900 10072
rect 46860 9625 46888 10066
rect 46846 9616 46902 9625
rect 46846 9551 46902 9560
rect 46676 9030 46796 9058
rect 46768 8974 46796 9030
rect 46756 8968 46808 8974
rect 46756 8910 46808 8916
rect 46388 8356 46440 8362
rect 46388 8298 46440 8304
rect 46386 7848 46442 7857
rect 46386 7783 46442 7792
rect 46400 7750 46428 7783
rect 46388 7744 46440 7750
rect 46388 7686 46440 7692
rect 46202 7375 46204 7384
rect 46256 7375 46258 7384
rect 46296 7404 46348 7410
rect 46204 7346 46256 7352
rect 46296 7346 46348 7352
rect 45926 6831 45982 6840
rect 46020 6860 46072 6866
rect 45940 6798 45968 6831
rect 46020 6802 46072 6808
rect 45928 6792 45980 6798
rect 45928 6734 45980 6740
rect 45940 6089 45968 6734
rect 46032 6662 46060 6802
rect 46020 6656 46072 6662
rect 46020 6598 46072 6604
rect 46018 6488 46074 6497
rect 46018 6423 46020 6432
rect 46072 6423 46074 6432
rect 46020 6394 46072 6400
rect 45926 6080 45982 6089
rect 45926 6015 45982 6024
rect 45928 5772 45980 5778
rect 45928 5714 45980 5720
rect 45836 5364 45888 5370
rect 45836 5306 45888 5312
rect 45848 4826 45876 5306
rect 45836 4820 45888 4826
rect 45836 4762 45888 4768
rect 45940 3058 45968 5714
rect 46216 4826 46244 7346
rect 46296 6860 46348 6866
rect 46296 6802 46348 6808
rect 46308 6322 46336 6802
rect 46296 6316 46348 6322
rect 46296 6258 46348 6264
rect 46204 4820 46256 4826
rect 46204 4762 46256 4768
rect 46308 4622 46336 6258
rect 46662 6216 46718 6225
rect 46388 6180 46440 6186
rect 46662 6151 46664 6160
rect 46388 6122 46440 6128
rect 46716 6151 46718 6160
rect 46664 6122 46716 6128
rect 46400 5642 46428 6122
rect 46572 5840 46624 5846
rect 46572 5782 46624 5788
rect 46584 5710 46612 5782
rect 46572 5704 46624 5710
rect 46572 5646 46624 5652
rect 46388 5636 46440 5642
rect 46388 5578 46440 5584
rect 46584 4758 46612 5646
rect 46768 4826 46796 8910
rect 46848 8424 46900 8430
rect 46848 8366 46900 8372
rect 46860 7993 46888 8366
rect 46846 7984 46902 7993
rect 46952 7970 46980 11698
rect 47044 8090 47072 11698
rect 47124 11552 47176 11558
rect 47124 11494 47176 11500
rect 47136 9500 47164 11494
rect 47228 9654 47256 12022
rect 47216 9648 47268 9654
rect 47216 9590 47268 9596
rect 47136 9472 47256 9500
rect 47124 9376 47176 9382
rect 47124 9318 47176 9324
rect 47032 8084 47084 8090
rect 47032 8026 47084 8032
rect 46952 7942 47072 7970
rect 46846 7919 46902 7928
rect 46940 7744 46992 7750
rect 46940 7686 46992 7692
rect 46848 6656 46900 6662
rect 46848 6598 46900 6604
rect 46860 6322 46888 6598
rect 46848 6316 46900 6322
rect 46848 6258 46900 6264
rect 46952 6254 46980 7686
rect 46940 6248 46992 6254
rect 46940 6190 46992 6196
rect 47044 5914 47072 7942
rect 47136 7886 47164 9318
rect 47124 7880 47176 7886
rect 47124 7822 47176 7828
rect 47228 7342 47256 9472
rect 47216 7336 47268 7342
rect 47216 7278 47268 7284
rect 47214 6760 47270 6769
rect 47124 6724 47176 6730
rect 47214 6695 47270 6704
rect 47124 6666 47176 6672
rect 47032 5908 47084 5914
rect 47032 5850 47084 5856
rect 46940 5704 46992 5710
rect 46940 5646 46992 5652
rect 46952 5370 46980 5646
rect 46940 5364 46992 5370
rect 46940 5306 46992 5312
rect 46756 4820 46808 4826
rect 46756 4762 46808 4768
rect 46572 4752 46624 4758
rect 46572 4694 46624 4700
rect 46296 4616 46348 4622
rect 46296 4558 46348 4564
rect 46664 4072 46716 4078
rect 46664 4014 46716 4020
rect 45744 3052 45796 3058
rect 45744 2994 45796 3000
rect 45928 3052 45980 3058
rect 45928 2994 45980 3000
rect 46676 1465 46704 4014
rect 47136 3534 47164 6666
rect 47228 6458 47256 6695
rect 47216 6452 47268 6458
rect 47216 6394 47268 6400
rect 47214 6352 47270 6361
rect 47214 6287 47270 6296
rect 47228 5914 47256 6287
rect 47216 5908 47268 5914
rect 47216 5850 47268 5856
rect 47320 4826 47348 12158
rect 47398 11384 47454 11393
rect 47398 11319 47400 11328
rect 47452 11319 47454 11328
rect 47400 11290 47452 11296
rect 47400 11144 47452 11150
rect 47400 11086 47452 11092
rect 47412 4826 47440 11086
rect 47504 9450 47532 13280
rect 47596 12889 47624 17546
rect 47688 16153 47716 21626
rect 47780 21418 47808 22578
rect 48412 22432 48464 22438
rect 48412 22374 48464 22380
rect 48320 22024 48372 22030
rect 48320 21966 48372 21972
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 47952 21480 48004 21486
rect 47952 21422 48004 21428
rect 47768 21412 47820 21418
rect 47768 21354 47820 21360
rect 47860 21140 47912 21146
rect 47860 21082 47912 21088
rect 47768 20528 47820 20534
rect 47768 20470 47820 20476
rect 47780 18057 47808 20470
rect 47872 19334 47900 21082
rect 47964 20874 47992 21422
rect 47952 20868 48004 20874
rect 47952 20810 48004 20816
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 48226 20496 48282 20505
rect 48226 20431 48282 20440
rect 48240 19836 48268 20431
rect 48332 19990 48360 21966
rect 48424 20777 48452 22374
rect 48504 22160 48556 22166
rect 48504 22102 48556 22108
rect 48516 20942 48544 22102
rect 48504 20936 48556 20942
rect 48504 20878 48556 20884
rect 48504 20800 48556 20806
rect 48410 20768 48466 20777
rect 48504 20742 48556 20748
rect 48410 20703 48466 20712
rect 48320 19984 48372 19990
rect 48320 19926 48372 19932
rect 48516 19854 48544 20742
rect 48412 19848 48464 19854
rect 48240 19808 48360 19836
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 47872 19306 47992 19334
rect 47860 19236 47912 19242
rect 47860 19178 47912 19184
rect 47872 18358 47900 19178
rect 47964 18737 47992 19306
rect 48228 19168 48280 19174
rect 48226 19136 48228 19145
rect 48280 19136 48282 19145
rect 48226 19071 48282 19080
rect 47950 18728 48006 18737
rect 47950 18663 48006 18672
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 47860 18352 47912 18358
rect 47860 18294 47912 18300
rect 47858 18184 47914 18193
rect 47858 18119 47914 18128
rect 47766 18048 47822 18057
rect 47766 17983 47822 17992
rect 47766 17912 47822 17921
rect 47766 17847 47822 17856
rect 47780 17066 47808 17847
rect 47768 17060 47820 17066
rect 47768 17002 47820 17008
rect 47674 16144 47730 16153
rect 47674 16079 47730 16088
rect 47768 15360 47820 15366
rect 47674 15328 47730 15337
rect 47768 15302 47820 15308
rect 47674 15263 47730 15272
rect 47688 15162 47716 15263
rect 47676 15156 47728 15162
rect 47676 15098 47728 15104
rect 47676 15020 47728 15026
rect 47676 14962 47728 14968
rect 47582 12880 47638 12889
rect 47688 12850 47716 14962
rect 47780 14414 47808 15302
rect 47872 15026 47900 18119
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 48332 16182 48360 19808
rect 48412 19790 48464 19796
rect 48504 19848 48556 19854
rect 48504 19790 48556 19796
rect 48424 18970 48452 19790
rect 48412 18964 48464 18970
rect 48412 18906 48464 18912
rect 48412 17672 48464 17678
rect 48412 17614 48464 17620
rect 48504 17672 48556 17678
rect 48504 17614 48556 17620
rect 48424 17338 48452 17614
rect 48412 17332 48464 17338
rect 48412 17274 48464 17280
rect 48412 16652 48464 16658
rect 48412 16594 48464 16600
rect 48320 16176 48372 16182
rect 48320 16118 48372 16124
rect 48320 15428 48372 15434
rect 48320 15370 48372 15376
rect 47950 15260 48258 15269
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 47860 15020 47912 15026
rect 47860 14962 47912 14968
rect 47768 14408 47820 14414
rect 47768 14350 47820 14356
rect 47766 14240 47822 14249
rect 47766 14175 47822 14184
rect 47780 14074 47808 14175
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 48332 14074 48360 15370
rect 47768 14068 47820 14074
rect 47768 14010 47820 14016
rect 48320 14068 48372 14074
rect 48320 14010 48372 14016
rect 47860 13932 47912 13938
rect 47860 13874 47912 13880
rect 47768 13728 47820 13734
rect 47768 13670 47820 13676
rect 47582 12815 47638 12824
rect 47676 12844 47728 12850
rect 47676 12786 47728 12792
rect 47780 12730 47808 13670
rect 47596 12702 47808 12730
rect 47492 9444 47544 9450
rect 47492 9386 47544 9392
rect 47596 9178 47624 12702
rect 47676 12640 47728 12646
rect 47676 12582 47728 12588
rect 47688 10810 47716 12582
rect 47676 10804 47728 10810
rect 47676 10746 47728 10752
rect 47676 10192 47728 10198
rect 47676 10134 47728 10140
rect 47584 9172 47636 9178
rect 47584 9114 47636 9120
rect 47688 6322 47716 10134
rect 47872 9654 47900 13874
rect 48318 13560 48374 13569
rect 48424 13530 48452 16594
rect 48516 16454 48544 17614
rect 48504 16448 48556 16454
rect 48504 16390 48556 16396
rect 48608 16266 48636 26200
rect 49240 25764 49292 25770
rect 49240 25706 49292 25712
rect 48962 25664 49018 25673
rect 48780 25628 48832 25634
rect 48962 25599 49018 25608
rect 48780 25570 48832 25576
rect 48792 24274 48820 25570
rect 48780 24268 48832 24274
rect 48780 24210 48832 24216
rect 48780 23316 48832 23322
rect 48780 23258 48832 23264
rect 48688 22704 48740 22710
rect 48688 22646 48740 22652
rect 48700 22030 48728 22646
rect 48688 22024 48740 22030
rect 48688 21966 48740 21972
rect 48688 21888 48740 21894
rect 48688 21830 48740 21836
rect 48516 16238 48636 16266
rect 48318 13495 48374 13504
rect 48412 13524 48464 13530
rect 48332 13394 48360 13495
rect 48412 13466 48464 13472
rect 48320 13388 48372 13394
rect 48320 13330 48372 13336
rect 48412 13388 48464 13394
rect 48412 13330 48464 13336
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 47950 11996 48258 12005
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 48424 10266 48452 13330
rect 48516 11286 48544 16238
rect 48596 15360 48648 15366
rect 48596 15302 48648 15308
rect 48608 15026 48636 15302
rect 48700 15094 48728 21830
rect 48792 17202 48820 23258
rect 48872 23112 48924 23118
rect 48872 23054 48924 23060
rect 48884 18306 48912 23054
rect 48976 18970 49004 25599
rect 49056 25356 49108 25362
rect 49056 25298 49108 25304
rect 49068 21690 49096 25298
rect 49148 23724 49200 23730
rect 49148 23666 49200 23672
rect 49160 22710 49188 23666
rect 49148 22704 49200 22710
rect 49148 22646 49200 22652
rect 49148 21888 49200 21894
rect 49148 21830 49200 21836
rect 49056 21684 49108 21690
rect 49056 21626 49108 21632
rect 49160 21622 49188 21830
rect 49148 21616 49200 21622
rect 49054 21584 49110 21593
rect 49148 21558 49200 21564
rect 49054 21519 49110 21528
rect 49068 20058 49096 21519
rect 49148 20392 49200 20398
rect 49148 20334 49200 20340
rect 49056 20052 49108 20058
rect 49056 19994 49108 20000
rect 49160 19938 49188 20334
rect 49068 19910 49188 19938
rect 48964 18964 49016 18970
rect 48964 18906 49016 18912
rect 48884 18278 49004 18306
rect 48872 18216 48924 18222
rect 48872 18158 48924 18164
rect 48780 17196 48832 17202
rect 48780 17138 48832 17144
rect 48780 16584 48832 16590
rect 48780 16526 48832 16532
rect 48792 16250 48820 16526
rect 48780 16244 48832 16250
rect 48780 16186 48832 16192
rect 48780 15904 48832 15910
rect 48780 15846 48832 15852
rect 48688 15088 48740 15094
rect 48688 15030 48740 15036
rect 48596 15020 48648 15026
rect 48596 14962 48648 14968
rect 48792 14906 48820 15846
rect 48700 14878 48820 14906
rect 48596 13932 48648 13938
rect 48596 13874 48648 13880
rect 48504 11280 48556 11286
rect 48504 11222 48556 11228
rect 48608 10742 48636 13874
rect 48700 13394 48728 14878
rect 48778 13424 48834 13433
rect 48688 13388 48740 13394
rect 48778 13359 48834 13368
rect 48688 13330 48740 13336
rect 48596 10736 48648 10742
rect 48596 10678 48648 10684
rect 48412 10260 48464 10266
rect 48412 10202 48464 10208
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 47860 9648 47912 9654
rect 47860 9590 47912 9596
rect 48318 9072 48374 9081
rect 48318 9007 48374 9016
rect 47860 8900 47912 8906
rect 47860 8842 47912 8848
rect 47768 8560 47820 8566
rect 47768 8502 47820 8508
rect 47780 6798 47808 8502
rect 47872 8498 47900 8842
rect 48332 8838 48360 9007
rect 48320 8832 48372 8838
rect 48320 8774 48372 8780
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 47860 8492 47912 8498
rect 47860 8434 47912 8440
rect 48320 7812 48372 7818
rect 48320 7754 48372 7760
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 47952 7404 48004 7410
rect 47952 7346 48004 7352
rect 47860 7268 47912 7274
rect 47860 7210 47912 7216
rect 47768 6792 47820 6798
rect 47768 6734 47820 6740
rect 47676 6316 47728 6322
rect 47676 6258 47728 6264
rect 47872 5234 47900 7210
rect 47964 7002 47992 7346
rect 47952 6996 48004 7002
rect 47952 6938 48004 6944
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 48332 5574 48360 7754
rect 48688 6724 48740 6730
rect 48688 6666 48740 6672
rect 48700 6361 48728 6666
rect 48686 6352 48742 6361
rect 48686 6287 48742 6296
rect 48320 5568 48372 5574
rect 48320 5510 48372 5516
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 47860 5228 47912 5234
rect 47860 5170 47912 5176
rect 48320 5160 48372 5166
rect 48320 5102 48372 5108
rect 47308 4820 47360 4826
rect 47308 4762 47360 4768
rect 47400 4820 47452 4826
rect 47400 4762 47452 4768
rect 48332 4729 48360 5102
rect 48318 4720 48374 4729
rect 48318 4655 48374 4664
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 47676 3596 47728 3602
rect 47676 3538 47728 3544
rect 47124 3528 47176 3534
rect 47124 3470 47176 3476
rect 46756 2984 46808 2990
rect 46756 2926 46808 2932
rect 46848 2984 46900 2990
rect 46848 2926 46900 2932
rect 46768 1873 46796 2926
rect 46860 2689 46888 2926
rect 46846 2680 46902 2689
rect 46846 2615 46902 2624
rect 46754 1864 46810 1873
rect 46754 1799 46810 1808
rect 46662 1456 46718 1465
rect 46662 1391 46718 1400
rect 47688 800 47716 3538
rect 48688 3460 48740 3466
rect 48688 3402 48740 3408
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 48700 3097 48728 3402
rect 48686 3088 48742 3097
rect 48686 3023 48742 3032
rect 48792 2774 48820 13359
rect 48884 10606 48912 18158
rect 48976 16658 49004 18278
rect 49068 17338 49096 19910
rect 49146 19408 49202 19417
rect 49146 19343 49148 19352
rect 49200 19343 49202 19352
rect 49148 19314 49200 19320
rect 49146 19000 49202 19009
rect 49146 18935 49202 18944
rect 49056 17332 49108 17338
rect 49056 17274 49108 17280
rect 49160 17270 49188 18935
rect 49252 18426 49280 25706
rect 49424 22976 49476 22982
rect 49424 22918 49476 22924
rect 49436 20534 49464 22918
rect 49424 20528 49476 20534
rect 49424 20470 49476 20476
rect 49528 20346 49556 26302
rect 49974 24712 50030 24721
rect 49974 24647 50030 24656
rect 49882 24304 49938 24313
rect 49882 24239 49938 24248
rect 49700 22024 49752 22030
rect 49700 21966 49752 21972
rect 49608 20460 49660 20466
rect 49608 20402 49660 20408
rect 49344 20318 49556 20346
rect 49240 18420 49292 18426
rect 49240 18362 49292 18368
rect 49238 18320 49294 18329
rect 49238 18255 49294 18264
rect 49148 17264 49200 17270
rect 49148 17206 49200 17212
rect 49056 17196 49108 17202
rect 49056 17138 49108 17144
rect 48964 16652 49016 16658
rect 48964 16594 49016 16600
rect 48964 16448 49016 16454
rect 48964 16390 49016 16396
rect 48872 10600 48924 10606
rect 48872 10542 48924 10548
rect 48976 4554 49004 16390
rect 49068 7954 49096 17138
rect 49252 16522 49280 18255
rect 49240 16516 49292 16522
rect 49240 16458 49292 16464
rect 49344 16232 49372 20318
rect 49516 20256 49568 20262
rect 49516 20198 49568 20204
rect 49422 19816 49478 19825
rect 49422 19751 49478 19760
rect 49160 16204 49372 16232
rect 49160 13938 49188 16204
rect 49240 16108 49292 16114
rect 49240 16050 49292 16056
rect 49252 15162 49280 16050
rect 49332 15496 49384 15502
rect 49332 15438 49384 15444
rect 49240 15156 49292 15162
rect 49240 15098 49292 15104
rect 49344 14618 49372 15438
rect 49332 14612 49384 14618
rect 49332 14554 49384 14560
rect 49148 13932 49200 13938
rect 49148 13874 49200 13880
rect 49148 13320 49200 13326
rect 49146 13288 49148 13297
rect 49200 13288 49202 13297
rect 49146 13223 49202 13232
rect 49146 12880 49202 12889
rect 49146 12815 49148 12824
rect 49200 12815 49202 12824
rect 49148 12786 49200 12792
rect 49146 12472 49202 12481
rect 49146 12407 49202 12416
rect 49160 12306 49188 12407
rect 49148 12300 49200 12306
rect 49148 12242 49200 12248
rect 49146 12064 49202 12073
rect 49146 11999 49202 12008
rect 49160 11830 49188 11999
rect 49148 11824 49200 11830
rect 49148 11766 49200 11772
rect 49146 11656 49202 11665
rect 49146 11591 49202 11600
rect 49160 11218 49188 11591
rect 49330 11248 49386 11257
rect 49148 11212 49200 11218
rect 49330 11183 49386 11192
rect 49148 11154 49200 11160
rect 49146 10840 49202 10849
rect 49146 10775 49202 10784
rect 49160 10130 49188 10775
rect 49344 10742 49372 11183
rect 49436 11082 49464 19751
rect 49424 11076 49476 11082
rect 49424 11018 49476 11024
rect 49332 10736 49384 10742
rect 49332 10678 49384 10684
rect 49422 10432 49478 10441
rect 49422 10367 49478 10376
rect 49148 10124 49200 10130
rect 49148 10066 49200 10072
rect 49238 10024 49294 10033
rect 49238 9959 49294 9968
rect 49146 9208 49202 9217
rect 49146 9143 49202 9152
rect 49160 8566 49188 9143
rect 49252 9042 49280 9959
rect 49436 9654 49464 10367
rect 49424 9648 49476 9654
rect 49424 9590 49476 9596
rect 49240 9036 49292 9042
rect 49240 8978 49292 8984
rect 49238 8800 49294 8809
rect 49238 8735 49294 8744
rect 49148 8560 49200 8566
rect 49148 8502 49200 8508
rect 49252 7954 49280 8735
rect 49330 8392 49386 8401
rect 49330 8327 49386 8336
rect 49056 7948 49108 7954
rect 49056 7890 49108 7896
rect 49240 7948 49292 7954
rect 49240 7890 49292 7896
rect 49146 7576 49202 7585
rect 49146 7511 49202 7520
rect 49160 6866 49188 7511
rect 49344 7478 49372 8327
rect 49332 7472 49384 7478
rect 49332 7414 49384 7420
rect 49238 7168 49294 7177
rect 49238 7103 49294 7112
rect 49148 6860 49200 6866
rect 49148 6802 49200 6808
rect 49252 6390 49280 7103
rect 49330 6760 49386 6769
rect 49330 6695 49386 6704
rect 49240 6384 49292 6390
rect 49240 6326 49292 6332
rect 49146 5944 49202 5953
rect 49146 5879 49202 5888
rect 49160 5302 49188 5879
rect 49344 5778 49372 6695
rect 49528 6633 49556 20198
rect 49620 15745 49648 20402
rect 49712 19786 49740 21966
rect 49790 21176 49846 21185
rect 49790 21111 49846 21120
rect 49700 19780 49752 19786
rect 49700 19722 49752 19728
rect 49804 18737 49832 21111
rect 49790 18728 49846 18737
rect 49700 18692 49752 18698
rect 49790 18663 49846 18672
rect 49700 18634 49752 18640
rect 49606 15736 49662 15745
rect 49606 15671 49662 15680
rect 49620 15366 49648 15671
rect 49608 15360 49660 15366
rect 49608 15302 49660 15308
rect 49712 14521 49740 18634
rect 49790 18592 49846 18601
rect 49790 18527 49846 18536
rect 49804 15450 49832 18527
rect 49896 17252 49924 24239
rect 49988 23338 50016 24647
rect 50066 23896 50122 23905
rect 50122 23854 50384 23882
rect 50066 23831 50122 23840
rect 49988 23310 50200 23338
rect 49974 23080 50030 23089
rect 49974 23015 50030 23024
rect 49988 17406 50016 23015
rect 50066 21856 50122 21865
rect 50066 21791 50122 21800
rect 50080 20738 50108 21791
rect 50068 20732 50120 20738
rect 50068 20674 50120 20680
rect 50066 20632 50122 20641
rect 50066 20567 50122 20576
rect 50080 19378 50108 20567
rect 50068 19372 50120 19378
rect 50068 19314 50120 19320
rect 50068 18284 50120 18290
rect 50068 18226 50120 18232
rect 49976 17400 50028 17406
rect 49976 17342 50028 17348
rect 49896 17224 50016 17252
rect 49884 17128 49936 17134
rect 49884 17070 49936 17076
rect 49896 15570 49924 17070
rect 49884 15564 49936 15570
rect 49884 15506 49936 15512
rect 49804 15422 49924 15450
rect 49792 15360 49844 15366
rect 49792 15302 49844 15308
rect 49698 14512 49754 14521
rect 49698 14447 49754 14456
rect 49514 6624 49570 6633
rect 49514 6559 49570 6568
rect 49332 5772 49384 5778
rect 49332 5714 49384 5720
rect 49422 5536 49478 5545
rect 49422 5471 49478 5480
rect 49148 5296 49200 5302
rect 49148 5238 49200 5244
rect 49238 5128 49294 5137
rect 49238 5063 49294 5072
rect 48964 4548 49016 4554
rect 48964 4490 49016 4496
rect 49146 4312 49202 4321
rect 49146 4247 49202 4256
rect 49160 3602 49188 4247
rect 49252 4146 49280 5063
rect 49436 4690 49464 5471
rect 49712 5370 49740 14447
rect 49700 5364 49752 5370
rect 49700 5306 49752 5312
rect 49424 4684 49476 4690
rect 49424 4626 49476 4632
rect 49240 4140 49292 4146
rect 49240 4082 49292 4088
rect 49804 4078 49832 15302
rect 49896 6905 49924 15422
rect 49988 7818 50016 17224
rect 50080 14929 50108 18226
rect 50066 14920 50122 14929
rect 50066 14855 50122 14864
rect 50066 14784 50122 14793
rect 50066 14719 50122 14728
rect 49976 7812 50028 7818
rect 49976 7754 50028 7760
rect 50080 7546 50108 14719
rect 50068 7540 50120 7546
rect 50068 7482 50120 7488
rect 50068 7336 50120 7342
rect 50066 7304 50068 7313
rect 50120 7304 50122 7313
rect 50066 7239 50122 7248
rect 49882 6896 49938 6905
rect 49882 6831 49938 6840
rect 50172 5914 50200 23310
rect 50252 20732 50304 20738
rect 50252 20674 50304 20680
rect 50264 6118 50292 20674
rect 50356 6798 50384 23854
rect 50528 22636 50580 22642
rect 50528 22578 50580 22584
rect 50436 20936 50488 20942
rect 50436 20878 50488 20884
rect 50448 15434 50476 20878
rect 50436 15428 50488 15434
rect 50436 15370 50488 15376
rect 50344 6792 50396 6798
rect 50344 6734 50396 6740
rect 50252 6112 50304 6118
rect 50252 6054 50304 6060
rect 50160 5908 50212 5914
rect 50160 5850 50212 5856
rect 50448 5846 50476 15370
rect 50540 7342 50568 22578
rect 50620 19712 50672 19718
rect 50620 19654 50672 19660
rect 50632 14006 50660 19654
rect 50804 19372 50856 19378
rect 50804 19314 50856 19320
rect 50712 17400 50764 17406
rect 50712 17342 50764 17348
rect 50620 14000 50672 14006
rect 50620 13942 50672 13948
rect 50724 12170 50752 17342
rect 50712 12164 50764 12170
rect 50712 12106 50764 12112
rect 50816 11694 50844 19314
rect 50896 14680 50948 14686
rect 50896 14622 50948 14628
rect 50804 11688 50856 11694
rect 50804 11630 50856 11636
rect 50528 7336 50580 7342
rect 50528 7278 50580 7284
rect 50908 6458 50936 14622
rect 50896 6452 50948 6458
rect 50896 6394 50948 6400
rect 50436 5840 50488 5846
rect 50436 5782 50488 5788
rect 49792 4072 49844 4078
rect 49792 4014 49844 4020
rect 49238 3904 49294 3913
rect 49238 3839 49294 3848
rect 49148 3596 49200 3602
rect 49148 3538 49200 3544
rect 49146 3496 49202 3505
rect 49146 3431 49202 3440
rect 48792 2746 48912 2774
rect 48884 2650 48912 2746
rect 48872 2644 48924 2650
rect 48872 2586 48924 2592
rect 49160 2514 49188 3431
rect 49252 3126 49280 3839
rect 49792 3664 49844 3670
rect 49792 3606 49844 3612
rect 49240 3120 49292 3126
rect 49240 3062 49292 3068
rect 49148 2508 49200 2514
rect 49148 2450 49200 2456
rect 48504 2372 48556 2378
rect 48504 2314 48556 2320
rect 48516 2281 48544 2314
rect 48502 2272 48558 2281
rect 47950 2204 48258 2213
rect 48502 2207 48558 2216
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 49804 800 49832 3606
rect 18156 734 18368 762
rect 20166 0 20222 800
rect 22282 0 22338 800
rect 24398 0 24454 800
rect 26514 0 26570 800
rect 28630 0 28686 800
rect 30746 0 30802 800
rect 32862 0 32918 800
rect 34978 0 35034 800
rect 37094 0 37150 800
rect 39210 0 39266 800
rect 41326 0 41382 800
rect 43442 0 43498 800
rect 45558 0 45614 800
rect 47674 0 47730 800
rect 49790 0 49846 800
<< via2 >>
rect 1766 21800 1822 21856
rect 1306 20712 1362 20768
rect 1214 17040 1270 17096
rect 1306 16632 1362 16688
rect 1306 16224 1362 16280
rect 1306 15816 1362 15872
rect 1306 15408 1362 15464
rect 1766 15272 1822 15328
rect 1306 15000 1362 15056
rect 1306 14592 1362 14648
rect 938 14184 994 14240
rect 1766 13232 1822 13288
rect 1306 12960 1362 13016
rect 1306 12144 1362 12200
rect 2042 18264 2098 18320
rect 2042 17448 2098 17504
rect 1306 10920 1362 10976
rect 2778 24384 2834 24440
rect 1214 10512 1270 10568
rect 1766 10532 1822 10568
rect 1766 10512 1768 10532
rect 1768 10512 1820 10532
rect 1820 10512 1822 10532
rect 1306 10104 1362 10160
rect 1582 9696 1638 9752
rect 1766 9444 1822 9480
rect 1766 9424 1768 9444
rect 1768 9424 1820 9444
rect 1820 9424 1822 9444
rect 1214 9288 1270 9344
rect 1306 8916 1308 8936
rect 1308 8916 1360 8936
rect 1360 8916 1362 8936
rect 1306 8880 1362 8916
rect 1766 8880 1822 8936
rect 1214 8508 1216 8528
rect 1216 8508 1268 8528
rect 1268 8508 1270 8528
rect 1214 8472 1270 8508
rect 1582 8064 1638 8120
rect 3422 25608 3478 25664
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 4066 25220 4122 25256
rect 4066 25200 4068 25220
rect 4068 25200 4120 25220
rect 4120 25200 4122 25220
rect 3698 24812 3754 24848
rect 3698 24792 3700 24812
rect 3700 24792 3752 24812
rect 3752 24792 3754 24812
rect 3330 23976 3386 24032
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 3238 23160 3294 23216
rect 2686 21528 2742 21584
rect 2778 21120 2834 21176
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 3238 21936 3294 21992
rect 3422 23196 3424 23216
rect 3424 23196 3476 23216
rect 3476 23196 3478 23216
rect 3422 23160 3478 23196
rect 3422 21836 3424 21856
rect 3424 21836 3476 21856
rect 3476 21836 3478 21856
rect 3422 21800 3478 21836
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2778 19080 2834 19136
rect 3330 19896 3386 19952
rect 2962 19488 3018 19544
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2870 18672 2926 18728
rect 2778 17856 2834 17912
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 3698 23588 3754 23624
rect 3698 23568 3700 23588
rect 3700 23568 3752 23588
rect 3752 23568 3754 23588
rect 3698 22752 3754 22808
rect 3514 20168 3570 20224
rect 3422 18536 3478 18592
rect 3606 18128 3662 18184
rect 3422 17620 3424 17640
rect 3424 17620 3476 17640
rect 3476 17620 3478 17640
rect 3422 17584 3478 17620
rect 3606 16108 3662 16144
rect 3606 16088 3608 16108
rect 3608 16088 3660 16108
rect 3660 16088 3662 16108
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2778 13776 2834 13832
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2870 13368 2926 13424
rect 3054 12860 3056 12880
rect 3056 12860 3108 12880
rect 3108 12860 3110 12880
rect 3054 12824 3110 12860
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 3422 13640 3478 13696
rect 3422 12300 3478 12336
rect 3422 12280 3424 12300
rect 3424 12280 3476 12300
rect 3476 12280 3478 12300
rect 3422 11192 3478 11248
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2870 9696 2926 9752
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 3882 20340 3884 20360
rect 3884 20340 3936 20360
rect 3936 20340 3938 20360
rect 3882 20304 3938 20340
rect 3882 16904 3938 16960
rect 4250 23432 4306 23488
rect 4618 23296 4674 23352
rect 4250 23060 4252 23080
rect 4252 23060 4304 23080
rect 4304 23060 4306 23080
rect 4250 23024 4306 23060
rect 4158 22072 4214 22128
rect 4158 20848 4214 20904
rect 3974 14492 3976 14512
rect 3976 14492 4028 14512
rect 4028 14492 4030 14512
rect 3974 14456 4030 14492
rect 3974 13252 4030 13288
rect 3974 13232 3976 13252
rect 3976 13232 4028 13252
rect 4028 13232 4030 13252
rect 3882 12980 3938 13016
rect 3882 12960 3884 12980
rect 3884 12960 3936 12980
rect 3936 12960 3938 12980
rect 3974 12688 4030 12744
rect 3882 11328 3938 11384
rect 3698 10512 3754 10568
rect 4158 11736 4214 11792
rect 4802 23568 4858 23624
rect 4710 17856 4766 17912
rect 5998 24656 6054 24712
rect 4802 15544 4858 15600
rect 4710 12552 4766 12608
rect 4618 11192 4674 11248
rect 5354 19352 5410 19408
rect 5814 21972 5816 21992
rect 5816 21972 5868 21992
rect 5868 21972 5870 21992
rect 5814 21936 5870 21972
rect 6550 25064 6606 25120
rect 5262 16532 5264 16552
rect 5264 16532 5316 16552
rect 5316 16532 5318 16552
rect 5262 16496 5318 16532
rect 5354 15700 5410 15736
rect 5354 15680 5356 15700
rect 5356 15680 5408 15700
rect 5408 15680 5410 15700
rect 5262 11620 5318 11656
rect 5262 11600 5264 11620
rect 5264 11600 5316 11620
rect 5316 11600 5318 11620
rect 5446 13640 5502 13696
rect 5722 20984 5778 21040
rect 5814 18264 5870 18320
rect 5998 14592 6054 14648
rect 6366 22072 6422 22128
rect 6182 18400 6238 18456
rect 6182 18128 6238 18184
rect 5722 11736 5778 11792
rect 5354 10920 5410 10976
rect 5170 10260 5226 10296
rect 5170 10240 5172 10260
rect 5172 10240 5224 10260
rect 5224 10240 5226 10260
rect 6182 12416 6238 12472
rect 5998 9288 6054 9344
rect 3514 8336 3570 8392
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 1306 7656 1362 7712
rect 6366 16632 6422 16688
rect 6826 26152 6882 26208
rect 6550 19116 6552 19136
rect 6552 19116 6604 19136
rect 6604 19116 6606 19136
rect 6550 19080 6606 19116
rect 6826 22652 6828 22672
rect 6828 22652 6880 22672
rect 6880 22652 6882 22672
rect 6826 22616 6882 22652
rect 6826 22108 6828 22128
rect 6828 22108 6880 22128
rect 6880 22108 6882 22128
rect 6826 22072 6882 22108
rect 6458 15816 6514 15872
rect 6366 13912 6422 13968
rect 6366 13776 6422 13832
rect 6734 15952 6790 16008
rect 6550 12416 6606 12472
rect 6734 12144 6790 12200
rect 7010 23432 7066 23488
rect 7654 24792 7710 24848
rect 7010 18808 7066 18864
rect 7010 17176 7066 17232
rect 7010 13776 7066 13832
rect 6642 9968 6698 10024
rect 1306 7248 1362 7304
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 1214 6840 1270 6896
rect 1306 6432 1362 6488
rect 1306 6024 1362 6080
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 1306 5652 1308 5672
rect 1308 5652 1360 5672
rect 1360 5652 1362 5672
rect 1306 5616 1362 5652
rect 2778 5208 2834 5264
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 1306 4820 1362 4856
rect 1306 4800 1308 4820
rect 1308 4800 1360 4820
rect 1360 4800 1362 4820
rect 1306 4392 1362 4448
rect 1306 3984 1362 4040
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 1214 3576 1270 3632
rect 1306 3188 1362 3224
rect 1306 3168 1308 3188
rect 1308 3168 1360 3188
rect 1360 3168 1362 3188
rect 1306 2760 1362 2816
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 1306 2388 1308 2408
rect 1308 2388 1360 2408
rect 1360 2388 1362 2408
rect 1306 2352 1362 2388
rect 1214 1944 1270 2000
rect 3238 1536 3294 1592
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7746 22480 7802 22536
rect 7470 18672 7526 18728
rect 7378 17176 7434 17232
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 8390 20476 8392 20496
rect 8392 20476 8444 20496
rect 8444 20476 8446 20496
rect 8390 20440 8446 20476
rect 8758 20304 8814 20360
rect 8298 19896 8354 19952
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 8206 19372 8262 19408
rect 8206 19352 8208 19372
rect 8208 19352 8260 19372
rect 8260 19352 8262 19372
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 8114 17212 8116 17232
rect 8116 17212 8168 17232
rect 8168 17212 8170 17232
rect 8114 17176 8170 17212
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 8022 15020 8078 15056
rect 8022 15000 8024 15020
rect 8024 15000 8076 15020
rect 8076 15000 8078 15020
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7378 10260 7434 10296
rect 7378 10240 7380 10260
rect 7380 10240 7432 10260
rect 7432 10240 7434 10260
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 8666 15544 8722 15600
rect 8390 9832 8446 9888
rect 7654 9560 7710 9616
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 9126 19660 9128 19680
rect 9128 19660 9180 19680
rect 9180 19660 9182 19680
rect 9126 19624 9182 19660
rect 9034 19216 9090 19272
rect 9402 23704 9458 23760
rect 9218 17604 9274 17640
rect 9218 17584 9220 17604
rect 9220 17584 9272 17604
rect 9272 17584 9274 17604
rect 9126 17448 9182 17504
rect 8942 15952 8998 16008
rect 8850 13368 8906 13424
rect 8482 8744 8538 8800
rect 8574 7656 8630 7712
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7470 3984 7526 4040
rect 8298 3576 8354 3632
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 9770 22344 9826 22400
rect 9770 21392 9826 21448
rect 11518 25200 11574 25256
rect 11058 22652 11060 22672
rect 11060 22652 11112 22672
rect 11112 22652 11114 22672
rect 11058 22616 11114 22652
rect 10138 21800 10194 21856
rect 11334 21664 11390 21720
rect 9862 19760 9918 19816
rect 9678 18808 9734 18864
rect 9586 17856 9642 17912
rect 9126 14728 9182 14784
rect 10046 15816 10102 15872
rect 10046 15564 10102 15600
rect 10046 15544 10048 15564
rect 10048 15544 10100 15564
rect 10100 15544 10102 15564
rect 9494 15428 9550 15464
rect 9494 15408 9496 15428
rect 9496 15408 9548 15428
rect 9548 15408 9550 15428
rect 9218 13640 9274 13696
rect 9310 12688 9366 12744
rect 9126 12552 9182 12608
rect 9126 10260 9182 10296
rect 9126 10240 9128 10260
rect 9128 10240 9180 10260
rect 9180 10240 9182 10260
rect 9402 10376 9458 10432
rect 9862 12008 9918 12064
rect 9862 10240 9918 10296
rect 9770 9560 9826 9616
rect 9494 7248 9550 7304
rect 11702 24132 11758 24168
rect 11702 24112 11704 24132
rect 11704 24112 11756 24132
rect 11756 24112 11758 24132
rect 11978 23568 12034 23624
rect 10506 18536 10562 18592
rect 10414 13368 10470 13424
rect 10230 12280 10286 12336
rect 10506 13096 10562 13152
rect 9954 8200 10010 8256
rect 10046 7948 10102 7984
rect 10046 7928 10048 7948
rect 10048 7928 10100 7948
rect 10100 7928 10102 7948
rect 11058 18964 11114 19000
rect 11058 18944 11060 18964
rect 11060 18944 11112 18964
rect 11112 18944 11114 18964
rect 10874 17720 10930 17776
rect 10966 16532 10968 16552
rect 10968 16532 11020 16552
rect 11020 16532 11022 16552
rect 10966 16496 11022 16532
rect 10966 15952 11022 16008
rect 10782 11736 10838 11792
rect 11058 14184 11114 14240
rect 11242 14048 11298 14104
rect 11058 12552 11114 12608
rect 11242 12416 11298 12472
rect 12162 23296 12218 23352
rect 12622 23296 12678 23352
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12806 23704 12862 23760
rect 12806 23432 12862 23488
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12622 23024 12678 23080
rect 12714 22072 12770 22128
rect 11886 20168 11942 20224
rect 11518 17720 11574 17776
rect 11794 18284 11850 18320
rect 11794 18264 11796 18284
rect 11796 18264 11848 18284
rect 11848 18264 11850 18284
rect 12070 18536 12126 18592
rect 11794 17720 11850 17776
rect 12070 17332 12126 17368
rect 12070 17312 12072 17332
rect 12072 17312 12124 17332
rect 12124 17312 12126 17332
rect 11794 17060 11850 17096
rect 11794 17040 11796 17060
rect 11796 17040 11848 17060
rect 11848 17040 11850 17060
rect 11978 16224 12034 16280
rect 11610 12960 11666 13016
rect 11978 15272 12034 15328
rect 13358 22344 13414 22400
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12990 20848 13046 20904
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 13634 21528 13690 21584
rect 13726 21256 13782 21312
rect 13542 20576 13598 20632
rect 12530 18808 12586 18864
rect 12530 18536 12586 18592
rect 12530 18148 12586 18184
rect 12530 18128 12532 18148
rect 12532 18128 12584 18148
rect 12584 18128 12586 18148
rect 12438 17856 12494 17912
rect 12346 17584 12402 17640
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12806 18400 12862 18456
rect 12438 17176 12494 17232
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 13634 19080 13690 19136
rect 13910 19488 13966 19544
rect 14462 22228 14518 22264
rect 14462 22208 14464 22228
rect 14464 22208 14516 22228
rect 14516 22208 14518 22228
rect 14646 22752 14702 22808
rect 14554 22072 14610 22128
rect 14094 20712 14150 20768
rect 14370 21120 14426 21176
rect 14738 21392 14794 21448
rect 14554 20032 14610 20088
rect 14554 19896 14610 19952
rect 13634 18264 13690 18320
rect 13542 17856 13598 17912
rect 12806 16904 12862 16960
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12990 15952 13046 16008
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12806 15564 12862 15600
rect 12806 15544 12808 15564
rect 12808 15544 12860 15564
rect 12860 15544 12862 15564
rect 12254 15000 12310 15056
rect 11978 13096 12034 13152
rect 11794 12008 11850 12064
rect 11702 11872 11758 11928
rect 11794 11328 11850 11384
rect 11242 11056 11298 11112
rect 11518 11056 11574 11112
rect 11610 10804 11666 10840
rect 11794 11056 11850 11112
rect 11610 10784 11612 10804
rect 11612 10784 11664 10804
rect 11664 10784 11666 10804
rect 11886 10376 11942 10432
rect 11610 10104 11666 10160
rect 11334 7540 11390 7576
rect 11334 7520 11336 7540
rect 11336 7520 11388 7540
rect 11388 7520 11390 7540
rect 11334 6840 11390 6896
rect 12346 13676 12348 13696
rect 12348 13676 12400 13696
rect 12400 13676 12402 13696
rect 12346 13640 12402 13676
rect 12438 12552 12494 12608
rect 13910 17312 13966 17368
rect 13542 16632 13598 16688
rect 12990 15272 13046 15328
rect 13634 15680 13690 15736
rect 13634 15308 13636 15328
rect 13636 15308 13688 15328
rect 13688 15308 13690 15328
rect 13634 15272 13690 15308
rect 13542 15020 13598 15056
rect 13542 15000 13544 15020
rect 13544 15000 13596 15020
rect 13596 15000 13598 15020
rect 12714 14728 12770 14784
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 13450 14592 13506 14648
rect 12622 12416 12678 12472
rect 12346 11872 12402 11928
rect 12070 9560 12126 9616
rect 11978 7404 12034 7440
rect 11978 7384 11980 7404
rect 11980 7384 12032 7404
rect 12032 7384 12034 7404
rect 12438 10376 12494 10432
rect 12530 10240 12586 10296
rect 12530 9696 12586 9752
rect 12346 6704 12402 6760
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 13174 13388 13230 13424
rect 13174 13368 13176 13388
rect 13176 13368 13228 13388
rect 13228 13368 13230 13388
rect 13266 12824 13322 12880
rect 13450 14320 13506 14376
rect 13450 14184 13506 14240
rect 13818 15952 13874 16008
rect 13726 14320 13782 14376
rect 13634 14220 13636 14240
rect 13636 14220 13688 14240
rect 13688 14220 13690 14240
rect 13634 14184 13690 14220
rect 13450 12844 13506 12880
rect 13450 12824 13452 12844
rect 13452 12824 13504 12844
rect 13504 12824 13506 12844
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12714 10804 12770 10840
rect 12714 10784 12716 10804
rect 12716 10784 12768 10804
rect 12768 10784 12770 10804
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 13542 12552 13598 12608
rect 13634 12008 13690 12064
rect 13358 9288 13414 9344
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 14278 17312 14334 17368
rect 14370 16088 14426 16144
rect 14370 15816 14426 15872
rect 14186 15000 14242 15056
rect 14094 13640 14150 13696
rect 14094 13504 14150 13560
rect 13910 11464 13966 11520
rect 15290 22752 15346 22808
rect 15014 20984 15070 21040
rect 14830 18028 14832 18048
rect 14832 18028 14884 18048
rect 14884 18028 14886 18048
rect 14830 17992 14886 18028
rect 15198 20984 15254 21040
rect 15382 20576 15438 20632
rect 15198 19796 15200 19816
rect 15200 19796 15252 19816
rect 15252 19796 15254 19816
rect 15198 19760 15254 19796
rect 16302 23704 16358 23760
rect 16946 24248 17002 24304
rect 16854 23724 16910 23760
rect 16854 23704 16856 23724
rect 16856 23704 16908 23724
rect 16908 23704 16910 23724
rect 16578 23160 16634 23216
rect 15658 20712 15714 20768
rect 16118 20460 16174 20496
rect 16118 20440 16120 20460
rect 16120 20440 16172 20460
rect 16172 20440 16174 20460
rect 16026 19760 16082 19816
rect 15106 18964 15162 19000
rect 15106 18944 15108 18964
rect 15108 18944 15160 18964
rect 15160 18944 15162 18964
rect 15014 18808 15070 18864
rect 14738 16768 14794 16824
rect 15106 16632 15162 16688
rect 14738 16108 14794 16144
rect 14738 16088 14740 16108
rect 14740 16088 14792 16108
rect 14792 16088 14794 16108
rect 15198 16360 15254 16416
rect 16026 19216 16082 19272
rect 16210 19080 16266 19136
rect 16026 18672 16082 18728
rect 15658 18400 15714 18456
rect 15566 17992 15622 18048
rect 14830 15000 14886 15056
rect 15014 14184 15070 14240
rect 15566 15952 15622 16008
rect 16302 18400 16358 18456
rect 16946 23432 17002 23488
rect 17130 23296 17186 23352
rect 16486 21664 16542 21720
rect 16762 21392 16818 21448
rect 16946 21392 17002 21448
rect 16946 20748 16948 20768
rect 16948 20748 17000 20768
rect 17000 20748 17002 20768
rect 16946 20712 17002 20748
rect 16486 20168 16542 20224
rect 16026 17076 16028 17096
rect 16028 17076 16080 17096
rect 16080 17076 16082 17096
rect 16026 17040 16082 17076
rect 16026 16360 16082 16416
rect 16026 16244 16082 16280
rect 16026 16224 16028 16244
rect 16028 16224 16080 16244
rect 16080 16224 16082 16244
rect 15934 15952 15990 16008
rect 16210 15680 16266 15736
rect 15842 15136 15898 15192
rect 14462 12008 14518 12064
rect 14370 11736 14426 11792
rect 13818 10104 13874 10160
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 13726 8472 13782 8528
rect 13726 6860 13782 6896
rect 13726 6840 13728 6860
rect 13728 6840 13780 6860
rect 13780 6840 13782 6860
rect 12346 6196 12348 6216
rect 12348 6196 12400 6216
rect 12400 6196 12402 6216
rect 12346 6160 12402 6196
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 14094 7792 14150 7848
rect 14646 12008 14702 12064
rect 14554 9560 14610 9616
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 14278 6704 14334 6760
rect 15198 12144 15254 12200
rect 14922 11756 14978 11792
rect 14922 11736 14924 11756
rect 14924 11736 14976 11756
rect 14976 11736 14978 11756
rect 15014 11464 15070 11520
rect 15566 13504 15622 13560
rect 15566 13368 15622 13424
rect 15382 10376 15438 10432
rect 15198 8608 15254 8664
rect 15106 7928 15162 7984
rect 16118 12416 16174 12472
rect 15842 11464 15898 11520
rect 15842 11056 15898 11112
rect 15842 10512 15898 10568
rect 16394 14728 16450 14784
rect 16118 11076 16174 11112
rect 16118 11056 16120 11076
rect 16120 11056 16172 11076
rect 16172 11056 16174 11076
rect 16026 9696 16082 9752
rect 16762 19352 16818 19408
rect 16578 15000 16634 15056
rect 17590 22072 17646 22128
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 18418 23296 18474 23352
rect 18694 23296 18750 23352
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17498 21836 17500 21856
rect 17500 21836 17552 21856
rect 17552 21836 17554 21856
rect 17498 21800 17554 21836
rect 18142 22616 18198 22672
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 18142 21564 18144 21584
rect 18144 21564 18196 21584
rect 18196 21564 18198 21584
rect 18142 21528 18198 21564
rect 18418 22616 18474 22672
rect 17130 19080 17186 19136
rect 16486 11056 16542 11112
rect 16210 8336 16266 8392
rect 17314 18128 17370 18184
rect 17222 17720 17278 17776
rect 17222 17448 17278 17504
rect 17314 16632 17370 16688
rect 17498 17312 17554 17368
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 19062 22888 19118 22944
rect 18970 22752 19026 22808
rect 18878 22480 18934 22536
rect 19062 22344 19118 22400
rect 19706 24132 19762 24168
rect 19706 24112 19708 24132
rect 19708 24112 19760 24132
rect 19760 24112 19762 24132
rect 19338 21664 19394 21720
rect 19154 20848 19210 20904
rect 18602 20168 18658 20224
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18786 20032 18842 20088
rect 18602 19624 18658 19680
rect 17774 19216 17830 19272
rect 17774 18536 17830 18592
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17958 18264 18014 18320
rect 17774 17992 17830 18048
rect 17130 15680 17186 15736
rect 17038 14864 17094 14920
rect 17222 14864 17278 14920
rect 17222 13912 17278 13968
rect 16670 8200 16726 8256
rect 16670 7112 16726 7168
rect 16946 11192 17002 11248
rect 17038 8472 17094 8528
rect 16670 6704 16726 6760
rect 17590 16496 17646 16552
rect 17590 15272 17646 15328
rect 17958 17584 18014 17640
rect 18326 17604 18382 17640
rect 18326 17584 18328 17604
rect 18328 17584 18380 17604
rect 18380 17584 18382 17604
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17958 16652 18014 16688
rect 18602 19080 18658 19136
rect 18510 17856 18566 17912
rect 18510 17448 18566 17504
rect 18786 17856 18842 17912
rect 17958 16632 17960 16652
rect 17960 16632 18012 16652
rect 18012 16632 18014 16652
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18326 16088 18382 16144
rect 17866 15680 17922 15736
rect 17222 8744 17278 8800
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18510 15136 18566 15192
rect 18418 14728 18474 14784
rect 18510 14048 18566 14104
rect 17590 10648 17646 10704
rect 17498 10376 17554 10432
rect 17406 10104 17462 10160
rect 17774 10920 17830 10976
rect 17774 10668 17830 10704
rect 17774 10648 17776 10668
rect 17776 10648 17828 10668
rect 17828 10648 17830 10668
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18694 15408 18750 15464
rect 18970 16652 19026 16688
rect 18970 16632 18972 16652
rect 18972 16632 19024 16652
rect 19024 16632 19026 16652
rect 18970 16496 19026 16552
rect 18878 15000 18934 15056
rect 19430 20748 19432 20768
rect 19432 20748 19484 20768
rect 19484 20748 19486 20768
rect 19430 20712 19486 20748
rect 19338 20324 19394 20360
rect 19338 20304 19340 20324
rect 19340 20304 19392 20324
rect 19392 20304 19394 20324
rect 19246 19352 19302 19408
rect 19246 18264 19302 18320
rect 19246 17992 19302 18048
rect 19522 17992 19578 18048
rect 19430 17720 19486 17776
rect 20074 24792 20130 24848
rect 19982 21256 20038 21312
rect 21086 23296 21142 23352
rect 21086 23044 21142 23080
rect 21086 23024 21088 23044
rect 21088 23024 21140 23044
rect 21140 23024 21142 23044
rect 20166 21664 20222 21720
rect 20258 20576 20314 20632
rect 19982 19760 20038 19816
rect 19982 19488 20038 19544
rect 20166 20168 20222 20224
rect 20166 19216 20222 19272
rect 20166 19080 20222 19136
rect 20258 18808 20314 18864
rect 20258 18536 20314 18592
rect 19798 17312 19854 17368
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17682 9288 17738 9344
rect 17590 8472 17646 8528
rect 18142 9968 18198 10024
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18602 11212 18658 11248
rect 18602 11192 18604 11212
rect 18604 11192 18656 11212
rect 18656 11192 18658 11212
rect 18786 11464 18842 11520
rect 18510 10920 18566 10976
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18050 8492 18106 8528
rect 18050 8472 18052 8492
rect 18052 8472 18104 8492
rect 18104 8472 18106 8492
rect 18694 9052 18696 9072
rect 18696 9052 18748 9072
rect 18748 9052 18750 9072
rect 18694 9016 18750 9052
rect 18418 8608 18474 8664
rect 18418 8336 18474 8392
rect 18142 8200 18198 8256
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17130 5208 17186 5264
rect 18970 10920 19026 10976
rect 18878 8744 18934 8800
rect 18878 8472 18934 8528
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 19246 13912 19302 13968
rect 19522 14900 19524 14920
rect 19524 14900 19576 14920
rect 19576 14900 19578 14920
rect 19522 14864 19578 14900
rect 19890 16088 19946 16144
rect 19890 15816 19946 15872
rect 19614 14592 19670 14648
rect 19338 12708 19394 12744
rect 19338 12688 19340 12708
rect 19340 12688 19392 12708
rect 19392 12688 19394 12708
rect 19246 11056 19302 11112
rect 19430 10920 19486 10976
rect 19430 10804 19486 10840
rect 19430 10784 19432 10804
rect 19432 10784 19484 10804
rect 19484 10784 19486 10804
rect 19154 10512 19210 10568
rect 19154 9968 19210 10024
rect 19430 9172 19486 9208
rect 19430 9152 19432 9172
rect 19432 9152 19484 9172
rect 19484 9152 19486 9172
rect 20626 20848 20682 20904
rect 20626 18536 20682 18592
rect 21638 24792 21694 24848
rect 21546 23432 21602 23488
rect 20994 20168 21050 20224
rect 21270 20204 21272 20224
rect 21272 20204 21324 20224
rect 21324 20204 21326 20224
rect 21270 20168 21326 20204
rect 21454 22208 21510 22264
rect 21454 20032 21510 20088
rect 21270 17720 21326 17776
rect 21362 17312 21418 17368
rect 21362 16224 21418 16280
rect 20534 14184 20590 14240
rect 20074 13912 20130 13968
rect 20350 13640 20406 13696
rect 20166 12144 20222 12200
rect 20442 11872 20498 11928
rect 20166 11056 20222 11112
rect 20350 10920 20406 10976
rect 18326 3576 18382 3632
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 21086 14340 21142 14376
rect 21086 14320 21088 14340
rect 21088 14320 21140 14340
rect 21140 14320 21142 14340
rect 22098 24248 22154 24304
rect 22558 25200 22614 25256
rect 22282 24656 22338 24712
rect 22098 21800 22154 21856
rect 22466 21800 22522 21856
rect 21730 19236 21786 19272
rect 21730 19216 21732 19236
rect 21732 19216 21784 19236
rect 21784 19216 21786 19236
rect 21638 16768 21694 16824
rect 21546 15680 21602 15736
rect 20166 9560 20222 9616
rect 20166 8472 20222 8528
rect 20718 8336 20774 8392
rect 20718 7248 20774 7304
rect 20902 7656 20958 7712
rect 21546 13640 21602 13696
rect 21362 10784 21418 10840
rect 21546 12960 21602 13016
rect 22466 20576 22522 20632
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 23202 23976 23258 24032
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22834 22752 22890 22808
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 23570 22888 23626 22944
rect 23846 23296 23902 23352
rect 23478 22344 23534 22400
rect 22742 22072 22798 22128
rect 22650 20884 22652 20904
rect 22652 20884 22704 20904
rect 22704 20884 22706 20904
rect 22650 20848 22706 20884
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22650 20576 22706 20632
rect 22558 20032 22614 20088
rect 22190 18944 22246 19000
rect 22834 20576 22890 20632
rect 22926 20340 22928 20360
rect 22928 20340 22980 20360
rect 22980 20340 22982 20360
rect 22926 20304 22982 20340
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 23662 22208 23718 22264
rect 23938 22208 23994 22264
rect 23754 21936 23810 21992
rect 23846 20712 23902 20768
rect 23478 19488 23534 19544
rect 23478 19372 23534 19408
rect 23478 19352 23480 19372
rect 23480 19352 23532 19372
rect 23532 19352 23534 19372
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22558 16632 22614 16688
rect 22466 16224 22522 16280
rect 22374 15680 22430 15736
rect 21914 14456 21970 14512
rect 22098 14456 22154 14512
rect 21822 14184 21878 14240
rect 22006 13776 22062 13832
rect 21730 11600 21786 11656
rect 21546 10784 21602 10840
rect 21730 8064 21786 8120
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 23294 16496 23350 16552
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22834 15272 22890 15328
rect 23110 15272 23166 15328
rect 23202 15000 23258 15056
rect 23938 19896 23994 19952
rect 23846 17584 23902 17640
rect 24214 23724 24270 23760
rect 24214 23704 24216 23724
rect 24216 23704 24268 23724
rect 24268 23704 24270 23724
rect 24122 23432 24178 23488
rect 24122 21664 24178 21720
rect 24306 21412 24362 21448
rect 24306 21392 24308 21412
rect 24308 21392 24360 21412
rect 24360 21392 24362 21412
rect 24490 20576 24546 20632
rect 24582 19780 24638 19816
rect 24582 19760 24584 19780
rect 24584 19760 24636 19780
rect 24636 19760 24638 19780
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22926 14456 22982 14512
rect 23386 14320 23442 14376
rect 22190 9868 22192 9888
rect 22192 9868 22244 9888
rect 22244 9868 22246 9888
rect 22190 9832 22246 9868
rect 22742 12960 22798 13016
rect 22374 9152 22430 9208
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 23018 13232 23074 13288
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 23478 13096 23534 13152
rect 23846 13912 23902 13968
rect 23386 10648 23442 10704
rect 22926 10512 22982 10568
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 23386 10124 23442 10160
rect 23386 10104 23388 10124
rect 23388 10104 23440 10124
rect 23440 10104 23442 10124
rect 23386 9560 23442 9616
rect 24030 16904 24086 16960
rect 24214 17176 24270 17232
rect 23938 11872 23994 11928
rect 22926 9424 22982 9480
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 23386 8880 23442 8936
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 24306 13368 24362 13424
rect 25502 26560 25558 26616
rect 25778 26288 25834 26344
rect 24766 21836 24768 21856
rect 24768 21836 24820 21856
rect 24820 21836 24822 21856
rect 24766 21800 24822 21836
rect 25134 22344 25190 22400
rect 24858 18944 24914 19000
rect 24950 18028 24952 18048
rect 24952 18028 25004 18048
rect 25004 18028 25006 18048
rect 24950 17992 25006 18028
rect 24766 16496 24822 16552
rect 24766 16108 24822 16144
rect 24766 16088 24768 16108
rect 24768 16088 24820 16108
rect 24820 16088 24822 16108
rect 25226 17448 25282 17504
rect 25686 23568 25742 23624
rect 25502 21956 25558 21992
rect 25502 21936 25504 21956
rect 25504 21936 25556 21956
rect 25556 21936 25558 21956
rect 24950 14456 25006 14512
rect 24122 10104 24178 10160
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 23754 3984 23810 4040
rect 24306 8472 24362 8528
rect 24582 8472 24638 8528
rect 25594 19216 25650 19272
rect 25962 20168 26018 20224
rect 25502 15952 25558 16008
rect 25778 16768 25834 16824
rect 25962 16904 26018 16960
rect 25686 15680 25742 15736
rect 25502 14592 25558 14648
rect 25318 13232 25374 13288
rect 25870 15544 25926 15600
rect 27342 23432 27398 23488
rect 26790 22208 26846 22264
rect 27158 22208 27214 22264
rect 26606 21392 26662 21448
rect 26514 20304 26570 20360
rect 26330 20168 26386 20224
rect 26514 18672 26570 18728
rect 26606 17992 26662 18048
rect 26882 19896 26938 19952
rect 27342 20168 27398 20224
rect 26882 18400 26938 18456
rect 27066 18420 27122 18456
rect 27066 18400 27068 18420
rect 27068 18400 27120 18420
rect 27120 18400 27122 18420
rect 27526 23976 27582 24032
rect 27342 19624 27398 19680
rect 27342 18400 27398 18456
rect 27066 17856 27122 17912
rect 26790 17332 26846 17368
rect 26790 17312 26792 17332
rect 26792 17312 26844 17332
rect 26844 17312 26846 17332
rect 26698 17076 26700 17096
rect 26700 17076 26752 17096
rect 26752 17076 26754 17096
rect 26698 17040 26754 17076
rect 26698 16108 26754 16144
rect 26698 16088 26700 16108
rect 26700 16088 26752 16108
rect 26752 16088 26754 16108
rect 26514 15272 26570 15328
rect 26606 15000 26662 15056
rect 26238 14728 26294 14784
rect 26054 11600 26110 11656
rect 24766 8628 24822 8664
rect 24766 8608 24768 8628
rect 24768 8608 24820 8628
rect 24820 8608 24822 8628
rect 25962 10124 26018 10160
rect 25962 10104 25964 10124
rect 25964 10104 26016 10124
rect 26016 10104 26018 10124
rect 25962 9832 26018 9888
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 24950 4020 24952 4040
rect 24952 4020 25004 4040
rect 25004 4020 25006 4040
rect 24950 3984 25006 4020
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 28354 23296 28410 23352
rect 28078 23060 28080 23080
rect 28080 23060 28132 23080
rect 28132 23060 28134 23080
rect 28078 23024 28134 23060
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 28538 23976 28594 24032
rect 28630 23432 28686 23488
rect 29182 24148 29184 24168
rect 29184 24148 29236 24168
rect 29236 24148 29238 24168
rect 29182 24112 29238 24148
rect 28722 23296 28778 23352
rect 28538 22752 28594 22808
rect 28722 23024 28778 23080
rect 28538 22344 28594 22400
rect 28538 22228 28594 22264
rect 28538 22208 28540 22228
rect 28540 22208 28592 22228
rect 28592 22208 28594 22228
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 27618 19760 27674 19816
rect 27342 18128 27398 18184
rect 27158 17040 27214 17096
rect 27710 19352 27766 19408
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 27158 16360 27214 16416
rect 27066 15544 27122 15600
rect 26974 15136 27030 15192
rect 26606 12144 26662 12200
rect 26422 10648 26478 10704
rect 27618 17720 27674 17776
rect 27802 18808 27858 18864
rect 27986 18672 28042 18728
rect 28262 19352 28318 19408
rect 28262 18944 28318 19000
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 28814 22072 28870 22128
rect 28906 21936 28962 21992
rect 29090 23180 29146 23216
rect 29090 23160 29092 23180
rect 29092 23160 29144 23180
rect 29144 23160 29146 23180
rect 29366 26152 29422 26208
rect 29090 22208 29146 22264
rect 28814 20984 28870 21040
rect 28446 17992 28502 18048
rect 27710 16904 27766 16960
rect 27526 16768 27582 16824
rect 27526 15580 27528 15600
rect 27528 15580 27580 15600
rect 27580 15580 27582 15600
rect 27526 15544 27582 15580
rect 27526 15272 27582 15328
rect 27526 14864 27582 14920
rect 27250 12824 27306 12880
rect 27250 12044 27252 12064
rect 27252 12044 27304 12064
rect 27304 12044 27306 12064
rect 27250 12008 27306 12044
rect 27342 9968 27398 10024
rect 28722 19216 28778 19272
rect 29090 20440 29146 20496
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 27986 17176 28042 17232
rect 27894 16632 27950 16688
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 27894 15680 27950 15736
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 27894 15000 27950 15056
rect 27986 14864 28042 14920
rect 28262 14864 28318 14920
rect 28262 14612 28318 14648
rect 28262 14592 28264 14612
rect 28264 14592 28316 14612
rect 28316 14592 28318 14612
rect 27710 14456 27766 14512
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 28446 15272 28502 15328
rect 28538 14764 28540 14784
rect 28540 14764 28592 14784
rect 28592 14764 28594 14784
rect 28538 14728 28594 14764
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 30746 25744 30802 25800
rect 29642 22072 29698 22128
rect 29918 23432 29974 23488
rect 29918 22072 29974 22128
rect 29274 20204 29276 20224
rect 29276 20204 29328 20224
rect 29328 20204 29330 20224
rect 29274 20168 29330 20204
rect 29274 20032 29330 20088
rect 29274 19372 29330 19408
rect 29274 19352 29276 19372
rect 29276 19352 29328 19372
rect 29328 19352 29330 19372
rect 29274 19236 29330 19272
rect 29274 19216 29276 19236
rect 29276 19216 29328 19236
rect 29328 19216 29330 19236
rect 29274 18944 29330 19000
rect 29182 16632 29238 16688
rect 28722 14592 28778 14648
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27618 11328 27674 11384
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27802 9968 27858 10024
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 28630 11636 28632 11656
rect 28632 11636 28684 11656
rect 28684 11636 28686 11656
rect 28630 11600 28686 11636
rect 28906 15000 28962 15056
rect 29090 15020 29146 15056
rect 29090 15000 29092 15020
rect 29092 15000 29144 15020
rect 29144 15000 29146 15020
rect 29182 14864 29238 14920
rect 29090 14184 29146 14240
rect 28906 13640 28962 13696
rect 28998 12280 29054 12336
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 29366 14764 29368 14784
rect 29368 14764 29420 14784
rect 29420 14764 29422 14784
rect 29366 14728 29422 14764
rect 30194 23296 30250 23352
rect 30286 21664 30342 21720
rect 29826 18944 29882 19000
rect 29826 18808 29882 18864
rect 30102 20440 30158 20496
rect 30654 23860 30710 23896
rect 30654 23840 30656 23860
rect 30656 23840 30708 23860
rect 30708 23840 30710 23860
rect 30470 19760 30526 19816
rect 30654 19760 30710 19816
rect 30562 19488 30618 19544
rect 30010 16652 30066 16688
rect 30010 16632 30012 16652
rect 30012 16632 30064 16652
rect 30064 16632 30066 16652
rect 29642 14728 29698 14784
rect 29826 14592 29882 14648
rect 30930 21392 30986 21448
rect 30470 18400 30526 18456
rect 29826 13640 29882 13696
rect 29366 12416 29422 12472
rect 29274 11328 29330 11384
rect 29182 9560 29238 9616
rect 30010 14340 30066 14376
rect 30010 14320 30012 14340
rect 30012 14320 30064 14340
rect 30064 14320 30066 14340
rect 29826 12280 29882 12336
rect 29550 7792 29606 7848
rect 30378 13776 30434 13832
rect 30470 13640 30526 13696
rect 30838 15136 30894 15192
rect 30194 12008 30250 12064
rect 30562 12144 30618 12200
rect 30470 11056 30526 11112
rect 30378 9832 30434 9888
rect 30562 10376 30618 10432
rect 30562 9696 30618 9752
rect 30194 7384 30250 7440
rect 31206 23432 31262 23488
rect 31022 13096 31078 13152
rect 31574 23432 31630 23488
rect 31482 23296 31538 23352
rect 31574 22636 31630 22672
rect 31574 22616 31576 22636
rect 31576 22616 31628 22636
rect 31628 22616 31630 22636
rect 31390 21800 31446 21856
rect 31666 22344 31722 22400
rect 31390 20748 31392 20768
rect 31392 20748 31444 20768
rect 31444 20748 31446 20768
rect 31390 20712 31446 20748
rect 32034 25336 32090 25392
rect 32034 23296 32090 23352
rect 32126 22480 32182 22536
rect 31850 22072 31906 22128
rect 31114 10648 31170 10704
rect 31390 19216 31446 19272
rect 31666 19080 31722 19136
rect 31758 18944 31814 19000
rect 32310 23704 32366 23760
rect 32310 22208 32366 22264
rect 32310 22072 32366 22128
rect 32770 25472 32826 25528
rect 32678 24792 32734 24848
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32862 24248 32918 24304
rect 32494 23432 32550 23488
rect 31942 19352 31998 19408
rect 31850 18808 31906 18864
rect 31482 16632 31538 16688
rect 31574 16360 31630 16416
rect 31666 15544 31722 15600
rect 31666 15136 31722 15192
rect 31574 15000 31630 15056
rect 31574 14184 31630 14240
rect 33046 23588 33102 23624
rect 33046 23568 33048 23588
rect 33048 23568 33100 23588
rect 33100 23568 33102 23588
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 33782 23432 33838 23488
rect 33322 23160 33378 23216
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 32770 21936 32826 21992
rect 32678 20576 32734 20632
rect 32862 21528 32918 21584
rect 32678 19896 32734 19952
rect 32218 17856 32274 17912
rect 31942 16632 31998 16688
rect 31942 15272 31998 15328
rect 31022 8744 31078 8800
rect 31206 9696 31262 9752
rect 31758 9696 31814 9752
rect 32218 12844 32274 12880
rect 32218 12824 32220 12844
rect 32220 12824 32272 12844
rect 32272 12824 32274 12844
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 33506 21528 33562 21584
rect 34702 25200 34758 25256
rect 34426 24792 34482 24848
rect 33966 24248 34022 24304
rect 33874 22752 33930 22808
rect 34150 23976 34206 24032
rect 34242 23296 34298 23352
rect 34150 22752 34206 22808
rect 33782 21836 33784 21856
rect 33784 21836 33836 21856
rect 33836 21836 33838 21856
rect 33782 21800 33838 21836
rect 33782 21140 33838 21176
rect 33782 21120 33784 21140
rect 33784 21120 33836 21140
rect 33836 21120 33838 21140
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 33230 19896 33286 19952
rect 33690 20848 33746 20904
rect 33598 19780 33654 19816
rect 32954 19352 33010 19408
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 32862 18808 32918 18864
rect 33046 18536 33102 18592
rect 33046 18264 33102 18320
rect 33598 19760 33600 19780
rect 33600 19760 33652 19780
rect 33652 19760 33654 19780
rect 33230 18164 33232 18184
rect 33232 18164 33284 18184
rect 33284 18164 33286 18184
rect 33230 18128 33286 18164
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 32862 17212 32864 17232
rect 32864 17212 32916 17232
rect 32916 17212 32918 17232
rect 32862 17176 32918 17212
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 33414 16496 33470 16552
rect 32862 16088 32918 16144
rect 32862 15952 32918 16008
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 32954 15308 32956 15328
rect 32956 15308 33008 15328
rect 33008 15308 33010 15328
rect 32954 15272 33010 15308
rect 32678 14728 32734 14784
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 32770 14592 32826 14648
rect 33598 19216 33654 19272
rect 33598 18672 33654 18728
rect 34058 21800 34114 21856
rect 33782 19236 33838 19272
rect 33782 19216 33784 19236
rect 33784 19216 33836 19236
rect 33836 19216 33838 19236
rect 33966 20440 34022 20496
rect 34518 22888 34574 22944
rect 34610 22480 34666 22536
rect 34702 21936 34758 21992
rect 34426 21664 34482 21720
rect 34426 20848 34482 20904
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 32862 13368 32918 13424
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 32770 11348 32826 11384
rect 32770 11328 32772 11348
rect 32772 11328 32824 11348
rect 32824 11328 32826 11348
rect 32586 9696 32642 9752
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 33690 15136 33746 15192
rect 34334 19252 34336 19272
rect 34336 19252 34388 19272
rect 34388 19252 34390 19272
rect 34334 19216 34390 19252
rect 34334 18692 34390 18728
rect 34334 18672 34336 18692
rect 34336 18672 34388 18692
rect 34388 18672 34390 18692
rect 34334 17856 34390 17912
rect 34702 19216 34758 19272
rect 34242 17584 34298 17640
rect 34334 16940 34336 16960
rect 34336 16940 34388 16960
rect 34388 16940 34390 16960
rect 34334 16904 34390 16940
rect 34058 16632 34114 16688
rect 33782 13912 33838 13968
rect 33782 12008 33838 12064
rect 33690 11872 33746 11928
rect 33690 11056 33746 11112
rect 33690 9832 33746 9888
rect 33046 8372 33048 8392
rect 33048 8372 33100 8392
rect 33100 8372 33102 8392
rect 33046 8336 33102 8372
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 33322 7828 33324 7848
rect 33324 7828 33376 7848
rect 33376 7828 33378 7848
rect 33322 7792 33378 7828
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 33966 13776 34022 13832
rect 34058 13524 34114 13560
rect 34058 13504 34060 13524
rect 34060 13504 34112 13524
rect 34112 13504 34114 13524
rect 34794 19080 34850 19136
rect 34702 18672 34758 18728
rect 34702 18300 34704 18320
rect 34704 18300 34756 18320
rect 34756 18300 34758 18320
rect 34702 18264 34758 18300
rect 34702 17040 34758 17096
rect 35254 21528 35310 21584
rect 35070 21392 35126 21448
rect 35070 20460 35126 20496
rect 35070 20440 35072 20460
rect 35072 20440 35124 20460
rect 35124 20440 35126 20460
rect 35162 20032 35218 20088
rect 35070 19896 35126 19952
rect 33966 12552 34022 12608
rect 33966 11464 34022 11520
rect 33782 9152 33838 9208
rect 33414 6024 33470 6080
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 34150 11092 34152 11112
rect 34152 11092 34204 11112
rect 34204 11092 34206 11112
rect 34150 11056 34206 11092
rect 34426 13676 34428 13696
rect 34428 13676 34480 13696
rect 34480 13676 34482 13696
rect 34426 13640 34482 13676
rect 34334 11464 34390 11520
rect 34334 10104 34390 10160
rect 34518 12144 34574 12200
rect 34518 10240 34574 10296
rect 34426 7928 34482 7984
rect 34886 13232 34942 13288
rect 35346 20984 35402 21040
rect 35346 20340 35348 20360
rect 35348 20340 35400 20360
rect 35400 20340 35402 20360
rect 35346 20304 35402 20340
rect 35254 18944 35310 19000
rect 35254 15952 35310 16008
rect 36082 26288 36138 26344
rect 35714 22208 35770 22264
rect 35530 22072 35586 22128
rect 35622 19624 35678 19680
rect 35438 18808 35494 18864
rect 35530 17992 35586 18048
rect 35898 21800 35954 21856
rect 35898 20576 35954 20632
rect 36174 25064 36230 25120
rect 36450 23840 36506 23896
rect 36358 23568 36414 23624
rect 36174 20712 36230 20768
rect 36082 20576 36138 20632
rect 35990 19760 36046 19816
rect 35898 19624 35954 19680
rect 35806 18128 35862 18184
rect 36818 23568 36874 23624
rect 36726 23296 36782 23352
rect 37002 23432 37058 23488
rect 36634 21256 36690 21312
rect 36542 20476 36544 20496
rect 36544 20476 36596 20496
rect 36596 20476 36598 20496
rect 36542 20440 36598 20476
rect 36082 18536 36138 18592
rect 36266 18128 36322 18184
rect 35714 17312 35770 17368
rect 35438 15272 35494 15328
rect 35346 14068 35402 14104
rect 35346 14048 35348 14068
rect 35348 14048 35400 14068
rect 35400 14048 35402 14068
rect 35530 15000 35586 15056
rect 35806 17040 35862 17096
rect 35990 15952 36046 16008
rect 35806 14728 35862 14784
rect 35254 11056 35310 11112
rect 36726 19896 36782 19952
rect 36450 19080 36506 19136
rect 36450 18400 36506 18456
rect 36726 18672 36782 18728
rect 36818 18400 36874 18456
rect 36450 17856 36506 17912
rect 36358 16768 36414 16824
rect 37462 20712 37518 20768
rect 37278 20576 37334 20632
rect 37002 19896 37058 19952
rect 36910 17720 36966 17776
rect 36726 17584 36782 17640
rect 36542 16904 36598 16960
rect 36266 13912 36322 13968
rect 36082 13776 36138 13832
rect 36174 13504 36230 13560
rect 36174 12416 36230 12472
rect 35162 9424 35218 9480
rect 35530 9460 35532 9480
rect 35532 9460 35584 9480
rect 35584 9460 35586 9480
rect 35530 9424 35586 9460
rect 36174 12008 36230 12064
rect 35806 11192 35862 11248
rect 36082 11192 36138 11248
rect 35898 9424 35954 9480
rect 35898 8880 35954 8936
rect 35898 8084 35954 8120
rect 35898 8064 35900 8084
rect 35900 8064 35952 8084
rect 35952 8064 35954 8084
rect 35806 6704 35862 6760
rect 36450 12008 36506 12064
rect 36910 16904 36966 16960
rect 36818 16360 36874 16416
rect 36818 15972 36874 16008
rect 36818 15952 36820 15972
rect 36820 15952 36872 15972
rect 36872 15952 36874 15972
rect 37002 16224 37058 16280
rect 37186 19488 37242 19544
rect 38290 26016 38346 26072
rect 37830 24928 37886 24984
rect 37738 23840 37794 23896
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 38382 23840 38438 23896
rect 37646 23432 37702 23488
rect 38566 23296 38622 23352
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 37738 22344 37794 22400
rect 38106 21936 38162 21992
rect 38934 23432 38990 23488
rect 38750 22888 38806 22944
rect 38658 22616 38714 22672
rect 37738 21664 37794 21720
rect 38382 21800 38438 21856
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 37830 21548 37886 21584
rect 37830 21528 37832 21548
rect 37832 21528 37884 21548
rect 37884 21528 37886 21548
rect 37646 21392 37702 21448
rect 37830 20984 37886 21040
rect 38566 21564 38568 21584
rect 38568 21564 38620 21584
rect 38620 21564 38622 21584
rect 38566 21528 38622 21564
rect 38934 23024 38990 23080
rect 38842 22108 38844 22128
rect 38844 22108 38896 22128
rect 38896 22108 38898 22128
rect 38842 22072 38898 22108
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 38474 20576 38530 20632
rect 37646 19352 37702 19408
rect 38382 20168 38438 20224
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 37278 18672 37334 18728
rect 37002 14864 37058 14920
rect 38198 19352 38254 19408
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 37646 17992 37702 18048
rect 38750 20168 38806 20224
rect 38474 19760 38530 19816
rect 38382 19352 38438 19408
rect 38750 18572 38752 18592
rect 38752 18572 38804 18592
rect 38804 18572 38806 18592
rect 38750 18536 38806 18572
rect 37462 16632 37518 16688
rect 37462 15680 37518 15736
rect 37370 13504 37426 13560
rect 37002 12280 37058 12336
rect 36910 11056 36966 11112
rect 36726 10920 36782 10976
rect 36542 10376 36598 10432
rect 36634 9868 36636 9888
rect 36636 9868 36688 9888
rect 36688 9868 36690 9888
rect 36634 9832 36690 9868
rect 35622 6432 35678 6488
rect 35898 5888 35954 5944
rect 35162 5208 35218 5264
rect 37462 11872 37518 11928
rect 37370 11328 37426 11384
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 38198 15000 38254 15056
rect 38750 17312 38806 17368
rect 39118 19896 39174 19952
rect 39118 18536 39174 18592
rect 38934 17448 38990 17504
rect 38658 16496 38714 16552
rect 38842 16360 38898 16416
rect 40958 26696 41014 26752
rect 39946 24384 40002 24440
rect 39394 20848 39450 20904
rect 39394 20576 39450 20632
rect 39578 20984 39634 21040
rect 39946 22616 40002 22672
rect 40038 22480 40094 22536
rect 39578 19216 39634 19272
rect 39486 18128 39542 18184
rect 40406 23432 40462 23488
rect 40314 22344 40370 22400
rect 40682 23160 40738 23216
rect 40498 23024 40554 23080
rect 40682 22752 40738 22808
rect 40406 22072 40462 22128
rect 40498 21664 40554 21720
rect 40222 20576 40278 20632
rect 40498 20848 40554 20904
rect 39854 20168 39910 20224
rect 40038 20204 40040 20224
rect 40040 20204 40092 20224
rect 40092 20204 40094 20224
rect 40038 20168 40094 20204
rect 39854 19896 39910 19952
rect 40406 20440 40462 20496
rect 40590 19896 40646 19952
rect 40498 19760 40554 19816
rect 38474 15408 38530 15464
rect 38290 14592 38346 14648
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 38842 15816 38898 15872
rect 38750 15272 38806 15328
rect 38934 15136 38990 15192
rect 38290 13812 38292 13832
rect 38292 13812 38344 13832
rect 38344 13812 38346 13832
rect 38290 13776 38346 13812
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 37738 12280 37794 12336
rect 37094 10804 37150 10840
rect 37094 10784 37096 10804
rect 37096 10784 37148 10804
rect 37148 10784 37150 10804
rect 37094 10376 37150 10432
rect 37002 9016 37058 9072
rect 36726 8880 36782 8936
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 37278 9696 37334 9752
rect 37186 9424 37242 9480
rect 37186 8744 37242 8800
rect 37462 11192 37518 11248
rect 37738 10920 37794 10976
rect 37462 9832 37518 9888
rect 37370 9152 37426 9208
rect 38382 12552 38438 12608
rect 38290 12280 38346 12336
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 38474 12280 38530 12336
rect 38934 13640 38990 13696
rect 38382 10920 38438 10976
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 37830 9424 37886 9480
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 40038 19216 40094 19272
rect 39854 18128 39910 18184
rect 40130 18400 40186 18456
rect 40314 18148 40370 18184
rect 40314 18128 40316 18148
rect 40316 18128 40368 18148
rect 40368 18128 40370 18148
rect 39762 16360 39818 16416
rect 40498 18128 40554 18184
rect 40590 16904 40646 16960
rect 40130 16224 40186 16280
rect 39670 15816 39726 15872
rect 39302 14492 39304 14512
rect 39304 14492 39356 14512
rect 39356 14492 39358 14512
rect 39302 14456 39358 14492
rect 39302 12824 39358 12880
rect 39118 11348 39174 11384
rect 39118 11328 39120 11348
rect 39120 11328 39172 11348
rect 39172 11328 39174 11348
rect 39026 9968 39082 10024
rect 38658 8880 38714 8936
rect 38842 9560 38898 9616
rect 38934 9424 38990 9480
rect 38750 8744 38806 8800
rect 39118 9424 39174 9480
rect 39578 15136 39634 15192
rect 39578 13912 39634 13968
rect 39762 14476 39818 14512
rect 39762 14456 39764 14476
rect 39764 14456 39816 14476
rect 39816 14456 39818 14476
rect 40498 16768 40554 16824
rect 40314 15136 40370 15192
rect 40222 14728 40278 14784
rect 40130 14340 40186 14376
rect 40130 14320 40132 14340
rect 40132 14320 40184 14340
rect 40184 14320 40186 14340
rect 39578 12588 39580 12608
rect 39580 12588 39632 12608
rect 39632 12588 39634 12608
rect 39578 12552 39634 12588
rect 40590 13912 40646 13968
rect 40498 13368 40554 13424
rect 40590 13232 40646 13288
rect 40498 12008 40554 12064
rect 39486 11192 39542 11248
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 38014 7404 38070 7440
rect 38014 7384 38016 7404
rect 38016 7384 38068 7404
rect 38068 7384 38070 7404
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 39210 8200 39266 8256
rect 39118 7248 39174 7304
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 38106 5228 38162 5264
rect 38106 5208 38108 5228
rect 38108 5208 38160 5228
rect 38160 5208 38162 5228
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 39578 9152 39634 9208
rect 39394 5616 39450 5672
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 39854 10376 39910 10432
rect 39854 9424 39910 9480
rect 40038 8508 40040 8528
rect 40040 8508 40092 8528
rect 40092 8508 40094 8528
rect 40038 8472 40094 8508
rect 40222 8064 40278 8120
rect 40130 7812 40186 7848
rect 40130 7792 40132 7812
rect 40132 7792 40184 7812
rect 40184 7792 40186 7812
rect 40038 6316 40094 6352
rect 40038 6296 40040 6316
rect 40040 6296 40092 6316
rect 40092 6296 40094 6316
rect 40958 21936 41014 21992
rect 40774 15816 40830 15872
rect 40958 21664 41014 21720
rect 41234 22516 41236 22536
rect 41236 22516 41288 22536
rect 41288 22516 41290 22536
rect 41234 22480 41290 22516
rect 41234 22344 41290 22400
rect 41234 22072 41290 22128
rect 41234 20848 41290 20904
rect 41142 20460 41198 20496
rect 41142 20440 41144 20460
rect 41144 20440 41196 20460
rect 41196 20440 41198 20460
rect 41418 21936 41474 21992
rect 41878 22208 41934 22264
rect 41602 21664 41658 21720
rect 41418 20304 41474 20360
rect 41326 20168 41382 20224
rect 40958 17332 41014 17368
rect 40958 17312 40960 17332
rect 40960 17312 41012 17332
rect 41012 17312 41014 17332
rect 40682 11192 40738 11248
rect 40866 15000 40922 15056
rect 40958 11056 41014 11112
rect 40958 10240 41014 10296
rect 41142 19388 41144 19408
rect 41144 19388 41196 19408
rect 41196 19388 41198 19408
rect 41142 19352 41198 19388
rect 41694 20848 41750 20904
rect 41878 20712 41934 20768
rect 42246 23976 42302 24032
rect 42430 23432 42486 23488
rect 42430 22636 42486 22672
rect 42430 22616 42432 22636
rect 42432 22616 42484 22636
rect 42484 22616 42486 22636
rect 42246 22208 42302 22264
rect 42246 21664 42302 21720
rect 41602 19080 41658 19136
rect 41510 18164 41512 18184
rect 41512 18164 41564 18184
rect 41564 18164 41566 18184
rect 41510 18128 41566 18164
rect 41234 17992 41290 18048
rect 41142 15272 41198 15328
rect 41326 16496 41382 16552
rect 41234 14728 41290 14784
rect 41326 13912 41382 13968
rect 41234 13640 41290 13696
rect 41418 9580 41474 9616
rect 41418 9560 41420 9580
rect 41420 9560 41472 9580
rect 41472 9560 41474 9580
rect 41694 16224 41750 16280
rect 41694 15816 41750 15872
rect 41602 10920 41658 10976
rect 41970 19252 41972 19272
rect 41972 19252 42024 19272
rect 42024 19252 42026 19272
rect 41970 19216 42026 19252
rect 41878 19080 41934 19136
rect 42062 18944 42118 19000
rect 42246 19116 42248 19136
rect 42248 19116 42300 19136
rect 42300 19116 42302 19136
rect 42246 19080 42302 19116
rect 41970 18400 42026 18456
rect 41970 17856 42026 17912
rect 42338 18672 42394 18728
rect 42246 18536 42302 18592
rect 42154 18400 42210 18456
rect 42154 18128 42210 18184
rect 42154 17584 42210 17640
rect 42338 17584 42394 17640
rect 42154 15272 42210 15328
rect 42062 13232 42118 13288
rect 42062 12144 42118 12200
rect 41786 8744 41842 8800
rect 41234 7792 41290 7848
rect 41510 8064 41566 8120
rect 42154 8608 42210 8664
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 42706 24248 42762 24304
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 42706 23296 42762 23352
rect 43258 23044 43314 23080
rect 43258 23024 43260 23044
rect 43260 23024 43312 23044
rect 43312 23024 43314 23044
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 43534 26016 43590 26072
rect 42798 21256 42854 21312
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 42706 21120 42762 21176
rect 42522 18808 42578 18864
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 44086 25200 44142 25256
rect 43902 23704 43958 23760
rect 43718 22752 43774 22808
rect 43442 19760 43498 19816
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 43350 17856 43406 17912
rect 42890 17312 42946 17368
rect 42798 17176 42854 17232
rect 43258 17076 43260 17096
rect 43260 17076 43312 17096
rect 43312 17076 43314 17096
rect 43258 17040 43314 17076
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 42798 16768 42854 16824
rect 42614 15952 42670 16008
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 42798 14612 42854 14648
rect 42798 14592 42800 14612
rect 42800 14592 42852 14612
rect 42852 14592 42854 14612
rect 43166 14476 43222 14512
rect 43166 14456 43168 14476
rect 43168 14456 43220 14476
rect 43220 14456 43222 14476
rect 42798 14048 42854 14104
rect 42706 13932 42762 13968
rect 42706 13912 42708 13932
rect 42708 13912 42760 13932
rect 42760 13912 42762 13932
rect 42430 11736 42486 11792
rect 42430 10784 42486 10840
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 42798 13524 42854 13560
rect 42798 13504 42800 13524
rect 42800 13504 42852 13524
rect 42852 13504 42854 13524
rect 42706 12824 42762 12880
rect 42614 11328 42670 11384
rect 42614 10104 42670 10160
rect 41602 6024 41658 6080
rect 41418 5208 41474 5264
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 43258 11192 43314 11248
rect 43718 19352 43774 19408
rect 44270 24928 44326 24984
rect 44086 22752 44142 22808
rect 44546 24656 44602 24712
rect 44454 23060 44456 23080
rect 44456 23060 44508 23080
rect 44508 23060 44510 23080
rect 44454 23024 44510 23060
rect 44362 20340 44364 20360
rect 44364 20340 44416 20360
rect 44416 20340 44418 20360
rect 44362 20304 44418 20340
rect 45650 26288 45706 26344
rect 45006 25472 45062 25528
rect 44822 22344 44878 22400
rect 44638 21392 44694 21448
rect 44638 21120 44694 21176
rect 44362 19488 44418 19544
rect 44270 18808 44326 18864
rect 45190 23568 45246 23624
rect 45374 23432 45430 23488
rect 45006 21800 45062 21856
rect 44914 20576 44970 20632
rect 44730 19080 44786 19136
rect 43902 18536 43958 18592
rect 43810 18128 43866 18184
rect 43810 16224 43866 16280
rect 44178 17992 44234 18048
rect 44086 17720 44142 17776
rect 44362 18284 44418 18320
rect 44362 18264 44364 18284
rect 44364 18264 44416 18284
rect 44416 18264 44418 18284
rect 44546 16360 44602 16416
rect 44086 14728 44142 14784
rect 43994 13368 44050 13424
rect 44730 16768 44786 16824
rect 43626 12552 43682 12608
rect 43534 12144 43590 12200
rect 43442 11192 43498 11248
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 43258 10104 43314 10160
rect 42890 9580 42946 9616
rect 42890 9560 42892 9580
rect 42892 9560 42944 9580
rect 42944 9560 42946 9580
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 42890 7928 42946 7984
rect 43534 8916 43536 8936
rect 43536 8916 43588 8936
rect 43588 8916 43590 8936
rect 43534 8880 43590 8916
rect 43442 8744 43498 8800
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 43350 6860 43406 6896
rect 43350 6840 43352 6860
rect 43352 6840 43404 6860
rect 43404 6840 43406 6860
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 43534 6976 43590 7032
rect 44362 11892 44418 11928
rect 44362 11872 44364 11892
rect 44364 11872 44416 11892
rect 44416 11872 44418 11892
rect 44178 11600 44234 11656
rect 44638 15444 44640 15464
rect 44640 15444 44692 15464
rect 44692 15444 44694 15464
rect 44638 15408 44694 15444
rect 44822 13640 44878 13696
rect 44546 11872 44602 11928
rect 44178 9560 44234 9616
rect 43902 8336 43958 8392
rect 44362 8472 44418 8528
rect 44730 11056 44786 11112
rect 44546 7656 44602 7712
rect 44454 7248 44510 7304
rect 44362 6704 44418 6760
rect 43442 5072 43498 5128
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 42706 4664 42762 4720
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 45282 19352 45338 19408
rect 45190 18400 45246 18456
rect 45098 16496 45154 16552
rect 44914 11756 44970 11792
rect 44914 11736 44916 11756
rect 44916 11736 44968 11756
rect 44968 11736 44970 11756
rect 45742 25880 45798 25936
rect 45926 25744 45982 25800
rect 45834 25064 45890 25120
rect 45650 20596 45706 20632
rect 45650 20576 45652 20596
rect 45652 20576 45704 20596
rect 45704 20576 45706 20596
rect 45558 19352 45614 19408
rect 45466 17448 45522 17504
rect 45650 17312 45706 17368
rect 45374 16360 45430 16416
rect 45466 15564 45522 15600
rect 45466 15544 45468 15564
rect 45468 15544 45520 15564
rect 45520 15544 45522 15564
rect 45374 15136 45430 15192
rect 45282 13776 45338 13832
rect 46662 25472 46718 25528
rect 46570 25336 46626 25392
rect 46018 23432 46074 23488
rect 46110 22616 46166 22672
rect 46294 22208 46350 22264
rect 46018 20576 46074 20632
rect 46202 21392 46258 21448
rect 46018 20168 46074 20224
rect 46110 19760 46166 19816
rect 46018 16904 46074 16960
rect 45834 15408 45890 15464
rect 45926 14864 45982 14920
rect 45190 9460 45192 9480
rect 45192 9460 45244 9480
rect 45244 9460 45246 9480
rect 45190 9424 45246 9460
rect 45006 7420 45008 7440
rect 45008 7420 45060 7440
rect 45060 7420 45062 7440
rect 45006 7384 45062 7420
rect 45190 7248 45246 7304
rect 45098 6060 45100 6080
rect 45100 6060 45152 6080
rect 45152 6060 45154 6080
rect 45098 6024 45154 6060
rect 45558 10104 45614 10160
rect 45466 6604 45468 6624
rect 45468 6604 45520 6624
rect 45520 6604 45522 6624
rect 45466 6568 45522 6604
rect 45006 5752 45062 5808
rect 45558 5616 45614 5672
rect 44730 4528 44786 4584
rect 45926 8200 45982 8256
rect 45926 6840 45982 6896
rect 46478 22072 46534 22128
rect 46662 24012 46664 24032
rect 46664 24012 46716 24032
rect 46716 24012 46718 24032
rect 46662 23976 46718 24012
rect 46386 20848 46442 20904
rect 46662 20984 46718 21040
rect 46294 17720 46350 17776
rect 46294 16360 46350 16416
rect 46570 17720 46626 17776
rect 46294 12688 46350 12744
rect 46110 11092 46112 11112
rect 46112 11092 46164 11112
rect 46164 11092 46166 11112
rect 46110 11056 46166 11092
rect 46110 10668 46166 10704
rect 46110 10648 46112 10668
rect 46112 10648 46164 10668
rect 46164 10648 46166 10668
rect 46202 10512 46258 10568
rect 46202 7404 46258 7440
rect 46938 24792 46994 24848
rect 46846 23432 46902 23488
rect 47030 24112 47086 24168
rect 47030 23568 47086 23624
rect 47214 23840 47270 23896
rect 47214 23568 47270 23624
rect 47030 22888 47086 22944
rect 46846 20984 46902 21040
rect 46938 20748 46940 20768
rect 46940 20748 46992 20768
rect 46992 20748 46994 20768
rect 46938 20712 46994 20748
rect 46938 19624 46994 19680
rect 46938 18808 46994 18864
rect 46754 16496 46810 16552
rect 47122 17992 47178 18048
rect 46938 16224 46994 16280
rect 46754 12300 46810 12336
rect 46754 12280 46756 12300
rect 46756 12280 46808 12300
rect 46808 12280 46810 12300
rect 47030 15952 47086 16008
rect 47214 16768 47270 16824
rect 47214 16668 47216 16688
rect 47216 16668 47268 16688
rect 47268 16668 47270 16688
rect 47214 16632 47270 16668
rect 47398 20576 47454 20632
rect 47398 18672 47454 18728
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 47306 13912 47362 13968
rect 47490 13404 47492 13424
rect 47492 13404 47544 13424
rect 47544 13404 47546 13424
rect 47490 13368 47546 13404
rect 47122 11892 47178 11928
rect 47122 11872 47124 11892
rect 47124 11872 47176 11892
rect 47176 11872 47178 11892
rect 46846 9560 46902 9616
rect 46386 7792 46442 7848
rect 46202 7384 46204 7404
rect 46204 7384 46256 7404
rect 46256 7384 46258 7404
rect 46018 6452 46074 6488
rect 46018 6432 46020 6452
rect 46020 6432 46072 6452
rect 46072 6432 46074 6452
rect 45926 6024 45982 6080
rect 46662 6180 46718 6216
rect 46662 6160 46664 6180
rect 46664 6160 46716 6180
rect 46716 6160 46718 6180
rect 46846 7928 46902 7984
rect 47214 6704 47270 6760
rect 47214 6296 47270 6352
rect 47398 11348 47454 11384
rect 47398 11328 47400 11348
rect 47400 11328 47452 11348
rect 47452 11328 47454 11348
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 48226 20440 48282 20496
rect 48410 20712 48466 20768
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 48226 19116 48228 19136
rect 48228 19116 48280 19136
rect 48280 19116 48282 19136
rect 48226 19080 48282 19116
rect 47950 18672 48006 18728
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 47858 18128 47914 18184
rect 47766 17992 47822 18048
rect 47766 17856 47822 17912
rect 47674 16088 47730 16144
rect 47674 15272 47730 15328
rect 47582 12824 47638 12880
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 47766 14184 47822 14240
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 48318 13504 48374 13560
rect 48962 25608 49018 25664
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 49054 21528 49110 21584
rect 48778 13368 48834 13424
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 48318 9016 48374 9072
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 48686 6296 48742 6352
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 48318 4664 48374 4720
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 46846 2624 46902 2680
rect 46754 1808 46810 1864
rect 46662 1400 46718 1456
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 48686 3032 48742 3088
rect 49146 19372 49202 19408
rect 49146 19352 49148 19372
rect 49148 19352 49200 19372
rect 49200 19352 49202 19372
rect 49146 18944 49202 19000
rect 49974 24656 50030 24712
rect 49882 24248 49938 24304
rect 49238 18264 49294 18320
rect 49422 19760 49478 19816
rect 49146 13268 49148 13288
rect 49148 13268 49200 13288
rect 49200 13268 49202 13288
rect 49146 13232 49202 13268
rect 49146 12844 49202 12880
rect 49146 12824 49148 12844
rect 49148 12824 49200 12844
rect 49200 12824 49202 12844
rect 49146 12416 49202 12472
rect 49146 12008 49202 12064
rect 49146 11600 49202 11656
rect 49330 11192 49386 11248
rect 49146 10784 49202 10840
rect 49422 10376 49478 10432
rect 49238 9968 49294 10024
rect 49146 9152 49202 9208
rect 49238 8744 49294 8800
rect 49330 8336 49386 8392
rect 49146 7520 49202 7576
rect 49238 7112 49294 7168
rect 49330 6704 49386 6760
rect 49146 5888 49202 5944
rect 49790 21120 49846 21176
rect 49790 18672 49846 18728
rect 49606 15680 49662 15736
rect 49790 18536 49846 18592
rect 50066 23840 50122 23896
rect 49974 23024 50030 23080
rect 50066 21800 50122 21856
rect 50066 20576 50122 20632
rect 49698 14456 49754 14512
rect 49514 6568 49570 6624
rect 49422 5480 49478 5536
rect 49238 5072 49294 5128
rect 49146 4256 49202 4312
rect 50066 14864 50122 14920
rect 50066 14728 50122 14784
rect 50066 7284 50068 7304
rect 50068 7284 50120 7304
rect 50120 7284 50122 7304
rect 50066 7248 50122 7284
rect 49882 6840 49938 6896
rect 49238 3848 49294 3904
rect 49146 3440 49202 3496
rect 48502 2216 48558 2272
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
<< metal3 >>
rect 24158 26692 24164 26756
rect 24228 26754 24234 26756
rect 40953 26754 41019 26757
rect 24228 26752 41019 26754
rect 24228 26696 40958 26752
rect 41014 26696 41019 26752
rect 24228 26694 41019 26696
rect 24228 26692 24234 26694
rect 40953 26691 41019 26694
rect 25497 26618 25563 26621
rect 47158 26618 47164 26620
rect 25497 26616 47164 26618
rect 25497 26560 25502 26616
rect 25558 26560 47164 26616
rect 25497 26558 47164 26560
rect 25497 26555 25563 26558
rect 47158 26556 47164 26558
rect 47228 26556 47234 26620
rect 25773 26346 25839 26349
rect 12390 26344 25839 26346
rect 12390 26288 25778 26344
rect 25834 26288 25839 26344
rect 12390 26286 25839 26288
rect 6821 26210 6887 26213
rect 12390 26210 12450 26286
rect 25773 26283 25839 26286
rect 36077 26346 36143 26349
rect 45645 26346 45711 26349
rect 36077 26344 45711 26346
rect 36077 26288 36082 26344
rect 36138 26288 45650 26344
rect 45706 26288 45711 26344
rect 36077 26286 45711 26288
rect 36077 26283 36143 26286
rect 45645 26283 45711 26286
rect 6821 26208 12450 26210
rect 6821 26152 6826 26208
rect 6882 26152 12450 26208
rect 6821 26150 12450 26152
rect 29361 26210 29427 26213
rect 46054 26210 46060 26212
rect 29361 26208 46060 26210
rect 29361 26152 29366 26208
rect 29422 26152 46060 26208
rect 29361 26150 46060 26152
rect 6821 26147 6887 26150
rect 29361 26147 29427 26150
rect 46054 26148 46060 26150
rect 46124 26148 46130 26212
rect 38285 26074 38351 26077
rect 43529 26074 43595 26077
rect 38285 26072 43595 26074
rect 38285 26016 38290 26072
rect 38346 26016 43534 26072
rect 43590 26016 43595 26072
rect 38285 26014 43595 26016
rect 38285 26011 38351 26014
rect 43529 26011 43595 26014
rect 30046 25876 30052 25940
rect 30116 25938 30122 25940
rect 45737 25938 45803 25941
rect 30116 25936 45803 25938
rect 30116 25880 45742 25936
rect 45798 25880 45803 25936
rect 30116 25878 45803 25880
rect 30116 25876 30122 25878
rect 45737 25875 45803 25878
rect 30741 25802 30807 25805
rect 45921 25802 45987 25805
rect 30741 25800 45987 25802
rect 30741 25744 30746 25800
rect 30802 25744 45926 25800
rect 45982 25744 45987 25800
rect 30741 25742 45987 25744
rect 30741 25739 30807 25742
rect 45921 25739 45987 25742
rect 0 25666 800 25696
rect 3417 25666 3483 25669
rect 0 25664 3483 25666
rect 0 25608 3422 25664
rect 3478 25608 3483 25664
rect 0 25606 3483 25608
rect 0 25576 800 25606
rect 3417 25603 3483 25606
rect 22502 25604 22508 25668
rect 22572 25666 22578 25668
rect 48957 25666 49023 25669
rect 22572 25664 49023 25666
rect 22572 25608 48962 25664
rect 49018 25608 49023 25664
rect 22572 25606 49023 25608
rect 22572 25604 22578 25606
rect 48957 25603 49023 25606
rect 32765 25530 32831 25533
rect 45001 25530 45067 25533
rect 32765 25528 45067 25530
rect 32765 25472 32770 25528
rect 32826 25472 45006 25528
rect 45062 25472 45067 25528
rect 32765 25470 45067 25472
rect 32765 25467 32831 25470
rect 45001 25467 45067 25470
rect 46657 25530 46723 25533
rect 50200 25530 51000 25560
rect 46657 25528 51000 25530
rect 46657 25472 46662 25528
rect 46718 25472 51000 25528
rect 46657 25470 51000 25472
rect 46657 25467 46723 25470
rect 50200 25440 51000 25470
rect 32029 25394 32095 25397
rect 46565 25394 46631 25397
rect 32029 25392 46631 25394
rect 32029 25336 32034 25392
rect 32090 25336 46570 25392
rect 46626 25336 46631 25392
rect 32029 25334 46631 25336
rect 32029 25331 32095 25334
rect 46565 25331 46631 25334
rect 0 25258 800 25288
rect 4061 25258 4127 25261
rect 0 25256 4127 25258
rect 0 25200 4066 25256
rect 4122 25200 4127 25256
rect 0 25198 4127 25200
rect 0 25168 800 25198
rect 4061 25195 4127 25198
rect 11513 25258 11579 25261
rect 22553 25258 22619 25261
rect 11513 25256 22619 25258
rect 11513 25200 11518 25256
rect 11574 25200 22558 25256
rect 22614 25200 22619 25256
rect 11513 25198 22619 25200
rect 11513 25195 11579 25198
rect 22553 25195 22619 25198
rect 34697 25258 34763 25261
rect 44081 25258 44147 25261
rect 34697 25256 44147 25258
rect 34697 25200 34702 25256
rect 34758 25200 44086 25256
rect 44142 25200 44147 25256
rect 34697 25198 44147 25200
rect 34697 25195 34763 25198
rect 44081 25195 44147 25198
rect 6545 25122 6611 25125
rect 19926 25122 19932 25124
rect 6545 25120 19932 25122
rect 6545 25064 6550 25120
rect 6606 25064 19932 25120
rect 6545 25062 19932 25064
rect 6545 25059 6611 25062
rect 19926 25060 19932 25062
rect 19996 25060 20002 25124
rect 36169 25122 36235 25125
rect 44214 25122 44220 25124
rect 36169 25120 44220 25122
rect 36169 25064 36174 25120
rect 36230 25064 44220 25120
rect 36169 25062 44220 25064
rect 36169 25059 36235 25062
rect 44214 25060 44220 25062
rect 44284 25060 44290 25124
rect 45829 25122 45895 25125
rect 50200 25122 51000 25152
rect 45829 25120 51000 25122
rect 45829 25064 45834 25120
rect 45890 25064 51000 25120
rect 45829 25062 51000 25064
rect 45829 25059 45895 25062
rect 50200 25032 51000 25062
rect 3366 24924 3372 24988
rect 3436 24986 3442 24988
rect 24894 24986 24900 24988
rect 3436 24926 24900 24986
rect 3436 24924 3442 24926
rect 24894 24924 24900 24926
rect 24964 24924 24970 24988
rect 37825 24986 37891 24989
rect 44265 24986 44331 24989
rect 37825 24984 44331 24986
rect 37825 24928 37830 24984
rect 37886 24928 44270 24984
rect 44326 24928 44331 24984
rect 37825 24926 44331 24928
rect 37825 24923 37891 24926
rect 44265 24923 44331 24926
rect 0 24850 800 24880
rect 3693 24850 3759 24853
rect 0 24848 3759 24850
rect 0 24792 3698 24848
rect 3754 24792 3759 24848
rect 0 24790 3759 24792
rect 0 24760 800 24790
rect 3693 24787 3759 24790
rect 7649 24850 7715 24853
rect 20069 24850 20135 24853
rect 7649 24848 20135 24850
rect 7649 24792 7654 24848
rect 7710 24792 20074 24848
rect 20130 24792 20135 24848
rect 7649 24790 20135 24792
rect 7649 24787 7715 24790
rect 20069 24787 20135 24790
rect 21633 24850 21699 24853
rect 32673 24850 32739 24853
rect 21633 24848 32739 24850
rect 21633 24792 21638 24848
rect 21694 24792 32678 24848
rect 32734 24792 32739 24848
rect 21633 24790 32739 24792
rect 21633 24787 21699 24790
rect 32673 24787 32739 24790
rect 34421 24850 34487 24853
rect 46933 24850 46999 24853
rect 34421 24848 46999 24850
rect 34421 24792 34426 24848
rect 34482 24792 46938 24848
rect 46994 24792 46999 24848
rect 34421 24790 46999 24792
rect 34421 24787 34487 24790
rect 46933 24787 46999 24790
rect 5993 24714 6059 24717
rect 22277 24714 22343 24717
rect 44541 24714 44607 24717
rect 5993 24712 22343 24714
rect 5993 24656 5998 24712
rect 6054 24656 22282 24712
rect 22338 24656 22343 24712
rect 5993 24654 22343 24656
rect 5993 24651 6059 24654
rect 22277 24651 22343 24654
rect 41370 24712 44607 24714
rect 41370 24656 44546 24712
rect 44602 24656 44607 24712
rect 41370 24654 44607 24656
rect 34646 24516 34652 24580
rect 34716 24578 34722 24580
rect 41370 24578 41430 24654
rect 44541 24651 44607 24654
rect 49969 24714 50035 24717
rect 50200 24714 51000 24744
rect 49969 24712 51000 24714
rect 49969 24656 49974 24712
rect 50030 24656 51000 24712
rect 49969 24654 51000 24656
rect 49969 24651 50035 24654
rect 50200 24624 51000 24654
rect 34716 24518 41430 24578
rect 34716 24516 34722 24518
rect 2946 24512 3262 24513
rect 0 24442 800 24472
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 2773 24442 2839 24445
rect 39941 24442 40007 24445
rect 0 24440 2839 24442
rect 0 24384 2778 24440
rect 2834 24384 2839 24440
rect 0 24382 2839 24384
rect 0 24352 800 24382
rect 2773 24379 2839 24382
rect 33366 24440 40007 24442
rect 33366 24384 39946 24440
rect 40002 24384 40007 24440
rect 33366 24382 40007 24384
rect 16941 24306 17007 24309
rect 22093 24306 22159 24309
rect 16941 24304 22159 24306
rect 16941 24248 16946 24304
rect 17002 24248 22098 24304
rect 22154 24248 22159 24304
rect 16941 24246 22159 24248
rect 16941 24243 17007 24246
rect 22093 24243 22159 24246
rect 32857 24306 32923 24309
rect 33366 24306 33426 24382
rect 39941 24379 40007 24382
rect 32857 24304 33426 24306
rect 32857 24248 32862 24304
rect 32918 24248 33426 24304
rect 32857 24246 33426 24248
rect 33961 24306 34027 24309
rect 42701 24306 42767 24309
rect 33961 24304 42767 24306
rect 33961 24248 33966 24304
rect 34022 24248 42706 24304
rect 42762 24248 42767 24304
rect 33961 24246 42767 24248
rect 32857 24243 32923 24246
rect 33961 24243 34027 24246
rect 42701 24243 42767 24246
rect 49877 24306 49943 24309
rect 50200 24306 51000 24336
rect 49877 24304 51000 24306
rect 49877 24248 49882 24304
rect 49938 24248 51000 24304
rect 49877 24246 51000 24248
rect 49877 24243 49943 24246
rect 50200 24216 51000 24246
rect 11697 24170 11763 24173
rect 19701 24170 19767 24173
rect 11697 24168 19767 24170
rect 11697 24112 11702 24168
rect 11758 24112 19706 24168
rect 19762 24112 19767 24168
rect 11697 24110 19767 24112
rect 11697 24107 11763 24110
rect 19701 24107 19767 24110
rect 29177 24170 29243 24173
rect 47025 24170 47091 24173
rect 29177 24168 47091 24170
rect 29177 24112 29182 24168
rect 29238 24112 47030 24168
rect 47086 24112 47091 24168
rect 29177 24110 47091 24112
rect 29177 24107 29243 24110
rect 47025 24107 47091 24110
rect 0 24034 800 24064
rect 3325 24034 3391 24037
rect 0 24032 3391 24034
rect 0 23976 3330 24032
rect 3386 23976 3391 24032
rect 0 23974 3391 23976
rect 0 23944 800 23974
rect 3325 23971 3391 23974
rect 23197 24034 23263 24037
rect 27521 24034 27587 24037
rect 23197 24032 27587 24034
rect 23197 23976 23202 24032
rect 23258 23976 27526 24032
rect 27582 23976 27587 24032
rect 23197 23974 27587 23976
rect 23197 23971 23263 23974
rect 27521 23971 27587 23974
rect 28533 24034 28599 24037
rect 34145 24034 34211 24037
rect 28533 24032 34211 24034
rect 28533 23976 28538 24032
rect 28594 23976 34150 24032
rect 34206 23976 34211 24032
rect 28533 23974 34211 23976
rect 28533 23971 28599 23974
rect 34145 23971 34211 23974
rect 40350 23972 40356 24036
rect 40420 24034 40426 24036
rect 42241 24034 42307 24037
rect 40420 24032 42307 24034
rect 40420 23976 42246 24032
rect 42302 23976 42307 24032
rect 40420 23974 42307 23976
rect 40420 23972 40426 23974
rect 42241 23971 42307 23974
rect 43662 23972 43668 24036
rect 43732 24034 43738 24036
rect 46657 24034 46723 24037
rect 43732 24032 46723 24034
rect 43732 23976 46662 24032
rect 46718 23976 46723 24032
rect 43732 23974 46723 23976
rect 43732 23972 43738 23974
rect 46657 23971 46723 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 30649 23898 30715 23901
rect 34462 23898 34468 23900
rect 30649 23896 34468 23898
rect 30649 23840 30654 23896
rect 30710 23840 34468 23896
rect 30649 23838 34468 23840
rect 30649 23835 30715 23838
rect 34462 23836 34468 23838
rect 34532 23836 34538 23900
rect 36445 23898 36511 23901
rect 37733 23898 37799 23901
rect 36445 23896 37799 23898
rect 36445 23840 36450 23896
rect 36506 23840 37738 23896
rect 37794 23840 37799 23896
rect 36445 23838 37799 23840
rect 36445 23835 36511 23838
rect 37733 23835 37799 23838
rect 38377 23898 38443 23901
rect 46974 23898 46980 23900
rect 38377 23896 46980 23898
rect 38377 23840 38382 23896
rect 38438 23840 46980 23896
rect 38377 23838 46980 23840
rect 38377 23835 38443 23838
rect 46974 23836 46980 23838
rect 47044 23898 47050 23900
rect 47209 23898 47275 23901
rect 47044 23896 47275 23898
rect 47044 23840 47214 23896
rect 47270 23840 47275 23896
rect 47044 23838 47275 23840
rect 47044 23836 47050 23838
rect 47209 23835 47275 23838
rect 50061 23898 50127 23901
rect 50200 23898 51000 23928
rect 50061 23896 51000 23898
rect 50061 23840 50066 23896
rect 50122 23840 51000 23896
rect 50061 23838 51000 23840
rect 50061 23835 50127 23838
rect 50200 23808 51000 23838
rect 3918 23700 3924 23764
rect 3988 23762 3994 23764
rect 9397 23762 9463 23765
rect 3988 23760 9463 23762
rect 3988 23704 9402 23760
rect 9458 23704 9463 23760
rect 3988 23702 9463 23704
rect 3988 23700 3994 23702
rect 9397 23699 9463 23702
rect 12801 23762 12867 23765
rect 16297 23762 16363 23765
rect 12801 23760 16363 23762
rect 12801 23704 12806 23760
rect 12862 23704 16302 23760
rect 16358 23704 16363 23760
rect 12801 23702 16363 23704
rect 12801 23699 12867 23702
rect 16297 23699 16363 23702
rect 16849 23762 16915 23765
rect 24209 23762 24275 23765
rect 16849 23760 24275 23762
rect 16849 23704 16854 23760
rect 16910 23704 24214 23760
rect 24270 23704 24275 23760
rect 16849 23702 24275 23704
rect 16849 23699 16915 23702
rect 24209 23699 24275 23702
rect 32305 23762 32371 23765
rect 43897 23762 43963 23765
rect 32305 23760 43963 23762
rect 32305 23704 32310 23760
rect 32366 23704 43902 23760
rect 43958 23704 43963 23760
rect 32305 23702 43963 23704
rect 32305 23699 32371 23702
rect 43897 23699 43963 23702
rect 0 23626 800 23656
rect 3693 23626 3759 23629
rect 0 23624 3759 23626
rect 0 23568 3698 23624
rect 3754 23568 3759 23624
rect 0 23566 3759 23568
rect 0 23536 800 23566
rect 3693 23563 3759 23566
rect 4797 23626 4863 23629
rect 7598 23626 7604 23628
rect 4797 23624 7604 23626
rect 4797 23568 4802 23624
rect 4858 23568 7604 23624
rect 4797 23566 7604 23568
rect 4797 23563 4863 23566
rect 7598 23564 7604 23566
rect 7668 23564 7674 23628
rect 11973 23626 12039 23629
rect 25681 23626 25747 23629
rect 11973 23624 25747 23626
rect 11973 23568 11978 23624
rect 12034 23568 25686 23624
rect 25742 23568 25747 23624
rect 11973 23566 25747 23568
rect 11973 23563 12039 23566
rect 25681 23563 25747 23566
rect 33041 23626 33107 23629
rect 34646 23626 34652 23628
rect 33041 23624 34652 23626
rect 33041 23568 33046 23624
rect 33102 23568 34652 23624
rect 33041 23566 34652 23568
rect 33041 23563 33107 23566
rect 34646 23564 34652 23566
rect 34716 23564 34722 23628
rect 36353 23626 36419 23629
rect 36486 23626 36492 23628
rect 36353 23624 36492 23626
rect 36353 23568 36358 23624
rect 36414 23568 36492 23624
rect 36353 23566 36492 23568
rect 36353 23563 36419 23566
rect 36486 23564 36492 23566
rect 36556 23564 36562 23628
rect 36813 23626 36879 23629
rect 45185 23626 45251 23629
rect 36813 23624 45251 23626
rect 36813 23568 36818 23624
rect 36874 23568 45190 23624
rect 45246 23568 45251 23624
rect 36813 23566 45251 23568
rect 36813 23563 36879 23566
rect 45185 23563 45251 23566
rect 47025 23626 47091 23629
rect 47209 23626 47275 23629
rect 47025 23624 47275 23626
rect 47025 23568 47030 23624
rect 47086 23568 47214 23624
rect 47270 23568 47275 23624
rect 47025 23566 47275 23568
rect 47025 23563 47091 23566
rect 47209 23563 47275 23566
rect 4245 23492 4311 23493
rect 4245 23488 4292 23492
rect 4356 23490 4362 23492
rect 7005 23490 7071 23493
rect 12801 23490 12867 23493
rect 4245 23432 4250 23488
rect 4245 23428 4292 23432
rect 4356 23430 4402 23490
rect 7005 23488 12867 23490
rect 7005 23432 7010 23488
rect 7066 23432 12806 23488
rect 12862 23432 12867 23488
rect 7005 23430 12867 23432
rect 4356 23428 4362 23430
rect 4245 23427 4311 23428
rect 7005 23427 7071 23430
rect 12801 23427 12867 23430
rect 16941 23490 17007 23493
rect 17166 23490 17172 23492
rect 16941 23488 17172 23490
rect 16941 23432 16946 23488
rect 17002 23432 17172 23488
rect 16941 23430 17172 23432
rect 16941 23427 17007 23430
rect 17166 23428 17172 23430
rect 17236 23428 17242 23492
rect 20662 23428 20668 23492
rect 20732 23490 20738 23492
rect 21541 23490 21607 23493
rect 20732 23488 21607 23490
rect 20732 23432 21546 23488
rect 21602 23432 21607 23488
rect 20732 23430 21607 23432
rect 20732 23428 20738 23430
rect 21541 23427 21607 23430
rect 23422 23428 23428 23492
rect 23492 23490 23498 23492
rect 24117 23490 24183 23493
rect 23492 23488 24183 23490
rect 23492 23432 24122 23488
rect 24178 23432 24183 23488
rect 23492 23430 24183 23432
rect 23492 23428 23498 23430
rect 24117 23427 24183 23430
rect 27337 23490 27403 23493
rect 27470 23490 27476 23492
rect 27337 23488 27476 23490
rect 27337 23432 27342 23488
rect 27398 23432 27476 23488
rect 27337 23430 27476 23432
rect 27337 23427 27403 23430
rect 27470 23428 27476 23430
rect 27540 23428 27546 23492
rect 28625 23490 28691 23493
rect 28758 23490 28764 23492
rect 28625 23488 28764 23490
rect 28625 23432 28630 23488
rect 28686 23432 28764 23488
rect 28625 23430 28764 23432
rect 28625 23427 28691 23430
rect 28758 23428 28764 23430
rect 28828 23428 28834 23492
rect 29913 23490 29979 23493
rect 30230 23490 30236 23492
rect 29913 23488 30236 23490
rect 29913 23432 29918 23488
rect 29974 23432 30236 23488
rect 29913 23430 30236 23432
rect 29913 23427 29979 23430
rect 30230 23428 30236 23430
rect 30300 23428 30306 23492
rect 30966 23428 30972 23492
rect 31036 23490 31042 23492
rect 31201 23490 31267 23493
rect 31569 23492 31635 23493
rect 32489 23492 32555 23493
rect 31518 23490 31524 23492
rect 31036 23488 31267 23490
rect 31036 23432 31206 23488
rect 31262 23432 31267 23488
rect 31036 23430 31267 23432
rect 31478 23430 31524 23490
rect 31588 23488 31635 23492
rect 32438 23490 32444 23492
rect 31630 23432 31635 23488
rect 31036 23428 31042 23430
rect 31201 23427 31267 23430
rect 31518 23428 31524 23430
rect 31588 23428 31635 23432
rect 32398 23430 32444 23490
rect 32508 23488 32555 23492
rect 32550 23432 32555 23488
rect 32438 23428 32444 23430
rect 32508 23428 32555 23432
rect 31569 23427 31635 23428
rect 32489 23427 32555 23428
rect 33777 23490 33843 23493
rect 34094 23490 34100 23492
rect 33777 23488 34100 23490
rect 33777 23432 33782 23488
rect 33838 23432 34100 23488
rect 33777 23430 34100 23432
rect 33777 23427 33843 23430
rect 34094 23428 34100 23430
rect 34164 23428 34170 23492
rect 36670 23428 36676 23492
rect 36740 23490 36746 23492
rect 36997 23490 37063 23493
rect 36740 23488 37063 23490
rect 36740 23432 37002 23488
rect 37058 23432 37063 23488
rect 36740 23430 37063 23432
rect 36740 23428 36746 23430
rect 36997 23427 37063 23430
rect 37641 23490 37707 23493
rect 38510 23490 38516 23492
rect 37641 23488 38516 23490
rect 37641 23432 37646 23488
rect 37702 23432 38516 23488
rect 37641 23430 38516 23432
rect 37641 23427 37707 23430
rect 38510 23428 38516 23430
rect 38580 23428 38586 23492
rect 38929 23490 38995 23493
rect 39430 23490 39436 23492
rect 38929 23488 39436 23490
rect 38929 23432 38934 23488
rect 38990 23432 39436 23488
rect 38929 23430 39436 23432
rect 38929 23427 38995 23430
rect 39430 23428 39436 23430
rect 39500 23428 39506 23492
rect 40401 23490 40467 23493
rect 40534 23490 40540 23492
rect 40401 23488 40540 23490
rect 40401 23432 40406 23488
rect 40462 23432 40540 23488
rect 40401 23430 40540 23432
rect 40401 23427 40467 23430
rect 40534 23428 40540 23430
rect 40604 23428 40610 23492
rect 42425 23490 42491 23493
rect 42558 23490 42564 23492
rect 42425 23488 42564 23490
rect 42425 23432 42430 23488
rect 42486 23432 42564 23488
rect 42425 23430 42564 23432
rect 42425 23427 42491 23430
rect 42558 23428 42564 23430
rect 42628 23428 42634 23492
rect 44950 23428 44956 23492
rect 45020 23490 45026 23492
rect 45369 23490 45435 23493
rect 45020 23488 45435 23490
rect 45020 23432 45374 23488
rect 45430 23432 45435 23488
rect 45020 23430 45435 23432
rect 45020 23428 45026 23430
rect 45369 23427 45435 23430
rect 46013 23490 46079 23493
rect 46841 23492 46907 23493
rect 46238 23490 46244 23492
rect 46013 23488 46244 23490
rect 46013 23432 46018 23488
rect 46074 23432 46244 23488
rect 46013 23430 46244 23432
rect 46013 23427 46079 23430
rect 46238 23428 46244 23430
rect 46308 23428 46314 23492
rect 46790 23490 46796 23492
rect 46750 23430 46796 23490
rect 46860 23488 46907 23492
rect 46902 23432 46907 23488
rect 46790 23428 46796 23430
rect 46860 23428 46907 23432
rect 48446 23428 48452 23492
rect 48516 23490 48522 23492
rect 50200 23490 51000 23520
rect 48516 23430 51000 23490
rect 48516 23428 48522 23430
rect 46841 23427 46907 23428
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 50200 23400 51000 23430
rect 42946 23359 43262 23360
rect 4613 23354 4679 23357
rect 12157 23354 12223 23357
rect 12617 23354 12683 23357
rect 17125 23354 17191 23357
rect 18413 23354 18479 23357
rect 4613 23352 12683 23354
rect 4613 23296 4618 23352
rect 4674 23296 12162 23352
rect 12218 23296 12622 23352
rect 12678 23296 12683 23352
rect 4613 23294 12683 23296
rect 4613 23291 4679 23294
rect 12157 23291 12223 23294
rect 12617 23291 12683 23294
rect 13494 23352 18479 23354
rect 13494 23296 17130 23352
rect 17186 23296 18418 23352
rect 18474 23296 18479 23352
rect 13494 23294 18479 23296
rect 0 23218 800 23248
rect 3233 23218 3299 23221
rect 0 23216 3299 23218
rect 0 23160 3238 23216
rect 3294 23160 3299 23216
rect 0 23158 3299 23160
rect 0 23128 800 23158
rect 3233 23155 3299 23158
rect 3417 23218 3483 23221
rect 13494 23218 13554 23294
rect 17125 23291 17191 23294
rect 18413 23291 18479 23294
rect 18689 23354 18755 23357
rect 21081 23354 21147 23357
rect 21214 23354 21220 23356
rect 18689 23352 21220 23354
rect 18689 23296 18694 23352
rect 18750 23296 21086 23352
rect 21142 23296 21220 23352
rect 18689 23294 21220 23296
rect 18689 23291 18755 23294
rect 21081 23291 21147 23294
rect 21214 23292 21220 23294
rect 21284 23292 21290 23356
rect 23841 23354 23907 23357
rect 28349 23354 28415 23357
rect 28717 23354 28783 23357
rect 23841 23352 28783 23354
rect 23841 23296 23846 23352
rect 23902 23296 28354 23352
rect 28410 23296 28722 23352
rect 28778 23296 28783 23352
rect 23841 23294 28783 23296
rect 23841 23291 23907 23294
rect 28349 23291 28415 23294
rect 28717 23291 28783 23294
rect 30046 23292 30052 23356
rect 30116 23354 30122 23356
rect 30189 23354 30255 23357
rect 30116 23352 30255 23354
rect 30116 23296 30194 23352
rect 30250 23296 30255 23352
rect 30116 23294 30255 23296
rect 30116 23292 30122 23294
rect 30189 23291 30255 23294
rect 31477 23354 31543 23357
rect 32029 23354 32095 23357
rect 31477 23352 32095 23354
rect 31477 23296 31482 23352
rect 31538 23296 32034 23352
rect 32090 23296 32095 23352
rect 31477 23294 32095 23296
rect 31477 23291 31543 23294
rect 32029 23291 32095 23294
rect 34237 23354 34303 23357
rect 36721 23354 36787 23357
rect 37406 23354 37412 23356
rect 34237 23352 35082 23354
rect 34237 23296 34242 23352
rect 34298 23296 35082 23352
rect 34237 23294 35082 23296
rect 34237 23291 34303 23294
rect 3417 23216 13554 23218
rect 3417 23160 3422 23216
rect 3478 23160 13554 23216
rect 3417 23158 13554 23160
rect 16573 23218 16639 23221
rect 29085 23218 29151 23221
rect 16573 23216 29151 23218
rect 16573 23160 16578 23216
rect 16634 23160 29090 23216
rect 29146 23160 29151 23216
rect 16573 23158 29151 23160
rect 3417 23155 3483 23158
rect 16573 23155 16639 23158
rect 29085 23155 29151 23158
rect 33317 23218 33383 23221
rect 34830 23218 34836 23220
rect 33317 23216 34836 23218
rect 33317 23160 33322 23216
rect 33378 23160 34836 23216
rect 33317 23158 34836 23160
rect 33317 23155 33383 23158
rect 34830 23156 34836 23158
rect 34900 23156 34906 23220
rect 35022 23218 35082 23294
rect 36721 23352 37412 23354
rect 36721 23296 36726 23352
rect 36782 23296 37412 23352
rect 36721 23294 37412 23296
rect 36721 23291 36787 23294
rect 37406 23292 37412 23294
rect 37476 23292 37482 23356
rect 38561 23354 38627 23357
rect 42701 23354 42767 23357
rect 38561 23352 42767 23354
rect 38561 23296 38566 23352
rect 38622 23296 42706 23352
rect 42762 23296 42767 23352
rect 38561 23294 42767 23296
rect 38561 23291 38627 23294
rect 42701 23291 42767 23294
rect 40677 23218 40743 23221
rect 35022 23216 40743 23218
rect 35022 23160 40682 23216
rect 40738 23160 40743 23216
rect 35022 23158 40743 23160
rect 40677 23155 40743 23158
rect 4245 23082 4311 23085
rect 5206 23082 5212 23084
rect 4245 23080 5212 23082
rect 4245 23024 4250 23080
rect 4306 23024 5212 23080
rect 4245 23022 5212 23024
rect 4245 23019 4311 23022
rect 5206 23020 5212 23022
rect 5276 23020 5282 23084
rect 12617 23082 12683 23085
rect 21081 23082 21147 23085
rect 28073 23082 28139 23085
rect 12617 23080 21147 23082
rect 12617 23024 12622 23080
rect 12678 23024 21086 23080
rect 21142 23024 21147 23080
rect 12617 23022 21147 23024
rect 12617 23019 12683 23022
rect 21081 23019 21147 23022
rect 21222 23080 28139 23082
rect 21222 23024 28078 23080
rect 28134 23024 28139 23080
rect 21222 23022 28139 23024
rect 19057 22946 19123 22949
rect 21222 22946 21282 23022
rect 28073 23019 28139 23022
rect 28717 23082 28783 23085
rect 38929 23082 38995 23085
rect 28717 23080 38995 23082
rect 28717 23024 28722 23080
rect 28778 23024 38934 23080
rect 38990 23024 38995 23080
rect 28717 23022 38995 23024
rect 28717 23019 28783 23022
rect 38929 23019 38995 23022
rect 40493 23082 40559 23085
rect 43253 23082 43319 23085
rect 40493 23080 43319 23082
rect 40493 23024 40498 23080
rect 40554 23024 43258 23080
rect 43314 23024 43319 23080
rect 40493 23022 43319 23024
rect 40493 23019 40559 23022
rect 43253 23019 43319 23022
rect 44030 23020 44036 23084
rect 44100 23082 44106 23084
rect 44449 23082 44515 23085
rect 44100 23080 44515 23082
rect 44100 23024 44454 23080
rect 44510 23024 44515 23080
rect 44100 23022 44515 23024
rect 44100 23020 44106 23022
rect 44449 23019 44515 23022
rect 49969 23082 50035 23085
rect 50200 23082 51000 23112
rect 49969 23080 51000 23082
rect 49969 23024 49974 23080
rect 50030 23024 51000 23080
rect 49969 23022 51000 23024
rect 49969 23019 50035 23022
rect 50200 22992 51000 23022
rect 23565 22946 23631 22949
rect 34513 22946 34579 22949
rect 19057 22944 21282 22946
rect 19057 22888 19062 22944
rect 19118 22888 21282 22944
rect 19057 22886 21282 22888
rect 21406 22944 23631 22946
rect 21406 22888 23570 22944
rect 23626 22888 23631 22944
rect 21406 22886 23631 22888
rect 19057 22883 19123 22886
rect 7946 22880 8262 22881
rect 0 22810 800 22840
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 3693 22810 3759 22813
rect 0 22808 3759 22810
rect 0 22752 3698 22808
rect 3754 22752 3759 22808
rect 0 22750 3759 22752
rect 0 22720 800 22750
rect 3693 22747 3759 22750
rect 9254 22748 9260 22812
rect 9324 22810 9330 22812
rect 14641 22810 14707 22813
rect 15285 22810 15351 22813
rect 9324 22808 15351 22810
rect 9324 22752 14646 22808
rect 14702 22752 15290 22808
rect 15346 22752 15351 22808
rect 9324 22750 15351 22752
rect 9324 22748 9330 22750
rect 14641 22747 14707 22750
rect 15285 22747 15351 22750
rect 18965 22810 19031 22813
rect 21406 22810 21466 22886
rect 23565 22883 23631 22886
rect 28398 22944 34579 22946
rect 28398 22888 34518 22944
rect 34574 22888 34579 22944
rect 28398 22886 34579 22888
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 18965 22808 21466 22810
rect 18965 22752 18970 22808
rect 19026 22752 21466 22808
rect 18965 22750 21466 22752
rect 18965 22747 19031 22750
rect 22134 22748 22140 22812
rect 22204 22810 22210 22812
rect 22829 22810 22895 22813
rect 22204 22808 22895 22810
rect 22204 22752 22834 22808
rect 22890 22752 22895 22808
rect 22204 22750 22895 22752
rect 22204 22748 22210 22750
rect 22829 22747 22895 22750
rect 5758 22612 5764 22676
rect 5828 22674 5834 22676
rect 6821 22674 6887 22677
rect 5828 22672 6887 22674
rect 5828 22616 6826 22672
rect 6882 22616 6887 22672
rect 5828 22614 6887 22616
rect 5828 22612 5834 22614
rect 6821 22611 6887 22614
rect 11053 22674 11119 22677
rect 18137 22674 18203 22677
rect 11053 22672 18203 22674
rect 11053 22616 11058 22672
rect 11114 22616 18142 22672
rect 18198 22616 18203 22672
rect 11053 22614 18203 22616
rect 11053 22611 11119 22614
rect 18137 22611 18203 22614
rect 18413 22674 18479 22677
rect 18413 22672 22110 22674
rect 18413 22616 18418 22672
rect 18474 22616 22110 22672
rect 18413 22614 22110 22616
rect 18413 22611 18479 22614
rect 7741 22538 7807 22541
rect 18873 22538 18939 22541
rect 7741 22536 18939 22538
rect 7741 22480 7746 22536
rect 7802 22480 18878 22536
rect 18934 22480 18939 22536
rect 7741 22478 18939 22480
rect 22050 22538 22110 22614
rect 27286 22612 27292 22676
rect 27356 22674 27362 22676
rect 28398 22674 28458 22886
rect 34513 22883 34579 22886
rect 38745 22946 38811 22949
rect 47025 22946 47091 22949
rect 38745 22944 47091 22946
rect 38745 22888 38750 22944
rect 38806 22888 47030 22944
rect 47086 22888 47091 22944
rect 38745 22886 47091 22888
rect 38745 22883 38811 22886
rect 47025 22883 47091 22886
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 47946 22815 48262 22816
rect 28533 22810 28599 22813
rect 33869 22810 33935 22813
rect 28533 22808 33935 22810
rect 28533 22752 28538 22808
rect 28594 22752 33874 22808
rect 33930 22752 33935 22808
rect 28533 22750 33935 22752
rect 28533 22747 28599 22750
rect 33869 22747 33935 22750
rect 34145 22810 34211 22813
rect 34278 22810 34284 22812
rect 34145 22808 34284 22810
rect 34145 22752 34150 22808
rect 34206 22752 34284 22808
rect 34145 22750 34284 22752
rect 34145 22747 34211 22750
rect 34278 22748 34284 22750
rect 34348 22748 34354 22812
rect 40677 22810 40743 22813
rect 43713 22810 43779 22813
rect 44081 22810 44147 22813
rect 40677 22808 44147 22810
rect 40677 22752 40682 22808
rect 40738 22752 43718 22808
rect 43774 22752 44086 22808
rect 44142 22752 44147 22808
rect 40677 22750 44147 22752
rect 40677 22747 40743 22750
rect 43713 22747 43779 22750
rect 44081 22747 44147 22750
rect 27356 22614 28458 22674
rect 31569 22674 31635 22677
rect 38653 22674 38719 22677
rect 31569 22672 38719 22674
rect 31569 22616 31574 22672
rect 31630 22616 38658 22672
rect 38714 22616 38719 22672
rect 31569 22614 38719 22616
rect 27356 22612 27362 22614
rect 31569 22611 31635 22614
rect 38653 22611 38719 22614
rect 39941 22674 40007 22677
rect 42425 22674 42491 22677
rect 39941 22672 42491 22674
rect 39941 22616 39946 22672
rect 40002 22616 42430 22672
rect 42486 22616 42491 22672
rect 39941 22614 42491 22616
rect 39941 22611 40007 22614
rect 42425 22611 42491 22614
rect 46105 22674 46171 22677
rect 50200 22674 51000 22704
rect 46105 22672 51000 22674
rect 46105 22616 46110 22672
rect 46166 22616 51000 22672
rect 46105 22614 51000 22616
rect 46105 22611 46171 22614
rect 50200 22584 51000 22614
rect 32121 22538 32187 22541
rect 34605 22538 34671 22541
rect 40033 22538 40099 22541
rect 22050 22536 32187 22538
rect 22050 22480 32126 22536
rect 32182 22480 32187 22536
rect 22050 22478 32187 22480
rect 7741 22475 7807 22478
rect 18873 22475 18939 22478
rect 32121 22475 32187 22478
rect 32814 22536 34671 22538
rect 32814 22480 34610 22536
rect 34666 22480 34671 22536
rect 32814 22478 34671 22480
rect 0 22402 800 22432
rect 9765 22404 9831 22405
rect 0 22342 2514 22402
rect 0 22312 800 22342
rect 2454 22130 2514 22342
rect 9765 22400 9812 22404
rect 9876 22402 9882 22404
rect 13353 22402 13419 22405
rect 19057 22402 19123 22405
rect 9765 22344 9770 22400
rect 9765 22340 9812 22344
rect 9876 22342 9922 22402
rect 13353 22400 19123 22402
rect 13353 22344 13358 22400
rect 13414 22344 19062 22400
rect 19118 22344 19123 22400
rect 13353 22342 19123 22344
rect 9876 22340 9882 22342
rect 9765 22339 9831 22340
rect 13353 22339 13419 22342
rect 19057 22339 19123 22342
rect 23473 22402 23539 22405
rect 25129 22402 25195 22405
rect 23473 22400 25195 22402
rect 23473 22344 23478 22400
rect 23534 22344 25134 22400
rect 25190 22344 25195 22400
rect 23473 22342 25195 22344
rect 23473 22339 23539 22342
rect 25129 22339 25195 22342
rect 25998 22340 26004 22404
rect 26068 22402 26074 22404
rect 28533 22402 28599 22405
rect 26068 22400 28599 22402
rect 26068 22344 28538 22400
rect 28594 22344 28599 22400
rect 26068 22342 28599 22344
rect 26068 22340 26074 22342
rect 28533 22339 28599 22342
rect 31661 22402 31727 22405
rect 32814 22402 32874 22478
rect 34605 22475 34671 22478
rect 34838 22536 40099 22538
rect 34838 22480 40038 22536
rect 40094 22480 40099 22536
rect 34838 22478 40099 22480
rect 31661 22400 32874 22402
rect 31661 22344 31666 22400
rect 31722 22344 32874 22400
rect 31661 22342 32874 22344
rect 31661 22339 31727 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 14457 22266 14523 22269
rect 21449 22266 21515 22269
rect 14457 22264 21515 22266
rect 14457 22208 14462 22264
rect 14518 22208 21454 22264
rect 21510 22208 21515 22264
rect 14457 22206 21515 22208
rect 14457 22203 14523 22206
rect 21449 22203 21515 22206
rect 23657 22266 23723 22269
rect 23790 22266 23796 22268
rect 23657 22264 23796 22266
rect 23657 22208 23662 22264
rect 23718 22208 23796 22264
rect 23657 22206 23796 22208
rect 23657 22203 23723 22206
rect 23790 22204 23796 22206
rect 23860 22204 23866 22268
rect 23933 22266 23999 22269
rect 26785 22266 26851 22269
rect 27153 22266 27219 22269
rect 23933 22264 27219 22266
rect 23933 22208 23938 22264
rect 23994 22208 26790 22264
rect 26846 22208 27158 22264
rect 27214 22208 27219 22264
rect 23933 22206 27219 22208
rect 23933 22203 23999 22206
rect 26785 22203 26851 22206
rect 27153 22203 27219 22206
rect 28533 22266 28599 22269
rect 29085 22266 29151 22269
rect 28533 22264 29151 22266
rect 28533 22208 28538 22264
rect 28594 22208 29090 22264
rect 29146 22208 29151 22264
rect 28533 22206 29151 22208
rect 28533 22203 28599 22206
rect 29085 22203 29151 22206
rect 29310 22204 29316 22268
rect 29380 22266 29386 22268
rect 32305 22266 32371 22269
rect 29380 22264 32371 22266
rect 29380 22208 32310 22264
rect 32366 22208 32371 22264
rect 29380 22206 32371 22208
rect 29380 22204 29386 22206
rect 32305 22203 32371 22206
rect 4153 22130 4219 22133
rect 2454 22128 4219 22130
rect 2454 22072 4158 22128
rect 4214 22072 4219 22128
rect 2454 22070 4219 22072
rect 4153 22067 4219 22070
rect 6361 22130 6427 22133
rect 6821 22130 6887 22133
rect 6361 22128 6887 22130
rect 6361 22072 6366 22128
rect 6422 22072 6826 22128
rect 6882 22072 6887 22128
rect 6361 22070 6887 22072
rect 6361 22067 6427 22070
rect 6821 22067 6887 22070
rect 11462 22068 11468 22132
rect 11532 22130 11538 22132
rect 12709 22130 12775 22133
rect 14549 22130 14615 22133
rect 11532 22128 12775 22130
rect 11532 22072 12714 22128
rect 12770 22072 12775 22128
rect 11532 22070 12775 22072
rect 11532 22068 11538 22070
rect 12709 22067 12775 22070
rect 14230 22128 14615 22130
rect 14230 22072 14554 22128
rect 14610 22072 14615 22128
rect 14230 22070 14615 22072
rect 0 21994 800 22024
rect 3233 21994 3299 21997
rect 0 21992 3299 21994
rect 0 21936 3238 21992
rect 3294 21936 3299 21992
rect 0 21934 3299 21936
rect 0 21904 800 21934
rect 3233 21931 3299 21934
rect 5574 21932 5580 21996
rect 5644 21994 5650 21996
rect 5809 21994 5875 21997
rect 14230 21994 14290 22070
rect 14549 22067 14615 22070
rect 17585 22130 17651 22133
rect 22737 22130 22803 22133
rect 17585 22128 22803 22130
rect 17585 22072 17590 22128
rect 17646 22072 22742 22128
rect 22798 22072 22803 22128
rect 17585 22070 22803 22072
rect 17585 22067 17651 22070
rect 22737 22067 22803 22070
rect 28809 22130 28875 22133
rect 29637 22130 29703 22133
rect 29913 22130 29979 22133
rect 28809 22128 29979 22130
rect 28809 22072 28814 22128
rect 28870 22072 29642 22128
rect 29698 22072 29918 22128
rect 29974 22072 29979 22128
rect 28809 22070 29979 22072
rect 28809 22067 28875 22070
rect 29637 22067 29703 22070
rect 29913 22067 29979 22070
rect 31334 22068 31340 22132
rect 31404 22130 31410 22132
rect 31845 22130 31911 22133
rect 31404 22128 31911 22130
rect 31404 22072 31850 22128
rect 31906 22072 31911 22128
rect 31404 22070 31911 22072
rect 31404 22068 31410 22070
rect 31845 22067 31911 22070
rect 32305 22130 32371 22133
rect 34838 22130 34898 22478
rect 40033 22475 40099 22478
rect 41086 22476 41092 22540
rect 41156 22538 41162 22540
rect 41229 22538 41295 22541
rect 41156 22536 41295 22538
rect 41156 22480 41234 22536
rect 41290 22480 41295 22536
rect 41156 22478 41295 22480
rect 41156 22476 41162 22478
rect 41229 22475 41295 22478
rect 41370 22478 43546 22538
rect 37590 22340 37596 22404
rect 37660 22402 37666 22404
rect 37733 22402 37799 22405
rect 37660 22400 37799 22402
rect 37660 22344 37738 22400
rect 37794 22344 37799 22400
rect 37660 22342 37799 22344
rect 37660 22340 37666 22342
rect 37733 22339 37799 22342
rect 40309 22402 40375 22405
rect 41229 22402 41295 22405
rect 40309 22400 41295 22402
rect 40309 22344 40314 22400
rect 40370 22344 41234 22400
rect 41290 22344 41295 22400
rect 40309 22342 41295 22344
rect 40309 22339 40375 22342
rect 41229 22339 41295 22342
rect 35709 22266 35775 22269
rect 35709 22264 39682 22266
rect 35709 22208 35714 22264
rect 35770 22208 39682 22264
rect 35709 22206 39682 22208
rect 35709 22203 35775 22206
rect 32305 22128 34898 22130
rect 32305 22072 32310 22128
rect 32366 22072 34898 22128
rect 32305 22070 34898 22072
rect 35525 22130 35591 22133
rect 38837 22130 38903 22133
rect 35525 22128 38903 22130
rect 35525 22072 35530 22128
rect 35586 22072 38842 22128
rect 38898 22072 38903 22128
rect 35525 22070 38903 22072
rect 39622 22130 39682 22206
rect 39798 22204 39804 22268
rect 39868 22266 39874 22268
rect 41370 22266 41430 22478
rect 43486 22402 43546 22478
rect 44817 22402 44883 22405
rect 45318 22402 45324 22404
rect 43486 22400 45324 22402
rect 43486 22344 44822 22400
rect 44878 22344 45324 22400
rect 43486 22342 45324 22344
rect 44817 22339 44883 22342
rect 45318 22340 45324 22342
rect 45388 22340 45394 22404
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 39868 22206 41430 22266
rect 41873 22266 41939 22269
rect 42241 22266 42307 22269
rect 41873 22264 42307 22266
rect 41873 22208 41878 22264
rect 41934 22208 42246 22264
rect 42302 22208 42307 22264
rect 41873 22206 42307 22208
rect 39868 22204 39874 22206
rect 41873 22203 41939 22206
rect 42241 22203 42307 22206
rect 46289 22266 46355 22269
rect 50200 22266 51000 22296
rect 46289 22264 51000 22266
rect 46289 22208 46294 22264
rect 46350 22208 51000 22264
rect 46289 22206 51000 22208
rect 46289 22203 46355 22206
rect 50200 22176 51000 22206
rect 40401 22130 40467 22133
rect 39622 22128 40467 22130
rect 39622 22072 40406 22128
rect 40462 22072 40467 22128
rect 39622 22070 40467 22072
rect 32305 22067 32371 22070
rect 35525 22067 35591 22070
rect 38837 22067 38903 22070
rect 40401 22067 40467 22070
rect 41229 22130 41295 22133
rect 46473 22130 46539 22133
rect 41229 22128 46539 22130
rect 41229 22072 41234 22128
rect 41290 22072 46478 22128
rect 46534 22072 46539 22128
rect 41229 22070 46539 22072
rect 41229 22067 41295 22070
rect 46473 22067 46539 22070
rect 23749 21994 23815 21997
rect 5644 21992 5875 21994
rect 5644 21936 5814 21992
rect 5870 21936 5875 21992
rect 5644 21934 5875 21936
rect 5644 21932 5650 21934
rect 5809 21931 5875 21934
rect 7790 21934 14290 21994
rect 17726 21992 23815 21994
rect 17726 21936 23754 21992
rect 23810 21936 23815 21992
rect 17726 21934 23815 21936
rect 1761 21858 1827 21861
rect 3417 21858 3483 21861
rect 7790 21858 7850 21934
rect 1761 21856 2790 21858
rect 1761 21800 1766 21856
rect 1822 21800 2790 21856
rect 1761 21798 2790 21800
rect 1761 21795 1827 21798
rect 2730 21722 2790 21798
rect 3417 21856 7850 21858
rect 3417 21800 3422 21856
rect 3478 21800 7850 21856
rect 3417 21798 7850 21800
rect 10133 21858 10199 21861
rect 17493 21858 17559 21861
rect 17726 21858 17786 21934
rect 23749 21931 23815 21934
rect 25497 21994 25563 21997
rect 28901 21996 28967 21997
rect 28901 21994 28948 21996
rect 25497 21992 28458 21994
rect 25497 21936 25502 21992
rect 25558 21936 28458 21992
rect 25497 21934 28458 21936
rect 28856 21992 28948 21994
rect 28856 21936 28906 21992
rect 28856 21934 28948 21936
rect 25497 21931 25563 21934
rect 10133 21856 16682 21858
rect 10133 21800 10138 21856
rect 10194 21800 16682 21856
rect 10133 21798 16682 21800
rect 3417 21795 3483 21798
rect 10133 21795 10199 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 7414 21722 7420 21724
rect 2730 21662 7420 21722
rect 7414 21660 7420 21662
rect 7484 21660 7490 21724
rect 11329 21722 11395 21725
rect 16481 21722 16547 21725
rect 11329 21720 16547 21722
rect 11329 21664 11334 21720
rect 11390 21664 16486 21720
rect 16542 21664 16547 21720
rect 11329 21662 16547 21664
rect 11329 21659 11395 21662
rect 16481 21659 16547 21662
rect 0 21586 800 21616
rect 2681 21586 2747 21589
rect 0 21584 2747 21586
rect 0 21528 2686 21584
rect 2742 21528 2747 21584
rect 0 21526 2747 21528
rect 0 21496 800 21526
rect 2681 21523 2747 21526
rect 13629 21586 13695 21589
rect 16622 21586 16682 21798
rect 17493 21856 17786 21858
rect 17493 21800 17498 21856
rect 17554 21800 17786 21856
rect 17493 21798 17786 21800
rect 22093 21858 22159 21861
rect 22318 21858 22324 21860
rect 22093 21856 22324 21858
rect 22093 21800 22098 21856
rect 22154 21800 22324 21856
rect 22093 21798 22324 21800
rect 17493 21795 17559 21798
rect 22093 21795 22159 21798
rect 22318 21796 22324 21798
rect 22388 21796 22394 21860
rect 22461 21858 22527 21861
rect 24761 21858 24827 21861
rect 22461 21856 24827 21858
rect 22461 21800 22466 21856
rect 22522 21800 24766 21856
rect 24822 21800 24827 21856
rect 22461 21798 24827 21800
rect 22461 21795 22527 21798
rect 24761 21795 24827 21798
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 19333 21722 19399 21725
rect 20161 21722 20227 21725
rect 24117 21724 24183 21725
rect 24117 21722 24164 21724
rect 19333 21720 24164 21722
rect 19333 21664 19338 21720
rect 19394 21664 20166 21720
rect 20222 21664 24122 21720
rect 19333 21662 24164 21664
rect 19333 21659 19399 21662
rect 20161 21659 20227 21662
rect 24117 21660 24164 21662
rect 24228 21660 24234 21724
rect 28398 21722 28458 21934
rect 28901 21932 28948 21934
rect 29012 21932 29018 21996
rect 32765 21994 32831 21997
rect 34697 21994 34763 21997
rect 32765 21992 34763 21994
rect 32765 21936 32770 21992
rect 32826 21936 34702 21992
rect 34758 21936 34763 21992
rect 32765 21934 34763 21936
rect 28901 21931 28967 21932
rect 32765 21931 32831 21934
rect 34697 21931 34763 21934
rect 35934 21932 35940 21996
rect 36004 21994 36010 21996
rect 38101 21994 38167 21997
rect 40953 21994 41019 21997
rect 41413 21994 41479 21997
rect 36004 21992 38167 21994
rect 36004 21936 38106 21992
rect 38162 21936 38167 21992
rect 36004 21934 38167 21936
rect 36004 21932 36010 21934
rect 38101 21931 38167 21934
rect 38932 21992 41019 21994
rect 38932 21936 40958 21992
rect 41014 21936 41019 21992
rect 38932 21934 41019 21936
rect 31385 21858 31451 21861
rect 33777 21858 33843 21861
rect 31385 21856 33843 21858
rect 31385 21800 31390 21856
rect 31446 21800 33782 21856
rect 33838 21800 33843 21856
rect 31385 21798 33843 21800
rect 31385 21795 31451 21798
rect 33777 21795 33843 21798
rect 34053 21858 34119 21861
rect 35893 21858 35959 21861
rect 34053 21856 35959 21858
rect 34053 21800 34058 21856
rect 34114 21800 35898 21856
rect 35954 21800 35959 21856
rect 34053 21798 35959 21800
rect 34053 21795 34119 21798
rect 35893 21795 35959 21798
rect 38377 21858 38443 21861
rect 38932 21858 38992 21934
rect 40953 21931 41019 21934
rect 41094 21992 41479 21994
rect 41094 21936 41418 21992
rect 41474 21936 41479 21992
rect 41094 21934 41479 21936
rect 38377 21856 38992 21858
rect 38377 21800 38382 21856
rect 38438 21800 38992 21856
rect 38377 21798 38992 21800
rect 38377 21795 38443 21798
rect 39062 21796 39068 21860
rect 39132 21858 39138 21860
rect 41094 21858 41154 21934
rect 41413 21931 41479 21934
rect 45001 21858 45067 21861
rect 39132 21798 41154 21858
rect 41370 21856 45067 21858
rect 41370 21800 45006 21856
rect 45062 21800 45067 21856
rect 41370 21798 45067 21800
rect 39132 21796 39138 21798
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 30281 21722 30347 21725
rect 34421 21722 34487 21725
rect 37733 21722 37799 21725
rect 40493 21722 40559 21725
rect 28398 21720 34487 21722
rect 28398 21664 30286 21720
rect 30342 21664 34426 21720
rect 34482 21664 34487 21720
rect 28398 21662 34487 21664
rect 24117 21659 24183 21660
rect 30281 21659 30347 21662
rect 34421 21659 34487 21662
rect 34838 21720 37799 21722
rect 34838 21664 37738 21720
rect 37794 21664 37799 21720
rect 34838 21662 37799 21664
rect 18137 21586 18203 21589
rect 32857 21586 32923 21589
rect 13629 21584 15026 21586
rect 13629 21528 13634 21584
rect 13690 21528 15026 21584
rect 13629 21526 15026 21528
rect 16622 21584 18203 21586
rect 16622 21528 18142 21584
rect 18198 21528 18203 21584
rect 16622 21526 18203 21528
rect 13629 21523 13695 21526
rect 9765 21450 9831 21453
rect 10174 21450 10180 21452
rect 9765 21448 10180 21450
rect 9765 21392 9770 21448
rect 9826 21392 10180 21448
rect 9765 21390 10180 21392
rect 9765 21387 9831 21390
rect 10174 21388 10180 21390
rect 10244 21450 10250 21452
rect 14733 21450 14799 21453
rect 10244 21448 14799 21450
rect 10244 21392 14738 21448
rect 14794 21392 14799 21448
rect 10244 21390 14799 21392
rect 14966 21450 15026 21526
rect 18137 21523 18203 21526
rect 18278 21584 32923 21586
rect 18278 21528 32862 21584
rect 32918 21528 32923 21584
rect 18278 21526 32923 21528
rect 16757 21450 16823 21453
rect 14966 21448 16823 21450
rect 14966 21392 16762 21448
rect 16818 21392 16823 21448
rect 14966 21390 16823 21392
rect 10244 21388 10250 21390
rect 14733 21387 14799 21390
rect 16757 21387 16823 21390
rect 16941 21450 17007 21453
rect 18278 21450 18338 21526
rect 32857 21523 32923 21526
rect 33501 21586 33567 21589
rect 34838 21586 34898 21662
rect 37733 21659 37799 21662
rect 38380 21720 40559 21722
rect 38380 21664 40498 21720
rect 40554 21664 40559 21720
rect 38380 21662 40559 21664
rect 33501 21584 34898 21586
rect 33501 21528 33506 21584
rect 33562 21528 34898 21584
rect 33501 21526 34898 21528
rect 35249 21586 35315 21589
rect 35750 21586 35756 21588
rect 35249 21584 35756 21586
rect 35249 21528 35254 21584
rect 35310 21528 35756 21584
rect 35249 21526 35756 21528
rect 33501 21523 33567 21526
rect 35249 21523 35315 21526
rect 35750 21524 35756 21526
rect 35820 21524 35826 21588
rect 37825 21586 37891 21589
rect 38380 21586 38440 21662
rect 40493 21659 40559 21662
rect 40953 21722 41019 21725
rect 41370 21722 41430 21798
rect 45001 21795 45067 21798
rect 50061 21858 50127 21861
rect 50200 21858 51000 21888
rect 50061 21856 51000 21858
rect 50061 21800 50066 21856
rect 50122 21800 51000 21856
rect 50061 21798 51000 21800
rect 50061 21795 50127 21798
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 50200 21768 51000 21798
rect 47946 21727 48262 21728
rect 40953 21720 41430 21722
rect 40953 21664 40958 21720
rect 41014 21664 41430 21720
rect 40953 21662 41430 21664
rect 41597 21722 41663 21725
rect 42241 21722 42307 21725
rect 41597 21720 42307 21722
rect 41597 21664 41602 21720
rect 41658 21664 42246 21720
rect 42302 21664 42307 21720
rect 41597 21662 42307 21664
rect 40953 21659 41019 21662
rect 41597 21659 41663 21662
rect 42241 21659 42307 21662
rect 37825 21584 38440 21586
rect 37825 21528 37830 21584
rect 37886 21528 38440 21584
rect 37825 21526 38440 21528
rect 38561 21586 38627 21589
rect 49049 21586 49115 21589
rect 38561 21584 49115 21586
rect 38561 21528 38566 21584
rect 38622 21528 49054 21584
rect 49110 21528 49115 21584
rect 38561 21526 49115 21528
rect 37825 21523 37891 21526
rect 38561 21523 38627 21526
rect 49049 21523 49115 21526
rect 24301 21450 24367 21453
rect 26601 21450 26667 21453
rect 16941 21448 18338 21450
rect 16941 21392 16946 21448
rect 17002 21392 18338 21448
rect 16941 21390 18338 21392
rect 22050 21390 23490 21450
rect 16941 21387 17007 21390
rect 13721 21314 13787 21317
rect 19977 21314 20043 21317
rect 13721 21312 20043 21314
rect 13721 21256 13726 21312
rect 13782 21256 19982 21312
rect 20038 21256 20043 21312
rect 13721 21254 20043 21256
rect 13721 21251 13787 21254
rect 19977 21251 20043 21254
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 0 21088 800 21118
rect 2773 21115 2839 21118
rect 14365 21178 14431 21181
rect 22050 21178 22110 21390
rect 23430 21314 23490 21390
rect 24301 21448 26667 21450
rect 24301 21392 24306 21448
rect 24362 21392 26606 21448
rect 26662 21392 26667 21448
rect 24301 21390 26667 21392
rect 24301 21387 24367 21390
rect 26601 21387 26667 21390
rect 30925 21450 30991 21453
rect 35065 21450 35131 21453
rect 30925 21448 35131 21450
rect 30925 21392 30930 21448
rect 30986 21392 35070 21448
rect 35126 21392 35131 21448
rect 30925 21390 35131 21392
rect 30925 21387 30991 21390
rect 35065 21387 35131 21390
rect 37641 21450 37707 21453
rect 44633 21450 44699 21453
rect 37641 21448 44699 21450
rect 37641 21392 37646 21448
rect 37702 21392 44638 21448
rect 44694 21392 44699 21448
rect 37641 21390 44699 21392
rect 37641 21387 37707 21390
rect 44633 21387 44699 21390
rect 46197 21450 46263 21453
rect 50200 21450 51000 21480
rect 46197 21448 51000 21450
rect 46197 21392 46202 21448
rect 46258 21392 51000 21448
rect 46197 21390 51000 21392
rect 46197 21387 46263 21390
rect 50200 21360 51000 21390
rect 26550 21314 26556 21316
rect 23430 21254 26556 21314
rect 26550 21252 26556 21254
rect 26620 21314 26626 21316
rect 36629 21314 36695 21317
rect 42793 21314 42859 21317
rect 26620 21254 31770 21314
rect 26620 21252 26626 21254
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 14365 21176 22110 21178
rect 14365 21120 14370 21176
rect 14426 21120 22110 21176
rect 14365 21118 22110 21120
rect 14365 21115 14431 21118
rect 5717 21042 5783 21045
rect 15009 21042 15075 21045
rect 5717 21040 15075 21042
rect 5717 20984 5722 21040
rect 5778 20984 15014 21040
rect 15070 20984 15075 21040
rect 5717 20982 15075 20984
rect 5717 20979 5783 20982
rect 15009 20979 15075 20982
rect 15193 21042 15259 21045
rect 28809 21042 28875 21045
rect 15193 21040 28875 21042
rect 15193 20984 15198 21040
rect 15254 20984 28814 21040
rect 28870 20984 28875 21040
rect 15193 20982 28875 20984
rect 31710 21042 31770 21254
rect 36629 21312 42859 21314
rect 36629 21256 36634 21312
rect 36690 21256 42798 21312
rect 42854 21256 42859 21312
rect 36629 21254 42859 21256
rect 36629 21251 36695 21254
rect 42793 21251 42859 21254
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 33777 21178 33843 21181
rect 42701 21178 42767 21181
rect 33777 21176 42767 21178
rect 33777 21120 33782 21176
rect 33838 21120 42706 21176
rect 42762 21120 42767 21176
rect 33777 21118 42767 21120
rect 33777 21115 33843 21118
rect 42701 21115 42767 21118
rect 44633 21178 44699 21181
rect 49785 21178 49851 21181
rect 44633 21176 49851 21178
rect 44633 21120 44638 21176
rect 44694 21120 49790 21176
rect 49846 21120 49851 21176
rect 44633 21118 49851 21120
rect 44633 21115 44699 21118
rect 49785 21115 49851 21118
rect 35341 21042 35407 21045
rect 37825 21042 37891 21045
rect 31710 21040 37891 21042
rect 31710 20984 35346 21040
rect 35402 20984 37830 21040
rect 37886 20984 37891 21040
rect 31710 20982 37891 20984
rect 15193 20979 15259 20982
rect 28809 20979 28875 20982
rect 35341 20979 35407 20982
rect 37825 20979 37891 20982
rect 39573 21042 39639 21045
rect 46657 21042 46723 21045
rect 39573 21040 46723 21042
rect 39573 20984 39578 21040
rect 39634 20984 46662 21040
rect 46718 20984 46723 21040
rect 39573 20982 46723 20984
rect 39573 20979 39639 20982
rect 46657 20979 46723 20982
rect 46841 21042 46907 21045
rect 50200 21042 51000 21072
rect 46841 21040 51000 21042
rect 46841 20984 46846 21040
rect 46902 20984 51000 21040
rect 46841 20982 51000 20984
rect 46841 20979 46907 20982
rect 50200 20952 51000 20982
rect 4153 20906 4219 20909
rect 4153 20904 9690 20906
rect 4153 20848 4158 20904
rect 4214 20848 9690 20904
rect 4153 20846 9690 20848
rect 4153 20843 4219 20846
rect 0 20770 800 20800
rect 1301 20770 1367 20773
rect 0 20768 1367 20770
rect 0 20712 1306 20768
rect 1362 20712 1367 20768
rect 0 20710 1367 20712
rect 0 20680 800 20710
rect 1301 20707 1367 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 9630 20634 9690 20846
rect 12566 20844 12572 20908
rect 12636 20906 12642 20908
rect 12985 20906 13051 20909
rect 19149 20906 19215 20909
rect 12636 20904 13051 20906
rect 12636 20848 12990 20904
rect 13046 20848 13051 20904
rect 12636 20846 13051 20848
rect 12636 20844 12642 20846
rect 12985 20843 13051 20846
rect 15518 20904 19215 20906
rect 15518 20848 19154 20904
rect 19210 20848 19215 20904
rect 15518 20846 19215 20848
rect 14089 20770 14155 20773
rect 15518 20770 15578 20846
rect 19149 20843 19215 20846
rect 20621 20906 20687 20909
rect 22645 20906 22711 20909
rect 33685 20906 33751 20909
rect 34421 20906 34487 20909
rect 39389 20906 39455 20909
rect 39614 20906 39620 20908
rect 20621 20904 22711 20906
rect 20621 20848 20626 20904
rect 20682 20848 22650 20904
rect 22706 20848 22711 20904
rect 20621 20846 22711 20848
rect 20621 20843 20687 20846
rect 22645 20843 22711 20846
rect 23844 20846 29010 20906
rect 23844 20773 23904 20846
rect 13310 20768 15578 20770
rect 13310 20712 14094 20768
rect 14150 20712 15578 20768
rect 13310 20710 15578 20712
rect 15653 20772 15719 20773
rect 16941 20772 17007 20773
rect 19425 20772 19491 20773
rect 15653 20768 15700 20772
rect 15764 20770 15770 20772
rect 15653 20712 15658 20768
rect 13310 20634 13370 20710
rect 14089 20707 14155 20710
rect 15653 20708 15700 20712
rect 15764 20710 15810 20770
rect 16941 20768 16988 20772
rect 17052 20770 17058 20772
rect 19374 20770 19380 20772
rect 16941 20712 16946 20768
rect 15764 20708 15770 20710
rect 16941 20708 16988 20712
rect 17052 20710 17098 20770
rect 19334 20710 19380 20770
rect 19444 20768 19491 20772
rect 19486 20712 19491 20768
rect 17052 20708 17058 20710
rect 19374 20708 19380 20710
rect 19444 20708 19491 20712
rect 15653 20707 15719 20708
rect 16941 20707 17007 20708
rect 19425 20707 19491 20708
rect 23841 20768 23907 20773
rect 23841 20712 23846 20768
rect 23902 20712 23907 20768
rect 23841 20707 23907 20712
rect 28950 20770 29010 20846
rect 33685 20904 34487 20906
rect 33685 20848 33690 20904
rect 33746 20848 34426 20904
rect 34482 20848 34487 20904
rect 33685 20846 34487 20848
rect 33685 20843 33751 20846
rect 34421 20843 34487 20846
rect 34654 20904 39620 20906
rect 34654 20848 39394 20904
rect 39450 20848 39620 20904
rect 34654 20846 39620 20848
rect 31385 20770 31451 20773
rect 34654 20770 34714 20846
rect 39389 20843 39455 20846
rect 39614 20844 39620 20846
rect 39684 20844 39690 20908
rect 40493 20906 40559 20909
rect 41229 20906 41295 20909
rect 40493 20904 41295 20906
rect 40493 20848 40498 20904
rect 40554 20848 41234 20904
rect 41290 20848 41295 20904
rect 40493 20846 41295 20848
rect 40493 20843 40559 20846
rect 41229 20843 41295 20846
rect 41689 20906 41755 20909
rect 41822 20906 41828 20908
rect 41689 20904 41828 20906
rect 41689 20848 41694 20904
rect 41750 20848 41828 20904
rect 41689 20846 41828 20848
rect 41689 20843 41755 20846
rect 41822 20844 41828 20846
rect 41892 20844 41898 20908
rect 45134 20844 45140 20908
rect 45204 20906 45210 20908
rect 46381 20906 46447 20909
rect 45204 20904 46447 20906
rect 45204 20848 46386 20904
rect 46442 20848 46447 20904
rect 45204 20846 46447 20848
rect 45204 20844 45210 20846
rect 46381 20843 46447 20846
rect 28950 20768 34714 20770
rect 28950 20712 31390 20768
rect 31446 20712 34714 20768
rect 28950 20710 34714 20712
rect 36169 20770 36235 20773
rect 37457 20770 37523 20773
rect 36169 20768 37523 20770
rect 36169 20712 36174 20768
rect 36230 20712 37462 20768
rect 37518 20712 37523 20768
rect 36169 20710 37523 20712
rect 31385 20707 31451 20710
rect 36169 20707 36235 20710
rect 37457 20707 37523 20710
rect 41873 20770 41939 20773
rect 46933 20770 46999 20773
rect 41873 20768 46999 20770
rect 41873 20712 41878 20768
rect 41934 20712 46938 20768
rect 46994 20712 46999 20768
rect 41873 20710 46999 20712
rect 41873 20707 41939 20710
rect 46933 20707 46999 20710
rect 48405 20770 48471 20773
rect 48630 20770 48636 20772
rect 48405 20768 48636 20770
rect 48405 20712 48410 20768
rect 48466 20712 48636 20768
rect 48405 20710 48636 20712
rect 48405 20707 48471 20710
rect 48630 20708 48636 20710
rect 48700 20708 48706 20772
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 9630 20574 13370 20634
rect 13537 20634 13603 20637
rect 15377 20634 15443 20637
rect 13537 20632 15443 20634
rect 13537 20576 13542 20632
rect 13598 20576 15382 20632
rect 15438 20576 15443 20632
rect 13537 20574 15443 20576
rect 13537 20571 13603 20574
rect 15377 20571 15443 20574
rect 20253 20634 20319 20637
rect 22461 20634 22527 20637
rect 22645 20634 22711 20637
rect 20253 20632 22711 20634
rect 20253 20576 20258 20632
rect 20314 20576 22466 20632
rect 22522 20576 22650 20632
rect 22706 20576 22711 20632
rect 20253 20574 22711 20576
rect 20253 20571 20319 20574
rect 22461 20571 22527 20574
rect 22645 20571 22711 20574
rect 22829 20634 22895 20637
rect 24485 20634 24551 20637
rect 22829 20632 24551 20634
rect 22829 20576 22834 20632
rect 22890 20576 24490 20632
rect 24546 20576 24551 20632
rect 22829 20574 24551 20576
rect 22829 20571 22895 20574
rect 24485 20571 24551 20574
rect 32673 20634 32739 20637
rect 35893 20634 35959 20637
rect 32673 20632 35959 20634
rect 32673 20576 32678 20632
rect 32734 20576 35898 20632
rect 35954 20576 35959 20632
rect 32673 20574 35959 20576
rect 32673 20571 32739 20574
rect 35893 20571 35959 20574
rect 36077 20634 36143 20637
rect 37273 20634 37339 20637
rect 36077 20632 37339 20634
rect 36077 20576 36082 20632
rect 36138 20576 37278 20632
rect 37334 20576 37339 20632
rect 36077 20574 37339 20576
rect 36077 20571 36143 20574
rect 37273 20571 37339 20574
rect 38469 20634 38535 20637
rect 39389 20634 39455 20637
rect 38469 20632 39455 20634
rect 38469 20576 38474 20632
rect 38530 20576 39394 20632
rect 39450 20576 39455 20632
rect 38469 20574 39455 20576
rect 38469 20571 38535 20574
rect 39389 20571 39455 20574
rect 40217 20634 40283 20637
rect 41270 20634 41276 20636
rect 40217 20632 41276 20634
rect 40217 20576 40222 20632
rect 40278 20576 41276 20632
rect 40217 20574 41276 20576
rect 40217 20571 40283 20574
rect 41270 20572 41276 20574
rect 41340 20572 41346 20636
rect 44909 20634 44975 20637
rect 45645 20634 45711 20637
rect 44909 20632 45711 20634
rect 44909 20576 44914 20632
rect 44970 20576 45650 20632
rect 45706 20576 45711 20632
rect 44909 20574 45711 20576
rect 44909 20571 44975 20574
rect 45645 20571 45711 20574
rect 46013 20634 46079 20637
rect 47393 20634 47459 20637
rect 46013 20632 47459 20634
rect 46013 20576 46018 20632
rect 46074 20576 47398 20632
rect 47454 20576 47459 20632
rect 46013 20574 47459 20576
rect 46013 20571 46079 20574
rect 47393 20571 47459 20574
rect 50061 20634 50127 20637
rect 50200 20634 51000 20664
rect 50061 20632 51000 20634
rect 50061 20576 50066 20632
rect 50122 20576 51000 20632
rect 50061 20574 51000 20576
rect 50061 20571 50127 20574
rect 50200 20544 51000 20574
rect 8385 20498 8451 20501
rect 16113 20498 16179 20501
rect 29085 20498 29151 20501
rect 8385 20496 29151 20498
rect 8385 20440 8390 20496
rect 8446 20440 16118 20496
rect 16174 20440 29090 20496
rect 29146 20440 29151 20496
rect 8385 20438 29151 20440
rect 8385 20435 8451 20438
rect 16113 20435 16179 20438
rect 29085 20435 29151 20438
rect 30097 20498 30163 20501
rect 33961 20498 34027 20501
rect 30097 20496 34027 20498
rect 30097 20440 30102 20496
rect 30158 20440 33966 20496
rect 34022 20440 34027 20496
rect 30097 20438 34027 20440
rect 30097 20435 30163 20438
rect 33961 20435 34027 20438
rect 34462 20436 34468 20500
rect 34532 20498 34538 20500
rect 35065 20498 35131 20501
rect 35198 20498 35204 20500
rect 34532 20496 35204 20498
rect 34532 20440 35070 20496
rect 35126 20440 35204 20496
rect 34532 20438 35204 20440
rect 34532 20436 34538 20438
rect 35065 20435 35131 20438
rect 35198 20436 35204 20438
rect 35268 20498 35274 20500
rect 36537 20498 36603 20501
rect 39798 20498 39804 20500
rect 35268 20438 36416 20498
rect 35268 20436 35274 20438
rect 0 20362 800 20392
rect 3877 20362 3943 20365
rect 0 20360 3943 20362
rect 0 20304 3882 20360
rect 3938 20304 3943 20360
rect 0 20302 3943 20304
rect 0 20272 800 20302
rect 3877 20299 3943 20302
rect 8753 20362 8819 20365
rect 8886 20362 8892 20364
rect 8753 20360 8892 20362
rect 8753 20304 8758 20360
rect 8814 20304 8892 20360
rect 8753 20302 8892 20304
rect 8753 20299 8819 20302
rect 8886 20300 8892 20302
rect 8956 20300 8962 20364
rect 19333 20362 19399 20365
rect 22921 20362 22987 20365
rect 26509 20362 26575 20365
rect 35341 20364 35407 20365
rect 12390 20360 26575 20362
rect 12390 20304 19338 20360
rect 19394 20304 22926 20360
rect 22982 20304 26514 20360
rect 26570 20304 26575 20360
rect 12390 20302 26575 20304
rect 3509 20226 3575 20229
rect 11881 20226 11947 20229
rect 3509 20224 11947 20226
rect 3509 20168 3514 20224
rect 3570 20168 11886 20224
rect 11942 20168 11947 20224
rect 3509 20166 11947 20168
rect 3509 20163 3575 20166
rect 11881 20163 11947 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 0 19954 800 19984
rect 3325 19954 3391 19957
rect 0 19952 3391 19954
rect 0 19896 3330 19952
rect 3386 19896 3391 19952
rect 0 19894 3391 19896
rect 0 19864 800 19894
rect 3325 19891 3391 19894
rect 8293 19954 8359 19957
rect 12390 19954 12450 20302
rect 19333 20299 19399 20302
rect 22921 20299 22987 20302
rect 26509 20299 26575 20302
rect 29318 20302 34576 20362
rect 29318 20229 29378 20302
rect 16481 20226 16547 20229
rect 18597 20226 18663 20229
rect 16481 20224 18663 20226
rect 16481 20168 16486 20224
rect 16542 20168 18602 20224
rect 18658 20168 18663 20224
rect 16481 20166 18663 20168
rect 16481 20163 16547 20166
rect 18597 20163 18663 20166
rect 20161 20226 20227 20229
rect 20989 20226 21055 20229
rect 21265 20226 21331 20229
rect 20161 20224 21331 20226
rect 20161 20168 20166 20224
rect 20222 20168 20994 20224
rect 21050 20168 21270 20224
rect 21326 20168 21331 20224
rect 20161 20166 21331 20168
rect 20161 20163 20227 20166
rect 20989 20163 21055 20166
rect 21265 20163 21331 20166
rect 25957 20226 26023 20229
rect 26325 20226 26391 20229
rect 25957 20224 26391 20226
rect 25957 20168 25962 20224
rect 26018 20168 26330 20224
rect 26386 20168 26391 20224
rect 25957 20166 26391 20168
rect 25957 20163 26023 20166
rect 26325 20163 26391 20166
rect 27337 20226 27403 20229
rect 29269 20226 29378 20229
rect 27337 20224 29378 20226
rect 27337 20168 27342 20224
rect 27398 20168 29274 20224
rect 29330 20168 29378 20224
rect 27337 20166 29378 20168
rect 34516 20226 34576 20302
rect 34646 20300 34652 20364
rect 34716 20362 34722 20364
rect 35341 20362 35388 20364
rect 34716 20360 35388 20362
rect 34716 20304 35346 20360
rect 34716 20302 35388 20304
rect 34716 20300 34722 20302
rect 35341 20300 35388 20302
rect 35452 20300 35458 20364
rect 36356 20362 36416 20438
rect 36537 20496 39804 20498
rect 36537 20440 36542 20496
rect 36598 20440 39804 20496
rect 36537 20438 39804 20440
rect 36537 20435 36603 20438
rect 39798 20436 39804 20438
rect 39868 20436 39874 20500
rect 40401 20498 40467 20501
rect 40718 20498 40724 20500
rect 40401 20496 40724 20498
rect 40401 20440 40406 20496
rect 40462 20440 40724 20496
rect 40401 20438 40724 20440
rect 40401 20435 40467 20438
rect 40718 20436 40724 20438
rect 40788 20436 40794 20500
rect 41137 20498 41203 20501
rect 48221 20498 48287 20501
rect 41137 20496 48287 20498
rect 41137 20440 41142 20496
rect 41198 20440 48226 20496
rect 48282 20440 48287 20496
rect 41137 20438 48287 20440
rect 41137 20435 41203 20438
rect 48221 20435 48287 20438
rect 40350 20362 40356 20364
rect 36356 20302 40356 20362
rect 40350 20300 40356 20302
rect 40420 20300 40426 20364
rect 41086 20362 41092 20364
rect 40496 20302 41092 20362
rect 35341 20299 35407 20300
rect 38377 20226 38443 20229
rect 34516 20224 38443 20226
rect 34516 20168 38382 20224
rect 38438 20168 38443 20224
rect 34516 20166 38443 20168
rect 27337 20163 27403 20166
rect 29269 20163 29335 20166
rect 38377 20163 38443 20166
rect 38745 20226 38811 20229
rect 39849 20226 39915 20229
rect 38745 20224 39915 20226
rect 38745 20168 38750 20224
rect 38806 20168 39854 20224
rect 39910 20168 39915 20224
rect 38745 20166 39915 20168
rect 38745 20163 38811 20166
rect 39849 20163 39915 20166
rect 40033 20226 40099 20229
rect 40496 20226 40556 20302
rect 41086 20300 41092 20302
rect 41156 20300 41162 20364
rect 41413 20362 41479 20365
rect 44357 20362 44423 20365
rect 41413 20360 44423 20362
rect 41413 20304 41418 20360
rect 41474 20304 44362 20360
rect 44418 20304 44423 20360
rect 41413 20302 44423 20304
rect 41413 20299 41479 20302
rect 44357 20299 44423 20302
rect 41321 20226 41387 20229
rect 42006 20226 42012 20228
rect 40033 20224 40556 20226
rect 40033 20168 40038 20224
rect 40094 20168 40556 20224
rect 40033 20166 40556 20168
rect 40680 20166 40970 20226
rect 40033 20163 40099 20166
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 14549 20090 14615 20093
rect 18781 20090 18847 20093
rect 14549 20088 18847 20090
rect 14549 20032 14554 20088
rect 14610 20032 18786 20088
rect 18842 20032 18847 20088
rect 14549 20030 18847 20032
rect 14549 20027 14615 20030
rect 18781 20027 18847 20030
rect 21449 20090 21515 20093
rect 22553 20090 22619 20093
rect 29269 20092 29335 20093
rect 29269 20090 29316 20092
rect 21449 20088 22619 20090
rect 21449 20032 21454 20088
rect 21510 20032 22558 20088
rect 22614 20032 22619 20088
rect 21449 20030 22619 20032
rect 29224 20088 29316 20090
rect 29224 20032 29274 20088
rect 29224 20030 29316 20032
rect 21449 20027 21515 20030
rect 22553 20027 22619 20030
rect 29269 20028 29316 20030
rect 29380 20028 29386 20092
rect 35157 20090 35223 20093
rect 40680 20090 40740 20166
rect 33366 20088 40740 20090
rect 33366 20032 35162 20088
rect 35218 20032 40740 20088
rect 33366 20030 40740 20032
rect 40910 20090 40970 20166
rect 41321 20224 42012 20226
rect 41321 20168 41326 20224
rect 41382 20168 42012 20224
rect 41321 20166 42012 20168
rect 41321 20163 41387 20166
rect 42006 20164 42012 20166
rect 42076 20164 42082 20228
rect 44214 20164 44220 20228
rect 44284 20226 44290 20228
rect 46013 20226 46079 20229
rect 44284 20224 46079 20226
rect 44284 20168 46018 20224
rect 46074 20168 46079 20224
rect 44284 20166 46079 20168
rect 44284 20164 44290 20166
rect 46013 20163 46079 20166
rect 46422 20164 46428 20228
rect 46492 20226 46498 20228
rect 50200 20226 51000 20256
rect 46492 20166 51000 20226
rect 46492 20164 46498 20166
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 50200 20136 51000 20166
rect 42946 20095 43262 20096
rect 42374 20090 42380 20092
rect 40910 20030 42380 20090
rect 29269 20027 29335 20028
rect 8293 19952 12450 19954
rect 8293 19896 8298 19952
rect 8354 19896 12450 19952
rect 8293 19894 12450 19896
rect 14549 19954 14615 19957
rect 23933 19954 23999 19957
rect 14549 19952 23999 19954
rect 14549 19896 14554 19952
rect 14610 19896 23938 19952
rect 23994 19896 23999 19952
rect 14549 19894 23999 19896
rect 8293 19891 8359 19894
rect 14549 19891 14615 19894
rect 23933 19891 23999 19894
rect 26877 19954 26943 19957
rect 32673 19954 32739 19957
rect 26877 19952 32739 19954
rect 26877 19896 26882 19952
rect 26938 19896 32678 19952
rect 32734 19896 32739 19952
rect 26877 19894 32739 19896
rect 26877 19891 26943 19894
rect 32673 19891 32739 19894
rect 33225 19954 33291 19957
rect 33366 19954 33426 20030
rect 35157 20027 35223 20030
rect 42374 20028 42380 20030
rect 42444 20028 42450 20092
rect 33225 19952 33426 19954
rect 33225 19896 33230 19952
rect 33286 19896 33426 19952
rect 33225 19894 33426 19896
rect 35065 19954 35131 19957
rect 36721 19954 36787 19957
rect 35065 19952 36787 19954
rect 35065 19896 35070 19952
rect 35126 19896 36726 19952
rect 36782 19896 36787 19952
rect 35065 19894 36787 19896
rect 33225 19891 33291 19894
rect 35065 19891 35131 19894
rect 36721 19891 36787 19894
rect 36997 19954 37063 19957
rect 38878 19954 38884 19956
rect 36997 19952 38884 19954
rect 36997 19896 37002 19952
rect 37058 19896 38884 19952
rect 36997 19894 38884 19896
rect 36997 19891 37063 19894
rect 38878 19892 38884 19894
rect 38948 19892 38954 19956
rect 39113 19954 39179 19957
rect 39849 19954 39915 19957
rect 40585 19954 40651 19957
rect 39113 19952 39915 19954
rect 39113 19896 39118 19952
rect 39174 19896 39854 19952
rect 39910 19896 39915 19952
rect 39113 19894 39915 19896
rect 39113 19891 39179 19894
rect 39849 19891 39915 19894
rect 40358 19952 40651 19954
rect 40358 19896 40590 19952
rect 40646 19896 40651 19952
rect 40358 19894 40651 19896
rect 9857 19818 9923 19821
rect 15193 19818 15259 19821
rect 9857 19816 15259 19818
rect 9857 19760 9862 19816
rect 9918 19760 15198 19816
rect 15254 19760 15259 19816
rect 9857 19758 15259 19760
rect 9857 19755 9923 19758
rect 15193 19755 15259 19758
rect 16021 19818 16087 19821
rect 19977 19818 20043 19821
rect 24577 19818 24643 19821
rect 16021 19816 18522 19818
rect 16021 19760 16026 19816
rect 16082 19760 18522 19816
rect 16021 19758 18522 19760
rect 16021 19755 16087 19758
rect 9121 19682 9187 19685
rect 15142 19682 15148 19684
rect 9121 19680 15148 19682
rect 9121 19624 9126 19680
rect 9182 19624 15148 19680
rect 9121 19622 15148 19624
rect 9121 19619 9187 19622
rect 15142 19620 15148 19622
rect 15212 19620 15218 19684
rect 7946 19616 8262 19617
rect 0 19546 800 19576
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 2957 19546 3023 19549
rect 0 19544 3023 19546
rect 0 19488 2962 19544
rect 3018 19488 3023 19544
rect 0 19486 3023 19488
rect 0 19456 800 19486
rect 2957 19483 3023 19486
rect 11094 19484 11100 19548
rect 11164 19546 11170 19548
rect 13905 19546 13971 19549
rect 11164 19544 13971 19546
rect 11164 19488 13910 19544
rect 13966 19488 13971 19544
rect 11164 19486 13971 19488
rect 18462 19546 18522 19758
rect 19977 19816 24643 19818
rect 19977 19760 19982 19816
rect 20038 19760 24582 19816
rect 24638 19760 24643 19816
rect 19977 19758 24643 19760
rect 19977 19755 20043 19758
rect 24577 19755 24643 19758
rect 27613 19818 27679 19821
rect 30465 19818 30531 19821
rect 27613 19816 30531 19818
rect 27613 19760 27618 19816
rect 27674 19760 30470 19816
rect 30526 19760 30531 19816
rect 27613 19758 30531 19760
rect 27613 19755 27679 19758
rect 30465 19755 30531 19758
rect 30649 19818 30715 19821
rect 33593 19818 33659 19821
rect 35985 19818 36051 19821
rect 38469 19818 38535 19821
rect 40358 19818 40418 19894
rect 40585 19891 40651 19894
rect 30649 19816 35818 19818
rect 30649 19760 30654 19816
rect 30710 19760 33598 19816
rect 33654 19760 35818 19816
rect 30649 19758 35818 19760
rect 30649 19755 30715 19758
rect 33593 19755 33659 19758
rect 18597 19682 18663 19685
rect 27337 19682 27403 19685
rect 35617 19682 35683 19685
rect 18597 19680 27403 19682
rect 18597 19624 18602 19680
rect 18658 19624 27342 19680
rect 27398 19624 27403 19680
rect 18597 19622 27403 19624
rect 18597 19619 18663 19622
rect 27337 19619 27403 19622
rect 28398 19680 35683 19682
rect 28398 19624 35622 19680
rect 35678 19624 35683 19680
rect 28398 19622 35683 19624
rect 35758 19682 35818 19758
rect 35985 19816 38394 19818
rect 35985 19760 35990 19816
rect 36046 19760 38394 19816
rect 35985 19758 38394 19760
rect 35985 19755 36051 19758
rect 35893 19682 35959 19685
rect 38334 19682 38394 19758
rect 38469 19816 40418 19818
rect 38469 19760 38474 19816
rect 38530 19760 40418 19816
rect 38469 19758 40418 19760
rect 40493 19818 40559 19821
rect 43437 19818 43503 19821
rect 40493 19816 43503 19818
rect 40493 19760 40498 19816
rect 40554 19760 43442 19816
rect 43498 19760 43503 19816
rect 40493 19758 43503 19760
rect 38469 19755 38535 19758
rect 40493 19755 40559 19758
rect 43437 19755 43503 19758
rect 46105 19818 46171 19821
rect 49417 19818 49483 19821
rect 50200 19818 51000 19848
rect 46105 19816 49250 19818
rect 46105 19760 46110 19816
rect 46166 19760 49250 19816
rect 46105 19758 49250 19760
rect 46105 19755 46171 19758
rect 46933 19682 46999 19685
rect 35758 19680 37842 19682
rect 35758 19624 35898 19680
rect 35954 19624 37842 19680
rect 35758 19622 37842 19624
rect 38334 19680 46999 19682
rect 38334 19624 46938 19680
rect 46994 19624 46999 19680
rect 38334 19622 46999 19624
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 19977 19546 20043 19549
rect 23473 19546 23539 19549
rect 18462 19544 23539 19546
rect 18462 19488 19982 19544
rect 20038 19488 23478 19544
rect 23534 19488 23539 19544
rect 18462 19486 23539 19488
rect 11164 19484 11170 19486
rect 13905 19483 13971 19486
rect 19977 19483 20043 19486
rect 23473 19483 23539 19486
rect 5349 19410 5415 19413
rect 8201 19410 8267 19413
rect 16757 19410 16823 19413
rect 19241 19410 19307 19413
rect 5349 19408 19307 19410
rect 5349 19352 5354 19408
rect 5410 19352 8206 19408
rect 8262 19352 16762 19408
rect 16818 19352 19246 19408
rect 19302 19352 19307 19408
rect 5349 19350 19307 19352
rect 5349 19347 5415 19350
rect 8201 19347 8267 19350
rect 16757 19347 16823 19350
rect 19241 19347 19307 19350
rect 22318 19348 22324 19412
rect 22388 19410 22394 19412
rect 23473 19410 23539 19413
rect 22388 19408 23539 19410
rect 22388 19352 23478 19408
rect 23534 19352 23539 19408
rect 22388 19350 23539 19352
rect 22388 19348 22394 19350
rect 23473 19347 23539 19350
rect 27705 19410 27771 19413
rect 28257 19410 28323 19413
rect 28398 19410 28458 19622
rect 35617 19619 35683 19622
rect 35893 19619 35959 19622
rect 30557 19546 30623 19549
rect 37181 19546 37247 19549
rect 30557 19544 37247 19546
rect 30557 19488 30562 19544
rect 30618 19488 37186 19544
rect 37242 19488 37247 19544
rect 30557 19486 37247 19488
rect 30557 19483 30623 19486
rect 37181 19483 37247 19486
rect 27705 19408 28458 19410
rect 27705 19352 27710 19408
rect 27766 19352 28262 19408
rect 28318 19352 28458 19408
rect 27705 19350 28458 19352
rect 29269 19410 29335 19413
rect 29494 19410 29500 19412
rect 29269 19408 29500 19410
rect 29269 19352 29274 19408
rect 29330 19352 29500 19408
rect 29269 19350 29500 19352
rect 27705 19347 27771 19350
rect 28257 19347 28323 19350
rect 29269 19347 29335 19350
rect 29494 19348 29500 19350
rect 29564 19348 29570 19412
rect 31937 19410 32003 19413
rect 32949 19410 33015 19413
rect 37641 19410 37707 19413
rect 31937 19408 37707 19410
rect 31937 19352 31942 19408
rect 31998 19352 32954 19408
rect 33010 19352 37646 19408
rect 37702 19352 37707 19408
rect 31937 19350 37707 19352
rect 37782 19410 37842 19622
rect 46933 19619 46999 19622
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 38878 19484 38884 19548
rect 38948 19546 38954 19548
rect 44357 19546 44423 19549
rect 38948 19544 44423 19546
rect 38948 19488 44362 19544
rect 44418 19488 44423 19544
rect 38948 19486 44423 19488
rect 49190 19546 49250 19758
rect 49417 19816 51000 19818
rect 49417 19760 49422 19816
rect 49478 19760 51000 19816
rect 49417 19758 51000 19760
rect 49417 19755 49483 19758
rect 50200 19728 51000 19758
rect 49190 19486 49434 19546
rect 38948 19484 38954 19486
rect 44357 19483 44423 19486
rect 38193 19410 38259 19413
rect 37782 19408 38259 19410
rect 37782 19352 38198 19408
rect 38254 19352 38259 19408
rect 37782 19350 38259 19352
rect 31937 19347 32003 19350
rect 32949 19347 33015 19350
rect 37641 19347 37707 19350
rect 38193 19347 38259 19350
rect 38377 19410 38443 19413
rect 41137 19410 41203 19413
rect 43713 19410 43779 19413
rect 38377 19408 43779 19410
rect 38377 19352 38382 19408
rect 38438 19352 41142 19408
rect 41198 19352 43718 19408
rect 43774 19352 43779 19408
rect 38377 19350 43779 19352
rect 38377 19347 38443 19350
rect 41137 19347 41203 19350
rect 43713 19347 43779 19350
rect 45277 19410 45343 19413
rect 45553 19410 45619 19413
rect 45277 19408 45619 19410
rect 45277 19352 45282 19408
rect 45338 19352 45558 19408
rect 45614 19352 45619 19408
rect 45277 19350 45619 19352
rect 45277 19347 45343 19350
rect 45553 19347 45619 19350
rect 49141 19412 49207 19413
rect 49141 19408 49188 19412
rect 49252 19410 49258 19412
rect 49374 19410 49434 19486
rect 50200 19410 51000 19440
rect 49141 19352 49146 19408
rect 49141 19348 49188 19352
rect 49252 19350 49298 19410
rect 49374 19350 51000 19410
rect 49252 19348 49258 19350
rect 49141 19347 49207 19348
rect 50200 19320 51000 19350
rect 9029 19274 9095 19277
rect 16021 19274 16087 19277
rect 9029 19272 16087 19274
rect 9029 19216 9034 19272
rect 9090 19216 16026 19272
rect 16082 19216 16087 19272
rect 9029 19214 16087 19216
rect 9029 19211 9095 19214
rect 16021 19211 16087 19214
rect 17769 19274 17835 19277
rect 20161 19274 20227 19277
rect 17769 19272 20227 19274
rect 17769 19216 17774 19272
rect 17830 19216 20166 19272
rect 20222 19216 20227 19272
rect 17769 19214 20227 19216
rect 17769 19211 17835 19214
rect 20161 19211 20227 19214
rect 21725 19274 21791 19277
rect 25589 19274 25655 19277
rect 28717 19274 28783 19277
rect 21725 19272 28783 19274
rect 21725 19216 21730 19272
rect 21786 19216 25594 19272
rect 25650 19216 28722 19272
rect 28778 19216 28783 19272
rect 21725 19214 28783 19216
rect 21725 19211 21791 19214
rect 25589 19211 25655 19214
rect 28717 19211 28783 19214
rect 29269 19274 29335 19277
rect 31385 19274 31451 19277
rect 33593 19274 33659 19277
rect 33777 19274 33843 19277
rect 29269 19272 30436 19274
rect 29269 19216 29274 19272
rect 29330 19216 30436 19272
rect 29269 19214 30436 19216
rect 29269 19211 29335 19214
rect 0 19138 800 19168
rect 2773 19138 2839 19141
rect 0 19136 2839 19138
rect 0 19080 2778 19136
rect 2834 19080 2839 19136
rect 0 19078 2839 19080
rect 0 19048 800 19078
rect 2773 19075 2839 19078
rect 6545 19138 6611 19141
rect 12198 19138 12204 19140
rect 6545 19136 12204 19138
rect 6545 19080 6550 19136
rect 6606 19080 12204 19136
rect 6545 19078 12204 19080
rect 6545 19075 6611 19078
rect 12198 19076 12204 19078
rect 12268 19138 12274 19140
rect 13629 19138 13695 19141
rect 16205 19138 16271 19141
rect 12268 19078 12818 19138
rect 12268 19076 12274 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 5574 18940 5580 19004
rect 5644 19002 5650 19004
rect 11053 19002 11119 19005
rect 5644 19000 11119 19002
rect 5644 18944 11058 19000
rect 11114 18944 11119 19000
rect 5644 18942 11119 18944
rect 5644 18940 5650 18942
rect 11053 18939 11119 18942
rect 7005 18866 7071 18869
rect 9673 18866 9739 18869
rect 12525 18866 12591 18869
rect 7005 18864 8586 18866
rect 7005 18808 7010 18864
rect 7066 18808 8586 18864
rect 7005 18806 8586 18808
rect 7005 18803 7071 18806
rect 0 18730 800 18760
rect 2865 18730 2931 18733
rect 0 18728 2931 18730
rect 0 18672 2870 18728
rect 2926 18672 2931 18728
rect 0 18670 2931 18672
rect 0 18640 800 18670
rect 2865 18667 2931 18670
rect 7465 18730 7531 18733
rect 8334 18730 8340 18732
rect 7465 18728 8340 18730
rect 7465 18672 7470 18728
rect 7526 18672 8340 18728
rect 7465 18670 8340 18672
rect 7465 18667 7531 18670
rect 8334 18668 8340 18670
rect 8404 18668 8410 18732
rect 8526 18730 8586 18806
rect 9673 18864 12591 18866
rect 9673 18808 9678 18864
rect 9734 18808 12530 18864
rect 12586 18808 12591 18864
rect 9673 18806 12591 18808
rect 12758 18866 12818 19078
rect 13629 19136 16271 19138
rect 13629 19080 13634 19136
rect 13690 19080 16210 19136
rect 16266 19080 16271 19136
rect 13629 19078 16271 19080
rect 13629 19075 13695 19078
rect 16205 19075 16271 19078
rect 17125 19138 17191 19141
rect 18597 19138 18663 19141
rect 17125 19136 18663 19138
rect 17125 19080 17130 19136
rect 17186 19080 18602 19136
rect 18658 19080 18663 19136
rect 17125 19078 18663 19080
rect 17125 19075 17191 19078
rect 18597 19075 18663 19078
rect 19926 19076 19932 19140
rect 19996 19138 20002 19140
rect 20161 19138 20227 19141
rect 19996 19136 20227 19138
rect 19996 19080 20166 19136
rect 20222 19080 20227 19136
rect 19996 19078 20227 19080
rect 30376 19138 30436 19214
rect 31385 19272 33426 19274
rect 31385 19216 31390 19272
rect 31446 19216 33426 19272
rect 31385 19214 33426 19216
rect 31385 19211 31451 19214
rect 31661 19138 31727 19141
rect 30376 19136 31727 19138
rect 30376 19080 31666 19136
rect 31722 19080 31727 19136
rect 30376 19078 31727 19080
rect 33366 19138 33426 19214
rect 33593 19272 33843 19274
rect 33593 19216 33598 19272
rect 33654 19216 33782 19272
rect 33838 19216 33843 19272
rect 33593 19214 33843 19216
rect 33593 19211 33659 19214
rect 33777 19211 33843 19214
rect 34329 19274 34395 19277
rect 34462 19274 34468 19276
rect 34329 19272 34468 19274
rect 34329 19216 34334 19272
rect 34390 19216 34468 19272
rect 34329 19214 34468 19216
rect 34329 19211 34395 19214
rect 34462 19212 34468 19214
rect 34532 19212 34538 19276
rect 34697 19274 34763 19277
rect 39573 19274 39639 19277
rect 34697 19272 39639 19274
rect 34697 19216 34702 19272
rect 34758 19216 39578 19272
rect 39634 19216 39639 19272
rect 34697 19214 39639 19216
rect 34697 19211 34763 19214
rect 39573 19211 39639 19214
rect 40033 19274 40099 19277
rect 41638 19274 41644 19276
rect 40033 19272 41644 19274
rect 40033 19216 40038 19272
rect 40094 19216 41644 19272
rect 40033 19214 41644 19216
rect 40033 19211 40099 19214
rect 41638 19212 41644 19214
rect 41708 19274 41714 19276
rect 41965 19274 42031 19277
rect 41708 19272 42031 19274
rect 41708 19216 41970 19272
rect 42026 19216 42031 19272
rect 41708 19214 42031 19216
rect 41708 19212 41714 19214
rect 41965 19211 42031 19214
rect 33542 19138 33548 19140
rect 33366 19078 33548 19138
rect 19996 19076 20002 19078
rect 20161 19075 20227 19078
rect 31661 19075 31727 19078
rect 33542 19076 33548 19078
rect 33612 19138 33618 19140
rect 34789 19138 34855 19141
rect 33612 19136 34855 19138
rect 33612 19080 34794 19136
rect 34850 19080 34855 19136
rect 33612 19078 34855 19080
rect 33612 19076 33618 19078
rect 34789 19075 34855 19078
rect 36445 19138 36511 19141
rect 41597 19138 41663 19141
rect 41873 19138 41939 19141
rect 36445 19136 41939 19138
rect 36445 19080 36450 19136
rect 36506 19080 41602 19136
rect 41658 19080 41878 19136
rect 41934 19080 41939 19136
rect 36445 19078 41939 19080
rect 36445 19075 36511 19078
rect 41597 19075 41663 19078
rect 41873 19075 41939 19078
rect 42241 19138 42307 19141
rect 44725 19140 44791 19141
rect 42374 19138 42380 19140
rect 42241 19136 42380 19138
rect 42241 19080 42246 19136
rect 42302 19080 42380 19136
rect 42241 19078 42380 19080
rect 42241 19075 42307 19078
rect 42374 19076 42380 19078
rect 42444 19076 42450 19140
rect 44725 19138 44772 19140
rect 44680 19136 44772 19138
rect 44680 19080 44730 19136
rect 44680 19078 44772 19080
rect 44725 19076 44772 19078
rect 44836 19076 44842 19140
rect 47158 19076 47164 19140
rect 47228 19138 47234 19140
rect 48221 19138 48287 19141
rect 48814 19138 48820 19140
rect 47228 19136 48820 19138
rect 47228 19080 48226 19136
rect 48282 19080 48820 19136
rect 47228 19078 48820 19080
rect 47228 19076 47234 19078
rect 44725 19075 44791 19076
rect 48221 19075 48287 19078
rect 48814 19076 48820 19078
rect 48884 19076 48890 19140
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 15101 19002 15167 19005
rect 22185 19002 22251 19005
rect 24853 19004 24919 19005
rect 24853 19002 24900 19004
rect 15101 19000 22251 19002
rect 15101 18944 15106 19000
rect 15162 18944 22190 19000
rect 22246 18944 22251 19000
rect 15101 18942 22251 18944
rect 24808 19000 24900 19002
rect 24808 18944 24858 19000
rect 24808 18942 24900 18944
rect 15101 18939 15167 18942
rect 22185 18939 22251 18942
rect 24853 18940 24900 18942
rect 24964 18940 24970 19004
rect 27654 18940 27660 19004
rect 27724 19002 27730 19004
rect 28257 19002 28323 19005
rect 27724 19000 28323 19002
rect 27724 18944 28262 19000
rect 28318 18944 28323 19000
rect 27724 18942 28323 18944
rect 27724 18940 27730 18942
rect 24853 18939 24919 18940
rect 28257 18939 28323 18942
rect 29269 19002 29335 19005
rect 29821 19002 29887 19005
rect 29269 19000 29887 19002
rect 29269 18944 29274 19000
rect 29330 18944 29826 19000
rect 29882 18944 29887 19000
rect 29269 18942 29887 18944
rect 29269 18939 29335 18942
rect 29821 18939 29887 18942
rect 31753 19002 31819 19005
rect 31886 19002 31892 19004
rect 31753 19000 31892 19002
rect 31753 18944 31758 19000
rect 31814 18944 31892 19000
rect 31753 18942 31892 18944
rect 31753 18939 31819 18942
rect 31886 18940 31892 18942
rect 31956 18940 31962 19004
rect 35249 19002 35315 19005
rect 42057 19002 42123 19005
rect 35249 19000 42123 19002
rect 35249 18944 35254 19000
rect 35310 18944 42062 19000
rect 42118 18944 42123 19000
rect 35249 18942 42123 18944
rect 35249 18939 35315 18942
rect 42057 18939 42123 18942
rect 49141 19002 49207 19005
rect 50200 19002 51000 19032
rect 49141 19000 51000 19002
rect 49141 18944 49146 19000
rect 49202 18944 51000 19000
rect 49141 18942 51000 18944
rect 49141 18939 49207 18942
rect 50200 18912 51000 18942
rect 15009 18866 15075 18869
rect 20253 18866 20319 18869
rect 12758 18864 15075 18866
rect 12758 18808 15014 18864
rect 15070 18808 15075 18864
rect 12758 18806 15075 18808
rect 9673 18803 9739 18806
rect 12525 18803 12591 18806
rect 15009 18803 15075 18806
rect 15886 18864 20319 18866
rect 15886 18808 20258 18864
rect 20314 18808 20319 18864
rect 15886 18806 20319 18808
rect 15886 18730 15946 18806
rect 20253 18803 20319 18806
rect 27102 18804 27108 18868
rect 27172 18866 27178 18868
rect 27797 18866 27863 18869
rect 27172 18864 27863 18866
rect 27172 18808 27802 18864
rect 27858 18808 27863 18864
rect 27172 18806 27863 18808
rect 27172 18804 27178 18806
rect 27797 18803 27863 18806
rect 29821 18866 29887 18869
rect 31845 18866 31911 18869
rect 29821 18864 31911 18866
rect 29821 18808 29826 18864
rect 29882 18808 31850 18864
rect 31906 18808 31911 18864
rect 29821 18806 31911 18808
rect 29821 18803 29887 18806
rect 31845 18803 31911 18806
rect 32857 18866 32923 18869
rect 35433 18866 35499 18869
rect 42517 18866 42583 18869
rect 44265 18868 44331 18869
rect 44214 18866 44220 18868
rect 32857 18864 42583 18866
rect 32857 18808 32862 18864
rect 32918 18808 35438 18864
rect 35494 18808 42522 18864
rect 42578 18808 42583 18864
rect 32857 18806 42583 18808
rect 44174 18806 44220 18866
rect 44284 18864 44331 18868
rect 46933 18868 46999 18869
rect 46933 18866 46980 18868
rect 44326 18808 44331 18864
rect 32857 18803 32923 18806
rect 35433 18803 35499 18806
rect 42517 18803 42583 18806
rect 44214 18804 44220 18806
rect 44284 18804 44331 18808
rect 46892 18864 46980 18866
rect 47044 18866 47050 18868
rect 49918 18866 49924 18868
rect 46892 18808 46938 18864
rect 46892 18806 46980 18808
rect 44265 18803 44331 18804
rect 46933 18804 46980 18806
rect 47044 18806 49924 18866
rect 47044 18804 47050 18806
rect 49918 18804 49924 18806
rect 49988 18804 49994 18868
rect 46933 18803 46999 18804
rect 8526 18670 15946 18730
rect 16021 18730 16087 18733
rect 26509 18730 26575 18733
rect 16021 18728 26575 18730
rect 16021 18672 16026 18728
rect 16082 18672 26514 18728
rect 26570 18672 26575 18728
rect 16021 18670 26575 18672
rect 16021 18667 16087 18670
rect 26509 18667 26575 18670
rect 27981 18730 28047 18733
rect 33593 18730 33659 18733
rect 27981 18728 33659 18730
rect 27981 18672 27986 18728
rect 28042 18672 33598 18728
rect 33654 18672 33659 18728
rect 27981 18670 33659 18672
rect 27981 18667 28047 18670
rect 33593 18667 33659 18670
rect 34329 18730 34395 18733
rect 34697 18730 34763 18733
rect 34329 18728 34763 18730
rect 34329 18672 34334 18728
rect 34390 18672 34702 18728
rect 34758 18672 34763 18728
rect 34329 18670 34763 18672
rect 34329 18667 34395 18670
rect 34697 18667 34763 18670
rect 36721 18730 36787 18733
rect 36854 18730 36860 18732
rect 36721 18728 36860 18730
rect 36721 18672 36726 18728
rect 36782 18672 36860 18728
rect 36721 18670 36860 18672
rect 36721 18667 36787 18670
rect 36854 18668 36860 18670
rect 36924 18668 36930 18732
rect 37273 18730 37339 18733
rect 42333 18730 42399 18733
rect 37273 18728 42399 18730
rect 37273 18672 37278 18728
rect 37334 18672 42338 18728
rect 42394 18672 42399 18728
rect 37273 18670 42399 18672
rect 37273 18667 37339 18670
rect 42333 18667 42399 18670
rect 47393 18730 47459 18733
rect 47945 18730 48011 18733
rect 49785 18730 49851 18733
rect 47393 18728 48011 18730
rect 47393 18672 47398 18728
rect 47454 18672 47950 18728
rect 48006 18672 48011 18728
rect 47393 18670 48011 18672
rect 47393 18667 47459 18670
rect 47945 18667 48011 18670
rect 49558 18728 49851 18730
rect 49558 18672 49790 18728
rect 49846 18672 49851 18728
rect 49558 18670 49851 18672
rect 3417 18596 3483 18597
rect 3366 18532 3372 18596
rect 3436 18594 3483 18596
rect 10501 18594 10567 18597
rect 12065 18594 12131 18597
rect 3436 18592 3528 18594
rect 3478 18536 3528 18592
rect 3436 18534 3528 18536
rect 10501 18592 12131 18594
rect 10501 18536 10506 18592
rect 10562 18536 12070 18592
rect 12126 18536 12131 18592
rect 10501 18534 12131 18536
rect 3436 18532 3483 18534
rect 3417 18531 3483 18532
rect 10501 18531 10567 18534
rect 12065 18531 12131 18534
rect 12525 18594 12591 18597
rect 17769 18594 17835 18597
rect 12525 18592 17835 18594
rect 12525 18536 12530 18592
rect 12586 18536 17774 18592
rect 17830 18536 17835 18592
rect 12525 18534 17835 18536
rect 12525 18531 12591 18534
rect 17769 18531 17835 18534
rect 20253 18594 20319 18597
rect 20621 18594 20687 18597
rect 20253 18592 20687 18594
rect 20253 18536 20258 18592
rect 20314 18536 20626 18592
rect 20682 18536 20687 18592
rect 20253 18534 20687 18536
rect 20253 18531 20319 18534
rect 20621 18531 20687 18534
rect 33041 18594 33107 18597
rect 36077 18594 36143 18597
rect 33041 18592 36143 18594
rect 33041 18536 33046 18592
rect 33102 18536 36082 18592
rect 36138 18536 36143 18592
rect 33041 18534 36143 18536
rect 33041 18531 33107 18534
rect 36077 18531 36143 18534
rect 38745 18594 38811 18597
rect 38878 18594 38884 18596
rect 38745 18592 38884 18594
rect 38745 18536 38750 18592
rect 38806 18536 38884 18592
rect 38745 18534 38884 18536
rect 38745 18531 38811 18534
rect 38878 18532 38884 18534
rect 38948 18532 38954 18596
rect 39113 18594 39179 18597
rect 42241 18594 42307 18597
rect 43897 18594 43963 18597
rect 39113 18592 43963 18594
rect 39113 18536 39118 18592
rect 39174 18536 42246 18592
rect 42302 18536 43902 18592
rect 43958 18536 43963 18592
rect 39113 18534 43963 18536
rect 39113 18531 39179 18534
rect 42241 18531 42307 18534
rect 43897 18531 43963 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 47946 18463 48262 18464
rect 6177 18458 6243 18461
rect 6310 18458 6316 18460
rect 6177 18456 6316 18458
rect 6177 18400 6182 18456
rect 6238 18400 6316 18456
rect 6177 18398 6316 18400
rect 6177 18395 6243 18398
rect 6310 18396 6316 18398
rect 6380 18396 6386 18460
rect 12801 18458 12867 18461
rect 15653 18458 15719 18461
rect 16297 18458 16363 18461
rect 26877 18458 26943 18461
rect 12801 18456 16363 18458
rect 12801 18400 12806 18456
rect 12862 18400 15658 18456
rect 15714 18400 16302 18456
rect 16358 18400 16363 18456
rect 12801 18398 16363 18400
rect 12801 18395 12867 18398
rect 15653 18395 15719 18398
rect 16297 18395 16363 18398
rect 18462 18456 26943 18458
rect 18462 18400 26882 18456
rect 26938 18400 26943 18456
rect 18462 18398 26943 18400
rect 0 18322 800 18352
rect 2037 18322 2103 18325
rect 0 18320 2103 18322
rect 0 18264 2042 18320
rect 2098 18264 2103 18320
rect 0 18262 2103 18264
rect 0 18232 800 18262
rect 2037 18259 2103 18262
rect 5809 18322 5875 18325
rect 11789 18322 11855 18325
rect 13629 18322 13695 18325
rect 5809 18320 11855 18322
rect 5809 18264 5814 18320
rect 5870 18264 11794 18320
rect 11850 18264 11855 18320
rect 5809 18262 11855 18264
rect 5809 18259 5875 18262
rect 11789 18259 11855 18262
rect 12390 18320 13695 18322
rect 12390 18264 13634 18320
rect 13690 18264 13695 18320
rect 12390 18262 13695 18264
rect 3601 18188 3667 18189
rect 3550 18124 3556 18188
rect 3620 18186 3667 18188
rect 6177 18186 6243 18189
rect 12390 18186 12450 18262
rect 13629 18259 13695 18262
rect 17953 18322 18019 18325
rect 18462 18322 18522 18398
rect 26877 18395 26943 18398
rect 27061 18458 27127 18461
rect 27337 18458 27403 18461
rect 27061 18456 27403 18458
rect 27061 18400 27066 18456
rect 27122 18400 27342 18456
rect 27398 18400 27403 18456
rect 27061 18398 27403 18400
rect 27061 18395 27127 18398
rect 27337 18395 27403 18398
rect 30465 18458 30531 18461
rect 36445 18458 36511 18461
rect 30465 18456 36511 18458
rect 30465 18400 30470 18456
rect 30526 18400 36450 18456
rect 36506 18400 36511 18456
rect 30465 18398 36511 18400
rect 30465 18395 30531 18398
rect 36445 18395 36511 18398
rect 36813 18458 36879 18461
rect 37038 18458 37044 18460
rect 36813 18456 37044 18458
rect 36813 18400 36818 18456
rect 36874 18400 37044 18456
rect 36813 18398 37044 18400
rect 36813 18395 36879 18398
rect 37038 18396 37044 18398
rect 37108 18396 37114 18460
rect 40125 18458 40191 18461
rect 41965 18458 42031 18461
rect 40125 18456 42031 18458
rect 40125 18400 40130 18456
rect 40186 18400 41970 18456
rect 42026 18400 42031 18456
rect 40125 18398 42031 18400
rect 40125 18395 40191 18398
rect 41965 18395 42031 18398
rect 42149 18458 42215 18461
rect 45185 18458 45251 18461
rect 42149 18456 45251 18458
rect 42149 18400 42154 18456
rect 42210 18400 45190 18456
rect 45246 18400 45251 18456
rect 42149 18398 45251 18400
rect 42149 18395 42215 18398
rect 45185 18395 45251 18398
rect 17953 18320 18522 18322
rect 17953 18264 17958 18320
rect 18014 18264 18522 18320
rect 17953 18262 18522 18264
rect 19241 18322 19307 18325
rect 33041 18322 33107 18325
rect 19241 18320 33107 18322
rect 19241 18264 19246 18320
rect 19302 18264 33046 18320
rect 33102 18264 33107 18320
rect 19241 18262 33107 18264
rect 17953 18259 18019 18262
rect 19241 18259 19307 18262
rect 33041 18259 33107 18262
rect 34697 18322 34763 18325
rect 44357 18322 44423 18325
rect 34697 18320 44423 18322
rect 34697 18264 34702 18320
rect 34758 18264 44362 18320
rect 44418 18264 44423 18320
rect 34697 18262 44423 18264
rect 34697 18259 34763 18262
rect 44357 18259 44423 18262
rect 49233 18322 49299 18325
rect 49558 18322 49618 18670
rect 49785 18667 49851 18670
rect 49785 18594 49851 18597
rect 50200 18594 51000 18624
rect 49785 18592 51000 18594
rect 49785 18536 49790 18592
rect 49846 18536 51000 18592
rect 49785 18534 51000 18536
rect 49785 18531 49851 18534
rect 50200 18504 51000 18534
rect 49233 18320 49618 18322
rect 49233 18264 49238 18320
rect 49294 18264 49618 18320
rect 49233 18262 49618 18264
rect 49233 18259 49299 18262
rect 3620 18184 3712 18186
rect 3662 18128 3712 18184
rect 3620 18126 3712 18128
rect 6177 18184 12450 18186
rect 6177 18128 6182 18184
rect 6238 18128 12450 18184
rect 6177 18126 12450 18128
rect 12525 18186 12591 18189
rect 17309 18186 17375 18189
rect 27337 18186 27403 18189
rect 12525 18184 27403 18186
rect 12525 18128 12530 18184
rect 12586 18128 17314 18184
rect 17370 18128 27342 18184
rect 27398 18128 27403 18184
rect 12525 18126 27403 18128
rect 3620 18124 3667 18126
rect 3601 18123 3667 18124
rect 6177 18123 6243 18126
rect 12525 18123 12591 18126
rect 17309 18123 17375 18126
rect 27337 18123 27403 18126
rect 33225 18186 33291 18189
rect 35801 18186 35867 18189
rect 33225 18184 35867 18186
rect 33225 18128 33230 18184
rect 33286 18128 35806 18184
rect 35862 18128 35867 18184
rect 33225 18126 35867 18128
rect 33225 18123 33291 18126
rect 35801 18123 35867 18126
rect 36261 18186 36327 18189
rect 39481 18186 39547 18189
rect 36261 18184 39547 18186
rect 36261 18128 36266 18184
rect 36322 18128 39486 18184
rect 39542 18128 39547 18184
rect 36261 18126 39547 18128
rect 36261 18123 36327 18126
rect 39481 18123 39547 18126
rect 39849 18186 39915 18189
rect 40309 18186 40375 18189
rect 39849 18184 40375 18186
rect 39849 18128 39854 18184
rect 39910 18128 40314 18184
rect 40370 18128 40375 18184
rect 39849 18126 40375 18128
rect 39849 18123 39915 18126
rect 40309 18123 40375 18126
rect 40493 18186 40559 18189
rect 41505 18186 41571 18189
rect 40493 18184 41571 18186
rect 40493 18128 40498 18184
rect 40554 18128 41510 18184
rect 41566 18128 41571 18184
rect 40493 18126 41571 18128
rect 40493 18123 40559 18126
rect 41505 18123 41571 18126
rect 42149 18186 42215 18189
rect 43805 18186 43871 18189
rect 42149 18184 43871 18186
rect 42149 18128 42154 18184
rect 42210 18128 43810 18184
rect 43866 18128 43871 18184
rect 42149 18126 43871 18128
rect 42149 18123 42215 18126
rect 43805 18123 43871 18126
rect 47853 18186 47919 18189
rect 50200 18186 51000 18216
rect 47853 18184 51000 18186
rect 47853 18128 47858 18184
rect 47914 18128 51000 18184
rect 47853 18126 51000 18128
rect 47853 18123 47919 18126
rect 50200 18096 51000 18126
rect 14825 18050 14891 18053
rect 14958 18050 14964 18052
rect 14825 18048 14964 18050
rect 14825 17992 14830 18048
rect 14886 17992 14964 18048
rect 14825 17990 14964 17992
rect 14825 17987 14891 17990
rect 14958 17988 14964 17990
rect 15028 17988 15034 18052
rect 15326 17988 15332 18052
rect 15396 18050 15402 18052
rect 15561 18050 15627 18053
rect 15396 18048 15627 18050
rect 15396 17992 15566 18048
rect 15622 17992 15627 18048
rect 15396 17990 15627 17992
rect 15396 17988 15402 17990
rect 15561 17987 15627 17990
rect 17769 18050 17835 18053
rect 19241 18050 19307 18053
rect 17769 18048 19307 18050
rect 17769 17992 17774 18048
rect 17830 17992 19246 18048
rect 19302 17992 19307 18048
rect 17769 17990 19307 17992
rect 17769 17987 17835 17990
rect 19241 17987 19307 17990
rect 19517 18052 19583 18053
rect 24945 18052 25011 18053
rect 26601 18052 26667 18053
rect 19517 18048 19564 18052
rect 19628 18050 19634 18052
rect 19517 17992 19522 18048
rect 19517 17988 19564 17992
rect 19628 17990 19674 18050
rect 19628 17988 19634 17990
rect 24894 17988 24900 18052
rect 24964 18050 25011 18052
rect 24964 18048 25056 18050
rect 25006 17992 25056 18048
rect 24964 17990 25056 17992
rect 24964 17988 25011 17990
rect 26550 17988 26556 18052
rect 26620 18050 26667 18052
rect 28441 18050 28507 18053
rect 26620 18048 26712 18050
rect 26662 17992 26712 18048
rect 26620 17990 26712 17992
rect 27340 18048 28507 18050
rect 27340 17992 28446 18048
rect 28502 17992 28507 18048
rect 27340 17990 28507 17992
rect 26620 17988 26667 17990
rect 19517 17987 19583 17988
rect 24945 17987 25011 17988
rect 26601 17987 26667 17988
rect 2946 17984 3262 17985
rect 0 17914 800 17944
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 2773 17914 2839 17917
rect 0 17912 2839 17914
rect 0 17856 2778 17912
rect 2834 17856 2839 17912
rect 0 17854 2839 17856
rect 0 17824 800 17854
rect 2773 17851 2839 17854
rect 4705 17914 4771 17917
rect 9581 17914 9647 17917
rect 4705 17912 9647 17914
rect 4705 17856 4710 17912
rect 4766 17856 9586 17912
rect 9642 17856 9647 17912
rect 4705 17854 9647 17856
rect 4705 17851 4771 17854
rect 9581 17851 9647 17854
rect 9990 17852 9996 17916
rect 10060 17914 10066 17916
rect 12433 17914 12499 17917
rect 10060 17912 12499 17914
rect 10060 17856 12438 17912
rect 12494 17856 12499 17912
rect 10060 17854 12499 17856
rect 10060 17852 10066 17854
rect 12433 17851 12499 17854
rect 13537 17914 13603 17917
rect 18505 17914 18571 17917
rect 13537 17912 18571 17914
rect 13537 17856 13542 17912
rect 13598 17856 18510 17912
rect 18566 17856 18571 17912
rect 13537 17854 18571 17856
rect 13537 17851 13603 17854
rect 18505 17851 18571 17854
rect 18781 17914 18847 17917
rect 27061 17914 27127 17917
rect 27340 17914 27400 17990
rect 28441 17987 28507 17990
rect 35525 18050 35591 18053
rect 37641 18050 37707 18053
rect 38326 18050 38332 18052
rect 35525 18048 37290 18050
rect 35525 17992 35530 18048
rect 35586 17992 37290 18048
rect 35525 17990 37290 17992
rect 35525 17987 35591 17990
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 18781 17912 22110 17914
rect 18781 17856 18786 17912
rect 18842 17856 22110 17912
rect 18781 17854 22110 17856
rect 18781 17851 18847 17854
rect 10869 17778 10935 17781
rect 11513 17778 11579 17781
rect 10869 17776 11579 17778
rect 10869 17720 10874 17776
rect 10930 17720 11518 17776
rect 11574 17720 11579 17776
rect 10869 17718 11579 17720
rect 10869 17715 10935 17718
rect 11513 17715 11579 17718
rect 11789 17778 11855 17781
rect 13670 17778 13676 17780
rect 11789 17776 13676 17778
rect 11789 17720 11794 17776
rect 11850 17720 13676 17776
rect 11789 17718 13676 17720
rect 11789 17715 11855 17718
rect 13670 17716 13676 17718
rect 13740 17716 13746 17780
rect 17217 17778 17283 17781
rect 19425 17778 19491 17781
rect 21265 17778 21331 17781
rect 17217 17776 18890 17778
rect 17217 17720 17222 17776
rect 17278 17720 18890 17776
rect 17217 17718 18890 17720
rect 17217 17715 17283 17718
rect 3417 17642 3483 17645
rect 9070 17642 9076 17644
rect 3417 17640 9076 17642
rect 3417 17584 3422 17640
rect 3478 17584 9076 17640
rect 3417 17582 9076 17584
rect 3417 17579 3483 17582
rect 9070 17580 9076 17582
rect 9140 17642 9146 17644
rect 9213 17642 9279 17645
rect 9140 17640 9279 17642
rect 9140 17584 9218 17640
rect 9274 17584 9279 17640
rect 9140 17582 9279 17584
rect 9140 17580 9146 17582
rect 9213 17579 9279 17582
rect 12341 17642 12407 17645
rect 17953 17642 18019 17645
rect 12341 17640 18019 17642
rect 12341 17584 12346 17640
rect 12402 17584 17958 17640
rect 18014 17584 18019 17640
rect 12341 17582 18019 17584
rect 12341 17579 12407 17582
rect 17953 17579 18019 17582
rect 18321 17642 18387 17645
rect 18454 17642 18460 17644
rect 18321 17640 18460 17642
rect 18321 17584 18326 17640
rect 18382 17584 18460 17640
rect 18321 17582 18460 17584
rect 18321 17579 18387 17582
rect 18454 17580 18460 17582
rect 18524 17580 18530 17644
rect 18830 17642 18890 17718
rect 19425 17776 21331 17778
rect 19425 17720 19430 17776
rect 19486 17720 21270 17776
rect 21326 17720 21331 17776
rect 19425 17718 21331 17720
rect 22050 17778 22110 17854
rect 27061 17912 27400 17914
rect 27061 17856 27066 17912
rect 27122 17856 27400 17912
rect 27061 17854 27400 17856
rect 27061 17851 27127 17854
rect 27470 17852 27476 17916
rect 27540 17914 27546 17916
rect 32213 17914 32279 17917
rect 32622 17914 32628 17916
rect 27540 17854 31770 17914
rect 27540 17852 27546 17854
rect 27613 17778 27679 17781
rect 22050 17776 27679 17778
rect 22050 17720 27618 17776
rect 27674 17720 27679 17776
rect 22050 17718 27679 17720
rect 31710 17778 31770 17854
rect 32213 17912 32628 17914
rect 32213 17856 32218 17912
rect 32274 17856 32628 17912
rect 32213 17854 32628 17856
rect 32213 17851 32279 17854
rect 32622 17852 32628 17854
rect 32692 17852 32698 17916
rect 34329 17914 34395 17917
rect 36445 17914 36511 17917
rect 34329 17912 36511 17914
rect 34329 17856 34334 17912
rect 34390 17856 36450 17912
rect 36506 17856 36511 17912
rect 34329 17854 36511 17856
rect 37230 17914 37290 17990
rect 37641 18048 38332 18050
rect 37641 17992 37646 18048
rect 37702 17992 38332 18048
rect 37641 17990 38332 17992
rect 37641 17987 37707 17990
rect 38326 17988 38332 17990
rect 38396 17988 38402 18052
rect 39798 17988 39804 18052
rect 39868 18050 39874 18052
rect 41229 18050 41295 18053
rect 39868 18048 41295 18050
rect 39868 17992 41234 18048
rect 41290 17992 41295 18048
rect 39868 17990 41295 17992
rect 39868 17988 39874 17990
rect 41229 17987 41295 17990
rect 44173 18050 44239 18053
rect 45318 18050 45324 18052
rect 44173 18048 45324 18050
rect 44173 17992 44178 18048
rect 44234 17992 45324 18048
rect 44173 17990 45324 17992
rect 44173 17987 44239 17990
rect 45318 17988 45324 17990
rect 45388 18050 45394 18052
rect 47117 18050 47183 18053
rect 47761 18052 47827 18053
rect 47710 18050 47716 18052
rect 45388 18048 47183 18050
rect 45388 17992 47122 18048
rect 47178 17992 47183 18048
rect 45388 17990 47183 17992
rect 47670 17990 47716 18050
rect 47780 18048 47827 18052
rect 47822 17992 47827 18048
rect 45388 17988 45394 17990
rect 47117 17987 47183 17990
rect 47710 17988 47716 17990
rect 47780 17988 47827 17992
rect 47761 17987 47827 17988
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 41965 17914 42031 17917
rect 37230 17912 42031 17914
rect 37230 17856 41970 17912
rect 42026 17856 42031 17912
rect 37230 17854 42031 17856
rect 34329 17851 34395 17854
rect 36445 17851 36511 17854
rect 41965 17851 42031 17854
rect 43345 17914 43411 17917
rect 46974 17914 46980 17916
rect 43345 17912 46980 17914
rect 43345 17856 43350 17912
rect 43406 17856 46980 17912
rect 43345 17854 46980 17856
rect 43345 17851 43411 17854
rect 46974 17852 46980 17854
rect 47044 17914 47050 17916
rect 47761 17914 47827 17917
rect 47044 17912 47827 17914
rect 47044 17856 47766 17912
rect 47822 17856 47827 17912
rect 47044 17854 47827 17856
rect 47044 17852 47050 17854
rect 47761 17851 47827 17854
rect 35934 17778 35940 17780
rect 31710 17718 35940 17778
rect 19425 17715 19491 17718
rect 21265 17715 21331 17718
rect 27613 17715 27679 17718
rect 35934 17716 35940 17718
rect 36004 17716 36010 17780
rect 36905 17778 36971 17781
rect 44081 17778 44147 17781
rect 36905 17776 44147 17778
rect 36905 17720 36910 17776
rect 36966 17720 44086 17776
rect 44142 17720 44147 17776
rect 36905 17718 44147 17720
rect 36905 17715 36971 17718
rect 44081 17715 44147 17718
rect 46289 17778 46355 17781
rect 46565 17778 46631 17781
rect 50200 17778 51000 17808
rect 46289 17776 51000 17778
rect 46289 17720 46294 17776
rect 46350 17720 46570 17776
rect 46626 17720 51000 17776
rect 46289 17718 51000 17720
rect 46289 17715 46355 17718
rect 46565 17715 46631 17718
rect 50200 17688 51000 17718
rect 23841 17642 23907 17645
rect 18830 17640 23907 17642
rect 18830 17584 23846 17640
rect 23902 17584 23907 17640
rect 18830 17582 23907 17584
rect 23841 17579 23907 17582
rect 26918 17580 26924 17644
rect 26988 17642 26994 17644
rect 34237 17642 34303 17645
rect 26988 17640 34303 17642
rect 26988 17584 34242 17640
rect 34298 17584 34303 17640
rect 26988 17582 34303 17584
rect 26988 17580 26994 17582
rect 34237 17579 34303 17582
rect 36721 17642 36787 17645
rect 42149 17642 42215 17645
rect 36721 17640 42215 17642
rect 36721 17584 36726 17640
rect 36782 17584 42154 17640
rect 42210 17584 42215 17640
rect 36721 17582 42215 17584
rect 36721 17579 36787 17582
rect 42149 17579 42215 17582
rect 42333 17642 42399 17645
rect 42333 17640 48514 17642
rect 42333 17584 42338 17640
rect 42394 17584 48514 17640
rect 42333 17582 48514 17584
rect 42333 17579 42399 17582
rect 0 17506 800 17536
rect 2037 17506 2103 17509
rect 0 17504 2103 17506
rect 0 17448 2042 17504
rect 2098 17448 2103 17504
rect 0 17446 2103 17448
rect 0 17416 800 17446
rect 2037 17443 2103 17446
rect 9121 17506 9187 17509
rect 9438 17506 9444 17508
rect 9121 17504 9444 17506
rect 9121 17448 9126 17504
rect 9182 17448 9444 17504
rect 9121 17446 9444 17448
rect 9121 17443 9187 17446
rect 9438 17444 9444 17446
rect 9508 17506 9514 17508
rect 17217 17506 17283 17509
rect 9508 17504 17283 17506
rect 9508 17448 17222 17504
rect 17278 17448 17283 17504
rect 9508 17446 17283 17448
rect 9508 17444 9514 17446
rect 17217 17443 17283 17446
rect 18505 17506 18571 17509
rect 25221 17506 25287 17509
rect 18505 17504 25287 17506
rect 18505 17448 18510 17504
rect 18566 17448 25226 17504
rect 25282 17448 25287 17504
rect 18505 17446 25287 17448
rect 18505 17443 18571 17446
rect 25221 17443 25287 17446
rect 38929 17506 38995 17509
rect 45318 17506 45324 17508
rect 38929 17504 45324 17506
rect 38929 17448 38934 17504
rect 38990 17448 45324 17504
rect 38929 17446 45324 17448
rect 38929 17443 38995 17446
rect 45318 17444 45324 17446
rect 45388 17506 45394 17508
rect 45461 17506 45527 17509
rect 45388 17504 45527 17506
rect 45388 17448 45466 17504
rect 45522 17448 45527 17504
rect 45388 17446 45527 17448
rect 45388 17444 45394 17446
rect 45461 17443 45527 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 12065 17370 12131 17373
rect 13905 17370 13971 17373
rect 12065 17368 13971 17370
rect 12065 17312 12070 17368
rect 12126 17312 13910 17368
rect 13966 17312 13971 17368
rect 12065 17310 13971 17312
rect 12065 17307 12131 17310
rect 13905 17307 13971 17310
rect 14273 17370 14339 17373
rect 17493 17370 17559 17373
rect 14273 17368 17559 17370
rect 14273 17312 14278 17368
rect 14334 17312 17498 17368
rect 17554 17312 17559 17368
rect 14273 17310 17559 17312
rect 14273 17307 14339 17310
rect 17493 17307 17559 17310
rect 19793 17370 19859 17373
rect 21357 17370 21423 17373
rect 19793 17368 21423 17370
rect 19793 17312 19798 17368
rect 19854 17312 21362 17368
rect 21418 17312 21423 17368
rect 19793 17310 21423 17312
rect 19793 17307 19859 17310
rect 21357 17307 21423 17310
rect 26785 17370 26851 17373
rect 27102 17370 27108 17372
rect 26785 17368 27108 17370
rect 26785 17312 26790 17368
rect 26846 17312 27108 17368
rect 26785 17310 27108 17312
rect 26785 17307 26851 17310
rect 27102 17308 27108 17310
rect 27172 17308 27178 17372
rect 35709 17370 35775 17373
rect 31710 17368 35775 17370
rect 31710 17312 35714 17368
rect 35770 17312 35775 17368
rect 31710 17310 35775 17312
rect 7005 17234 7071 17237
rect 7373 17234 7439 17237
rect 7005 17232 7439 17234
rect 7005 17176 7010 17232
rect 7066 17176 7378 17232
rect 7434 17176 7439 17232
rect 7005 17174 7439 17176
rect 7005 17171 7071 17174
rect 7373 17171 7439 17174
rect 8109 17234 8175 17237
rect 12433 17234 12499 17237
rect 24209 17234 24275 17237
rect 8109 17232 24275 17234
rect 8109 17176 8114 17232
rect 8170 17176 12438 17232
rect 12494 17176 24214 17232
rect 24270 17176 24275 17232
rect 8109 17174 24275 17176
rect 8109 17171 8175 17174
rect 12433 17171 12499 17174
rect 24209 17171 24275 17174
rect 27981 17234 28047 17237
rect 31710 17234 31770 17310
rect 35709 17307 35775 17310
rect 38745 17370 38811 17373
rect 40953 17370 41019 17373
rect 38745 17368 41019 17370
rect 38745 17312 38750 17368
rect 38806 17312 40958 17368
rect 41014 17312 41019 17368
rect 38745 17310 41019 17312
rect 38745 17307 38811 17310
rect 40953 17307 41019 17310
rect 42885 17370 42951 17373
rect 45645 17370 45711 17373
rect 42885 17368 45711 17370
rect 42885 17312 42890 17368
rect 42946 17312 45650 17368
rect 45706 17312 45711 17368
rect 42885 17310 45711 17312
rect 48454 17370 48514 17582
rect 50200 17370 51000 17400
rect 48454 17310 51000 17370
rect 42885 17307 42951 17310
rect 45645 17307 45711 17310
rect 50200 17280 51000 17310
rect 27981 17232 31770 17234
rect 27981 17176 27986 17232
rect 28042 17176 31770 17232
rect 27981 17174 31770 17176
rect 32857 17234 32923 17237
rect 42793 17234 42859 17237
rect 32857 17232 42859 17234
rect 32857 17176 32862 17232
rect 32918 17176 42798 17232
rect 42854 17176 42859 17232
rect 32857 17174 42859 17176
rect 27981 17171 28047 17174
rect 32857 17171 32923 17174
rect 42793 17171 42859 17174
rect 0 17098 800 17128
rect 1209 17098 1275 17101
rect 0 17096 1275 17098
rect 0 17040 1214 17096
rect 1270 17040 1275 17096
rect 0 17038 1275 17040
rect 0 17008 800 17038
rect 1209 17035 1275 17038
rect 11789 17098 11855 17101
rect 16021 17098 16087 17101
rect 26693 17098 26759 17101
rect 11789 17096 26759 17098
rect 11789 17040 11794 17096
rect 11850 17040 16026 17096
rect 16082 17040 26698 17096
rect 26754 17040 26759 17096
rect 11789 17038 26759 17040
rect 11789 17035 11855 17038
rect 16021 17035 16087 17038
rect 26693 17035 26759 17038
rect 27153 17098 27219 17101
rect 33358 17098 33364 17100
rect 27153 17096 33364 17098
rect 27153 17040 27158 17096
rect 27214 17040 33364 17096
rect 27153 17038 33364 17040
rect 27153 17035 27219 17038
rect 33358 17036 33364 17038
rect 33428 17098 33434 17100
rect 34697 17098 34763 17101
rect 33428 17096 34763 17098
rect 33428 17040 34702 17096
rect 34758 17040 34763 17096
rect 33428 17038 34763 17040
rect 33428 17036 33434 17038
rect 34697 17035 34763 17038
rect 35801 17098 35867 17101
rect 43253 17098 43319 17101
rect 35801 17096 43319 17098
rect 35801 17040 35806 17096
rect 35862 17040 43258 17096
rect 43314 17040 43319 17096
rect 35801 17038 43319 17040
rect 35801 17035 35867 17038
rect 43253 17035 43319 17038
rect 3877 16962 3943 16965
rect 12801 16962 12867 16965
rect 3877 16960 12867 16962
rect 3877 16904 3882 16960
rect 3938 16904 12806 16960
rect 12862 16904 12867 16960
rect 3877 16902 12867 16904
rect 3877 16899 3943 16902
rect 12801 16899 12867 16902
rect 13670 16900 13676 16964
rect 13740 16962 13746 16964
rect 18638 16962 18644 16964
rect 13740 16902 18644 16962
rect 13740 16900 13746 16902
rect 18638 16900 18644 16902
rect 18708 16900 18714 16964
rect 24025 16962 24091 16965
rect 25957 16962 26023 16965
rect 27705 16964 27771 16965
rect 27654 16962 27660 16964
rect 24025 16960 26023 16962
rect 24025 16904 24030 16960
rect 24086 16904 25962 16960
rect 26018 16904 26023 16960
rect 24025 16902 26023 16904
rect 27614 16902 27660 16962
rect 27724 16960 27771 16964
rect 27766 16904 27771 16960
rect 24025 16899 24091 16902
rect 25957 16899 26023 16902
rect 27654 16900 27660 16902
rect 27724 16900 27771 16904
rect 27705 16899 27771 16900
rect 34329 16962 34395 16965
rect 34462 16962 34468 16964
rect 34329 16960 34468 16962
rect 34329 16904 34334 16960
rect 34390 16904 34468 16960
rect 34329 16902 34468 16904
rect 34329 16899 34395 16902
rect 34462 16900 34468 16902
rect 34532 16962 34538 16964
rect 36537 16962 36603 16965
rect 36905 16964 36971 16965
rect 36854 16962 36860 16964
rect 34532 16960 36603 16962
rect 34532 16904 36542 16960
rect 36598 16904 36603 16960
rect 34532 16902 36603 16904
rect 36814 16902 36860 16962
rect 36924 16962 36971 16964
rect 40585 16962 40651 16965
rect 36924 16960 40651 16962
rect 36966 16904 40590 16960
rect 40646 16904 40651 16960
rect 34532 16900 34538 16902
rect 36537 16899 36603 16902
rect 36854 16900 36860 16902
rect 36924 16902 40651 16904
rect 36924 16900 36971 16902
rect 36905 16899 36971 16900
rect 40585 16899 40651 16902
rect 46013 16962 46079 16965
rect 50200 16962 51000 16992
rect 46013 16960 51000 16962
rect 46013 16904 46018 16960
rect 46074 16904 51000 16960
rect 46013 16902 51000 16904
rect 46013 16899 46079 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 50200 16872 51000 16902
rect 42946 16831 43262 16832
rect 14733 16826 14799 16829
rect 21633 16826 21699 16829
rect 14733 16824 21699 16826
rect 14733 16768 14738 16824
rect 14794 16768 21638 16824
rect 21694 16768 21699 16824
rect 14733 16766 21699 16768
rect 14733 16763 14799 16766
rect 21633 16763 21699 16766
rect 25773 16826 25839 16829
rect 27521 16826 27587 16829
rect 25773 16824 27587 16826
rect 25773 16768 25778 16824
rect 25834 16768 27526 16824
rect 27582 16768 27587 16824
rect 25773 16766 27587 16768
rect 25773 16763 25839 16766
rect 27521 16763 27587 16766
rect 36353 16826 36419 16829
rect 38694 16826 38700 16828
rect 36353 16824 38700 16826
rect 36353 16768 36358 16824
rect 36414 16768 38700 16824
rect 36353 16766 38700 16768
rect 36353 16763 36419 16766
rect 38694 16764 38700 16766
rect 38764 16826 38770 16828
rect 40493 16826 40559 16829
rect 42793 16826 42859 16829
rect 38764 16824 42859 16826
rect 38764 16768 40498 16824
rect 40554 16768 42798 16824
rect 42854 16768 42859 16824
rect 38764 16766 42859 16768
rect 38764 16764 38770 16766
rect 40493 16763 40559 16766
rect 42793 16763 42859 16766
rect 44725 16826 44791 16829
rect 47209 16826 47275 16829
rect 44725 16824 47275 16826
rect 44725 16768 44730 16824
rect 44786 16768 47214 16824
rect 47270 16768 47275 16824
rect 44725 16766 47275 16768
rect 44725 16763 44791 16766
rect 47209 16763 47275 16766
rect 0 16690 800 16720
rect 1301 16690 1367 16693
rect 0 16688 1367 16690
rect 0 16632 1306 16688
rect 1362 16632 1367 16688
rect 0 16630 1367 16632
rect 0 16600 800 16630
rect 1301 16627 1367 16630
rect 6361 16690 6427 16693
rect 13537 16690 13603 16693
rect 6361 16688 13603 16690
rect 6361 16632 6366 16688
rect 6422 16632 13542 16688
rect 13598 16632 13603 16688
rect 6361 16630 13603 16632
rect 6361 16627 6427 16630
rect 13537 16627 13603 16630
rect 14774 16628 14780 16692
rect 14844 16690 14850 16692
rect 15101 16690 15167 16693
rect 14844 16688 15167 16690
rect 14844 16632 15106 16688
rect 15162 16632 15167 16688
rect 14844 16630 15167 16632
rect 14844 16628 14850 16630
rect 15101 16627 15167 16630
rect 17309 16692 17375 16693
rect 17309 16688 17356 16692
rect 17420 16690 17426 16692
rect 17953 16690 18019 16693
rect 18965 16690 19031 16693
rect 22553 16690 22619 16693
rect 27889 16690 27955 16693
rect 29177 16690 29243 16693
rect 17309 16632 17314 16688
rect 17309 16628 17356 16632
rect 17420 16630 17466 16690
rect 17953 16688 19031 16690
rect 17953 16632 17958 16688
rect 18014 16632 18970 16688
rect 19026 16632 19031 16688
rect 17953 16630 19031 16632
rect 17420 16628 17426 16630
rect 17309 16627 17375 16628
rect 17953 16627 18019 16630
rect 18965 16627 19031 16630
rect 22050 16688 29243 16690
rect 22050 16632 22558 16688
rect 22614 16632 27894 16688
rect 27950 16632 29182 16688
rect 29238 16632 29243 16688
rect 22050 16630 29243 16632
rect 5257 16554 5323 16557
rect 10961 16554 11027 16557
rect 17585 16554 17651 16557
rect 5257 16552 8402 16554
rect 5257 16496 5262 16552
rect 5318 16496 8402 16552
rect 5257 16494 8402 16496
rect 5257 16491 5323 16494
rect 8342 16418 8402 16494
rect 10961 16552 17651 16554
rect 10961 16496 10966 16552
rect 11022 16496 17590 16552
rect 17646 16496 17651 16552
rect 10961 16494 17651 16496
rect 10961 16491 11027 16494
rect 17585 16491 17651 16494
rect 18965 16554 19031 16557
rect 22050 16554 22110 16630
rect 22553 16627 22619 16630
rect 27889 16627 27955 16630
rect 29177 16627 29243 16630
rect 30005 16690 30071 16693
rect 31477 16690 31543 16693
rect 30005 16688 31543 16690
rect 30005 16632 30010 16688
rect 30066 16632 31482 16688
rect 31538 16632 31543 16688
rect 30005 16630 31543 16632
rect 30005 16627 30071 16630
rect 31477 16627 31543 16630
rect 31937 16690 32003 16693
rect 34053 16690 34119 16693
rect 31937 16688 34119 16690
rect 31937 16632 31942 16688
rect 31998 16632 34058 16688
rect 34114 16632 34119 16688
rect 31937 16630 34119 16632
rect 31937 16627 32003 16630
rect 34053 16627 34119 16630
rect 35750 16628 35756 16692
rect 35820 16690 35826 16692
rect 37457 16690 37523 16693
rect 35820 16688 37523 16690
rect 35820 16632 37462 16688
rect 37518 16632 37523 16688
rect 35820 16630 37523 16632
rect 35820 16628 35826 16630
rect 37457 16627 37523 16630
rect 47209 16690 47275 16693
rect 47342 16690 47348 16692
rect 47209 16688 47348 16690
rect 47209 16632 47214 16688
rect 47270 16632 47348 16688
rect 47209 16630 47348 16632
rect 47209 16627 47275 16630
rect 47342 16628 47348 16630
rect 47412 16628 47418 16692
rect 18965 16552 22110 16554
rect 18965 16496 18970 16552
rect 19026 16496 22110 16552
rect 18965 16494 22110 16496
rect 23289 16554 23355 16557
rect 24761 16554 24827 16557
rect 23289 16552 23490 16554
rect 23289 16496 23294 16552
rect 23350 16496 23490 16552
rect 23289 16494 23490 16496
rect 18965 16491 19031 16494
rect 23289 16491 23355 16494
rect 15193 16418 15259 16421
rect 8342 16416 15259 16418
rect 8342 16360 15198 16416
rect 15254 16360 15259 16416
rect 8342 16358 15259 16360
rect 15193 16355 15259 16358
rect 16021 16420 16087 16421
rect 16021 16416 16068 16420
rect 16132 16418 16138 16420
rect 23430 16418 23490 16494
rect 24761 16552 28458 16554
rect 24761 16496 24766 16552
rect 24822 16496 28458 16552
rect 24761 16494 28458 16496
rect 24761 16491 24827 16494
rect 27153 16418 27219 16421
rect 16021 16360 16026 16416
rect 16021 16356 16068 16360
rect 16132 16358 16178 16418
rect 23430 16416 27219 16418
rect 23430 16360 27158 16416
rect 27214 16360 27219 16416
rect 23430 16358 27219 16360
rect 28398 16418 28458 16494
rect 29494 16492 29500 16556
rect 29564 16554 29570 16556
rect 33409 16554 33475 16557
rect 29564 16552 33475 16554
rect 29564 16496 33414 16552
rect 33470 16496 33475 16552
rect 29564 16494 33475 16496
rect 29564 16492 29570 16494
rect 33409 16491 33475 16494
rect 34278 16492 34284 16556
rect 34348 16554 34354 16556
rect 38653 16554 38719 16557
rect 41321 16554 41387 16557
rect 34348 16552 41387 16554
rect 34348 16496 38658 16552
rect 38714 16496 41326 16552
rect 41382 16496 41387 16552
rect 34348 16494 41387 16496
rect 34348 16492 34354 16494
rect 38653 16491 38719 16494
rect 41321 16491 41387 16494
rect 45093 16554 45159 16557
rect 46749 16554 46815 16557
rect 50200 16554 51000 16584
rect 45093 16552 46815 16554
rect 45093 16496 45098 16552
rect 45154 16496 46754 16552
rect 46810 16496 46815 16552
rect 45093 16494 46815 16496
rect 45093 16491 45159 16494
rect 46749 16491 46815 16494
rect 47718 16494 51000 16554
rect 31569 16418 31635 16421
rect 28398 16416 31635 16418
rect 28398 16360 31574 16416
rect 31630 16360 31635 16416
rect 28398 16358 31635 16360
rect 16132 16356 16138 16358
rect 16021 16355 16087 16356
rect 27153 16355 27219 16358
rect 31569 16355 31635 16358
rect 31886 16356 31892 16420
rect 31956 16418 31962 16420
rect 36813 16418 36879 16421
rect 31956 16416 36879 16418
rect 31956 16360 36818 16416
rect 36874 16360 36879 16416
rect 31956 16358 36879 16360
rect 31956 16356 31962 16358
rect 36813 16355 36879 16358
rect 38837 16416 38903 16421
rect 38837 16360 38842 16416
rect 38898 16360 38903 16416
rect 38837 16355 38903 16360
rect 39757 16418 39823 16421
rect 44541 16418 44607 16421
rect 45369 16420 45435 16421
rect 45318 16418 45324 16420
rect 39757 16416 44607 16418
rect 39757 16360 39762 16416
rect 39818 16360 44546 16416
rect 44602 16360 44607 16416
rect 39757 16358 44607 16360
rect 45278 16358 45324 16418
rect 45388 16416 45435 16420
rect 45430 16360 45435 16416
rect 39757 16355 39823 16358
rect 44541 16355 44607 16358
rect 45318 16356 45324 16358
rect 45388 16356 45435 16360
rect 45502 16356 45508 16420
rect 45572 16418 45578 16420
rect 46289 16418 46355 16421
rect 45572 16416 46355 16418
rect 45572 16360 46294 16416
rect 46350 16360 46355 16416
rect 45572 16358 46355 16360
rect 45572 16356 45578 16358
rect 45369 16355 45435 16356
rect 46289 16355 46355 16358
rect 46790 16356 46796 16420
rect 46860 16418 46866 16420
rect 47718 16418 47778 16494
rect 50200 16464 51000 16494
rect 46860 16358 47778 16418
rect 46860 16356 46866 16358
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 1301 16282 1367 16285
rect 0 16280 1367 16282
rect 0 16224 1306 16280
rect 1362 16224 1367 16280
rect 0 16222 1367 16224
rect 0 16192 800 16222
rect 1301 16219 1367 16222
rect 11973 16282 12039 16285
rect 16021 16282 16087 16285
rect 11973 16280 16087 16282
rect 11973 16224 11978 16280
rect 12034 16224 16026 16280
rect 16082 16224 16087 16280
rect 11973 16222 16087 16224
rect 11973 16219 12039 16222
rect 16021 16219 16087 16222
rect 18638 16220 18644 16284
rect 18708 16282 18714 16284
rect 21357 16282 21423 16285
rect 22461 16284 22527 16285
rect 22461 16282 22508 16284
rect 18708 16280 22508 16282
rect 18708 16224 21362 16280
rect 21418 16224 22466 16280
rect 18708 16222 22508 16224
rect 18708 16220 18714 16222
rect 21357 16219 21423 16222
rect 22461 16220 22508 16222
rect 22572 16220 22578 16284
rect 36997 16282 37063 16285
rect 32630 16280 37063 16282
rect 32630 16224 37002 16280
rect 37058 16224 37063 16280
rect 32630 16222 37063 16224
rect 38840 16282 38900 16355
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 40125 16282 40191 16285
rect 38840 16280 40191 16282
rect 38840 16224 40130 16280
rect 40186 16224 40191 16280
rect 38840 16222 40191 16224
rect 22461 16219 22527 16220
rect 3601 16146 3667 16149
rect 14365 16146 14431 16149
rect 14733 16146 14799 16149
rect 3601 16144 14799 16146
rect 3601 16088 3606 16144
rect 3662 16088 14370 16144
rect 14426 16088 14738 16144
rect 14794 16088 14799 16144
rect 3601 16086 14799 16088
rect 3601 16083 3667 16086
rect 14365 16083 14431 16086
rect 14733 16083 14799 16086
rect 15142 16084 15148 16148
rect 15212 16146 15218 16148
rect 18321 16146 18387 16149
rect 15212 16144 18387 16146
rect 15212 16088 18326 16144
rect 18382 16088 18387 16144
rect 15212 16086 18387 16088
rect 15212 16084 15218 16086
rect 18321 16083 18387 16086
rect 19885 16146 19951 16149
rect 24761 16146 24827 16149
rect 19885 16144 24827 16146
rect 19885 16088 19890 16144
rect 19946 16088 24766 16144
rect 24822 16088 24827 16144
rect 19885 16086 24827 16088
rect 19885 16083 19951 16086
rect 24761 16083 24827 16086
rect 26693 16146 26759 16149
rect 32630 16146 32690 16222
rect 36997 16219 37063 16222
rect 40125 16219 40191 16222
rect 41689 16282 41755 16285
rect 43805 16282 43871 16285
rect 46933 16282 46999 16285
rect 41689 16280 43871 16282
rect 41689 16224 41694 16280
rect 41750 16224 43810 16280
rect 43866 16224 43871 16280
rect 41689 16222 43871 16224
rect 41689 16219 41755 16222
rect 43805 16219 43871 16222
rect 45510 16280 46999 16282
rect 45510 16224 46938 16280
rect 46994 16224 46999 16280
rect 45510 16222 46999 16224
rect 32857 16148 32923 16149
rect 26693 16144 32690 16146
rect 26693 16088 26698 16144
rect 26754 16088 32690 16144
rect 26693 16086 32690 16088
rect 26693 16083 26759 16086
rect 32806 16084 32812 16148
rect 32876 16146 32923 16148
rect 45510 16146 45570 16222
rect 46933 16219 46999 16222
rect 47669 16146 47735 16149
rect 50200 16146 51000 16176
rect 32876 16144 32968 16146
rect 32918 16088 32968 16144
rect 32876 16086 32968 16088
rect 33044 16086 45570 16146
rect 47350 16144 51000 16146
rect 47350 16088 47674 16144
rect 47730 16088 51000 16144
rect 47350 16086 51000 16088
rect 32876 16084 32923 16086
rect 32857 16083 32923 16084
rect 6729 16010 6795 16013
rect 8937 16010 9003 16013
rect 6729 16008 9003 16010
rect 6729 15952 6734 16008
rect 6790 15952 8942 16008
rect 8998 15952 9003 16008
rect 6729 15950 9003 15952
rect 6729 15947 6795 15950
rect 8937 15947 9003 15950
rect 10961 16010 11027 16013
rect 12985 16010 13051 16013
rect 10961 16008 13051 16010
rect 10961 15952 10966 16008
rect 11022 15952 12990 16008
rect 13046 15952 13051 16008
rect 10961 15950 13051 15952
rect 10961 15947 11027 15950
rect 12985 15947 13051 15950
rect 13813 16010 13879 16013
rect 14038 16010 14044 16012
rect 13813 16008 14044 16010
rect 13813 15952 13818 16008
rect 13874 15952 14044 16008
rect 13813 15950 14044 15952
rect 13813 15947 13879 15950
rect 14038 15948 14044 15950
rect 14108 16010 14114 16012
rect 15561 16010 15627 16013
rect 14108 16008 15627 16010
rect 14108 15952 15566 16008
rect 15622 15952 15627 16008
rect 14108 15950 15627 15952
rect 14108 15948 14114 15950
rect 15561 15947 15627 15950
rect 15929 16010 15995 16013
rect 25497 16010 25563 16013
rect 15929 16008 25563 16010
rect 15929 15952 15934 16008
rect 15990 15952 25502 16008
rect 25558 15952 25563 16008
rect 15929 15950 25563 15952
rect 15929 15947 15995 15950
rect 25497 15947 25563 15950
rect 32857 16010 32923 16013
rect 33044 16010 33104 16086
rect 32857 16008 33104 16010
rect 32857 15952 32862 16008
rect 32918 15952 33104 16008
rect 32857 15950 33104 15952
rect 35249 16010 35315 16013
rect 35985 16010 36051 16013
rect 36813 16010 36879 16013
rect 42609 16010 42675 16013
rect 47025 16010 47091 16013
rect 35249 16008 42675 16010
rect 35249 15952 35254 16008
rect 35310 15952 35990 16008
rect 36046 15952 36818 16008
rect 36874 15952 42614 16008
rect 42670 15952 42675 16008
rect 35249 15950 42675 15952
rect 32857 15947 32923 15950
rect 35249 15947 35315 15950
rect 35985 15947 36051 15950
rect 36813 15947 36879 15950
rect 42609 15947 42675 15950
rect 42750 16008 47091 16010
rect 42750 15952 47030 16008
rect 47086 15952 47091 16008
rect 42750 15950 47091 15952
rect 0 15874 800 15904
rect 1301 15874 1367 15877
rect 0 15872 1367 15874
rect 0 15816 1306 15872
rect 1362 15816 1367 15872
rect 0 15814 1367 15816
rect 0 15784 800 15814
rect 1301 15811 1367 15814
rect 6453 15874 6519 15877
rect 10041 15874 10107 15877
rect 6453 15872 10107 15874
rect 6453 15816 6458 15872
rect 6514 15816 10046 15872
rect 10102 15816 10107 15872
rect 6453 15814 10107 15816
rect 6453 15811 6519 15814
rect 10041 15811 10107 15814
rect 14365 15874 14431 15877
rect 19885 15874 19951 15877
rect 14365 15872 19951 15874
rect 14365 15816 14370 15872
rect 14426 15816 19890 15872
rect 19946 15816 19951 15872
rect 14365 15814 19951 15816
rect 14365 15811 14431 15814
rect 19885 15811 19951 15814
rect 38837 15874 38903 15877
rect 39665 15874 39731 15877
rect 40769 15874 40835 15877
rect 41689 15874 41755 15877
rect 38837 15872 41755 15874
rect 38837 15816 38842 15872
rect 38898 15816 39670 15872
rect 39726 15816 40774 15872
rect 40830 15816 41694 15872
rect 41750 15816 41755 15872
rect 38837 15814 41755 15816
rect 38837 15811 38903 15814
rect 39665 15811 39731 15814
rect 40769 15811 40835 15814
rect 41689 15811 41755 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 5349 15738 5415 15741
rect 11094 15738 11100 15740
rect 5349 15736 11100 15738
rect 5349 15680 5354 15736
rect 5410 15680 11100 15736
rect 5349 15678 11100 15680
rect 5349 15675 5415 15678
rect 11094 15676 11100 15678
rect 11164 15676 11170 15740
rect 13629 15738 13695 15741
rect 16205 15738 16271 15741
rect 13629 15736 16271 15738
rect 13629 15680 13634 15736
rect 13690 15680 16210 15736
rect 16266 15680 16271 15736
rect 13629 15678 16271 15680
rect 13629 15675 13695 15678
rect 16205 15675 16271 15678
rect 17125 15738 17191 15741
rect 17861 15738 17927 15741
rect 17125 15736 17927 15738
rect 17125 15680 17130 15736
rect 17186 15680 17866 15736
rect 17922 15680 17927 15736
rect 17125 15678 17927 15680
rect 17125 15675 17191 15678
rect 17861 15675 17927 15678
rect 21541 15738 21607 15741
rect 22369 15738 22435 15741
rect 21541 15736 22435 15738
rect 21541 15680 21546 15736
rect 21602 15680 22374 15736
rect 22430 15680 22435 15736
rect 21541 15678 22435 15680
rect 21541 15675 21607 15678
rect 22369 15675 22435 15678
rect 25681 15738 25747 15741
rect 27889 15738 27955 15741
rect 25681 15736 27955 15738
rect 25681 15680 25686 15736
rect 25742 15680 27894 15736
rect 27950 15680 27955 15736
rect 25681 15678 27955 15680
rect 25681 15675 25747 15678
rect 27889 15675 27955 15678
rect 37457 15738 37523 15741
rect 42750 15738 42810 15950
rect 47025 15947 47091 15950
rect 44398 15812 44404 15876
rect 44468 15874 44474 15876
rect 47350 15874 47410 16086
rect 47669 16083 47735 16086
rect 50200 16056 51000 16086
rect 44468 15814 47410 15874
rect 44468 15812 44474 15814
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 37457 15736 42810 15738
rect 37457 15680 37462 15736
rect 37518 15680 42810 15736
rect 37457 15678 42810 15680
rect 49601 15738 49667 15741
rect 50200 15738 51000 15768
rect 49601 15736 51000 15738
rect 49601 15680 49606 15736
rect 49662 15680 51000 15736
rect 49601 15678 51000 15680
rect 37457 15675 37523 15678
rect 49601 15675 49667 15678
rect 50200 15648 51000 15678
rect 4797 15602 4863 15605
rect 8661 15602 8727 15605
rect 4797 15600 8727 15602
rect 4797 15544 4802 15600
rect 4858 15544 8666 15600
rect 8722 15544 8727 15600
rect 4797 15542 8727 15544
rect 4797 15539 4863 15542
rect 8661 15539 8727 15542
rect 10041 15602 10107 15605
rect 12801 15602 12867 15605
rect 25865 15602 25931 15605
rect 10041 15600 25931 15602
rect 10041 15544 10046 15600
rect 10102 15544 12806 15600
rect 12862 15544 25870 15600
rect 25926 15544 25931 15600
rect 10041 15542 25931 15544
rect 10041 15539 10107 15542
rect 12801 15539 12867 15542
rect 25865 15539 25931 15542
rect 27061 15602 27127 15605
rect 27521 15602 27587 15605
rect 27061 15600 27587 15602
rect 27061 15544 27066 15600
rect 27122 15544 27526 15600
rect 27582 15544 27587 15600
rect 27061 15542 27587 15544
rect 27061 15539 27127 15542
rect 27521 15539 27587 15542
rect 31661 15602 31727 15605
rect 45461 15602 45527 15605
rect 31661 15600 45527 15602
rect 31661 15544 31666 15600
rect 31722 15544 45466 15600
rect 45522 15544 45527 15600
rect 31661 15542 45527 15544
rect 31661 15539 31727 15542
rect 45461 15539 45527 15542
rect 0 15466 800 15496
rect 1301 15466 1367 15469
rect 0 15464 1367 15466
rect 0 15408 1306 15464
rect 1362 15408 1367 15464
rect 0 15406 1367 15408
rect 0 15376 800 15406
rect 1301 15403 1367 15406
rect 9489 15466 9555 15469
rect 18689 15466 18755 15469
rect 38469 15466 38535 15469
rect 44633 15466 44699 15469
rect 9489 15464 18522 15466
rect 9489 15408 9494 15464
rect 9550 15408 18522 15464
rect 9489 15406 18522 15408
rect 9489 15403 9555 15406
rect 1761 15330 1827 15333
rect 11973 15330 12039 15333
rect 12985 15330 13051 15333
rect 1761 15328 7666 15330
rect 1761 15272 1766 15328
rect 1822 15272 7666 15328
rect 1761 15270 7666 15272
rect 1761 15267 1827 15270
rect 0 15058 800 15088
rect 1301 15058 1367 15061
rect 0 15056 1367 15058
rect 0 15000 1306 15056
rect 1362 15000 1367 15056
rect 0 14998 1367 15000
rect 0 14968 800 14998
rect 1301 14995 1367 14998
rect 7606 14922 7666 15270
rect 11973 15328 13051 15330
rect 11973 15272 11978 15328
rect 12034 15272 12990 15328
rect 13046 15272 13051 15328
rect 11973 15270 13051 15272
rect 11973 15267 12039 15270
rect 12985 15267 13051 15270
rect 13629 15330 13695 15333
rect 17585 15330 17651 15333
rect 13629 15328 17651 15330
rect 13629 15272 13634 15328
rect 13690 15272 17590 15328
rect 17646 15272 17651 15328
rect 13629 15270 17651 15272
rect 18462 15330 18522 15406
rect 18689 15464 38394 15466
rect 18689 15408 18694 15464
rect 18750 15408 38394 15464
rect 18689 15406 38394 15408
rect 18689 15403 18755 15406
rect 22829 15330 22895 15333
rect 23105 15330 23171 15333
rect 18462 15328 23171 15330
rect 18462 15272 22834 15328
rect 22890 15272 23110 15328
rect 23166 15272 23171 15328
rect 18462 15270 23171 15272
rect 13629 15267 13695 15270
rect 17585 15267 17651 15270
rect 22829 15267 22895 15270
rect 23105 15267 23171 15270
rect 26509 15330 26575 15333
rect 27521 15330 27587 15333
rect 26509 15328 27587 15330
rect 26509 15272 26514 15328
rect 26570 15272 27526 15328
rect 27582 15272 27587 15328
rect 26509 15270 27587 15272
rect 26509 15267 26575 15270
rect 27521 15267 27587 15270
rect 28441 15330 28507 15333
rect 31937 15330 32003 15333
rect 28441 15328 32003 15330
rect 28441 15272 28446 15328
rect 28502 15272 31942 15328
rect 31998 15272 32003 15328
rect 28441 15270 32003 15272
rect 28441 15267 28507 15270
rect 31937 15267 32003 15270
rect 32949 15330 33015 15333
rect 35433 15330 35499 15333
rect 32949 15328 35499 15330
rect 32949 15272 32954 15328
rect 33010 15272 35438 15328
rect 35494 15272 35499 15328
rect 32949 15270 35499 15272
rect 38334 15330 38394 15406
rect 38469 15464 44699 15466
rect 38469 15408 38474 15464
rect 38530 15408 44638 15464
rect 44694 15408 44699 15464
rect 38469 15406 44699 15408
rect 38469 15403 38535 15406
rect 44633 15403 44699 15406
rect 45829 15466 45895 15469
rect 45829 15464 48514 15466
rect 45829 15408 45834 15464
rect 45890 15408 48514 15464
rect 45829 15406 48514 15408
rect 45829 15403 45895 15406
rect 38745 15330 38811 15333
rect 38334 15328 38811 15330
rect 38334 15272 38750 15328
rect 38806 15272 38811 15328
rect 38334 15270 38811 15272
rect 32949 15267 33015 15270
rect 35433 15267 35499 15270
rect 38745 15267 38811 15270
rect 40350 15268 40356 15332
rect 40420 15330 40426 15332
rect 41137 15330 41203 15333
rect 40420 15328 41203 15330
rect 40420 15272 41142 15328
rect 41198 15272 41203 15328
rect 40420 15270 41203 15272
rect 40420 15268 40426 15270
rect 41137 15267 41203 15270
rect 41270 15268 41276 15332
rect 41340 15330 41346 15332
rect 42149 15330 42215 15333
rect 41340 15328 42215 15330
rect 41340 15272 42154 15328
rect 42210 15272 42215 15328
rect 41340 15270 42215 15272
rect 41340 15268 41346 15270
rect 42149 15267 42215 15270
rect 46054 15268 46060 15332
rect 46124 15330 46130 15332
rect 47669 15330 47735 15333
rect 46124 15328 47735 15330
rect 46124 15272 47674 15328
rect 47730 15272 47735 15328
rect 46124 15270 47735 15272
rect 48454 15330 48514 15406
rect 50200 15330 51000 15360
rect 48454 15270 51000 15330
rect 46124 15268 46130 15270
rect 47669 15267 47735 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 50200 15240 51000 15270
rect 47946 15199 48262 15200
rect 15837 15194 15903 15197
rect 10228 15192 15903 15194
rect 10228 15136 15842 15192
rect 15898 15136 15903 15192
rect 10228 15134 15903 15136
rect 8017 15058 8083 15061
rect 10228 15058 10288 15134
rect 15837 15131 15903 15134
rect 18505 15194 18571 15197
rect 26969 15194 27035 15197
rect 30833 15194 30899 15197
rect 31150 15194 31156 15196
rect 18505 15192 18890 15194
rect 18505 15136 18510 15192
rect 18566 15136 18890 15192
rect 18505 15134 18890 15136
rect 18505 15131 18571 15134
rect 18830 15061 18890 15134
rect 26969 15192 27722 15194
rect 26969 15136 26974 15192
rect 27030 15136 27722 15192
rect 26969 15134 27722 15136
rect 26969 15131 27035 15134
rect 8017 15056 10288 15058
rect 8017 15000 8022 15056
rect 8078 15000 10288 15056
rect 8017 14998 10288 15000
rect 8017 14995 8083 14998
rect 12014 14996 12020 15060
rect 12084 15058 12090 15060
rect 12249 15058 12315 15061
rect 12084 15056 12315 15058
rect 12084 15000 12254 15056
rect 12310 15000 12315 15056
rect 12084 14998 12315 15000
rect 12084 14996 12090 14998
rect 12249 14995 12315 14998
rect 13537 15058 13603 15061
rect 14181 15058 14247 15061
rect 13537 15056 14247 15058
rect 13537 15000 13542 15056
rect 13598 15000 14186 15056
rect 14242 15000 14247 15056
rect 13537 14998 14247 15000
rect 13537 14995 13603 14998
rect 14181 14995 14247 14998
rect 14825 15058 14891 15061
rect 16573 15058 16639 15061
rect 14825 15056 16639 15058
rect 14825 15000 14830 15056
rect 14886 15000 16578 15056
rect 16634 15000 16639 15056
rect 14825 14998 16639 15000
rect 18830 15056 18939 15061
rect 18830 15000 18878 15056
rect 18934 15000 18939 15056
rect 18830 14998 18939 15000
rect 14825 14995 14891 14998
rect 16573 14995 16639 14998
rect 18873 14995 18939 14998
rect 23197 15058 23263 15061
rect 26601 15058 26667 15061
rect 27662 15058 27722 15134
rect 30833 15192 31156 15194
rect 30833 15136 30838 15192
rect 30894 15136 31156 15192
rect 30833 15134 31156 15136
rect 30833 15131 30899 15134
rect 31150 15132 31156 15134
rect 31220 15132 31226 15196
rect 31661 15194 31727 15197
rect 33685 15194 33751 15197
rect 38929 15196 38995 15197
rect 38878 15194 38884 15196
rect 31661 15192 33751 15194
rect 31661 15136 31666 15192
rect 31722 15136 33690 15192
rect 33746 15136 33751 15192
rect 31661 15134 33751 15136
rect 38838 15134 38884 15194
rect 38948 15192 38995 15196
rect 38990 15136 38995 15192
rect 31661 15131 31727 15134
rect 33685 15131 33751 15134
rect 38878 15132 38884 15134
rect 38948 15132 38995 15136
rect 38929 15131 38995 15132
rect 39573 15194 39639 15197
rect 40309 15194 40375 15197
rect 45369 15194 45435 15197
rect 39573 15192 45435 15194
rect 39573 15136 39578 15192
rect 39634 15136 40314 15192
rect 40370 15136 45374 15192
rect 45430 15136 45435 15192
rect 39573 15134 45435 15136
rect 39573 15131 39639 15134
rect 40309 15131 40375 15134
rect 45369 15131 45435 15134
rect 27889 15058 27955 15061
rect 28901 15058 28967 15061
rect 23197 15056 27584 15058
rect 23197 15000 23202 15056
rect 23258 15000 26606 15056
rect 26662 15000 27584 15056
rect 23197 14998 27584 15000
rect 27662 15056 28967 15058
rect 27662 15000 27894 15056
rect 27950 15000 28906 15056
rect 28962 15000 28967 15056
rect 27662 14998 28967 15000
rect 23197 14995 23263 14998
rect 26601 14995 26667 14998
rect 27524 14925 27584 14998
rect 27889 14995 27955 14998
rect 28901 14995 28967 14998
rect 29085 15058 29151 15061
rect 31569 15058 31635 15061
rect 29085 15056 31635 15058
rect 29085 15000 29090 15056
rect 29146 15000 31574 15056
rect 31630 15000 31635 15056
rect 29085 14998 31635 15000
rect 29085 14995 29151 14998
rect 31569 14995 31635 14998
rect 35525 15058 35591 15061
rect 38193 15058 38259 15061
rect 35525 15056 38259 15058
rect 35525 15000 35530 15056
rect 35586 15000 38198 15056
rect 38254 15000 38259 15056
rect 35525 14998 38259 15000
rect 35525 14995 35591 14998
rect 38193 14995 38259 14998
rect 40861 15058 40927 15061
rect 41638 15058 41644 15060
rect 40861 15056 41644 15058
rect 40861 15000 40866 15056
rect 40922 15000 41644 15056
rect 40861 14998 41644 15000
rect 40861 14995 40927 14998
rect 41638 14996 41644 14998
rect 41708 14996 41714 15060
rect 17033 14922 17099 14925
rect 7606 14920 17099 14922
rect 7606 14864 17038 14920
rect 17094 14864 17099 14920
rect 7606 14862 17099 14864
rect 17033 14859 17099 14862
rect 17217 14922 17283 14925
rect 18454 14922 18460 14924
rect 17217 14920 18460 14922
rect 17217 14864 17222 14920
rect 17278 14864 18460 14920
rect 17217 14862 18460 14864
rect 17217 14859 17283 14862
rect 18454 14860 18460 14862
rect 18524 14860 18530 14924
rect 19517 14922 19583 14925
rect 26734 14922 26740 14924
rect 19517 14920 26740 14922
rect 19517 14864 19522 14920
rect 19578 14864 26740 14920
rect 19517 14862 26740 14864
rect 19517 14859 19583 14862
rect 26734 14860 26740 14862
rect 26804 14860 26810 14924
rect 27521 14922 27587 14925
rect 27981 14922 28047 14925
rect 27430 14920 28047 14922
rect 27430 14864 27526 14920
rect 27582 14864 27986 14920
rect 28042 14864 28047 14920
rect 27430 14862 28047 14864
rect 27521 14859 27587 14862
rect 27981 14859 28047 14862
rect 28257 14922 28323 14925
rect 29177 14922 29243 14925
rect 36997 14922 37063 14925
rect 28257 14920 28826 14922
rect 28257 14864 28262 14920
rect 28318 14864 28826 14920
rect 28257 14862 28826 14864
rect 28257 14859 28323 14862
rect 9121 14786 9187 14789
rect 12709 14786 12775 14789
rect 16389 14788 16455 14789
rect 16389 14786 16436 14788
rect 9121 14784 12775 14786
rect 9121 14728 9126 14784
rect 9182 14728 12714 14784
rect 12770 14728 12775 14784
rect 9121 14726 12775 14728
rect 16344 14784 16436 14786
rect 16500 14786 16506 14788
rect 18413 14786 18479 14789
rect 16500 14784 18479 14786
rect 16344 14728 16394 14784
rect 16500 14728 18418 14784
rect 18474 14728 18479 14784
rect 16344 14726 16436 14728
rect 9121 14723 9187 14726
rect 12709 14723 12775 14726
rect 16389 14724 16436 14726
rect 16500 14726 18479 14728
rect 16500 14724 16506 14726
rect 16389 14723 16455 14724
rect 18413 14723 18479 14726
rect 26233 14786 26299 14789
rect 28533 14786 28599 14789
rect 26233 14784 28599 14786
rect 26233 14728 26238 14784
rect 26294 14728 28538 14784
rect 28594 14728 28599 14784
rect 26233 14726 28599 14728
rect 28766 14786 28826 14862
rect 29177 14920 37063 14922
rect 29177 14864 29182 14920
rect 29238 14864 37002 14920
rect 37058 14864 37063 14920
rect 29177 14862 37063 14864
rect 29177 14859 29243 14862
rect 36997 14859 37063 14862
rect 37590 14860 37596 14924
rect 37660 14922 37666 14924
rect 45921 14922 45987 14925
rect 50061 14922 50127 14925
rect 50200 14922 51000 14952
rect 37660 14862 44098 14922
rect 37660 14860 37666 14862
rect 44038 14789 44098 14862
rect 45921 14920 51000 14922
rect 45921 14864 45926 14920
rect 45982 14864 50066 14920
rect 50122 14864 51000 14920
rect 45921 14862 51000 14864
rect 45921 14859 45987 14862
rect 50061 14859 50127 14862
rect 50200 14832 51000 14862
rect 29361 14786 29427 14789
rect 28766 14784 29427 14786
rect 28766 14728 29366 14784
rect 29422 14728 29427 14784
rect 28766 14726 29427 14728
rect 26233 14723 26299 14726
rect 28533 14723 28599 14726
rect 29361 14723 29427 14726
rect 29637 14786 29703 14789
rect 32673 14786 32739 14789
rect 29637 14784 32739 14786
rect 29637 14728 29642 14784
rect 29698 14728 32678 14784
rect 32734 14728 32739 14784
rect 29637 14726 32739 14728
rect 29637 14723 29703 14726
rect 32673 14723 32739 14726
rect 35801 14786 35867 14789
rect 40217 14786 40283 14789
rect 35801 14784 40283 14786
rect 35801 14728 35806 14784
rect 35862 14728 40222 14784
rect 40278 14728 40283 14784
rect 35801 14726 40283 14728
rect 35801 14723 35867 14726
rect 40217 14723 40283 14726
rect 40902 14724 40908 14788
rect 40972 14786 40978 14788
rect 41229 14786 41295 14789
rect 40972 14784 41295 14786
rect 40972 14728 41234 14784
rect 41290 14728 41295 14784
rect 40972 14726 41295 14728
rect 44038 14784 44147 14789
rect 44038 14728 44086 14784
rect 44142 14728 44147 14784
rect 44038 14726 44147 14728
rect 40972 14724 40978 14726
rect 41229 14723 41295 14726
rect 44081 14723 44147 14726
rect 49918 14724 49924 14788
rect 49988 14786 49994 14788
rect 50061 14786 50127 14789
rect 49988 14784 50127 14786
rect 49988 14728 50066 14784
rect 50122 14728 50127 14784
rect 49988 14726 50127 14728
rect 49988 14724 49994 14726
rect 50061 14723 50127 14726
rect 2946 14720 3262 14721
rect 0 14650 800 14680
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 1301 14650 1367 14653
rect 0 14648 1367 14650
rect 0 14592 1306 14648
rect 1362 14592 1367 14648
rect 0 14590 1367 14592
rect 0 14560 800 14590
rect 1301 14587 1367 14590
rect 5993 14650 6059 14653
rect 9254 14650 9260 14652
rect 5993 14648 9260 14650
rect 5993 14592 5998 14648
rect 6054 14592 9260 14648
rect 5993 14590 9260 14592
rect 5993 14587 6059 14590
rect 9254 14588 9260 14590
rect 9324 14588 9330 14652
rect 13445 14650 13511 14653
rect 19609 14650 19675 14653
rect 13445 14648 19675 14650
rect 13445 14592 13450 14648
rect 13506 14592 19614 14648
rect 19670 14592 19675 14648
rect 13445 14590 19675 14592
rect 13445 14587 13511 14590
rect 19609 14587 19675 14590
rect 25497 14650 25563 14653
rect 28257 14650 28323 14653
rect 28717 14650 28783 14653
rect 25497 14648 28323 14650
rect 25497 14592 25502 14648
rect 25558 14592 28262 14648
rect 28318 14592 28323 14648
rect 25497 14590 28323 14592
rect 25497 14587 25563 14590
rect 28257 14587 28323 14590
rect 28398 14648 28783 14650
rect 28398 14592 28722 14648
rect 28778 14592 28783 14648
rect 28398 14590 28783 14592
rect 3969 14514 4035 14517
rect 21909 14514 21975 14517
rect 3969 14512 21975 14514
rect 3969 14456 3974 14512
rect 4030 14456 21914 14512
rect 21970 14456 21975 14512
rect 3969 14454 21975 14456
rect 3969 14451 4035 14454
rect 21909 14451 21975 14454
rect 22093 14514 22159 14517
rect 22921 14514 22987 14517
rect 22093 14512 22987 14514
rect 22093 14456 22098 14512
rect 22154 14456 22926 14512
rect 22982 14456 22987 14512
rect 22093 14454 22987 14456
rect 22093 14451 22159 14454
rect 22921 14451 22987 14454
rect 24945 14514 25011 14517
rect 27705 14514 27771 14517
rect 24945 14512 27771 14514
rect 24945 14456 24950 14512
rect 25006 14456 27710 14512
rect 27766 14456 27771 14512
rect 24945 14454 27771 14456
rect 24945 14451 25011 14454
rect 27705 14451 27771 14454
rect 6310 14316 6316 14380
rect 6380 14378 6386 14380
rect 13445 14378 13511 14381
rect 6380 14376 13511 14378
rect 6380 14320 13450 14376
rect 13506 14320 13511 14376
rect 6380 14318 13511 14320
rect 6380 14316 6386 14318
rect 13445 14315 13511 14318
rect 13721 14378 13787 14381
rect 21081 14378 21147 14381
rect 13721 14376 21147 14378
rect 13721 14320 13726 14376
rect 13782 14320 21086 14376
rect 21142 14320 21147 14376
rect 13721 14318 21147 14320
rect 13721 14315 13787 14318
rect 21081 14315 21147 14318
rect 23381 14378 23447 14381
rect 28398 14378 28458 14590
rect 28717 14587 28783 14590
rect 29821 14650 29887 14653
rect 32765 14650 32831 14653
rect 29821 14648 32831 14650
rect 29821 14592 29826 14648
rect 29882 14592 32770 14648
rect 32826 14592 32831 14648
rect 29821 14590 32831 14592
rect 29821 14587 29887 14590
rect 32765 14587 32831 14590
rect 38285 14650 38351 14653
rect 42793 14650 42859 14653
rect 38285 14648 42859 14650
rect 38285 14592 38290 14648
rect 38346 14592 42798 14648
rect 42854 14592 42859 14648
rect 38285 14590 42859 14592
rect 38285 14587 38351 14590
rect 42793 14587 42859 14590
rect 31518 14452 31524 14516
rect 31588 14514 31594 14516
rect 39297 14514 39363 14517
rect 31588 14512 39363 14514
rect 31588 14456 39302 14512
rect 39358 14456 39363 14512
rect 31588 14454 39363 14456
rect 31588 14452 31594 14454
rect 39297 14451 39363 14454
rect 39757 14514 39823 14517
rect 43161 14514 43227 14517
rect 39757 14512 43227 14514
rect 39757 14456 39762 14512
rect 39818 14456 43166 14512
rect 43222 14456 43227 14512
rect 39757 14454 43227 14456
rect 39757 14451 39823 14454
rect 43161 14451 43227 14454
rect 49693 14514 49759 14517
rect 50200 14514 51000 14544
rect 49693 14512 51000 14514
rect 49693 14456 49698 14512
rect 49754 14456 51000 14512
rect 49693 14454 51000 14456
rect 49693 14451 49759 14454
rect 50200 14424 51000 14454
rect 23381 14376 28458 14378
rect 23381 14320 23386 14376
rect 23442 14320 28458 14376
rect 23381 14318 28458 14320
rect 30005 14378 30071 14381
rect 40125 14378 40191 14381
rect 30005 14376 40191 14378
rect 30005 14320 30010 14376
rect 30066 14320 40130 14376
rect 40186 14320 40191 14376
rect 30005 14318 40191 14320
rect 23381 14315 23447 14318
rect 30005 14315 30071 14318
rect 40125 14315 40191 14318
rect 0 14242 800 14272
rect 933 14242 999 14245
rect 0 14240 999 14242
rect 0 14184 938 14240
rect 994 14184 999 14240
rect 0 14182 999 14184
rect 0 14152 800 14182
rect 933 14179 999 14182
rect 11053 14242 11119 14245
rect 13445 14242 13511 14245
rect 11053 14240 13511 14242
rect 11053 14184 11058 14240
rect 11114 14184 13450 14240
rect 13506 14184 13511 14240
rect 11053 14182 13511 14184
rect 11053 14179 11119 14182
rect 13445 14179 13511 14182
rect 13629 14242 13695 14245
rect 13854 14242 13860 14244
rect 13629 14240 13860 14242
rect 13629 14184 13634 14240
rect 13690 14184 13860 14240
rect 13629 14182 13860 14184
rect 13629 14179 13695 14182
rect 13854 14180 13860 14182
rect 13924 14242 13930 14244
rect 15009 14242 15075 14245
rect 13924 14240 15075 14242
rect 13924 14184 15014 14240
rect 15070 14184 15075 14240
rect 13924 14182 15075 14184
rect 13924 14180 13930 14182
rect 15009 14179 15075 14182
rect 20529 14242 20595 14245
rect 21817 14242 21883 14245
rect 20529 14240 21883 14242
rect 20529 14184 20534 14240
rect 20590 14184 21822 14240
rect 21878 14184 21883 14240
rect 20529 14182 21883 14184
rect 20529 14179 20595 14182
rect 21817 14179 21883 14182
rect 29085 14242 29151 14245
rect 31569 14242 31635 14245
rect 29085 14240 31635 14242
rect 29085 14184 29090 14240
rect 29146 14184 31574 14240
rect 31630 14184 31635 14240
rect 29085 14182 31635 14184
rect 29085 14179 29151 14182
rect 31569 14179 31635 14182
rect 38326 14180 38332 14244
rect 38396 14242 38402 14244
rect 47761 14242 47827 14245
rect 38396 14240 47827 14242
rect 38396 14184 47766 14240
rect 47822 14184 47827 14240
rect 38396 14182 47827 14184
rect 38396 14180 38402 14182
rect 47761 14179 47827 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 11237 14106 11303 14109
rect 18505 14106 18571 14109
rect 11237 14104 17832 14106
rect 11237 14048 11242 14104
rect 11298 14048 17832 14104
rect 11237 14046 17832 14048
rect 11237 14043 11303 14046
rect 6361 13970 6427 13973
rect 17217 13970 17283 13973
rect 6361 13968 17283 13970
rect 6361 13912 6366 13968
rect 6422 13912 17222 13968
rect 17278 13912 17283 13968
rect 6361 13910 17283 13912
rect 17772 13970 17832 14046
rect 18505 14104 26986 14106
rect 18505 14048 18510 14104
rect 18566 14048 26986 14104
rect 18505 14046 26986 14048
rect 18505 14043 18571 14046
rect 19241 13970 19307 13973
rect 17772 13968 19307 13970
rect 17772 13912 19246 13968
rect 19302 13912 19307 13968
rect 17772 13910 19307 13912
rect 6361 13907 6427 13910
rect 17217 13907 17283 13910
rect 19241 13907 19307 13910
rect 20069 13970 20135 13973
rect 23841 13970 23907 13973
rect 20069 13968 23907 13970
rect 20069 13912 20074 13968
rect 20130 13912 23846 13968
rect 23902 13912 23907 13968
rect 20069 13910 23907 13912
rect 26926 13970 26986 14046
rect 28942 14044 28948 14108
rect 29012 14106 29018 14108
rect 35341 14106 35407 14109
rect 29012 14104 35407 14106
rect 29012 14048 35346 14104
rect 35402 14048 35407 14104
rect 29012 14046 35407 14048
rect 29012 14044 29018 14046
rect 35341 14043 35407 14046
rect 40718 14044 40724 14108
rect 40788 14106 40794 14108
rect 42793 14106 42859 14109
rect 40788 14104 42859 14106
rect 40788 14048 42798 14104
rect 42854 14048 42859 14104
rect 40788 14046 42859 14048
rect 40788 14044 40794 14046
rect 42793 14043 42859 14046
rect 49182 14044 49188 14108
rect 49252 14106 49258 14108
rect 50200 14106 51000 14136
rect 49252 14046 51000 14106
rect 49252 14044 49258 14046
rect 33542 13970 33548 13972
rect 26926 13910 33548 13970
rect 20069 13907 20135 13910
rect 23841 13907 23907 13910
rect 33542 13908 33548 13910
rect 33612 13970 33618 13972
rect 33777 13970 33843 13973
rect 33612 13968 33843 13970
rect 33612 13912 33782 13968
rect 33838 13912 33843 13968
rect 33612 13910 33843 13912
rect 33612 13908 33618 13910
rect 33777 13907 33843 13910
rect 36261 13970 36327 13973
rect 39573 13970 39639 13973
rect 36261 13968 39639 13970
rect 36261 13912 36266 13968
rect 36322 13912 39578 13968
rect 39634 13912 39639 13968
rect 36261 13910 39639 13912
rect 36261 13907 36327 13910
rect 39573 13907 39639 13910
rect 40585 13970 40651 13973
rect 41321 13970 41387 13973
rect 42701 13970 42767 13973
rect 40585 13968 42767 13970
rect 40585 13912 40590 13968
rect 40646 13912 41326 13968
rect 41382 13912 42706 13968
rect 42762 13912 42767 13968
rect 40585 13910 42767 13912
rect 40585 13907 40651 13910
rect 41321 13907 41387 13910
rect 42701 13907 42767 13910
rect 47301 13970 47367 13973
rect 49190 13970 49250 14044
rect 50200 14016 51000 14046
rect 47301 13968 49250 13970
rect 47301 13912 47306 13968
rect 47362 13912 49250 13968
rect 47301 13910 49250 13912
rect 47301 13907 47367 13910
rect 0 13834 800 13864
rect 2773 13834 2839 13837
rect 6361 13836 6427 13837
rect 0 13832 2839 13834
rect 0 13776 2778 13832
rect 2834 13776 2839 13832
rect 0 13774 2839 13776
rect 0 13744 800 13774
rect 2773 13771 2839 13774
rect 6310 13772 6316 13836
rect 6380 13834 6427 13836
rect 7005 13834 7071 13837
rect 22001 13834 22067 13837
rect 6380 13832 6472 13834
rect 6422 13776 6472 13832
rect 6380 13774 6472 13776
rect 7005 13832 22067 13834
rect 7005 13776 7010 13832
rect 7066 13776 22006 13832
rect 22062 13776 22067 13832
rect 7005 13774 22067 13776
rect 6380 13772 6427 13774
rect 6361 13771 6427 13772
rect 7005 13771 7071 13774
rect 22001 13771 22067 13774
rect 24894 13772 24900 13836
rect 24964 13834 24970 13836
rect 30373 13834 30439 13837
rect 24964 13832 30439 13834
rect 24964 13776 30378 13832
rect 30434 13776 30439 13832
rect 24964 13774 30439 13776
rect 24964 13772 24970 13774
rect 30373 13771 30439 13774
rect 31150 13772 31156 13836
rect 31220 13834 31226 13836
rect 33961 13834 34027 13837
rect 31220 13832 34027 13834
rect 31220 13776 33966 13832
rect 34022 13776 34027 13832
rect 31220 13774 34027 13776
rect 31220 13772 31226 13774
rect 33961 13771 34027 13774
rect 36077 13834 36143 13837
rect 38285 13834 38351 13837
rect 36077 13832 38351 13834
rect 36077 13776 36082 13832
rect 36138 13776 38290 13832
rect 38346 13776 38351 13832
rect 36077 13774 38351 13776
rect 36077 13771 36143 13774
rect 38285 13771 38351 13774
rect 44766 13772 44772 13836
rect 44836 13834 44842 13836
rect 45277 13834 45343 13837
rect 44836 13832 45343 13834
rect 44836 13776 45282 13832
rect 45338 13776 45343 13832
rect 44836 13774 45343 13776
rect 44836 13772 44842 13774
rect 45277 13771 45343 13774
rect 3417 13700 3483 13701
rect 3366 13636 3372 13700
rect 3436 13698 3483 13700
rect 5441 13698 5507 13701
rect 5574 13698 5580 13700
rect 3436 13696 3528 13698
rect 3478 13640 3528 13696
rect 3436 13638 3528 13640
rect 5441 13696 5580 13698
rect 5441 13640 5446 13696
rect 5502 13640 5580 13696
rect 5441 13638 5580 13640
rect 3436 13636 3483 13638
rect 3417 13635 3483 13636
rect 5441 13635 5507 13638
rect 5574 13636 5580 13638
rect 5644 13636 5650 13700
rect 9213 13698 9279 13701
rect 12341 13698 12407 13701
rect 9213 13696 12407 13698
rect 9213 13640 9218 13696
rect 9274 13640 12346 13696
rect 12402 13640 12407 13696
rect 9213 13638 12407 13640
rect 9213 13635 9279 13638
rect 12341 13635 12407 13638
rect 13486 13636 13492 13700
rect 13556 13698 13562 13700
rect 14089 13698 14155 13701
rect 13556 13696 14155 13698
rect 13556 13640 14094 13696
rect 14150 13640 14155 13696
rect 13556 13638 14155 13640
rect 13556 13636 13562 13638
rect 14089 13635 14155 13638
rect 20345 13698 20411 13701
rect 21541 13698 21607 13701
rect 20345 13696 21607 13698
rect 20345 13640 20350 13696
rect 20406 13640 21546 13696
rect 21602 13640 21607 13696
rect 20345 13638 21607 13640
rect 20345 13635 20411 13638
rect 21541 13635 21607 13638
rect 28901 13698 28967 13701
rect 29821 13698 29887 13701
rect 30465 13698 30531 13701
rect 28901 13696 30531 13698
rect 28901 13640 28906 13696
rect 28962 13640 29826 13696
rect 29882 13640 30470 13696
rect 30526 13640 30531 13696
rect 28901 13638 30531 13640
rect 28901 13635 28967 13638
rect 29821 13635 29887 13638
rect 30465 13635 30531 13638
rect 34421 13698 34487 13701
rect 38929 13698 38995 13701
rect 34421 13696 38995 13698
rect 34421 13640 34426 13696
rect 34482 13640 38934 13696
rect 38990 13640 38995 13696
rect 34421 13638 38995 13640
rect 34421 13635 34487 13638
rect 38929 13635 38995 13638
rect 41086 13636 41092 13700
rect 41156 13698 41162 13700
rect 41229 13698 41295 13701
rect 41156 13696 41295 13698
rect 41156 13640 41234 13696
rect 41290 13640 41295 13696
rect 41156 13638 41295 13640
rect 41156 13636 41162 13638
rect 41229 13635 41295 13638
rect 44817 13698 44883 13701
rect 50200 13698 51000 13728
rect 44817 13696 51000 13698
rect 44817 13640 44822 13696
rect 44878 13640 51000 13696
rect 44817 13638 51000 13640
rect 44817 13635 44883 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 50200 13608 51000 13638
rect 42946 13567 43262 13568
rect 4286 13500 4292 13564
rect 4356 13562 4362 13564
rect 11646 13562 11652 13564
rect 4356 13502 11652 13562
rect 4356 13500 4362 13502
rect 11646 13500 11652 13502
rect 11716 13500 11722 13564
rect 14089 13562 14155 13565
rect 15561 13562 15627 13565
rect 14089 13560 15627 13562
rect 14089 13504 14094 13560
rect 14150 13504 15566 13560
rect 15622 13504 15627 13560
rect 14089 13502 15627 13504
rect 14089 13499 14155 13502
rect 15561 13499 15627 13502
rect 34053 13562 34119 13565
rect 36169 13562 36235 13565
rect 34053 13560 36235 13562
rect 34053 13504 34058 13560
rect 34114 13504 36174 13560
rect 36230 13504 36235 13560
rect 34053 13502 36235 13504
rect 34053 13499 34119 13502
rect 36169 13499 36235 13502
rect 37365 13562 37431 13565
rect 42793 13562 42859 13565
rect 37365 13560 42859 13562
rect 37365 13504 37370 13560
rect 37426 13504 42798 13560
rect 42854 13504 42859 13560
rect 37365 13502 42859 13504
rect 37365 13499 37431 13502
rect 42793 13499 42859 13502
rect 43662 13500 43668 13564
rect 43732 13562 43738 13564
rect 45686 13562 45692 13564
rect 43732 13502 45692 13562
rect 43732 13500 43738 13502
rect 45686 13500 45692 13502
rect 45756 13500 45762 13564
rect 48313 13562 48379 13565
rect 48630 13562 48636 13564
rect 48313 13560 48636 13562
rect 48313 13504 48318 13560
rect 48374 13504 48636 13560
rect 48313 13502 48636 13504
rect 48313 13499 48379 13502
rect 48630 13500 48636 13502
rect 48700 13500 48706 13564
rect 0 13426 800 13456
rect 2865 13426 2931 13429
rect 8845 13426 8911 13429
rect 0 13424 2931 13426
rect 0 13368 2870 13424
rect 2926 13368 2931 13424
rect 0 13366 2931 13368
rect 0 13336 800 13366
rect 2865 13363 2931 13366
rect 3742 13424 8911 13426
rect 3742 13368 8850 13424
rect 8906 13368 8911 13424
rect 3742 13366 8911 13368
rect 1761 13290 1827 13293
rect 3742 13290 3802 13366
rect 8845 13363 8911 13366
rect 10409 13426 10475 13429
rect 13169 13426 13235 13429
rect 10409 13424 13235 13426
rect 10409 13368 10414 13424
rect 10470 13368 13174 13424
rect 13230 13368 13235 13424
rect 10409 13366 13235 13368
rect 10409 13363 10475 13366
rect 13169 13363 13235 13366
rect 15561 13426 15627 13429
rect 24301 13426 24367 13429
rect 15561 13424 24367 13426
rect 15561 13368 15566 13424
rect 15622 13368 24306 13424
rect 24362 13368 24367 13424
rect 15561 13366 24367 13368
rect 15561 13363 15627 13366
rect 24301 13363 24367 13366
rect 32857 13426 32923 13429
rect 40493 13426 40559 13429
rect 32857 13424 40559 13426
rect 32857 13368 32862 13424
rect 32918 13368 40498 13424
rect 40554 13368 40559 13424
rect 32857 13366 40559 13368
rect 32857 13363 32923 13366
rect 40493 13363 40559 13366
rect 43662 13364 43668 13428
rect 43732 13426 43738 13428
rect 43989 13426 44055 13429
rect 43732 13424 44055 13426
rect 43732 13368 43994 13424
rect 44050 13368 44055 13424
rect 43732 13366 44055 13368
rect 43732 13364 43738 13366
rect 43989 13363 44055 13366
rect 47485 13426 47551 13429
rect 47710 13426 47716 13428
rect 47485 13424 47716 13426
rect 47485 13368 47490 13424
rect 47546 13368 47716 13424
rect 47485 13366 47716 13368
rect 47485 13363 47551 13366
rect 47710 13364 47716 13366
rect 47780 13426 47786 13428
rect 48773 13426 48839 13429
rect 47780 13424 48839 13426
rect 47780 13368 48778 13424
rect 48834 13368 48839 13424
rect 47780 13366 48839 13368
rect 47780 13364 47786 13366
rect 48773 13363 48839 13366
rect 1761 13288 3802 13290
rect 1761 13232 1766 13288
rect 1822 13232 3802 13288
rect 1761 13230 3802 13232
rect 3969 13290 4035 13293
rect 3969 13288 12450 13290
rect 3969 13232 3974 13288
rect 4030 13232 12450 13288
rect 3969 13230 12450 13232
rect 1761 13227 1827 13230
rect 3969 13227 4035 13230
rect 10501 13154 10567 13157
rect 11973 13154 12039 13157
rect 10501 13152 12039 13154
rect 10501 13096 10506 13152
rect 10562 13096 11978 13152
rect 12034 13096 12039 13152
rect 10501 13094 12039 13096
rect 12390 13154 12450 13230
rect 16246 13228 16252 13292
rect 16316 13290 16322 13292
rect 23013 13290 23079 13293
rect 25313 13290 25379 13293
rect 16316 13288 25379 13290
rect 16316 13232 23018 13288
rect 23074 13232 25318 13288
rect 25374 13232 25379 13288
rect 16316 13230 25379 13232
rect 16316 13228 16322 13230
rect 23013 13227 23079 13230
rect 25313 13227 25379 13230
rect 34881 13290 34947 13293
rect 35014 13290 35020 13292
rect 34881 13288 35020 13290
rect 34881 13232 34886 13288
rect 34942 13232 35020 13288
rect 34881 13230 35020 13232
rect 34881 13227 34947 13230
rect 35014 13228 35020 13230
rect 35084 13228 35090 13292
rect 40585 13290 40651 13293
rect 37782 13288 40651 13290
rect 37782 13232 40590 13288
rect 40646 13232 40651 13288
rect 37782 13230 40651 13232
rect 15142 13154 15148 13156
rect 12390 13094 15148 13154
rect 10501 13091 10567 13094
rect 11973 13091 12039 13094
rect 15142 13092 15148 13094
rect 15212 13092 15218 13156
rect 23473 13154 23539 13157
rect 22050 13152 23539 13154
rect 22050 13096 23478 13152
rect 23534 13096 23539 13152
rect 22050 13094 23539 13096
rect 7946 13088 8262 13089
rect 0 13018 800 13048
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 1301 13018 1367 13021
rect 3877 13020 3943 13021
rect 3877 13018 3924 13020
rect 0 13016 1367 13018
rect 0 12960 1306 13016
rect 1362 12960 1367 13016
rect 0 12958 1367 12960
rect 3832 13016 3924 13018
rect 3832 12960 3882 13016
rect 3832 12958 3924 12960
rect 0 12928 800 12958
rect 1301 12955 1367 12958
rect 3877 12956 3924 12958
rect 3988 12956 3994 13020
rect 11605 13018 11671 13021
rect 16246 13018 16252 13020
rect 11605 13016 16252 13018
rect 11605 12960 11610 13016
rect 11666 12960 16252 13016
rect 11605 12958 16252 12960
rect 3877 12955 3943 12956
rect 11605 12955 11671 12958
rect 16246 12956 16252 12958
rect 16316 12956 16322 13020
rect 21541 13018 21607 13021
rect 22050 13018 22110 13094
rect 23473 13091 23539 13094
rect 31017 13154 31083 13157
rect 37782 13154 37842 13230
rect 40585 13227 40651 13230
rect 42057 13290 42123 13293
rect 46422 13290 46428 13292
rect 42057 13288 46428 13290
rect 42057 13232 42062 13288
rect 42118 13232 46428 13288
rect 42057 13230 46428 13232
rect 42057 13227 42123 13230
rect 46422 13228 46428 13230
rect 46492 13228 46498 13292
rect 49141 13290 49207 13293
rect 50200 13290 51000 13320
rect 49141 13288 51000 13290
rect 49141 13232 49146 13288
rect 49202 13232 51000 13288
rect 49141 13230 51000 13232
rect 49141 13227 49207 13230
rect 50200 13200 51000 13230
rect 31017 13152 37842 13154
rect 31017 13096 31022 13152
rect 31078 13096 37842 13152
rect 31017 13094 37842 13096
rect 31017 13091 31083 13094
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 21541 13016 22110 13018
rect 21541 12960 21546 13016
rect 21602 12960 22110 13016
rect 21541 12958 22110 12960
rect 22737 13018 22803 13021
rect 22737 13016 27538 13018
rect 22737 12960 22742 13016
rect 22798 12960 27538 13016
rect 22737 12958 27538 12960
rect 21541 12955 21607 12958
rect 22737 12955 22803 12958
rect 3049 12882 3115 12885
rect 3550 12882 3556 12884
rect 3049 12880 3556 12882
rect 3049 12824 3054 12880
rect 3110 12824 3556 12880
rect 3049 12822 3556 12824
rect 3049 12819 3115 12822
rect 3550 12820 3556 12822
rect 3620 12882 3626 12884
rect 13261 12882 13327 12885
rect 3620 12880 13327 12882
rect 3620 12824 13266 12880
rect 13322 12824 13327 12880
rect 3620 12822 13327 12824
rect 3620 12820 3626 12822
rect 13261 12819 13327 12822
rect 13445 12882 13511 12885
rect 27245 12882 27311 12885
rect 13445 12880 27311 12882
rect 13445 12824 13450 12880
rect 13506 12824 27250 12880
rect 27306 12824 27311 12880
rect 13445 12822 27311 12824
rect 27478 12882 27538 12958
rect 32213 12882 32279 12885
rect 39297 12882 39363 12885
rect 27478 12822 31770 12882
rect 13445 12819 13511 12822
rect 27245 12819 27311 12822
rect 3969 12746 4035 12749
rect 2454 12744 4035 12746
rect 2454 12688 3974 12744
rect 4030 12688 4035 12744
rect 2454 12686 4035 12688
rect 0 12610 800 12640
rect 2454 12610 2514 12686
rect 3969 12683 4035 12686
rect 9070 12684 9076 12748
rect 9140 12746 9146 12748
rect 9305 12746 9371 12749
rect 9140 12744 11346 12746
rect 9140 12688 9310 12744
rect 9366 12688 11346 12744
rect 9140 12686 11346 12688
rect 9140 12684 9146 12686
rect 9305 12683 9371 12686
rect 0 12550 2514 12610
rect 0 12520 800 12550
rect 4286 12548 4292 12612
rect 4356 12610 4362 12612
rect 4705 12610 4771 12613
rect 4356 12608 4771 12610
rect 4356 12552 4710 12608
rect 4766 12552 4771 12608
rect 4356 12550 4771 12552
rect 4356 12548 4362 12550
rect 4705 12547 4771 12550
rect 9121 12610 9187 12613
rect 11053 12610 11119 12613
rect 9121 12608 11119 12610
rect 9121 12552 9126 12608
rect 9182 12552 11058 12608
rect 11114 12552 11119 12608
rect 9121 12550 11119 12552
rect 11286 12610 11346 12686
rect 11646 12684 11652 12748
rect 11716 12746 11722 12748
rect 19333 12746 19399 12749
rect 11716 12744 19399 12746
rect 11716 12688 19338 12744
rect 19394 12688 19399 12744
rect 11716 12686 19399 12688
rect 31710 12746 31770 12822
rect 32213 12880 39363 12882
rect 32213 12824 32218 12880
rect 32274 12824 39302 12880
rect 39358 12824 39363 12880
rect 32213 12822 39363 12824
rect 32213 12819 32279 12822
rect 39297 12819 39363 12822
rect 42701 12882 42767 12885
rect 47577 12882 47643 12885
rect 42701 12880 47643 12882
rect 42701 12824 42706 12880
rect 42762 12824 47582 12880
rect 47638 12824 47643 12880
rect 42701 12822 47643 12824
rect 42701 12819 42767 12822
rect 47577 12819 47643 12822
rect 49141 12882 49207 12885
rect 50200 12882 51000 12912
rect 49141 12880 51000 12882
rect 49141 12824 49146 12880
rect 49202 12824 51000 12880
rect 49141 12822 51000 12824
rect 49141 12819 49207 12822
rect 50200 12792 51000 12822
rect 46289 12746 46355 12749
rect 31710 12744 46355 12746
rect 31710 12688 46294 12744
rect 46350 12688 46355 12744
rect 31710 12686 46355 12688
rect 11716 12684 11722 12686
rect 19333 12683 19399 12686
rect 46289 12683 46355 12686
rect 12433 12610 12499 12613
rect 11286 12608 12499 12610
rect 11286 12552 12438 12608
rect 12494 12552 12499 12608
rect 11286 12550 12499 12552
rect 9121 12547 9187 12550
rect 11053 12547 11119 12550
rect 12433 12547 12499 12550
rect 13537 12608 13603 12613
rect 13537 12552 13542 12608
rect 13598 12552 13603 12608
rect 13537 12547 13603 12552
rect 33961 12610 34027 12613
rect 38377 12610 38443 12613
rect 33961 12608 38443 12610
rect 33961 12552 33966 12608
rect 34022 12552 38382 12608
rect 38438 12552 38443 12608
rect 33961 12550 38443 12552
rect 33961 12547 34027 12550
rect 38377 12547 38443 12550
rect 39573 12608 39639 12613
rect 39573 12552 39578 12608
rect 39634 12552 39639 12608
rect 39573 12547 39639 12552
rect 43478 12548 43484 12612
rect 43548 12610 43554 12612
rect 43621 12610 43687 12613
rect 43548 12608 43687 12610
rect 43548 12552 43626 12608
rect 43682 12552 43687 12608
rect 43548 12550 43687 12552
rect 43548 12548 43554 12550
rect 43621 12547 43687 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 6177 12474 6243 12477
rect 6545 12474 6611 12477
rect 6177 12472 6611 12474
rect 6177 12416 6182 12472
rect 6238 12416 6550 12472
rect 6606 12416 6611 12472
rect 6177 12414 6611 12416
rect 6177 12411 6243 12414
rect 6545 12411 6611 12414
rect 11237 12474 11303 12477
rect 12617 12474 12683 12477
rect 11237 12472 12683 12474
rect 11237 12416 11242 12472
rect 11298 12416 12622 12472
rect 12678 12416 12683 12472
rect 11237 12414 12683 12416
rect 13540 12474 13600 12547
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 13670 12474 13676 12476
rect 13540 12414 13676 12474
rect 11237 12411 11303 12414
rect 12617 12411 12683 12414
rect 13670 12412 13676 12414
rect 13740 12474 13746 12476
rect 16113 12474 16179 12477
rect 29361 12474 29427 12477
rect 13740 12472 16179 12474
rect 13740 12416 16118 12472
rect 16174 12416 16179 12472
rect 13740 12414 16179 12416
rect 13740 12412 13746 12414
rect 16113 12411 16179 12414
rect 29318 12472 29427 12474
rect 29318 12416 29366 12472
rect 29422 12416 29427 12472
rect 29318 12411 29427 12416
rect 36169 12474 36235 12477
rect 39576 12474 39636 12547
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 36169 12472 39636 12474
rect 36169 12416 36174 12472
rect 36230 12416 39636 12472
rect 36169 12414 39636 12416
rect 49141 12474 49207 12477
rect 50200 12474 51000 12504
rect 49141 12472 51000 12474
rect 49141 12416 49146 12472
rect 49202 12416 51000 12472
rect 49141 12414 51000 12416
rect 36169 12411 36235 12414
rect 49141 12411 49207 12414
rect 3417 12338 3483 12341
rect 9806 12338 9812 12340
rect 3417 12336 9812 12338
rect 3417 12280 3422 12336
rect 3478 12280 9812 12336
rect 3417 12278 9812 12280
rect 3417 12275 3483 12278
rect 9806 12276 9812 12278
rect 9876 12276 9882 12340
rect 10225 12338 10291 12341
rect 26918 12338 26924 12340
rect 10225 12336 26924 12338
rect 10225 12280 10230 12336
rect 10286 12280 26924 12336
rect 10225 12278 26924 12280
rect 10225 12275 10291 12278
rect 26918 12276 26924 12278
rect 26988 12276 26994 12340
rect 28993 12338 29059 12341
rect 29318 12338 29378 12411
rect 50200 12384 51000 12414
rect 28993 12336 29378 12338
rect 28993 12280 28998 12336
rect 29054 12280 29378 12336
rect 28993 12278 29378 12280
rect 29821 12338 29887 12341
rect 29821 12336 34714 12338
rect 29821 12280 29826 12336
rect 29882 12280 34714 12336
rect 29821 12278 34714 12280
rect 28993 12275 29059 12278
rect 29821 12275 29887 12278
rect 0 12202 800 12232
rect 1301 12202 1367 12205
rect 0 12200 1367 12202
rect 0 12144 1306 12200
rect 1362 12144 1367 12200
rect 0 12142 1367 12144
rect 0 12112 800 12142
rect 1301 12139 1367 12142
rect 6729 12202 6795 12205
rect 15193 12202 15259 12205
rect 6729 12200 15259 12202
rect 6729 12144 6734 12200
rect 6790 12144 15198 12200
rect 15254 12144 15259 12200
rect 6729 12142 15259 12144
rect 6729 12139 6795 12142
rect 15193 12139 15259 12142
rect 16430 12140 16436 12204
rect 16500 12202 16506 12204
rect 20161 12202 20227 12205
rect 16500 12200 20227 12202
rect 16500 12144 20166 12200
rect 20222 12144 20227 12200
rect 16500 12142 20227 12144
rect 16500 12140 16506 12142
rect 20161 12139 20227 12142
rect 26601 12202 26667 12205
rect 30557 12202 30623 12205
rect 34513 12202 34579 12205
rect 26601 12200 29010 12202
rect 26601 12144 26606 12200
rect 26662 12144 29010 12200
rect 26601 12142 29010 12144
rect 26601 12139 26667 12142
rect 9857 12066 9923 12069
rect 11789 12066 11855 12069
rect 9857 12064 11855 12066
rect 9857 12008 9862 12064
rect 9918 12008 11794 12064
rect 11850 12008 11855 12064
rect 9857 12006 11855 12008
rect 9857 12003 9923 12006
rect 11789 12003 11855 12006
rect 13629 12066 13695 12069
rect 13854 12066 13860 12068
rect 13629 12064 13860 12066
rect 13629 12008 13634 12064
rect 13690 12008 13860 12064
rect 13629 12006 13860 12008
rect 13629 12003 13695 12006
rect 13854 12004 13860 12006
rect 13924 12004 13930 12068
rect 14457 12066 14523 12069
rect 14641 12066 14707 12069
rect 14457 12064 14707 12066
rect 14457 12008 14462 12064
rect 14518 12008 14646 12064
rect 14702 12008 14707 12064
rect 14457 12006 14707 12008
rect 14457 12003 14523 12006
rect 14641 12003 14707 12006
rect 26734 12004 26740 12068
rect 26804 12066 26810 12068
rect 27102 12066 27108 12068
rect 26804 12006 27108 12066
rect 26804 12004 26810 12006
rect 27102 12004 27108 12006
rect 27172 12066 27178 12068
rect 27245 12066 27311 12069
rect 27172 12064 27311 12066
rect 27172 12008 27250 12064
rect 27306 12008 27311 12064
rect 27172 12006 27311 12008
rect 28950 12066 29010 12142
rect 30557 12200 34579 12202
rect 30557 12144 30562 12200
rect 30618 12144 34518 12200
rect 34574 12144 34579 12200
rect 30557 12142 34579 12144
rect 34654 12202 34714 12278
rect 35198 12276 35204 12340
rect 35268 12338 35274 12340
rect 36997 12338 37063 12341
rect 35268 12336 37063 12338
rect 35268 12280 37002 12336
rect 37058 12280 37063 12336
rect 35268 12278 37063 12280
rect 35268 12276 35274 12278
rect 36997 12275 37063 12278
rect 37222 12276 37228 12340
rect 37292 12338 37298 12340
rect 37733 12338 37799 12341
rect 38285 12340 38351 12341
rect 38285 12338 38332 12340
rect 37292 12336 37799 12338
rect 37292 12280 37738 12336
rect 37794 12280 37799 12336
rect 37292 12278 37799 12280
rect 38240 12336 38332 12338
rect 38240 12280 38290 12336
rect 38240 12278 38332 12280
rect 37292 12276 37298 12278
rect 37733 12275 37799 12278
rect 38285 12276 38332 12278
rect 38396 12276 38402 12340
rect 38469 12338 38535 12341
rect 46749 12338 46815 12341
rect 38469 12336 46815 12338
rect 38469 12280 38474 12336
rect 38530 12280 46754 12336
rect 46810 12280 46815 12336
rect 38469 12278 46815 12280
rect 38285 12275 38351 12276
rect 38469 12275 38535 12278
rect 46749 12275 46815 12278
rect 42057 12202 42123 12205
rect 34654 12200 42123 12202
rect 34654 12144 42062 12200
rect 42118 12144 42123 12200
rect 34654 12142 42123 12144
rect 30557 12139 30623 12142
rect 34513 12139 34579 12142
rect 42057 12139 42123 12142
rect 43529 12202 43595 12205
rect 44398 12202 44404 12204
rect 43529 12200 44404 12202
rect 43529 12144 43534 12200
rect 43590 12144 44404 12200
rect 43529 12142 44404 12144
rect 43529 12139 43595 12142
rect 44398 12140 44404 12142
rect 44468 12140 44474 12204
rect 30189 12066 30255 12069
rect 28950 12064 30255 12066
rect 28950 12008 30194 12064
rect 30250 12008 30255 12064
rect 28950 12006 30255 12008
rect 27172 12004 27178 12006
rect 27245 12003 27311 12006
rect 30189 12003 30255 12006
rect 33777 12066 33843 12069
rect 34278 12066 34284 12068
rect 33777 12064 34284 12066
rect 33777 12008 33782 12064
rect 33838 12008 34284 12064
rect 33777 12006 34284 12008
rect 33777 12003 33843 12006
rect 34278 12004 34284 12006
rect 34348 12004 34354 12068
rect 36169 12066 36235 12069
rect 36445 12066 36511 12069
rect 36169 12064 36511 12066
rect 36169 12008 36174 12064
rect 36230 12008 36450 12064
rect 36506 12008 36511 12064
rect 36169 12006 36511 12008
rect 36169 12003 36235 12006
rect 36445 12003 36511 12006
rect 38326 12004 38332 12068
rect 38396 12066 38402 12068
rect 40493 12066 40559 12069
rect 38396 12064 40559 12066
rect 38396 12008 40498 12064
rect 40554 12008 40559 12064
rect 38396 12006 40559 12008
rect 38396 12004 38402 12006
rect 40493 12003 40559 12006
rect 49141 12066 49207 12069
rect 50200 12066 51000 12096
rect 49141 12064 51000 12066
rect 49141 12008 49146 12064
rect 49202 12008 51000 12064
rect 49141 12006 51000 12008
rect 49141 12003 49207 12006
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 50200 11976 51000 12006
rect 47946 11935 48262 11936
rect 11697 11930 11763 11933
rect 12341 11930 12407 11933
rect 11697 11928 12407 11930
rect 11697 11872 11702 11928
rect 11758 11872 12346 11928
rect 12402 11872 12407 11928
rect 11697 11870 12407 11872
rect 11697 11867 11763 11870
rect 12341 11867 12407 11870
rect 20437 11930 20503 11933
rect 23933 11930 23999 11933
rect 20437 11928 23999 11930
rect 20437 11872 20442 11928
rect 20498 11872 23938 11928
rect 23994 11872 23999 11928
rect 20437 11870 23999 11872
rect 20437 11867 20503 11870
rect 23933 11867 23999 11870
rect 33685 11930 33751 11933
rect 37457 11930 37523 11933
rect 33685 11928 37523 11930
rect 33685 11872 33690 11928
rect 33746 11872 37462 11928
rect 37518 11872 37523 11928
rect 33685 11870 37523 11872
rect 33685 11867 33751 11870
rect 37457 11867 37523 11870
rect 39614 11868 39620 11932
rect 39684 11930 39690 11932
rect 44357 11930 44423 11933
rect 39684 11928 44423 11930
rect 39684 11872 44362 11928
rect 44418 11872 44423 11928
rect 39684 11870 44423 11872
rect 39684 11868 39690 11870
rect 44357 11867 44423 11870
rect 44541 11930 44607 11933
rect 44766 11930 44772 11932
rect 44541 11928 44772 11930
rect 44541 11872 44546 11928
rect 44602 11872 44772 11928
rect 44541 11870 44772 11872
rect 44541 11867 44607 11870
rect 44766 11868 44772 11870
rect 44836 11868 44842 11932
rect 46974 11868 46980 11932
rect 47044 11930 47050 11932
rect 47117 11930 47183 11933
rect 47044 11928 47183 11930
rect 47044 11872 47122 11928
rect 47178 11872 47183 11928
rect 47044 11870 47183 11872
rect 47044 11868 47050 11870
rect 47117 11867 47183 11870
rect 0 11794 800 11824
rect 4153 11794 4219 11797
rect 0 11792 4219 11794
rect 0 11736 4158 11792
rect 4214 11736 4219 11792
rect 0 11734 4219 11736
rect 0 11704 800 11734
rect 4153 11731 4219 11734
rect 5717 11796 5783 11797
rect 5717 11792 5764 11796
rect 5828 11794 5834 11796
rect 10777 11794 10843 11797
rect 13670 11794 13676 11796
rect 5717 11736 5722 11792
rect 5717 11732 5764 11736
rect 5828 11734 5874 11794
rect 10777 11792 13676 11794
rect 10777 11736 10782 11792
rect 10838 11736 13676 11792
rect 10777 11734 13676 11736
rect 5828 11732 5834 11734
rect 5717 11731 5783 11732
rect 10777 11731 10843 11734
rect 13670 11732 13676 11734
rect 13740 11732 13746 11796
rect 14365 11794 14431 11797
rect 14917 11794 14983 11797
rect 38694 11794 38700 11796
rect 14365 11792 38700 11794
rect 14365 11736 14370 11792
rect 14426 11736 14922 11792
rect 14978 11736 38700 11792
rect 14365 11734 38700 11736
rect 14365 11731 14431 11734
rect 14917 11731 14983 11734
rect 38694 11732 38700 11734
rect 38764 11732 38770 11796
rect 41822 11732 41828 11796
rect 41892 11794 41898 11796
rect 42425 11794 42491 11797
rect 41892 11792 42491 11794
rect 41892 11736 42430 11792
rect 42486 11736 42491 11792
rect 41892 11734 42491 11736
rect 41892 11732 41898 11734
rect 42425 11731 42491 11734
rect 44909 11796 44975 11797
rect 44909 11792 44956 11796
rect 45020 11794 45026 11796
rect 44909 11736 44914 11792
rect 44909 11732 44956 11736
rect 45020 11734 45066 11794
rect 45020 11732 45026 11734
rect 44909 11731 44975 11732
rect 5257 11658 5323 11661
rect 21725 11658 21791 11661
rect 5257 11656 21791 11658
rect 5257 11600 5262 11656
rect 5318 11600 21730 11656
rect 21786 11600 21791 11656
rect 5257 11598 21791 11600
rect 5257 11595 5323 11598
rect 21725 11595 21791 11598
rect 26049 11658 26115 11661
rect 28625 11658 28691 11661
rect 26049 11656 28691 11658
rect 26049 11600 26054 11656
rect 26110 11600 28630 11656
rect 28686 11600 28691 11656
rect 26049 11598 28691 11600
rect 26049 11595 26115 11598
rect 28625 11595 28691 11598
rect 32622 11596 32628 11660
rect 32692 11658 32698 11660
rect 44173 11658 44239 11661
rect 32692 11656 44239 11658
rect 32692 11600 44178 11656
rect 44234 11600 44239 11656
rect 32692 11598 44239 11600
rect 32692 11596 32698 11598
rect 44173 11595 44239 11598
rect 49141 11658 49207 11661
rect 50200 11658 51000 11688
rect 49141 11656 51000 11658
rect 49141 11600 49146 11656
rect 49202 11600 51000 11656
rect 49141 11598 51000 11600
rect 49141 11595 49207 11598
rect 50200 11568 51000 11598
rect 13905 11522 13971 11525
rect 15009 11522 15075 11525
rect 13905 11520 15075 11522
rect 13905 11464 13910 11520
rect 13966 11464 15014 11520
rect 15070 11464 15075 11520
rect 13905 11462 15075 11464
rect 13905 11459 13971 11462
rect 15009 11459 15075 11462
rect 15837 11522 15903 11525
rect 18454 11522 18460 11524
rect 15837 11520 18460 11522
rect 15837 11464 15842 11520
rect 15898 11464 18460 11520
rect 15837 11462 18460 11464
rect 15837 11459 15903 11462
rect 18454 11460 18460 11462
rect 18524 11522 18530 11524
rect 18781 11522 18847 11525
rect 18524 11520 18847 11522
rect 18524 11464 18786 11520
rect 18842 11464 18847 11520
rect 18524 11462 18847 11464
rect 18524 11460 18530 11462
rect 18781 11459 18847 11462
rect 27286 11460 27292 11524
rect 27356 11522 27362 11524
rect 32254 11522 32260 11524
rect 27356 11462 32260 11522
rect 27356 11460 27362 11462
rect 32254 11460 32260 11462
rect 32324 11460 32330 11524
rect 33961 11522 34027 11525
rect 34329 11522 34395 11525
rect 33961 11520 34395 11522
rect 33961 11464 33966 11520
rect 34022 11464 34334 11520
rect 34390 11464 34395 11520
rect 33961 11462 34395 11464
rect 33961 11459 34027 11462
rect 34329 11459 34395 11462
rect 35014 11460 35020 11524
rect 35084 11522 35090 11524
rect 39062 11522 39068 11524
rect 35084 11462 39068 11522
rect 35084 11460 35090 11462
rect 39062 11460 39068 11462
rect 39132 11460 39138 11524
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 3877 11386 3943 11389
rect 11789 11386 11855 11389
rect 0 11326 2790 11386
rect 0 11296 800 11326
rect 2730 11250 2790 11326
rect 3877 11384 11855 11386
rect 3877 11328 3882 11384
rect 3938 11328 11794 11384
rect 11850 11328 11855 11384
rect 3877 11326 11855 11328
rect 3877 11323 3943 11326
rect 11789 11323 11855 11326
rect 27286 11324 27292 11388
rect 27356 11386 27362 11388
rect 27613 11386 27679 11389
rect 29269 11386 29335 11389
rect 32765 11388 32831 11389
rect 32765 11386 32812 11388
rect 27356 11384 29335 11386
rect 27356 11328 27618 11384
rect 27674 11328 29274 11384
rect 29330 11328 29335 11384
rect 27356 11326 29335 11328
rect 32720 11384 32812 11386
rect 32720 11328 32770 11384
rect 32720 11326 32812 11328
rect 27356 11324 27362 11326
rect 27613 11323 27679 11326
rect 29269 11323 29335 11326
rect 32765 11324 32812 11326
rect 32876 11324 32882 11388
rect 33358 11324 33364 11388
rect 33428 11386 33434 11388
rect 37365 11386 37431 11389
rect 39113 11386 39179 11389
rect 33428 11326 37290 11386
rect 33428 11324 33434 11326
rect 32765 11323 32831 11324
rect 3417 11250 3483 11253
rect 2730 11248 3483 11250
rect 2730 11192 3422 11248
rect 3478 11192 3483 11248
rect 2730 11190 3483 11192
rect 3417 11187 3483 11190
rect 4613 11250 4679 11253
rect 16941 11250 17007 11253
rect 18597 11252 18663 11253
rect 18597 11250 18644 11252
rect 4613 11248 17007 11250
rect 4613 11192 4618 11248
rect 4674 11192 16946 11248
rect 17002 11192 17007 11248
rect 4613 11190 17007 11192
rect 18552 11248 18644 11250
rect 18552 11192 18602 11248
rect 18552 11190 18644 11192
rect 4613 11187 4679 11190
rect 16941 11187 17007 11190
rect 18597 11188 18644 11190
rect 18708 11188 18714 11252
rect 32438 11188 32444 11252
rect 32508 11250 32514 11252
rect 34462 11250 34468 11252
rect 32508 11190 34468 11250
rect 32508 11188 32514 11190
rect 34462 11188 34468 11190
rect 34532 11188 34538 11252
rect 35801 11250 35867 11253
rect 36077 11250 36143 11253
rect 35801 11248 36143 11250
rect 35801 11192 35806 11248
rect 35862 11192 36082 11248
rect 36138 11192 36143 11248
rect 35801 11190 36143 11192
rect 18597 11187 18663 11188
rect 35801 11187 35867 11190
rect 36077 11187 36143 11190
rect 7790 11054 8402 11114
rect 0 10978 800 11008
rect 1301 10978 1367 10981
rect 0 10976 1367 10978
rect 0 10920 1306 10976
rect 1362 10920 1367 10976
rect 0 10918 1367 10920
rect 0 10888 800 10918
rect 1301 10915 1367 10918
rect 5349 10978 5415 10981
rect 7790 10978 7850 11054
rect 5349 10976 7850 10978
rect 5349 10920 5354 10976
rect 5410 10920 7850 10976
rect 5349 10918 7850 10920
rect 8342 10978 8402 11054
rect 8886 11052 8892 11116
rect 8956 11114 8962 11116
rect 9622 11114 9628 11116
rect 8956 11054 9628 11114
rect 8956 11052 8962 11054
rect 9622 11052 9628 11054
rect 9692 11052 9698 11116
rect 11237 11114 11303 11117
rect 11513 11114 11579 11117
rect 11237 11112 11579 11114
rect 11237 11056 11242 11112
rect 11298 11056 11518 11112
rect 11574 11056 11579 11112
rect 11237 11054 11579 11056
rect 11237 11051 11303 11054
rect 11513 11051 11579 11054
rect 11789 11114 11855 11117
rect 15837 11114 15903 11117
rect 11789 11112 15903 11114
rect 11789 11056 11794 11112
rect 11850 11056 15842 11112
rect 15898 11056 15903 11112
rect 11789 11054 15903 11056
rect 11789 11051 11855 11054
rect 15837 11051 15903 11054
rect 16113 11114 16179 11117
rect 16246 11114 16252 11116
rect 16113 11112 16252 11114
rect 16113 11056 16118 11112
rect 16174 11056 16252 11112
rect 16113 11054 16252 11056
rect 16113 11051 16179 11054
rect 16246 11052 16252 11054
rect 16316 11052 16322 11116
rect 16481 11114 16547 11117
rect 19241 11114 19307 11117
rect 16481 11112 19307 11114
rect 16481 11056 16486 11112
rect 16542 11056 19246 11112
rect 19302 11056 19307 11112
rect 16481 11054 19307 11056
rect 16481 11051 16547 11054
rect 19241 11051 19307 11054
rect 20161 11114 20227 11117
rect 30465 11114 30531 11117
rect 33685 11114 33751 11117
rect 20161 11112 33751 11114
rect 20161 11056 20166 11112
rect 20222 11056 30470 11112
rect 30526 11056 33690 11112
rect 33746 11056 33751 11112
rect 20161 11054 33751 11056
rect 20161 11051 20227 11054
rect 30465 11051 30531 11054
rect 33685 11051 33751 11054
rect 34145 11114 34211 11117
rect 34278 11114 34284 11116
rect 34145 11112 34284 11114
rect 34145 11056 34150 11112
rect 34206 11056 34284 11112
rect 34145 11054 34284 11056
rect 34145 11051 34211 11054
rect 34278 11052 34284 11054
rect 34348 11052 34354 11116
rect 35249 11114 35315 11117
rect 36905 11114 36971 11117
rect 35249 11112 36971 11114
rect 35249 11056 35254 11112
rect 35310 11056 36910 11112
rect 36966 11056 36971 11112
rect 35249 11054 36971 11056
rect 37230 11114 37290 11326
rect 37365 11384 39179 11386
rect 37365 11328 37370 11384
rect 37426 11328 39118 11384
rect 39174 11328 39179 11384
rect 37365 11326 39179 11328
rect 37365 11323 37431 11326
rect 39113 11323 39179 11326
rect 39430 11324 39436 11388
rect 39500 11386 39506 11388
rect 42609 11386 42675 11389
rect 47393 11388 47459 11389
rect 39500 11384 42675 11386
rect 39500 11328 42614 11384
rect 42670 11328 42675 11384
rect 39500 11326 42675 11328
rect 39500 11324 39506 11326
rect 42609 11323 42675 11326
rect 47342 11324 47348 11388
rect 47412 11386 47459 11388
rect 47412 11384 47504 11386
rect 47454 11328 47504 11384
rect 47412 11326 47504 11328
rect 47412 11324 47459 11326
rect 47393 11323 47459 11324
rect 37457 11250 37523 11253
rect 39481 11250 39547 11253
rect 37457 11248 39547 11250
rect 37457 11192 37462 11248
rect 37518 11192 39486 11248
rect 39542 11192 39547 11248
rect 37457 11190 39547 11192
rect 37457 11187 37523 11190
rect 39481 11187 39547 11190
rect 40677 11250 40743 11253
rect 43253 11250 43319 11253
rect 43437 11252 43503 11253
rect 43437 11250 43484 11252
rect 40677 11248 43319 11250
rect 40677 11192 40682 11248
rect 40738 11192 43258 11248
rect 43314 11192 43319 11248
rect 40677 11190 43319 11192
rect 43392 11248 43484 11250
rect 43392 11192 43442 11248
rect 43392 11190 43484 11192
rect 40677 11187 40743 11190
rect 43253 11187 43319 11190
rect 43437 11188 43484 11190
rect 43548 11188 43554 11252
rect 49325 11250 49391 11253
rect 50200 11250 51000 11280
rect 49325 11248 51000 11250
rect 49325 11192 49330 11248
rect 49386 11192 51000 11248
rect 49325 11190 51000 11192
rect 43437 11187 43503 11188
rect 49325 11187 49391 11190
rect 50200 11160 51000 11190
rect 39982 11114 39988 11116
rect 37230 11054 39988 11114
rect 35249 11051 35315 11054
rect 36905 11051 36971 11054
rect 39982 11052 39988 11054
rect 40052 11114 40058 11116
rect 40953 11114 41019 11117
rect 40052 11112 41019 11114
rect 40052 11056 40958 11112
rect 41014 11056 41019 11112
rect 40052 11054 41019 11056
rect 40052 11052 40058 11054
rect 40953 11051 41019 11054
rect 43846 11052 43852 11116
rect 43916 11114 43922 11116
rect 44725 11114 44791 11117
rect 43916 11112 44791 11114
rect 43916 11056 44730 11112
rect 44786 11056 44791 11112
rect 43916 11054 44791 11056
rect 43916 11052 43922 11054
rect 44725 11051 44791 11054
rect 46105 11114 46171 11117
rect 46974 11114 46980 11116
rect 46105 11112 46980 11114
rect 46105 11056 46110 11112
rect 46166 11056 46980 11112
rect 46105 11054 46980 11056
rect 46105 11051 46171 11054
rect 46974 11052 46980 11054
rect 47044 11052 47050 11116
rect 17769 10978 17835 10981
rect 8342 10976 17835 10978
rect 8342 10920 17774 10976
rect 17830 10920 17835 10976
rect 8342 10918 17835 10920
rect 5349 10915 5415 10918
rect 17769 10915 17835 10918
rect 18505 10978 18571 10981
rect 18965 10978 19031 10981
rect 18505 10976 19031 10978
rect 18505 10920 18510 10976
rect 18566 10920 18970 10976
rect 19026 10920 19031 10976
rect 18505 10918 19031 10920
rect 18505 10915 18571 10918
rect 18965 10915 19031 10918
rect 19425 10978 19491 10981
rect 20345 10978 20411 10981
rect 19425 10976 20411 10978
rect 19425 10920 19430 10976
rect 19486 10920 20350 10976
rect 20406 10920 20411 10976
rect 19425 10918 20411 10920
rect 19425 10915 19491 10918
rect 20345 10915 20411 10918
rect 30966 10916 30972 10980
rect 31036 10978 31042 10980
rect 36721 10978 36787 10981
rect 37733 10978 37799 10981
rect 31036 10976 36787 10978
rect 31036 10920 36726 10976
rect 36782 10920 36787 10976
rect 31036 10918 36787 10920
rect 31036 10916 31042 10918
rect 36721 10915 36787 10918
rect 36862 10976 37799 10978
rect 36862 10920 37738 10976
rect 37794 10920 37799 10976
rect 36862 10918 37799 10920
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 11605 10842 11671 10845
rect 12709 10842 12775 10845
rect 11605 10840 12775 10842
rect 11605 10784 11610 10840
rect 11666 10784 12714 10840
rect 12770 10784 12775 10840
rect 11605 10782 12775 10784
rect 11605 10779 11671 10782
rect 12709 10779 12775 10782
rect 19425 10842 19491 10845
rect 21357 10842 21423 10845
rect 21541 10842 21607 10845
rect 36862 10842 36922 10918
rect 37733 10915 37799 10918
rect 38377 10978 38443 10981
rect 41597 10978 41663 10981
rect 41822 10978 41828 10980
rect 38377 10976 41828 10978
rect 38377 10920 38382 10976
rect 38438 10920 41602 10976
rect 41658 10920 41828 10976
rect 38377 10918 41828 10920
rect 38377 10915 38443 10918
rect 41597 10915 41663 10918
rect 41822 10916 41828 10918
rect 41892 10916 41898 10980
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 37089 10844 37155 10845
rect 42425 10844 42491 10845
rect 19425 10840 21607 10842
rect 19425 10784 19430 10840
rect 19486 10784 21362 10840
rect 21418 10784 21546 10840
rect 21602 10784 21607 10840
rect 19425 10782 21607 10784
rect 19425 10779 19491 10782
rect 21357 10779 21423 10782
rect 21541 10779 21607 10782
rect 28950 10782 36922 10842
rect 17585 10706 17651 10709
rect 2730 10704 17651 10706
rect 2730 10648 17590 10704
rect 17646 10648 17651 10704
rect 2730 10646 17651 10648
rect 0 10570 800 10600
rect 1209 10570 1275 10573
rect 0 10568 1275 10570
rect 0 10512 1214 10568
rect 1270 10512 1275 10568
rect 0 10510 1275 10512
rect 0 10480 800 10510
rect 1209 10507 1275 10510
rect 1761 10570 1827 10573
rect 2730 10570 2790 10646
rect 17585 10643 17651 10646
rect 17769 10706 17835 10709
rect 23381 10706 23447 10709
rect 17769 10704 23447 10706
rect 17769 10648 17774 10704
rect 17830 10648 23386 10704
rect 23442 10648 23447 10704
rect 17769 10646 23447 10648
rect 17769 10643 17835 10646
rect 23381 10643 23447 10646
rect 26417 10706 26483 10709
rect 28950 10706 29010 10782
rect 37038 10780 37044 10844
rect 37108 10842 37155 10844
rect 42374 10842 42380 10844
rect 37108 10840 37200 10842
rect 37150 10784 37200 10840
rect 37108 10782 37200 10784
rect 42334 10782 42380 10842
rect 42444 10840 42491 10844
rect 42486 10784 42491 10840
rect 37108 10780 37155 10782
rect 42374 10780 42380 10782
rect 42444 10780 42491 10784
rect 37089 10779 37155 10780
rect 42425 10779 42491 10780
rect 49141 10842 49207 10845
rect 50200 10842 51000 10872
rect 49141 10840 51000 10842
rect 49141 10784 49146 10840
rect 49202 10784 51000 10840
rect 49141 10782 51000 10784
rect 49141 10779 49207 10782
rect 50200 10752 51000 10782
rect 26417 10704 29010 10706
rect 26417 10648 26422 10704
rect 26478 10648 29010 10704
rect 26417 10646 29010 10648
rect 31109 10706 31175 10709
rect 46105 10706 46171 10709
rect 31109 10704 46171 10706
rect 31109 10648 31114 10704
rect 31170 10648 46110 10704
rect 46166 10648 46171 10704
rect 31109 10646 46171 10648
rect 26417 10643 26483 10646
rect 31109 10643 31175 10646
rect 46105 10643 46171 10646
rect 1761 10568 2790 10570
rect 1761 10512 1766 10568
rect 1822 10512 2790 10568
rect 1761 10510 2790 10512
rect 3693 10570 3759 10573
rect 13486 10570 13492 10572
rect 3693 10568 13492 10570
rect 3693 10512 3698 10568
rect 3754 10512 13492 10568
rect 3693 10510 13492 10512
rect 1761 10507 1827 10510
rect 3693 10507 3759 10510
rect 13486 10508 13492 10510
rect 13556 10508 13562 10572
rect 15837 10570 15903 10573
rect 19149 10570 19215 10573
rect 15837 10568 19215 10570
rect 15837 10512 15842 10568
rect 15898 10512 19154 10568
rect 19210 10512 19215 10568
rect 15837 10510 19215 10512
rect 15837 10507 15903 10510
rect 19149 10507 19215 10510
rect 22921 10570 22987 10573
rect 22921 10568 23490 10570
rect 22921 10512 22926 10568
rect 22982 10512 23490 10568
rect 22921 10510 23490 10512
rect 22921 10507 22987 10510
rect 8334 10372 8340 10436
rect 8404 10434 8410 10436
rect 9397 10434 9463 10437
rect 8404 10432 9463 10434
rect 8404 10376 9402 10432
rect 9458 10376 9463 10432
rect 8404 10374 9463 10376
rect 8404 10372 8410 10374
rect 9397 10371 9463 10374
rect 11881 10434 11947 10437
rect 12433 10434 12499 10437
rect 11881 10432 12499 10434
rect 11881 10376 11886 10432
rect 11942 10376 12438 10432
rect 12494 10376 12499 10432
rect 11881 10374 12499 10376
rect 11881 10371 11947 10374
rect 12433 10371 12499 10374
rect 15377 10434 15443 10437
rect 17493 10434 17559 10437
rect 15377 10432 17559 10434
rect 15377 10376 15382 10432
rect 15438 10376 17498 10432
rect 17554 10376 17559 10432
rect 15377 10374 17559 10376
rect 23430 10434 23490 10510
rect 25998 10508 26004 10572
rect 26068 10570 26074 10572
rect 46197 10570 46263 10573
rect 26068 10568 46263 10570
rect 26068 10512 46202 10568
rect 46258 10512 46263 10568
rect 26068 10510 46263 10512
rect 26068 10508 26074 10510
rect 46197 10507 46263 10510
rect 30557 10434 30623 10437
rect 23430 10432 30623 10434
rect 23430 10376 30562 10432
rect 30618 10376 30623 10432
rect 23430 10374 30623 10376
rect 15377 10371 15443 10374
rect 17493 10371 17559 10374
rect 30557 10371 30623 10374
rect 36537 10434 36603 10437
rect 37089 10434 37155 10437
rect 39849 10434 39915 10437
rect 36537 10432 39915 10434
rect 36537 10376 36542 10432
rect 36598 10376 37094 10432
rect 37150 10376 39854 10432
rect 39910 10376 39915 10432
rect 36537 10374 39915 10376
rect 36537 10371 36603 10374
rect 37089 10371 37155 10374
rect 39849 10371 39915 10374
rect 49417 10434 49483 10437
rect 50200 10434 51000 10464
rect 49417 10432 51000 10434
rect 49417 10376 49422 10432
rect 49478 10376 51000 10432
rect 49417 10374 51000 10376
rect 49417 10371 49483 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 50200 10344 51000 10374
rect 42946 10303 43262 10304
rect 5165 10300 5231 10301
rect 7373 10300 7439 10301
rect 5165 10298 5212 10300
rect 5120 10296 5212 10298
rect 5120 10240 5170 10296
rect 5120 10238 5212 10240
rect 5165 10236 5212 10238
rect 5276 10236 5282 10300
rect 7373 10298 7420 10300
rect 7328 10296 7420 10298
rect 7328 10240 7378 10296
rect 7328 10238 7420 10240
rect 7373 10236 7420 10238
rect 7484 10236 7490 10300
rect 9121 10298 9187 10301
rect 9438 10298 9444 10300
rect 9121 10296 9444 10298
rect 9121 10240 9126 10296
rect 9182 10240 9444 10296
rect 9121 10238 9444 10240
rect 5165 10235 5231 10236
rect 7373 10235 7439 10236
rect 9121 10235 9187 10238
rect 9438 10236 9444 10238
rect 9508 10236 9514 10300
rect 9857 10298 9923 10301
rect 12525 10298 12591 10301
rect 9857 10296 12591 10298
rect 9857 10240 9862 10296
rect 9918 10240 12530 10296
rect 12586 10240 12591 10296
rect 9857 10238 12591 10240
rect 9857 10235 9923 10238
rect 12525 10235 12591 10238
rect 16614 10236 16620 10300
rect 16684 10298 16690 10300
rect 19374 10298 19380 10300
rect 16684 10238 19380 10298
rect 16684 10236 16690 10238
rect 19374 10236 19380 10238
rect 19444 10236 19450 10300
rect 34513 10298 34579 10301
rect 40953 10298 41019 10301
rect 34513 10296 41019 10298
rect 34513 10240 34518 10296
rect 34574 10240 40958 10296
rect 41014 10240 41019 10296
rect 34513 10238 41019 10240
rect 34513 10235 34579 10238
rect 40953 10235 41019 10238
rect 0 10162 800 10192
rect 1301 10162 1367 10165
rect 0 10160 1367 10162
rect 0 10104 1306 10160
rect 1362 10104 1367 10160
rect 0 10102 1367 10104
rect 0 10072 800 10102
rect 1301 10099 1367 10102
rect 11605 10162 11671 10165
rect 13813 10162 13879 10165
rect 11605 10160 13879 10162
rect 11605 10104 11610 10160
rect 11666 10104 13818 10160
rect 13874 10104 13879 10160
rect 11605 10102 13879 10104
rect 11605 10099 11671 10102
rect 13813 10099 13879 10102
rect 17401 10162 17467 10165
rect 23381 10162 23447 10165
rect 24117 10162 24183 10165
rect 17401 10160 23306 10162
rect 17401 10104 17406 10160
rect 17462 10104 23306 10160
rect 17401 10102 23306 10104
rect 17401 10099 17467 10102
rect 6637 10026 6703 10029
rect 18137 10026 18203 10029
rect 6637 10024 18203 10026
rect 6637 9968 6642 10024
rect 6698 9968 18142 10024
rect 18198 9968 18203 10024
rect 6637 9966 18203 9968
rect 6637 9963 6703 9966
rect 18137 9963 18203 9966
rect 19149 10026 19215 10029
rect 23246 10026 23306 10102
rect 23381 10160 24183 10162
rect 23381 10104 23386 10160
rect 23442 10104 24122 10160
rect 24178 10104 24183 10160
rect 23381 10102 24183 10104
rect 23381 10099 23447 10102
rect 24117 10099 24183 10102
rect 25957 10162 26023 10165
rect 34329 10162 34395 10165
rect 25957 10160 34395 10162
rect 25957 10104 25962 10160
rect 26018 10104 34334 10160
rect 34390 10104 34395 10160
rect 25957 10102 34395 10104
rect 25957 10099 26023 10102
rect 34329 10099 34395 10102
rect 34462 10100 34468 10164
rect 34532 10162 34538 10164
rect 42609 10162 42675 10165
rect 34532 10160 42675 10162
rect 34532 10104 42614 10160
rect 42670 10104 42675 10160
rect 34532 10102 42675 10104
rect 34532 10100 34538 10102
rect 42609 10099 42675 10102
rect 43253 10162 43319 10165
rect 44214 10162 44220 10164
rect 43253 10160 44220 10162
rect 43253 10104 43258 10160
rect 43314 10104 44220 10160
rect 43253 10102 44220 10104
rect 43253 10099 43319 10102
rect 44214 10100 44220 10102
rect 44284 10100 44290 10164
rect 45553 10162 45619 10165
rect 46238 10162 46244 10164
rect 45553 10160 46244 10162
rect 45553 10104 45558 10160
rect 45614 10104 46244 10160
rect 45553 10102 46244 10104
rect 45553 10099 45619 10102
rect 46238 10100 46244 10102
rect 46308 10100 46314 10164
rect 27337 10026 27403 10029
rect 19149 10024 22110 10026
rect 19149 9968 19154 10024
rect 19210 9968 22110 10024
rect 19149 9966 22110 9968
rect 23246 10024 27403 10026
rect 23246 9968 27342 10024
rect 27398 9968 27403 10024
rect 23246 9966 27403 9968
rect 19149 9963 19215 9966
rect 8385 9890 8451 9893
rect 16062 9890 16068 9892
rect 8385 9888 16068 9890
rect 8385 9832 8390 9888
rect 8446 9832 16068 9888
rect 8385 9830 16068 9832
rect 8385 9827 8451 9830
rect 16062 9828 16068 9830
rect 16132 9828 16138 9892
rect 22050 9890 22110 9966
rect 27337 9963 27403 9966
rect 27797 10026 27863 10029
rect 39021 10026 39087 10029
rect 27797 10024 39087 10026
rect 27797 9968 27802 10024
rect 27858 9968 39026 10024
rect 39082 9968 39087 10024
rect 27797 9966 39087 9968
rect 27797 9963 27863 9966
rect 39021 9963 39087 9966
rect 49233 10026 49299 10029
rect 50200 10026 51000 10056
rect 49233 10024 51000 10026
rect 49233 9968 49238 10024
rect 49294 9968 51000 10024
rect 49233 9966 51000 9968
rect 49233 9963 49299 9966
rect 50200 9936 51000 9966
rect 22185 9890 22251 9893
rect 25957 9890 26023 9893
rect 22050 9888 26023 9890
rect 22050 9832 22190 9888
rect 22246 9832 25962 9888
rect 26018 9832 26023 9888
rect 22050 9830 26023 9832
rect 22185 9827 22251 9830
rect 25957 9827 26023 9830
rect 30373 9890 30439 9893
rect 33685 9890 33751 9893
rect 30373 9888 33751 9890
rect 30373 9832 30378 9888
rect 30434 9832 33690 9888
rect 33746 9832 33751 9888
rect 30373 9830 33751 9832
rect 30373 9827 30439 9830
rect 33685 9827 33751 9830
rect 36629 9890 36695 9893
rect 37457 9890 37523 9893
rect 36629 9888 37523 9890
rect 36629 9832 36634 9888
rect 36690 9832 37462 9888
rect 37518 9832 37523 9888
rect 36629 9830 37523 9832
rect 36629 9827 36695 9830
rect 37457 9827 37523 9830
rect 7946 9824 8262 9825
rect 0 9754 800 9784
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 1577 9754 1643 9757
rect 2865 9754 2931 9757
rect 12525 9754 12591 9757
rect 14038 9754 14044 9756
rect 0 9752 2931 9754
rect 0 9696 1582 9752
rect 1638 9696 2870 9752
rect 2926 9696 2931 9752
rect 0 9694 2931 9696
rect 0 9664 800 9694
rect 1577 9691 1643 9694
rect 2865 9691 2931 9694
rect 11838 9694 12266 9754
rect 7649 9620 7715 9621
rect 7598 9618 7604 9620
rect 7558 9558 7604 9618
rect 7668 9616 7715 9620
rect 7710 9560 7715 9616
rect 7598 9556 7604 9558
rect 7668 9556 7715 9560
rect 7649 9555 7715 9556
rect 9765 9618 9831 9621
rect 11838 9618 11898 9694
rect 12065 9620 12131 9621
rect 12014 9618 12020 9620
rect 9765 9616 11898 9618
rect 9765 9560 9770 9616
rect 9826 9560 11898 9616
rect 9765 9558 11898 9560
rect 11974 9558 12020 9618
rect 12084 9616 12131 9620
rect 12126 9560 12131 9616
rect 9765 9555 9831 9558
rect 12014 9556 12020 9558
rect 12084 9556 12131 9560
rect 12206 9618 12266 9694
rect 12525 9752 14044 9754
rect 12525 9696 12530 9752
rect 12586 9696 14044 9752
rect 12525 9694 14044 9696
rect 12525 9691 12591 9694
rect 14038 9692 14044 9694
rect 14108 9692 14114 9756
rect 16021 9754 16087 9757
rect 16982 9754 16988 9756
rect 16021 9752 16988 9754
rect 16021 9696 16026 9752
rect 16082 9696 16988 9752
rect 16021 9694 16988 9696
rect 16021 9691 16087 9694
rect 16982 9692 16988 9694
rect 17052 9692 17058 9756
rect 27286 9754 27292 9756
rect 23430 9694 27292 9754
rect 23430 9621 23490 9694
rect 27286 9692 27292 9694
rect 27356 9692 27362 9756
rect 30557 9754 30623 9757
rect 31201 9754 31267 9757
rect 30557 9752 31267 9754
rect 30557 9696 30562 9752
rect 30618 9696 31206 9752
rect 31262 9696 31267 9752
rect 30557 9694 31267 9696
rect 30557 9691 30623 9694
rect 31201 9691 31267 9694
rect 31753 9754 31819 9757
rect 32581 9754 32647 9757
rect 37273 9754 37339 9757
rect 31753 9752 37339 9754
rect 31753 9696 31758 9752
rect 31814 9696 32586 9752
rect 32642 9696 37278 9752
rect 37334 9696 37339 9752
rect 31753 9694 37339 9696
rect 31753 9691 31819 9694
rect 32581 9691 32647 9694
rect 37273 9691 37339 9694
rect 14549 9618 14615 9621
rect 20161 9618 20227 9621
rect 12206 9616 20227 9618
rect 12206 9560 14554 9616
rect 14610 9560 20166 9616
rect 20222 9560 20227 9616
rect 12206 9558 20227 9560
rect 12065 9555 12131 9556
rect 14549 9555 14615 9558
rect 20161 9555 20227 9558
rect 23381 9616 23490 9621
rect 23381 9560 23386 9616
rect 23442 9560 23490 9616
rect 23381 9558 23490 9560
rect 29177 9618 29243 9621
rect 29177 9616 32138 9618
rect 29177 9560 29182 9616
rect 29238 9560 32138 9616
rect 29177 9558 32138 9560
rect 23381 9555 23447 9558
rect 29177 9555 29243 9558
rect 1761 9482 1827 9485
rect 22921 9482 22987 9485
rect 1761 9480 22110 9482
rect 1761 9424 1766 9480
rect 1822 9424 22110 9480
rect 1761 9422 22110 9424
rect 1761 9419 1827 9422
rect 0 9346 800 9376
rect 1209 9346 1275 9349
rect 0 9344 1275 9346
rect 0 9288 1214 9344
rect 1270 9288 1275 9344
rect 0 9286 1275 9288
rect 0 9256 800 9286
rect 1209 9283 1275 9286
rect 5993 9346 6059 9349
rect 12566 9346 12572 9348
rect 5993 9344 12572 9346
rect 5993 9288 5998 9344
rect 6054 9288 12572 9344
rect 5993 9286 12572 9288
rect 5993 9283 6059 9286
rect 12566 9284 12572 9286
rect 12636 9284 12642 9348
rect 13353 9346 13419 9349
rect 17677 9346 17743 9349
rect 13353 9344 17743 9346
rect 13353 9288 13358 9344
rect 13414 9288 17682 9344
rect 17738 9288 17743 9344
rect 13353 9286 17743 9288
rect 13353 9283 13419 9286
rect 17677 9283 17743 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 18638 9148 18644 9212
rect 18708 9210 18714 9212
rect 19425 9210 19491 9213
rect 18708 9208 19491 9210
rect 18708 9152 19430 9208
rect 19486 9152 19491 9208
rect 18708 9150 19491 9152
rect 18708 9148 18714 9150
rect 19425 9147 19491 9150
rect 9622 9012 9628 9076
rect 9692 9074 9698 9076
rect 18689 9074 18755 9077
rect 9692 9072 18755 9074
rect 9692 9016 18694 9072
rect 18750 9016 18755 9072
rect 9692 9014 18755 9016
rect 22050 9074 22110 9422
rect 22510 9480 22987 9482
rect 22510 9424 22926 9480
rect 22982 9424 22987 9480
rect 22510 9422 22987 9424
rect 32078 9482 32138 9558
rect 34278 9556 34284 9620
rect 34348 9618 34354 9620
rect 38837 9618 38903 9621
rect 34348 9616 38903 9618
rect 34348 9560 38842 9616
rect 38898 9560 38903 9616
rect 34348 9558 38903 9560
rect 34348 9556 34354 9558
rect 38837 9555 38903 9558
rect 39062 9556 39068 9620
rect 39132 9618 39138 9620
rect 41413 9618 41479 9621
rect 39132 9616 41479 9618
rect 39132 9560 41418 9616
rect 41474 9560 41479 9616
rect 39132 9558 41479 9560
rect 39132 9556 39138 9558
rect 41413 9555 41479 9558
rect 42885 9618 42951 9621
rect 43662 9618 43668 9620
rect 42885 9616 43668 9618
rect 42885 9560 42890 9616
rect 42946 9560 43668 9616
rect 42885 9558 43668 9560
rect 42885 9555 42951 9558
rect 43662 9556 43668 9558
rect 43732 9556 43738 9620
rect 44030 9556 44036 9620
rect 44100 9618 44106 9620
rect 44173 9618 44239 9621
rect 44100 9616 44239 9618
rect 44100 9560 44178 9616
rect 44234 9560 44239 9616
rect 44100 9558 44239 9560
rect 44100 9556 44106 9558
rect 44173 9555 44239 9558
rect 46841 9618 46907 9621
rect 50200 9618 51000 9648
rect 46841 9616 51000 9618
rect 46841 9560 46846 9616
rect 46902 9560 51000 9616
rect 46841 9558 51000 9560
rect 46841 9555 46907 9558
rect 50200 9528 51000 9558
rect 35157 9482 35223 9485
rect 35525 9482 35591 9485
rect 32078 9480 35591 9482
rect 32078 9424 35162 9480
rect 35218 9424 35530 9480
rect 35586 9424 35591 9480
rect 32078 9422 35591 9424
rect 22369 9210 22435 9213
rect 22510 9210 22570 9422
rect 22921 9419 22987 9422
rect 35157 9419 35223 9422
rect 35525 9419 35591 9422
rect 35893 9482 35959 9485
rect 37181 9482 37247 9485
rect 35893 9480 37247 9482
rect 35893 9424 35898 9480
rect 35954 9424 37186 9480
rect 37242 9424 37247 9480
rect 35893 9422 37247 9424
rect 35893 9419 35959 9422
rect 37181 9419 37247 9422
rect 37825 9482 37891 9485
rect 38929 9482 38995 9485
rect 37825 9480 38995 9482
rect 37825 9424 37830 9480
rect 37886 9424 38934 9480
rect 38990 9424 38995 9480
rect 37825 9422 38995 9424
rect 37825 9419 37891 9422
rect 38929 9419 38995 9422
rect 39113 9482 39179 9485
rect 39849 9482 39915 9485
rect 45185 9482 45251 9485
rect 39113 9480 39915 9482
rect 39113 9424 39118 9480
rect 39174 9424 39854 9480
rect 39910 9424 39915 9480
rect 39113 9422 39915 9424
rect 39113 9419 39179 9422
rect 39849 9419 39915 9422
rect 41370 9480 45251 9482
rect 41370 9424 45190 9480
rect 45246 9424 45251 9480
rect 41370 9422 45251 9424
rect 34830 9284 34836 9348
rect 34900 9346 34906 9348
rect 41370 9346 41430 9422
rect 45185 9419 45251 9422
rect 34900 9286 41430 9346
rect 34900 9284 34906 9286
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 22369 9208 22570 9210
rect 22369 9152 22374 9208
rect 22430 9152 22570 9208
rect 22369 9150 22570 9152
rect 33777 9210 33843 9213
rect 37365 9210 37431 9213
rect 39573 9210 39639 9213
rect 33777 9208 39639 9210
rect 33777 9152 33782 9208
rect 33838 9152 37370 9208
rect 37426 9152 39578 9208
rect 39634 9152 39639 9208
rect 33777 9150 39639 9152
rect 22369 9147 22435 9150
rect 33777 9147 33843 9150
rect 37365 9147 37431 9150
rect 39573 9147 39639 9150
rect 49141 9210 49207 9213
rect 50200 9210 51000 9240
rect 49141 9208 51000 9210
rect 49141 9152 49146 9208
rect 49202 9152 51000 9208
rect 49141 9150 51000 9152
rect 49141 9147 49207 9150
rect 50200 9120 51000 9150
rect 36997 9074 37063 9077
rect 22050 9072 37063 9074
rect 22050 9016 37002 9072
rect 37058 9016 37063 9072
rect 22050 9014 37063 9016
rect 9692 9012 9698 9014
rect 18689 9011 18755 9014
rect 36997 9011 37063 9014
rect 37406 9012 37412 9076
rect 37476 9074 37482 9076
rect 46974 9074 46980 9076
rect 37476 9014 46980 9074
rect 37476 9012 37482 9014
rect 46974 9012 46980 9014
rect 47044 9012 47050 9076
rect 48313 9074 48379 9077
rect 48814 9074 48820 9076
rect 48313 9072 48820 9074
rect 48313 9016 48318 9072
rect 48374 9016 48820 9072
rect 48313 9014 48820 9016
rect 48313 9011 48379 9014
rect 48814 9012 48820 9014
rect 48884 9012 48890 9076
rect 0 8938 800 8968
rect 1301 8938 1367 8941
rect 0 8936 1367 8938
rect 0 8880 1306 8936
rect 1362 8880 1367 8936
rect 0 8878 1367 8880
rect 0 8848 800 8878
rect 1301 8875 1367 8878
rect 1761 8938 1827 8941
rect 23381 8938 23447 8941
rect 1761 8936 23447 8938
rect 1761 8880 1766 8936
rect 1822 8880 23386 8936
rect 23442 8880 23447 8936
rect 1761 8878 23447 8880
rect 1761 8875 1827 8878
rect 23381 8875 23447 8878
rect 32254 8876 32260 8940
rect 32324 8938 32330 8940
rect 35893 8938 35959 8941
rect 32324 8936 35959 8938
rect 32324 8880 35898 8936
rect 35954 8880 35959 8936
rect 32324 8878 35959 8880
rect 32324 8876 32330 8878
rect 35893 8875 35959 8878
rect 36721 8938 36787 8941
rect 38653 8938 38719 8941
rect 43529 8938 43595 8941
rect 36721 8936 38394 8938
rect 36721 8880 36726 8936
rect 36782 8880 38394 8936
rect 36721 8878 38394 8880
rect 36721 8875 36787 8878
rect 8477 8802 8543 8805
rect 17217 8802 17283 8805
rect 8477 8800 17283 8802
rect 8477 8744 8482 8800
rect 8538 8744 17222 8800
rect 17278 8744 17283 8800
rect 8477 8742 17283 8744
rect 8477 8739 8543 8742
rect 17217 8739 17283 8742
rect 18638 8740 18644 8804
rect 18708 8802 18714 8804
rect 18873 8802 18939 8805
rect 18708 8800 18939 8802
rect 18708 8744 18878 8800
rect 18934 8744 18939 8800
rect 18708 8742 18939 8744
rect 18708 8740 18714 8742
rect 18873 8739 18939 8742
rect 31017 8802 31083 8805
rect 37181 8802 37247 8805
rect 31017 8800 37247 8802
rect 31017 8744 31022 8800
rect 31078 8744 37186 8800
rect 37242 8744 37247 8800
rect 31017 8742 37247 8744
rect 31017 8739 31083 8742
rect 37181 8739 37247 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 15193 8666 15259 8669
rect 17350 8666 17356 8668
rect 15193 8664 17356 8666
rect 15193 8608 15198 8664
rect 15254 8608 17356 8664
rect 15193 8606 17356 8608
rect 15193 8603 15259 8606
rect 17350 8604 17356 8606
rect 17420 8604 17426 8668
rect 18413 8666 18479 8669
rect 24761 8666 24827 8669
rect 18413 8664 24827 8666
rect 18413 8608 18418 8664
rect 18474 8608 24766 8664
rect 24822 8608 24827 8664
rect 18413 8606 24827 8608
rect 38334 8666 38394 8878
rect 38653 8936 43595 8938
rect 38653 8880 38658 8936
rect 38714 8880 43534 8936
rect 43590 8880 43595 8936
rect 38653 8878 43595 8880
rect 38653 8875 38719 8878
rect 43529 8875 43595 8878
rect 38745 8804 38811 8805
rect 38694 8802 38700 8804
rect 38654 8742 38700 8802
rect 38764 8800 38811 8804
rect 38806 8744 38811 8800
rect 38694 8740 38700 8742
rect 38764 8740 38811 8744
rect 38745 8739 38811 8740
rect 41781 8802 41847 8805
rect 43437 8802 43503 8805
rect 41781 8800 43503 8802
rect 41781 8744 41786 8800
rect 41842 8744 43442 8800
rect 43498 8744 43503 8800
rect 41781 8742 43503 8744
rect 41781 8739 41847 8742
rect 43437 8739 43503 8742
rect 49233 8802 49299 8805
rect 50200 8802 51000 8832
rect 49233 8800 51000 8802
rect 49233 8744 49238 8800
rect 49294 8744 51000 8800
rect 49233 8742 51000 8744
rect 49233 8739 49299 8742
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 50200 8712 51000 8742
rect 47946 8671 48262 8672
rect 42149 8666 42215 8669
rect 38334 8664 42215 8666
rect 38334 8608 42154 8664
rect 42210 8608 42215 8664
rect 38334 8606 42215 8608
rect 18413 8603 18479 8606
rect 24761 8603 24827 8606
rect 42149 8603 42215 8606
rect 0 8530 800 8560
rect 1209 8530 1275 8533
rect 0 8528 1275 8530
rect 0 8472 1214 8528
rect 1270 8472 1275 8528
rect 0 8470 1275 8472
rect 0 8440 800 8470
rect 1209 8467 1275 8470
rect 13721 8530 13787 8533
rect 17033 8530 17099 8533
rect 17585 8530 17651 8533
rect 13721 8528 17651 8530
rect 13721 8472 13726 8528
rect 13782 8472 17038 8528
rect 17094 8472 17590 8528
rect 17646 8472 17651 8528
rect 13721 8470 17651 8472
rect 13721 8467 13787 8470
rect 17033 8467 17099 8470
rect 17585 8467 17651 8470
rect 18045 8530 18111 8533
rect 18454 8530 18460 8532
rect 18045 8528 18460 8530
rect 18045 8472 18050 8528
rect 18106 8472 18460 8528
rect 18045 8470 18460 8472
rect 18045 8467 18111 8470
rect 18454 8468 18460 8470
rect 18524 8530 18530 8532
rect 18873 8530 18939 8533
rect 18524 8528 18939 8530
rect 18524 8472 18878 8528
rect 18934 8472 18939 8528
rect 18524 8470 18939 8472
rect 18524 8468 18530 8470
rect 18873 8467 18939 8470
rect 20161 8530 20227 8533
rect 24301 8530 24367 8533
rect 20161 8528 24367 8530
rect 20161 8472 20166 8528
rect 20222 8472 24306 8528
rect 24362 8472 24367 8528
rect 20161 8470 24367 8472
rect 20161 8467 20227 8470
rect 24301 8467 24367 8470
rect 24577 8530 24643 8533
rect 40033 8530 40099 8533
rect 24577 8528 40099 8530
rect 24577 8472 24582 8528
rect 24638 8472 40038 8528
rect 40094 8472 40099 8528
rect 24577 8470 40099 8472
rect 24577 8467 24643 8470
rect 40033 8467 40099 8470
rect 42558 8468 42564 8532
rect 42628 8530 42634 8532
rect 44357 8530 44423 8533
rect 42628 8528 44423 8530
rect 42628 8472 44362 8528
rect 44418 8472 44423 8528
rect 42628 8470 44423 8472
rect 42628 8468 42634 8470
rect 44357 8467 44423 8470
rect 3509 8394 3575 8397
rect 15694 8394 15700 8396
rect 3509 8392 15700 8394
rect 3509 8336 3514 8392
rect 3570 8336 15700 8392
rect 3509 8334 15700 8336
rect 3509 8331 3575 8334
rect 15694 8332 15700 8334
rect 15764 8332 15770 8396
rect 16205 8394 16271 8397
rect 18413 8394 18479 8397
rect 16205 8392 18479 8394
rect 16205 8336 16210 8392
rect 16266 8336 18418 8392
rect 18474 8336 18479 8392
rect 16205 8334 18479 8336
rect 16205 8331 16271 8334
rect 18413 8331 18479 8334
rect 20713 8394 20779 8397
rect 22134 8394 22140 8396
rect 20713 8392 22140 8394
rect 20713 8336 20718 8392
rect 20774 8336 22140 8392
rect 20713 8334 22140 8336
rect 20713 8331 20779 8334
rect 22134 8332 22140 8334
rect 22204 8332 22210 8396
rect 33041 8394 33107 8397
rect 33041 8392 33426 8394
rect 33041 8336 33046 8392
rect 33102 8336 33426 8392
rect 33041 8334 33426 8336
rect 33041 8331 33107 8334
rect 9949 8260 10015 8261
rect 9949 8256 9996 8260
rect 10060 8258 10066 8260
rect 9949 8200 9954 8256
rect 9949 8196 9996 8200
rect 10060 8198 10106 8258
rect 10060 8196 10066 8198
rect 16246 8196 16252 8260
rect 16316 8258 16322 8260
rect 16665 8258 16731 8261
rect 16316 8256 16731 8258
rect 16316 8200 16670 8256
rect 16726 8200 16731 8256
rect 16316 8198 16731 8200
rect 16316 8196 16322 8198
rect 9949 8195 10015 8196
rect 16665 8195 16731 8198
rect 18137 8258 18203 8261
rect 18638 8258 18644 8260
rect 18137 8256 18644 8258
rect 18137 8200 18142 8256
rect 18198 8200 18644 8256
rect 18137 8198 18644 8200
rect 18137 8195 18203 8198
rect 18638 8196 18644 8198
rect 18708 8196 18714 8260
rect 33366 8258 33426 8334
rect 34094 8332 34100 8396
rect 34164 8394 34170 8396
rect 43897 8394 43963 8397
rect 34164 8392 43963 8394
rect 34164 8336 43902 8392
rect 43958 8336 43963 8392
rect 34164 8334 43963 8336
rect 34164 8332 34170 8334
rect 43897 8331 43963 8334
rect 49325 8394 49391 8397
rect 50200 8394 51000 8424
rect 49325 8392 51000 8394
rect 49325 8336 49330 8392
rect 49386 8336 51000 8392
rect 49325 8334 51000 8336
rect 49325 8331 49391 8334
rect 50200 8304 51000 8334
rect 39205 8258 39271 8261
rect 33366 8256 39271 8258
rect 33366 8200 39210 8256
rect 39266 8200 39271 8256
rect 33366 8198 39271 8200
rect 39205 8195 39271 8198
rect 45921 8258 45987 8261
rect 48446 8258 48452 8260
rect 45921 8256 48452 8258
rect 45921 8200 45926 8256
rect 45982 8200 48452 8256
rect 45921 8198 48452 8200
rect 45921 8195 45987 8198
rect 48446 8196 48452 8198
rect 48516 8196 48522 8260
rect 2946 8192 3262 8193
rect 0 8122 800 8152
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 1577 8122 1643 8125
rect 0 8120 1643 8122
rect 0 8064 1582 8120
rect 1638 8064 1643 8120
rect 0 8062 1643 8064
rect 0 8032 800 8062
rect 1577 8059 1643 8062
rect 14774 8060 14780 8124
rect 14844 8122 14850 8124
rect 21725 8122 21791 8125
rect 14844 8120 21791 8122
rect 14844 8064 21730 8120
rect 21786 8064 21791 8120
rect 14844 8062 21791 8064
rect 14844 8060 14850 8062
rect 21725 8059 21791 8062
rect 35893 8122 35959 8125
rect 40217 8122 40283 8125
rect 35893 8120 40283 8122
rect 35893 8064 35898 8120
rect 35954 8064 40222 8120
rect 40278 8064 40283 8120
rect 35893 8062 40283 8064
rect 35893 8059 35959 8062
rect 40217 8059 40283 8062
rect 40534 8060 40540 8124
rect 40604 8122 40610 8124
rect 41505 8122 41571 8125
rect 40604 8120 41571 8122
rect 40604 8064 41510 8120
rect 41566 8064 41571 8120
rect 40604 8062 41571 8064
rect 40604 8060 40610 8062
rect 41505 8059 41571 8062
rect 10041 7986 10107 7989
rect 10174 7986 10180 7988
rect 10041 7984 10180 7986
rect 10041 7928 10046 7984
rect 10102 7928 10180 7984
rect 10041 7926 10180 7928
rect 10041 7923 10107 7926
rect 10174 7924 10180 7926
rect 10244 7924 10250 7988
rect 15101 7986 15167 7989
rect 16430 7986 16436 7988
rect 15101 7984 16436 7986
rect 15101 7928 15106 7984
rect 15162 7928 16436 7984
rect 15101 7926 16436 7928
rect 15101 7923 15167 7926
rect 16430 7924 16436 7926
rect 16500 7924 16506 7988
rect 34421 7986 34487 7989
rect 38694 7986 38700 7988
rect 34421 7984 38700 7986
rect 34421 7928 34426 7984
rect 34482 7928 38700 7984
rect 34421 7926 38700 7928
rect 34421 7923 34487 7926
rect 38694 7924 38700 7926
rect 38764 7924 38770 7988
rect 42006 7924 42012 7988
rect 42076 7986 42082 7988
rect 42885 7986 42951 7989
rect 42076 7984 42951 7986
rect 42076 7928 42890 7984
rect 42946 7928 42951 7984
rect 42076 7926 42951 7928
rect 42076 7924 42082 7926
rect 42885 7923 42951 7926
rect 46841 7986 46907 7989
rect 50200 7986 51000 8016
rect 46841 7984 51000 7986
rect 46841 7928 46846 7984
rect 46902 7928 51000 7984
rect 46841 7926 51000 7928
rect 46841 7923 46907 7926
rect 50200 7896 51000 7926
rect 14089 7850 14155 7853
rect 23422 7850 23428 7852
rect 14089 7848 23428 7850
rect 14089 7792 14094 7848
rect 14150 7792 23428 7848
rect 14089 7790 23428 7792
rect 14089 7787 14155 7790
rect 23422 7788 23428 7790
rect 23492 7788 23498 7852
rect 29545 7850 29611 7853
rect 33317 7850 33383 7853
rect 40125 7850 40191 7853
rect 29545 7848 40191 7850
rect 29545 7792 29550 7848
rect 29606 7792 33322 7848
rect 33378 7792 40130 7848
rect 40186 7792 40191 7848
rect 29545 7790 40191 7792
rect 29545 7787 29611 7790
rect 33317 7787 33383 7790
rect 40125 7787 40191 7790
rect 41229 7850 41295 7853
rect 46381 7850 46447 7853
rect 41229 7848 46447 7850
rect 41229 7792 41234 7848
rect 41290 7792 46386 7848
rect 46442 7792 46447 7848
rect 41229 7790 46447 7792
rect 41229 7787 41295 7790
rect 46381 7787 46447 7790
rect 0 7714 800 7744
rect 1301 7714 1367 7717
rect 0 7712 1367 7714
rect 0 7656 1306 7712
rect 1362 7656 1367 7712
rect 0 7654 1367 7656
rect 0 7624 800 7654
rect 1301 7651 1367 7654
rect 8569 7714 8635 7717
rect 14958 7714 14964 7716
rect 8569 7712 14964 7714
rect 8569 7656 8574 7712
rect 8630 7656 14964 7712
rect 8569 7654 14964 7656
rect 8569 7651 8635 7654
rect 14958 7652 14964 7654
rect 15028 7652 15034 7716
rect 20897 7714 20963 7717
rect 24894 7714 24900 7716
rect 20897 7712 24900 7714
rect 20897 7656 20902 7712
rect 20958 7656 24900 7712
rect 20897 7654 24900 7656
rect 20897 7651 20963 7654
rect 24894 7652 24900 7654
rect 24964 7652 24970 7716
rect 38510 7652 38516 7716
rect 38580 7714 38586 7716
rect 44541 7714 44607 7717
rect 38580 7712 44607 7714
rect 38580 7656 44546 7712
rect 44602 7656 44607 7712
rect 38580 7654 44607 7656
rect 38580 7652 38586 7654
rect 44541 7651 44607 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 11329 7578 11395 7581
rect 16614 7578 16620 7580
rect 11329 7576 16620 7578
rect 11329 7520 11334 7576
rect 11390 7520 16620 7576
rect 11329 7518 16620 7520
rect 11329 7515 11395 7518
rect 16614 7516 16620 7518
rect 16684 7516 16690 7580
rect 49141 7578 49207 7581
rect 50200 7578 51000 7608
rect 49141 7576 51000 7578
rect 49141 7520 49146 7576
rect 49202 7520 51000 7576
rect 49141 7518 51000 7520
rect 49141 7515 49207 7518
rect 50200 7488 51000 7518
rect 11973 7442 12039 7445
rect 23790 7442 23796 7444
rect 11973 7440 23796 7442
rect 11973 7384 11978 7440
rect 12034 7384 23796 7440
rect 11973 7382 23796 7384
rect 11973 7379 12039 7382
rect 23790 7380 23796 7382
rect 23860 7380 23866 7444
rect 30189 7442 30255 7445
rect 38009 7442 38075 7445
rect 30189 7440 38075 7442
rect 30189 7384 30194 7440
rect 30250 7384 38014 7440
rect 38070 7384 38075 7440
rect 30189 7382 38075 7384
rect 30189 7379 30255 7382
rect 38009 7379 38075 7382
rect 39982 7380 39988 7444
rect 40052 7442 40058 7444
rect 45001 7442 45067 7445
rect 40052 7440 45067 7442
rect 40052 7384 45006 7440
rect 45062 7384 45067 7440
rect 40052 7382 45067 7384
rect 40052 7380 40058 7382
rect 45001 7379 45067 7382
rect 45134 7380 45140 7444
rect 45204 7442 45210 7444
rect 46197 7442 46263 7445
rect 45204 7440 46263 7442
rect 45204 7384 46202 7440
rect 46258 7384 46263 7440
rect 45204 7382 46263 7384
rect 45204 7380 45210 7382
rect 46197 7379 46263 7382
rect 0 7306 800 7336
rect 1301 7306 1367 7309
rect 0 7304 1367 7306
rect 0 7248 1306 7304
rect 1362 7248 1367 7304
rect 0 7246 1367 7248
rect 0 7216 800 7246
rect 1301 7243 1367 7246
rect 9489 7306 9555 7309
rect 20713 7306 20779 7309
rect 9489 7304 20779 7306
rect 9489 7248 9494 7304
rect 9550 7248 20718 7304
rect 20774 7248 20779 7304
rect 9489 7246 20779 7248
rect 9489 7243 9555 7246
rect 20713 7243 20779 7246
rect 30230 7244 30236 7308
rect 30300 7306 30306 7308
rect 39113 7306 39179 7309
rect 30300 7304 39179 7306
rect 30300 7248 39118 7304
rect 39174 7248 39179 7304
rect 30300 7246 39179 7248
rect 30300 7244 30306 7246
rect 39113 7243 39179 7246
rect 44449 7306 44515 7309
rect 45185 7306 45251 7309
rect 50061 7306 50127 7309
rect 44449 7304 50127 7306
rect 44449 7248 44454 7304
rect 44510 7248 45190 7304
rect 45246 7248 50066 7304
rect 50122 7248 50127 7304
rect 44449 7246 50127 7248
rect 44449 7243 44515 7246
rect 45185 7243 45251 7246
rect 50061 7243 50127 7246
rect 16665 7170 16731 7173
rect 19558 7170 19564 7172
rect 16665 7168 19564 7170
rect 16665 7112 16670 7168
rect 16726 7112 19564 7168
rect 16665 7110 19564 7112
rect 16665 7107 16731 7110
rect 19558 7108 19564 7110
rect 19628 7108 19634 7172
rect 49233 7170 49299 7173
rect 50200 7170 51000 7200
rect 49233 7168 51000 7170
rect 49233 7112 49238 7168
rect 49294 7112 51000 7168
rect 49233 7110 51000 7112
rect 49233 7107 49299 7110
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 50200 7080 51000 7110
rect 42946 7039 43262 7040
rect 43529 7034 43595 7037
rect 45686 7034 45692 7036
rect 43529 7032 45692 7034
rect 43529 6976 43534 7032
rect 43590 6976 45692 7032
rect 43529 6974 45692 6976
rect 43529 6971 43595 6974
rect 45686 6972 45692 6974
rect 45756 6972 45762 7036
rect 0 6898 800 6928
rect 1209 6898 1275 6901
rect 0 6896 1275 6898
rect 0 6840 1214 6896
rect 1270 6840 1275 6896
rect 0 6838 1275 6840
rect 0 6808 800 6838
rect 1209 6835 1275 6838
rect 11329 6898 11395 6901
rect 11462 6898 11468 6900
rect 11329 6896 11468 6898
rect 11329 6840 11334 6896
rect 11390 6840 11468 6896
rect 11329 6838 11468 6840
rect 11329 6835 11395 6838
rect 11462 6836 11468 6838
rect 11532 6836 11538 6900
rect 13721 6898 13787 6901
rect 29494 6898 29500 6900
rect 13721 6896 29500 6898
rect 13721 6840 13726 6896
rect 13782 6840 29500 6896
rect 13721 6838 29500 6840
rect 13721 6835 13787 6838
rect 29494 6836 29500 6838
rect 29564 6836 29570 6900
rect 43345 6898 43411 6901
rect 43846 6898 43852 6900
rect 43345 6896 43852 6898
rect 43345 6840 43350 6896
rect 43406 6840 43852 6896
rect 43345 6838 43852 6840
rect 43345 6835 43411 6838
rect 43846 6836 43852 6838
rect 43916 6836 43922 6900
rect 45921 6898 45987 6901
rect 49877 6898 49943 6901
rect 44222 6838 45754 6898
rect 12198 6700 12204 6764
rect 12268 6762 12274 6764
rect 12341 6762 12407 6765
rect 12268 6760 12407 6762
rect 12268 6704 12346 6760
rect 12402 6704 12407 6760
rect 12268 6702 12407 6704
rect 12268 6700 12274 6702
rect 12341 6699 12407 6702
rect 14273 6762 14339 6765
rect 16665 6762 16731 6765
rect 14273 6760 16731 6762
rect 14273 6704 14278 6760
rect 14334 6704 16670 6760
rect 16726 6704 16731 6760
rect 14273 6702 16731 6704
rect 14273 6699 14339 6702
rect 16665 6699 16731 6702
rect 35801 6762 35867 6765
rect 44222 6762 44282 6838
rect 35801 6760 44282 6762
rect 35801 6704 35806 6760
rect 35862 6704 44282 6760
rect 35801 6702 44282 6704
rect 44357 6762 44423 6765
rect 45502 6762 45508 6764
rect 44357 6760 45508 6762
rect 44357 6704 44362 6760
rect 44418 6704 45508 6760
rect 44357 6702 45508 6704
rect 35801 6699 35867 6702
rect 44357 6699 44423 6702
rect 45502 6700 45508 6702
rect 45572 6700 45578 6764
rect 39798 6564 39804 6628
rect 39868 6626 39874 6628
rect 45461 6626 45527 6629
rect 39868 6624 45527 6626
rect 39868 6568 45466 6624
rect 45522 6568 45527 6624
rect 39868 6566 45527 6568
rect 45694 6626 45754 6838
rect 45921 6896 49943 6898
rect 45921 6840 45926 6896
rect 45982 6840 49882 6896
rect 49938 6840 49943 6896
rect 45921 6838 49943 6840
rect 45921 6835 45987 6838
rect 49877 6835 49943 6838
rect 46974 6700 46980 6764
rect 47044 6762 47050 6764
rect 47209 6762 47275 6765
rect 49325 6762 49391 6765
rect 50200 6762 51000 6792
rect 47044 6760 47275 6762
rect 47044 6704 47214 6760
rect 47270 6704 47275 6760
rect 47044 6702 47275 6704
rect 47044 6700 47050 6702
rect 47209 6699 47275 6702
rect 47350 6702 48514 6762
rect 47350 6626 47410 6702
rect 45694 6566 47410 6626
rect 48454 6626 48514 6702
rect 49325 6760 51000 6762
rect 49325 6704 49330 6760
rect 49386 6704 51000 6760
rect 49325 6702 51000 6704
rect 49325 6699 49391 6702
rect 50200 6672 51000 6702
rect 49509 6626 49575 6629
rect 48454 6624 49575 6626
rect 48454 6568 49514 6624
rect 49570 6568 49575 6624
rect 48454 6566 49575 6568
rect 39868 6564 39874 6566
rect 45461 6563 45527 6566
rect 49509 6563 49575 6566
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 1301 6490 1367 6493
rect 0 6488 1367 6490
rect 0 6432 1306 6488
rect 1362 6432 1367 6488
rect 0 6430 1367 6432
rect 0 6400 800 6430
rect 1301 6427 1367 6430
rect 28758 6428 28764 6492
rect 28828 6490 28834 6492
rect 35617 6490 35683 6493
rect 28828 6488 35683 6490
rect 28828 6432 35622 6488
rect 35678 6432 35683 6488
rect 28828 6430 35683 6432
rect 28828 6428 28834 6430
rect 35617 6427 35683 6430
rect 44766 6428 44772 6492
rect 44836 6490 44842 6492
rect 46013 6490 46079 6493
rect 44836 6488 46079 6490
rect 44836 6432 46018 6488
rect 46074 6432 46079 6488
rect 44836 6430 46079 6432
rect 44836 6428 44842 6430
rect 46013 6427 46079 6430
rect 21214 6292 21220 6356
rect 21284 6354 21290 6356
rect 40033 6354 40099 6357
rect 21284 6352 40099 6354
rect 21284 6296 40038 6352
rect 40094 6296 40099 6352
rect 21284 6294 40099 6296
rect 21284 6292 21290 6294
rect 40033 6291 40099 6294
rect 40350 6292 40356 6356
rect 40420 6354 40426 6356
rect 47209 6354 47275 6357
rect 40420 6352 47275 6354
rect 40420 6296 47214 6352
rect 47270 6296 47275 6352
rect 40420 6294 47275 6296
rect 40420 6292 40426 6294
rect 47209 6291 47275 6294
rect 48681 6354 48747 6357
rect 50200 6354 51000 6384
rect 48681 6352 51000 6354
rect 48681 6296 48686 6352
rect 48742 6296 51000 6352
rect 48681 6294 51000 6296
rect 48681 6291 48747 6294
rect 50200 6264 51000 6294
rect 12341 6218 12407 6221
rect 20662 6218 20668 6220
rect 12341 6216 20668 6218
rect 12341 6160 12346 6216
rect 12402 6160 20668 6216
rect 12341 6158 20668 6160
rect 12341 6155 12407 6158
rect 20662 6156 20668 6158
rect 20732 6156 20738 6220
rect 40902 6156 40908 6220
rect 40972 6218 40978 6220
rect 46657 6218 46723 6221
rect 40972 6216 46723 6218
rect 40972 6160 46662 6216
rect 46718 6160 46723 6216
rect 40972 6158 46723 6160
rect 40972 6156 40978 6158
rect 46657 6155 46723 6158
rect 0 6082 800 6112
rect 1301 6082 1367 6085
rect 0 6080 1367 6082
rect 0 6024 1306 6080
rect 1362 6024 1367 6080
rect 0 6022 1367 6024
rect 0 5992 800 6022
rect 1301 6019 1367 6022
rect 33409 6082 33475 6085
rect 41597 6082 41663 6085
rect 33409 6080 41663 6082
rect 33409 6024 33414 6080
rect 33470 6024 41602 6080
rect 41658 6024 41663 6080
rect 33409 6022 41663 6024
rect 33409 6019 33475 6022
rect 41597 6019 41663 6022
rect 45093 6082 45159 6085
rect 45921 6082 45987 6085
rect 45093 6080 45987 6082
rect 45093 6024 45098 6080
rect 45154 6024 45926 6080
rect 45982 6024 45987 6080
rect 45093 6022 45987 6024
rect 45093 6019 45159 6022
rect 45921 6019 45987 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 35893 5946 35959 5949
rect 37222 5946 37228 5948
rect 35893 5944 37228 5946
rect 35893 5888 35898 5944
rect 35954 5888 37228 5944
rect 35893 5886 37228 5888
rect 35893 5883 35959 5886
rect 37222 5884 37228 5886
rect 37292 5884 37298 5948
rect 49141 5946 49207 5949
rect 50200 5946 51000 5976
rect 49141 5944 51000 5946
rect 49141 5888 49146 5944
rect 49202 5888 51000 5944
rect 49141 5886 51000 5888
rect 49141 5883 49207 5886
rect 50200 5856 51000 5886
rect 27470 5748 27476 5812
rect 27540 5810 27546 5812
rect 45001 5810 45067 5813
rect 27540 5808 45067 5810
rect 27540 5752 45006 5808
rect 45062 5752 45067 5808
rect 27540 5750 45067 5752
rect 27540 5748 27546 5750
rect 45001 5747 45067 5750
rect 0 5674 800 5704
rect 1301 5674 1367 5677
rect 0 5672 1367 5674
rect 0 5616 1306 5672
rect 1362 5616 1367 5672
rect 0 5614 1367 5616
rect 0 5584 800 5614
rect 1301 5611 1367 5614
rect 27102 5612 27108 5676
rect 27172 5674 27178 5676
rect 39389 5674 39455 5677
rect 27172 5672 39455 5674
rect 27172 5616 39394 5672
rect 39450 5616 39455 5672
rect 27172 5614 39455 5616
rect 27172 5612 27178 5614
rect 39389 5611 39455 5614
rect 45553 5674 45619 5677
rect 46790 5674 46796 5676
rect 45553 5672 46796 5674
rect 45553 5616 45558 5672
rect 45614 5616 46796 5672
rect 45553 5614 46796 5616
rect 45553 5611 45619 5614
rect 46790 5612 46796 5614
rect 46860 5612 46866 5676
rect 49417 5538 49483 5541
rect 50200 5538 51000 5568
rect 49417 5536 51000 5538
rect 49417 5480 49422 5536
rect 49478 5480 51000 5536
rect 49417 5478 51000 5480
rect 49417 5475 49483 5478
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 50200 5448 51000 5478
rect 47946 5407 48262 5408
rect 0 5266 800 5296
rect 2773 5266 2839 5269
rect 17125 5268 17191 5269
rect 17125 5266 17172 5268
rect 0 5264 2839 5266
rect 0 5208 2778 5264
rect 2834 5208 2839 5264
rect 0 5206 2839 5208
rect 17080 5264 17172 5266
rect 17080 5208 17130 5264
rect 17080 5206 17172 5208
rect 0 5176 800 5206
rect 2773 5203 2839 5206
rect 17125 5204 17172 5206
rect 17236 5204 17242 5268
rect 35157 5266 35223 5269
rect 38101 5266 38167 5269
rect 41413 5266 41479 5269
rect 35157 5264 38167 5266
rect 35157 5208 35162 5264
rect 35218 5208 38106 5264
rect 38162 5208 38167 5264
rect 35157 5206 38167 5208
rect 17125 5203 17191 5204
rect 35157 5203 35223 5206
rect 38101 5203 38167 5206
rect 38380 5264 41479 5266
rect 38380 5208 41418 5264
rect 41474 5208 41479 5264
rect 38380 5206 41479 5208
rect 36670 5068 36676 5132
rect 36740 5130 36746 5132
rect 38380 5130 38440 5206
rect 41413 5203 41479 5206
rect 43437 5130 43503 5133
rect 36740 5070 38440 5130
rect 41370 5128 43503 5130
rect 41370 5072 43442 5128
rect 43498 5072 43503 5128
rect 41370 5070 43503 5072
rect 36740 5068 36746 5070
rect 36486 4932 36492 4996
rect 36556 4994 36562 4996
rect 41370 4994 41430 5070
rect 43437 5067 43503 5070
rect 49233 5130 49299 5133
rect 50200 5130 51000 5160
rect 49233 5128 51000 5130
rect 49233 5072 49238 5128
rect 49294 5072 51000 5128
rect 49233 5070 51000 5072
rect 49233 5067 49299 5070
rect 50200 5040 51000 5070
rect 36556 4934 41430 4994
rect 36556 4932 36562 4934
rect 2946 4928 3262 4929
rect 0 4858 800 4888
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 31334 4660 31340 4724
rect 31404 4722 31410 4724
rect 42701 4722 42767 4725
rect 31404 4720 42767 4722
rect 31404 4664 42706 4720
rect 42762 4664 42767 4720
rect 31404 4662 42767 4664
rect 31404 4660 31410 4662
rect 42701 4659 42767 4662
rect 48313 4722 48379 4725
rect 50200 4722 51000 4752
rect 48313 4720 51000 4722
rect 48313 4664 48318 4720
rect 48374 4664 51000 4720
rect 48313 4662 51000 4664
rect 48313 4659 48379 4662
rect 50200 4632 51000 4662
rect 35382 4524 35388 4588
rect 35452 4586 35458 4588
rect 44725 4586 44791 4589
rect 35452 4584 44791 4586
rect 35452 4528 44730 4584
rect 44786 4528 44791 4584
rect 35452 4526 44791 4528
rect 35452 4524 35458 4526
rect 44725 4523 44791 4526
rect 0 4450 800 4480
rect 1301 4450 1367 4453
rect 0 4448 1367 4450
rect 0 4392 1306 4448
rect 1362 4392 1367 4448
rect 0 4390 1367 4392
rect 0 4360 800 4390
rect 1301 4387 1367 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 49141 4314 49207 4317
rect 50200 4314 51000 4344
rect 49141 4312 51000 4314
rect 49141 4256 49146 4312
rect 49202 4256 51000 4312
rect 49141 4254 51000 4256
rect 49141 4251 49207 4254
rect 50200 4224 51000 4254
rect 0 4042 800 4072
rect 1301 4042 1367 4045
rect 0 4040 1367 4042
rect 0 3984 1306 4040
rect 1362 3984 1367 4040
rect 0 3982 1367 3984
rect 0 3952 800 3982
rect 1301 3979 1367 3982
rect 7465 4042 7531 4045
rect 23749 4042 23815 4045
rect 24945 4042 25011 4045
rect 7465 4040 25011 4042
rect 7465 3984 7470 4040
rect 7526 3984 23754 4040
rect 23810 3984 24950 4040
rect 25006 3984 25011 4040
rect 7465 3982 25011 3984
rect 7465 3979 7531 3982
rect 23749 3979 23815 3982
rect 24945 3979 25011 3982
rect 49233 3906 49299 3909
rect 50200 3906 51000 3936
rect 49233 3904 51000 3906
rect 49233 3848 49238 3904
rect 49294 3848 51000 3904
rect 49233 3846 51000 3848
rect 49233 3843 49299 3846
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 50200 3816 51000 3846
rect 42946 3775 43262 3776
rect 0 3634 800 3664
rect 1209 3634 1275 3637
rect 0 3632 1275 3634
rect 0 3576 1214 3632
rect 1270 3576 1275 3632
rect 0 3574 1275 3576
rect 0 3544 800 3574
rect 1209 3571 1275 3574
rect 8293 3634 8359 3637
rect 18321 3634 18387 3637
rect 8293 3632 18387 3634
rect 8293 3576 8298 3632
rect 8354 3576 18326 3632
rect 18382 3576 18387 3632
rect 8293 3574 18387 3576
rect 8293 3571 8359 3574
rect 18321 3571 18387 3574
rect 49141 3498 49207 3501
rect 50200 3498 51000 3528
rect 49141 3496 51000 3498
rect 49141 3440 49146 3496
rect 49202 3440 51000 3496
rect 49141 3438 51000 3440
rect 49141 3435 49207 3438
rect 50200 3408 51000 3438
rect 7946 3296 8262 3297
rect 0 3226 800 3256
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 1301 3226 1367 3229
rect 0 3224 1367 3226
rect 0 3168 1306 3224
rect 1362 3168 1367 3224
rect 0 3166 1367 3168
rect 0 3136 800 3166
rect 1301 3163 1367 3166
rect 48681 3090 48747 3093
rect 50200 3090 51000 3120
rect 48681 3088 51000 3090
rect 48681 3032 48686 3088
rect 48742 3032 51000 3088
rect 48681 3030 51000 3032
rect 48681 3027 48747 3030
rect 50200 3000 51000 3030
rect 0 2818 800 2848
rect 1301 2818 1367 2821
rect 0 2816 1367 2818
rect 0 2760 1306 2816
rect 1362 2760 1367 2816
rect 0 2758 1367 2760
rect 0 2728 800 2758
rect 1301 2755 1367 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 46841 2682 46907 2685
rect 50200 2682 51000 2712
rect 46841 2680 51000 2682
rect 46841 2624 46846 2680
rect 46902 2624 51000 2680
rect 46841 2622 51000 2624
rect 46841 2619 46907 2622
rect 50200 2592 51000 2622
rect 0 2410 800 2440
rect 1301 2410 1367 2413
rect 0 2408 1367 2410
rect 0 2352 1306 2408
rect 1362 2352 1367 2408
rect 0 2350 1367 2352
rect 0 2320 800 2350
rect 1301 2347 1367 2350
rect 48497 2274 48563 2277
rect 50200 2274 51000 2304
rect 48497 2272 51000 2274
rect 48497 2216 48502 2272
rect 48558 2216 51000 2272
rect 48497 2214 51000 2216
rect 48497 2211 48563 2214
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 50200 2184 51000 2214
rect 47946 2143 48262 2144
rect 0 2002 800 2032
rect 1209 2002 1275 2005
rect 0 2000 1275 2002
rect 0 1944 1214 2000
rect 1270 1944 1275 2000
rect 0 1942 1275 1944
rect 0 1912 800 1942
rect 1209 1939 1275 1942
rect 46749 1866 46815 1869
rect 50200 1866 51000 1896
rect 46749 1864 51000 1866
rect 46749 1808 46754 1864
rect 46810 1808 51000 1864
rect 46749 1806 51000 1808
rect 46749 1803 46815 1806
rect 50200 1776 51000 1806
rect 0 1594 800 1624
rect 3233 1594 3299 1597
rect 0 1592 3299 1594
rect 0 1536 3238 1592
rect 3294 1536 3299 1592
rect 0 1534 3299 1536
rect 0 1504 800 1534
rect 3233 1531 3299 1534
rect 46657 1458 46723 1461
rect 50200 1458 51000 1488
rect 46657 1456 51000 1458
rect 46657 1400 46662 1456
rect 46718 1400 51000 1456
rect 46657 1398 51000 1400
rect 46657 1395 46723 1398
rect 50200 1368 51000 1398
<< via3 >>
rect 24164 26692 24228 26756
rect 47164 26556 47228 26620
rect 46060 26148 46124 26212
rect 30052 25876 30116 25940
rect 22508 25604 22572 25668
rect 19932 25060 19996 25124
rect 44220 25060 44284 25124
rect 3372 24924 3436 24988
rect 24900 24924 24964 24988
rect 34652 24516 34716 24580
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 40356 23972 40420 24036
rect 43668 23972 43732 24036
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 34468 23836 34532 23900
rect 46980 23836 47044 23900
rect 3924 23700 3988 23764
rect 7604 23564 7668 23628
rect 34652 23564 34716 23628
rect 36492 23564 36556 23628
rect 4292 23488 4356 23492
rect 4292 23432 4306 23488
rect 4306 23432 4356 23488
rect 4292 23428 4356 23432
rect 17172 23428 17236 23492
rect 20668 23428 20732 23492
rect 23428 23428 23492 23492
rect 27476 23428 27540 23492
rect 28764 23428 28828 23492
rect 30236 23428 30300 23492
rect 30972 23428 31036 23492
rect 31524 23488 31588 23492
rect 31524 23432 31574 23488
rect 31574 23432 31588 23488
rect 31524 23428 31588 23432
rect 32444 23488 32508 23492
rect 32444 23432 32494 23488
rect 32494 23432 32508 23488
rect 32444 23428 32508 23432
rect 34100 23428 34164 23492
rect 36676 23428 36740 23492
rect 38516 23428 38580 23492
rect 39436 23428 39500 23492
rect 40540 23428 40604 23492
rect 42564 23428 42628 23492
rect 44956 23428 45020 23492
rect 46244 23428 46308 23492
rect 46796 23488 46860 23492
rect 46796 23432 46846 23488
rect 46846 23432 46860 23488
rect 46796 23428 46860 23432
rect 48452 23428 48516 23492
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 21220 23292 21284 23356
rect 30052 23292 30116 23356
rect 34836 23156 34900 23220
rect 37412 23292 37476 23356
rect 5212 23020 5276 23084
rect 44036 23020 44100 23084
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 9260 22748 9324 22812
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 22140 22748 22204 22812
rect 5764 22612 5828 22676
rect 27292 22612 27356 22676
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 34284 22748 34348 22812
rect 9812 22400 9876 22404
rect 9812 22344 9826 22400
rect 9826 22344 9876 22400
rect 9812 22340 9876 22344
rect 26004 22340 26068 22404
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 23796 22204 23860 22268
rect 29316 22204 29380 22268
rect 11468 22068 11532 22132
rect 5580 21932 5644 21996
rect 31340 22068 31404 22132
rect 41092 22476 41156 22540
rect 37596 22340 37660 22404
rect 39804 22204 39868 22268
rect 45324 22340 45388 22404
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 28948 21992 29012 21996
rect 28948 21936 28962 21992
rect 28962 21936 29012 21992
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 7420 21660 7484 21724
rect 22324 21796 22388 21860
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 24164 21720 24228 21724
rect 24164 21664 24178 21720
rect 24178 21664 24228 21720
rect 24164 21660 24228 21664
rect 28948 21932 29012 21936
rect 35940 21932 36004 21996
rect 39068 21796 39132 21860
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 10180 21388 10244 21452
rect 35756 21524 35820 21588
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 26556 21252 26620 21316
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 12572 20844 12636 20908
rect 15700 20768 15764 20772
rect 15700 20712 15714 20768
rect 15714 20712 15764 20768
rect 15700 20708 15764 20712
rect 16988 20768 17052 20772
rect 16988 20712 17002 20768
rect 17002 20712 17052 20768
rect 16988 20708 17052 20712
rect 19380 20768 19444 20772
rect 19380 20712 19430 20768
rect 19430 20712 19444 20768
rect 19380 20708 19444 20712
rect 39620 20844 39684 20908
rect 41828 20844 41892 20908
rect 45140 20844 45204 20908
rect 48636 20708 48700 20772
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 41276 20572 41340 20636
rect 34468 20436 34532 20500
rect 35204 20436 35268 20500
rect 8892 20300 8956 20364
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 34652 20300 34716 20364
rect 35388 20360 35452 20364
rect 35388 20304 35402 20360
rect 35402 20304 35452 20360
rect 35388 20300 35452 20304
rect 39804 20436 39868 20500
rect 40724 20436 40788 20500
rect 40356 20300 40420 20364
rect 41092 20300 41156 20364
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 29316 20088 29380 20092
rect 29316 20032 29330 20088
rect 29330 20032 29380 20088
rect 29316 20028 29380 20032
rect 42012 20164 42076 20228
rect 44220 20164 44284 20228
rect 46428 20164 46492 20228
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 42380 20028 42444 20092
rect 38884 19892 38948 19956
rect 15148 19620 15212 19684
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 11100 19484 11164 19548
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 22324 19348 22388 19412
rect 29500 19348 29564 19412
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 38884 19484 38948 19548
rect 49188 19408 49252 19412
rect 49188 19352 49202 19408
rect 49202 19352 49252 19408
rect 49188 19348 49252 19352
rect 12204 19076 12268 19140
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 5580 18940 5644 19004
rect 8340 18668 8404 18732
rect 19932 19076 19996 19140
rect 34468 19212 34532 19276
rect 41644 19212 41708 19276
rect 33548 19076 33612 19140
rect 42380 19076 42444 19140
rect 44772 19136 44836 19140
rect 44772 19080 44786 19136
rect 44786 19080 44836 19136
rect 44772 19076 44836 19080
rect 47164 19076 47228 19140
rect 48820 19076 48884 19140
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 24900 19000 24964 19004
rect 24900 18944 24914 19000
rect 24914 18944 24964 19000
rect 24900 18940 24964 18944
rect 27660 18940 27724 19004
rect 31892 18940 31956 19004
rect 27108 18804 27172 18868
rect 44220 18864 44284 18868
rect 44220 18808 44270 18864
rect 44270 18808 44284 18864
rect 44220 18804 44284 18808
rect 46980 18864 47044 18868
rect 46980 18808 46994 18864
rect 46994 18808 47044 18864
rect 46980 18804 47044 18808
rect 49924 18804 49988 18868
rect 36860 18668 36924 18732
rect 3372 18592 3436 18596
rect 3372 18536 3422 18592
rect 3422 18536 3436 18592
rect 3372 18532 3436 18536
rect 38884 18532 38948 18596
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 6316 18396 6380 18460
rect 3556 18184 3620 18188
rect 37044 18396 37108 18460
rect 3556 18128 3606 18184
rect 3606 18128 3620 18184
rect 3556 18124 3620 18128
rect 14964 17988 15028 18052
rect 15332 17988 15396 18052
rect 19564 18048 19628 18052
rect 19564 17992 19578 18048
rect 19578 17992 19628 18048
rect 19564 17988 19628 17992
rect 24900 18048 24964 18052
rect 24900 17992 24950 18048
rect 24950 17992 24964 18048
rect 24900 17988 24964 17992
rect 26556 18048 26620 18052
rect 26556 17992 26606 18048
rect 26606 17992 26620 18048
rect 26556 17988 26620 17992
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 9996 17852 10060 17916
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 13676 17716 13740 17780
rect 9076 17580 9140 17644
rect 18460 17580 18524 17644
rect 27476 17852 27540 17916
rect 32628 17852 32692 17916
rect 38332 17988 38396 18052
rect 39804 17988 39868 18052
rect 45324 17988 45388 18052
rect 47716 18048 47780 18052
rect 47716 17992 47766 18048
rect 47766 17992 47780 18048
rect 47716 17988 47780 17992
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 46980 17852 47044 17916
rect 35940 17716 36004 17780
rect 26924 17580 26988 17644
rect 9444 17444 9508 17508
rect 45324 17444 45388 17508
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 27108 17308 27172 17372
rect 33364 17036 33428 17100
rect 13676 16900 13740 16964
rect 18644 16900 18708 16964
rect 27660 16960 27724 16964
rect 27660 16904 27710 16960
rect 27710 16904 27724 16960
rect 27660 16900 27724 16904
rect 34468 16900 34532 16964
rect 36860 16960 36924 16964
rect 36860 16904 36910 16960
rect 36910 16904 36924 16960
rect 36860 16900 36924 16904
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 38700 16764 38764 16828
rect 14780 16628 14844 16692
rect 17356 16688 17420 16692
rect 17356 16632 17370 16688
rect 17370 16632 17420 16688
rect 17356 16628 17420 16632
rect 35756 16628 35820 16692
rect 47348 16628 47412 16692
rect 16068 16416 16132 16420
rect 16068 16360 16082 16416
rect 16082 16360 16132 16416
rect 16068 16356 16132 16360
rect 29500 16492 29564 16556
rect 34284 16492 34348 16556
rect 31892 16356 31956 16420
rect 45324 16416 45388 16420
rect 45324 16360 45374 16416
rect 45374 16360 45388 16416
rect 45324 16356 45388 16360
rect 45508 16356 45572 16420
rect 46796 16356 46860 16420
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 18644 16220 18708 16284
rect 22508 16280 22572 16284
rect 22508 16224 22522 16280
rect 22522 16224 22572 16280
rect 22508 16220 22572 16224
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 15148 16084 15212 16148
rect 32812 16144 32876 16148
rect 32812 16088 32862 16144
rect 32862 16088 32876 16144
rect 32812 16084 32876 16088
rect 14044 15948 14108 16012
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 11100 15676 11164 15740
rect 44404 15812 44468 15876
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 40356 15268 40420 15332
rect 41276 15268 41340 15332
rect 46060 15268 46124 15332
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 12020 14996 12084 15060
rect 31156 15132 31220 15196
rect 38884 15192 38948 15196
rect 38884 15136 38934 15192
rect 38934 15136 38948 15192
rect 38884 15132 38948 15136
rect 41644 14996 41708 15060
rect 18460 14860 18524 14924
rect 26740 14860 26804 14924
rect 16436 14784 16500 14788
rect 16436 14728 16450 14784
rect 16450 14728 16500 14784
rect 16436 14724 16500 14728
rect 37596 14860 37660 14924
rect 40908 14724 40972 14788
rect 49924 14724 49988 14788
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 9260 14588 9324 14652
rect 6316 14316 6380 14380
rect 31524 14452 31588 14516
rect 13860 14180 13924 14244
rect 38332 14180 38396 14244
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 28948 14044 29012 14108
rect 40724 14044 40788 14108
rect 49188 14044 49252 14108
rect 33548 13908 33612 13972
rect 6316 13832 6380 13836
rect 6316 13776 6366 13832
rect 6366 13776 6380 13832
rect 6316 13772 6380 13776
rect 24900 13772 24964 13836
rect 31156 13772 31220 13836
rect 44772 13772 44836 13836
rect 3372 13696 3436 13700
rect 3372 13640 3422 13696
rect 3422 13640 3436 13696
rect 3372 13636 3436 13640
rect 5580 13636 5644 13700
rect 13492 13636 13556 13700
rect 41092 13636 41156 13700
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 4292 13500 4356 13564
rect 11652 13500 11716 13564
rect 43668 13500 43732 13564
rect 45692 13500 45756 13564
rect 48636 13500 48700 13564
rect 43668 13364 43732 13428
rect 47716 13364 47780 13428
rect 16252 13228 16316 13292
rect 35020 13228 35084 13292
rect 15148 13092 15212 13156
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 3924 13016 3988 13020
rect 3924 12960 3938 13016
rect 3938 12960 3988 13016
rect 3924 12956 3988 12960
rect 16252 12956 16316 13020
rect 46428 13228 46492 13292
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 3556 12820 3620 12884
rect 9076 12684 9140 12748
rect 4292 12548 4356 12612
rect 11652 12684 11716 12748
rect 43484 12548 43548 12612
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 13676 12412 13740 12476
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 9812 12276 9876 12340
rect 26924 12276 26988 12340
rect 16436 12140 16500 12204
rect 13860 12004 13924 12068
rect 26740 12004 26804 12068
rect 27108 12004 27172 12068
rect 35204 12276 35268 12340
rect 37228 12276 37292 12340
rect 38332 12336 38396 12340
rect 38332 12280 38346 12336
rect 38346 12280 38396 12336
rect 38332 12276 38396 12280
rect 44404 12140 44468 12204
rect 34284 12004 34348 12068
rect 38332 12004 38396 12068
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 39620 11868 39684 11932
rect 44772 11868 44836 11932
rect 46980 11868 47044 11932
rect 5764 11792 5828 11796
rect 5764 11736 5778 11792
rect 5778 11736 5828 11792
rect 5764 11732 5828 11736
rect 13676 11732 13740 11796
rect 38700 11732 38764 11796
rect 41828 11732 41892 11796
rect 44956 11792 45020 11796
rect 44956 11736 44970 11792
rect 44970 11736 45020 11792
rect 44956 11732 45020 11736
rect 32628 11596 32692 11660
rect 18460 11460 18524 11524
rect 27292 11460 27356 11524
rect 32260 11460 32324 11524
rect 35020 11460 35084 11524
rect 39068 11460 39132 11524
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 27292 11324 27356 11388
rect 32812 11384 32876 11388
rect 32812 11328 32826 11384
rect 32826 11328 32876 11384
rect 32812 11324 32876 11328
rect 33364 11324 33428 11388
rect 18644 11248 18708 11252
rect 18644 11192 18658 11248
rect 18658 11192 18708 11248
rect 18644 11188 18708 11192
rect 32444 11188 32508 11252
rect 34468 11188 34532 11252
rect 8892 11052 8956 11116
rect 9628 11052 9692 11116
rect 16252 11052 16316 11116
rect 34284 11052 34348 11116
rect 39436 11324 39500 11388
rect 47348 11384 47412 11388
rect 47348 11328 47398 11384
rect 47398 11328 47412 11384
rect 47348 11324 47412 11328
rect 43484 11248 43548 11252
rect 43484 11192 43498 11248
rect 43498 11192 43548 11248
rect 43484 11188 43548 11192
rect 39988 11052 40052 11116
rect 43852 11052 43916 11116
rect 46980 11052 47044 11116
rect 30972 10916 31036 10980
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 41828 10916 41892 10980
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 37044 10840 37108 10844
rect 37044 10784 37094 10840
rect 37094 10784 37108 10840
rect 37044 10780 37108 10784
rect 42380 10840 42444 10844
rect 42380 10784 42430 10840
rect 42430 10784 42444 10840
rect 42380 10780 42444 10784
rect 13492 10508 13556 10572
rect 8340 10372 8404 10436
rect 26004 10508 26068 10572
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 5212 10296 5276 10300
rect 5212 10240 5226 10296
rect 5226 10240 5276 10296
rect 5212 10236 5276 10240
rect 7420 10296 7484 10300
rect 7420 10240 7434 10296
rect 7434 10240 7484 10296
rect 7420 10236 7484 10240
rect 9444 10236 9508 10300
rect 16620 10236 16684 10300
rect 19380 10236 19444 10300
rect 34468 10100 34532 10164
rect 44220 10100 44284 10164
rect 46244 10100 46308 10164
rect 16068 9828 16132 9892
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 7604 9616 7668 9620
rect 7604 9560 7654 9616
rect 7654 9560 7668 9616
rect 7604 9556 7668 9560
rect 12020 9616 12084 9620
rect 12020 9560 12070 9616
rect 12070 9560 12084 9616
rect 12020 9556 12084 9560
rect 14044 9692 14108 9756
rect 16988 9692 17052 9756
rect 27292 9692 27356 9756
rect 12572 9284 12636 9348
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 18644 9148 18708 9212
rect 9628 9012 9692 9076
rect 34284 9556 34348 9620
rect 39068 9556 39132 9620
rect 43668 9556 43732 9620
rect 44036 9556 44100 9620
rect 34836 9284 34900 9348
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 37412 9012 37476 9076
rect 46980 9012 47044 9076
rect 48820 9012 48884 9076
rect 32260 8876 32324 8940
rect 18644 8740 18708 8804
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 17356 8604 17420 8668
rect 38700 8800 38764 8804
rect 38700 8744 38750 8800
rect 38750 8744 38764 8800
rect 38700 8740 38764 8744
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 18460 8468 18524 8532
rect 42564 8468 42628 8532
rect 15700 8332 15764 8396
rect 22140 8332 22204 8396
rect 9996 8256 10060 8260
rect 9996 8200 10010 8256
rect 10010 8200 10060 8256
rect 9996 8196 10060 8200
rect 16252 8196 16316 8260
rect 18644 8196 18708 8260
rect 34100 8332 34164 8396
rect 48452 8196 48516 8260
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 14780 8060 14844 8124
rect 40540 8060 40604 8124
rect 10180 7924 10244 7988
rect 16436 7924 16500 7988
rect 38700 7924 38764 7988
rect 42012 7924 42076 7988
rect 23428 7788 23492 7852
rect 14964 7652 15028 7716
rect 24900 7652 24964 7716
rect 38516 7652 38580 7716
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 16620 7516 16684 7580
rect 23796 7380 23860 7444
rect 39988 7380 40052 7444
rect 45140 7380 45204 7444
rect 30236 7244 30300 7308
rect 19564 7108 19628 7172
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 45692 6972 45756 7036
rect 11468 6836 11532 6900
rect 29500 6836 29564 6900
rect 43852 6836 43916 6900
rect 12204 6700 12268 6764
rect 45508 6700 45572 6764
rect 39804 6564 39868 6628
rect 46980 6700 47044 6764
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 28764 6428 28828 6492
rect 44772 6428 44836 6492
rect 21220 6292 21284 6356
rect 40356 6292 40420 6356
rect 20668 6156 20732 6220
rect 40908 6156 40972 6220
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 37228 5884 37292 5948
rect 27476 5748 27540 5812
rect 27108 5612 27172 5676
rect 46796 5612 46860 5676
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 17172 5264 17236 5268
rect 17172 5208 17186 5264
rect 17186 5208 17236 5264
rect 17172 5204 17236 5208
rect 36676 5068 36740 5132
rect 36492 4932 36556 4996
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 31340 4660 31404 4724
rect 35388 4524 35452 4588
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 24163 26756 24229 26757
rect 24163 26692 24164 26756
rect 24228 26692 24229 26756
rect 24163 26691 24229 26692
rect 22507 25668 22573 25669
rect 22507 25604 22508 25668
rect 22572 25604 22573 25668
rect 22507 25603 22573 25604
rect 19931 25124 19997 25125
rect 19931 25060 19932 25124
rect 19996 25060 19997 25124
rect 19931 25059 19997 25060
rect 3371 24988 3437 24989
rect 3371 24924 3372 24988
rect 3436 24924 3437 24988
rect 3371 24923 3437 24924
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 3374 18597 3434 24923
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 3923 23764 3989 23765
rect 3923 23700 3924 23764
rect 3988 23700 3989 23764
rect 3923 23699 3989 23700
rect 3371 18596 3437 18597
rect 3371 18532 3372 18596
rect 3436 18532 3437 18596
rect 3371 18531 3437 18532
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 3374 13701 3434 18531
rect 3555 18188 3621 18189
rect 3555 18124 3556 18188
rect 3620 18124 3621 18188
rect 3555 18123 3621 18124
rect 3371 13700 3437 13701
rect 3371 13636 3372 13700
rect 3436 13636 3437 13700
rect 3371 13635 3437 13636
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 3558 12885 3618 18123
rect 3926 13021 3986 23699
rect 7603 23628 7669 23629
rect 7603 23564 7604 23628
rect 7668 23564 7669 23628
rect 7603 23563 7669 23564
rect 4291 23492 4357 23493
rect 4291 23428 4292 23492
rect 4356 23428 4357 23492
rect 4291 23427 4357 23428
rect 4294 13565 4354 23427
rect 5211 23084 5277 23085
rect 5211 23020 5212 23084
rect 5276 23020 5277 23084
rect 5211 23019 5277 23020
rect 4291 13564 4357 13565
rect 4291 13500 4292 13564
rect 4356 13500 4357 13564
rect 4291 13499 4357 13500
rect 3923 13020 3989 13021
rect 3923 12956 3924 13020
rect 3988 12956 3989 13020
rect 3923 12955 3989 12956
rect 3555 12884 3621 12885
rect 3555 12820 3556 12884
rect 3620 12820 3621 12884
rect 3555 12819 3621 12820
rect 4294 12613 4354 13499
rect 4291 12612 4357 12613
rect 4291 12548 4292 12612
rect 4356 12548 4357 12612
rect 4291 12547 4357 12548
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 5214 10301 5274 23019
rect 5763 22676 5829 22677
rect 5763 22612 5764 22676
rect 5828 22612 5829 22676
rect 5763 22611 5829 22612
rect 5579 21996 5645 21997
rect 5579 21932 5580 21996
rect 5644 21932 5645 21996
rect 5579 21931 5645 21932
rect 5582 19005 5642 21931
rect 5579 19004 5645 19005
rect 5579 18940 5580 19004
rect 5644 18940 5645 19004
rect 5579 18939 5645 18940
rect 5582 13701 5642 18939
rect 5579 13700 5645 13701
rect 5579 13636 5580 13700
rect 5644 13636 5645 13700
rect 5579 13635 5645 13636
rect 5766 11797 5826 22611
rect 7419 21724 7485 21725
rect 7419 21660 7420 21724
rect 7484 21660 7485 21724
rect 7419 21659 7485 21660
rect 6315 18460 6381 18461
rect 6315 18396 6316 18460
rect 6380 18396 6381 18460
rect 6315 18395 6381 18396
rect 6318 14381 6378 18395
rect 6315 14380 6381 14381
rect 6315 14316 6316 14380
rect 6380 14316 6381 14380
rect 6315 14315 6381 14316
rect 6318 13837 6378 14315
rect 6315 13836 6381 13837
rect 6315 13772 6316 13836
rect 6380 13772 6381 13836
rect 6315 13771 6381 13772
rect 5763 11796 5829 11797
rect 5763 11732 5764 11796
rect 5828 11732 5829 11796
rect 5763 11731 5829 11732
rect 7422 10301 7482 21659
rect 5211 10300 5277 10301
rect 5211 10236 5212 10300
rect 5276 10236 5277 10300
rect 5211 10235 5277 10236
rect 7419 10300 7485 10301
rect 7419 10236 7420 10300
rect 7484 10236 7485 10300
rect 7419 10235 7485 10236
rect 7606 9621 7666 23563
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 17944 23968 18264 24528
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17171 23492 17237 23493
rect 17171 23428 17172 23492
rect 17236 23428 17237 23492
rect 17171 23427 17237 23428
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 9259 22812 9325 22813
rect 9259 22748 9260 22812
rect 9324 22748 9325 22812
rect 9259 22747 9325 22748
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 8891 20364 8957 20365
rect 8891 20300 8892 20364
rect 8956 20300 8957 20364
rect 8891 20299 8957 20300
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 8339 18732 8405 18733
rect 8339 18668 8340 18732
rect 8404 18668 8405 18732
rect 8339 18667 8405 18668
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 8342 10437 8402 18667
rect 8894 11117 8954 20299
rect 9075 17644 9141 17645
rect 9075 17580 9076 17644
rect 9140 17580 9141 17644
rect 9075 17579 9141 17580
rect 9078 12749 9138 17579
rect 9262 14653 9322 22747
rect 9811 22404 9877 22405
rect 9811 22340 9812 22404
rect 9876 22340 9877 22404
rect 9811 22339 9877 22340
rect 9443 17508 9509 17509
rect 9443 17444 9444 17508
rect 9508 17444 9509 17508
rect 9443 17443 9509 17444
rect 9259 14652 9325 14653
rect 9259 14588 9260 14652
rect 9324 14588 9325 14652
rect 9259 14587 9325 14588
rect 9075 12748 9141 12749
rect 9075 12684 9076 12748
rect 9140 12684 9141 12748
rect 9075 12683 9141 12684
rect 8891 11116 8957 11117
rect 8891 11052 8892 11116
rect 8956 11052 8957 11116
rect 8891 11051 8957 11052
rect 8339 10436 8405 10437
rect 8339 10372 8340 10436
rect 8404 10372 8405 10436
rect 8339 10371 8405 10372
rect 9446 10301 9506 17443
rect 9814 12341 9874 22339
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 11467 22132 11533 22133
rect 11467 22068 11468 22132
rect 11532 22068 11533 22132
rect 11467 22067 11533 22068
rect 10179 21452 10245 21453
rect 10179 21388 10180 21452
rect 10244 21388 10245 21452
rect 10179 21387 10245 21388
rect 9995 17916 10061 17917
rect 9995 17852 9996 17916
rect 10060 17852 10061 17916
rect 9995 17851 10061 17852
rect 9811 12340 9877 12341
rect 9811 12276 9812 12340
rect 9876 12276 9877 12340
rect 9811 12275 9877 12276
rect 9627 11116 9693 11117
rect 9627 11052 9628 11116
rect 9692 11052 9693 11116
rect 9627 11051 9693 11052
rect 9443 10300 9509 10301
rect 9443 10236 9444 10300
rect 9508 10236 9509 10300
rect 9443 10235 9509 10236
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7603 9620 7669 9621
rect 7603 9556 7604 9620
rect 7668 9556 7669 9620
rect 7603 9555 7669 9556
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 8736 8264 9760
rect 9630 9077 9690 11051
rect 9627 9076 9693 9077
rect 9627 9012 9628 9076
rect 9692 9012 9693 9076
rect 9627 9011 9693 9012
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 9998 8261 10058 17851
rect 9995 8260 10061 8261
rect 9995 8196 9996 8260
rect 10060 8196 10061 8260
rect 9995 8195 10061 8196
rect 10182 7989 10242 21387
rect 11099 19548 11165 19549
rect 11099 19484 11100 19548
rect 11164 19484 11165 19548
rect 11099 19483 11165 19484
rect 11102 15741 11162 19483
rect 11099 15740 11165 15741
rect 11099 15676 11100 15740
rect 11164 15676 11165 15740
rect 11099 15675 11165 15676
rect 10179 7988 10245 7989
rect 10179 7924 10180 7988
rect 10244 7924 10245 7988
rect 10179 7923 10245 7924
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 11470 6901 11530 22067
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12571 20908 12637 20909
rect 12571 20844 12572 20908
rect 12636 20844 12637 20908
rect 12571 20843 12637 20844
rect 12203 19140 12269 19141
rect 12203 19076 12204 19140
rect 12268 19076 12269 19140
rect 12203 19075 12269 19076
rect 12019 15060 12085 15061
rect 12019 14996 12020 15060
rect 12084 14996 12085 15060
rect 12019 14995 12085 14996
rect 11651 13564 11717 13565
rect 11651 13500 11652 13564
rect 11716 13500 11717 13564
rect 11651 13499 11717 13500
rect 11654 12749 11714 13499
rect 11651 12748 11717 12749
rect 11651 12684 11652 12748
rect 11716 12684 11717 12748
rect 11651 12683 11717 12684
rect 12022 9621 12082 14995
rect 12019 9620 12085 9621
rect 12019 9556 12020 9620
rect 12084 9556 12085 9620
rect 12019 9555 12085 9556
rect 11467 6900 11533 6901
rect 11467 6836 11468 6900
rect 11532 6836 11533 6900
rect 11467 6835 11533 6836
rect 12206 6765 12266 19075
rect 12574 9349 12634 20843
rect 12944 20160 13264 21184
rect 15699 20772 15765 20773
rect 15699 20708 15700 20772
rect 15764 20708 15765 20772
rect 15699 20707 15765 20708
rect 16987 20772 17053 20773
rect 16987 20708 16988 20772
rect 17052 20708 17053 20772
rect 16987 20707 17053 20708
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 15147 19684 15213 19685
rect 15147 19620 15148 19684
rect 15212 19620 15213 19684
rect 15147 19619 15213 19620
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 14963 18052 15029 18053
rect 14963 17988 14964 18052
rect 15028 17988 15029 18052
rect 14963 17987 15029 17988
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 13675 17780 13741 17781
rect 13675 17716 13676 17780
rect 13740 17716 13741 17780
rect 13675 17715 13741 17716
rect 13678 16965 13738 17715
rect 13675 16964 13741 16965
rect 13675 16900 13676 16964
rect 13740 16900 13741 16964
rect 13675 16899 13741 16900
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 14779 16692 14845 16693
rect 14779 16628 14780 16692
rect 14844 16628 14845 16692
rect 14779 16627 14845 16628
rect 14043 16012 14109 16013
rect 14043 15948 14044 16012
rect 14108 15948 14109 16012
rect 14043 15947 14109 15948
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 13859 14244 13925 14245
rect 13859 14180 13860 14244
rect 13924 14180 13925 14244
rect 13859 14179 13925 14180
rect 13491 13700 13557 13701
rect 13491 13636 13492 13700
rect 13556 13636 13557 13700
rect 13491 13635 13557 13636
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 13494 10573 13554 13635
rect 13675 12476 13741 12477
rect 13675 12412 13676 12476
rect 13740 12412 13741 12476
rect 13675 12411 13741 12412
rect 13678 11797 13738 12411
rect 13862 12069 13922 14179
rect 13859 12068 13925 12069
rect 13859 12004 13860 12068
rect 13924 12004 13925 12068
rect 13859 12003 13925 12004
rect 13675 11796 13741 11797
rect 13675 11732 13676 11796
rect 13740 11732 13741 11796
rect 13675 11731 13741 11732
rect 13491 10572 13557 10573
rect 13491 10508 13492 10572
rect 13556 10508 13557 10572
rect 13491 10507 13557 10508
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12571 9348 12637 9349
rect 12571 9284 12572 9348
rect 12636 9284 12637 9348
rect 12571 9283 12637 9284
rect 12944 9280 13264 10304
rect 14046 9757 14106 15947
rect 14043 9756 14109 9757
rect 14043 9692 14044 9756
rect 14108 9692 14109 9756
rect 14043 9691 14109 9692
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 14782 8125 14842 16627
rect 14779 8124 14845 8125
rect 14779 8060 14780 8124
rect 14844 8060 14845 8124
rect 14779 8059 14845 8060
rect 14966 7717 15026 17987
rect 15150 16149 15210 19619
rect 15331 18052 15397 18053
rect 15331 17988 15332 18052
rect 15396 17988 15397 18052
rect 15331 17987 15397 17988
rect 15147 16148 15213 16149
rect 15147 16084 15148 16148
rect 15212 16084 15213 16148
rect 15147 16083 15213 16084
rect 15334 13970 15394 17987
rect 15150 13910 15394 13970
rect 15150 13157 15210 13910
rect 15147 13156 15213 13157
rect 15147 13092 15148 13156
rect 15212 13092 15213 13156
rect 15147 13091 15213 13092
rect 15702 8397 15762 20707
rect 16067 16420 16133 16421
rect 16067 16356 16068 16420
rect 16132 16356 16133 16420
rect 16067 16355 16133 16356
rect 16070 9893 16130 16355
rect 16435 14788 16501 14789
rect 16435 14724 16436 14788
rect 16500 14724 16501 14788
rect 16435 14723 16501 14724
rect 16251 13292 16317 13293
rect 16251 13228 16252 13292
rect 16316 13228 16317 13292
rect 16251 13227 16317 13228
rect 16254 13021 16314 13227
rect 16251 13020 16317 13021
rect 16251 12956 16252 13020
rect 16316 12956 16317 13020
rect 16251 12955 16317 12956
rect 16254 11117 16314 12955
rect 16438 12205 16498 14723
rect 16435 12204 16501 12205
rect 16435 12140 16436 12204
rect 16500 12140 16501 12204
rect 16435 12139 16501 12140
rect 16251 11116 16317 11117
rect 16251 11052 16252 11116
rect 16316 11052 16317 11116
rect 16251 11051 16317 11052
rect 16067 9892 16133 9893
rect 16067 9828 16068 9892
rect 16132 9828 16133 9892
rect 16067 9827 16133 9828
rect 15699 8396 15765 8397
rect 15699 8332 15700 8396
rect 15764 8332 15765 8396
rect 15699 8331 15765 8332
rect 16254 8261 16314 11051
rect 16251 8260 16317 8261
rect 16251 8196 16252 8260
rect 16316 8196 16317 8260
rect 16251 8195 16317 8196
rect 16438 7989 16498 12139
rect 16619 10300 16685 10301
rect 16619 10236 16620 10300
rect 16684 10236 16685 10300
rect 16619 10235 16685 10236
rect 16435 7988 16501 7989
rect 16435 7924 16436 7988
rect 16500 7924 16501 7988
rect 16435 7923 16501 7924
rect 14963 7716 15029 7717
rect 14963 7652 14964 7716
rect 15028 7652 15029 7716
rect 14963 7651 15029 7652
rect 16622 7581 16682 10235
rect 16990 9757 17050 20707
rect 16987 9756 17053 9757
rect 16987 9692 16988 9756
rect 17052 9692 17053 9756
rect 16987 9691 17053 9692
rect 16619 7580 16685 7581
rect 16619 7516 16620 7580
rect 16684 7516 16685 7580
rect 16619 7515 16685 7516
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12203 6764 12269 6765
rect 12203 6700 12204 6764
rect 12268 6700 12269 6764
rect 12203 6699 12269 6700
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 17174 5269 17234 23427
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 19379 20772 19445 20773
rect 19379 20708 19380 20772
rect 19444 20708 19445 20772
rect 19379 20707 19445 20708
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 18459 17644 18525 17645
rect 18459 17580 18460 17644
rect 18524 17580 18525 17644
rect 18459 17579 18525 17580
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17355 16692 17421 16693
rect 17355 16628 17356 16692
rect 17420 16628 17421 16692
rect 17355 16627 17421 16628
rect 17358 8669 17418 16627
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 18462 14925 18522 17579
rect 18643 16964 18709 16965
rect 18643 16900 18644 16964
rect 18708 16900 18709 16964
rect 18643 16899 18709 16900
rect 18646 16285 18706 16899
rect 18643 16284 18709 16285
rect 18643 16220 18644 16284
rect 18708 16220 18709 16284
rect 18643 16219 18709 16220
rect 18459 14924 18525 14925
rect 18459 14860 18460 14924
rect 18524 14860 18525 14924
rect 18459 14859 18525 14860
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 18459 11524 18525 11525
rect 18459 11460 18460 11524
rect 18524 11460 18525 11524
rect 18459 11459 18525 11460
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17355 8668 17421 8669
rect 17355 8604 17356 8668
rect 17420 8604 17421 8668
rect 17355 8603 17421 8604
rect 17944 7648 18264 8672
rect 18462 8533 18522 11459
rect 18646 11253 18706 16219
rect 18643 11252 18709 11253
rect 18643 11188 18644 11252
rect 18708 11188 18709 11252
rect 18643 11187 18709 11188
rect 18646 9213 18706 11187
rect 19382 10301 19442 20707
rect 19934 19141 19994 25059
rect 20667 23492 20733 23493
rect 20667 23428 20668 23492
rect 20732 23428 20733 23492
rect 20667 23427 20733 23428
rect 19931 19140 19997 19141
rect 19931 19076 19932 19140
rect 19996 19076 19997 19140
rect 19931 19075 19997 19076
rect 19563 18052 19629 18053
rect 19563 17988 19564 18052
rect 19628 17988 19629 18052
rect 19563 17987 19629 17988
rect 19379 10300 19445 10301
rect 19379 10236 19380 10300
rect 19444 10236 19445 10300
rect 19379 10235 19445 10236
rect 18643 9212 18709 9213
rect 18643 9148 18644 9212
rect 18708 9148 18709 9212
rect 18643 9147 18709 9148
rect 18643 8804 18709 8805
rect 18643 8740 18644 8804
rect 18708 8740 18709 8804
rect 18643 8739 18709 8740
rect 18459 8532 18525 8533
rect 18459 8468 18460 8532
rect 18524 8468 18525 8532
rect 18459 8467 18525 8468
rect 18646 8261 18706 8739
rect 18643 8260 18709 8261
rect 18643 8196 18644 8260
rect 18708 8196 18709 8260
rect 18643 8195 18709 8196
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 19566 7173 19626 17987
rect 19563 7172 19629 7173
rect 19563 7108 19564 7172
rect 19628 7108 19629 7172
rect 19563 7107 19629 7108
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 20670 6221 20730 23427
rect 21219 23356 21285 23357
rect 21219 23292 21220 23356
rect 21284 23292 21285 23356
rect 21219 23291 21285 23292
rect 21222 6357 21282 23291
rect 22139 22812 22205 22813
rect 22139 22748 22140 22812
rect 22204 22748 22205 22812
rect 22139 22747 22205 22748
rect 22142 8397 22202 22747
rect 22323 21860 22389 21861
rect 22323 21796 22324 21860
rect 22388 21796 22389 21860
rect 22323 21795 22389 21796
rect 22326 19413 22386 21795
rect 22323 19412 22389 19413
rect 22323 19348 22324 19412
rect 22388 19348 22389 19412
rect 22323 19347 22389 19348
rect 22510 16285 22570 25603
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 23427 23492 23493 23493
rect 23427 23428 23428 23492
rect 23492 23428 23493 23492
rect 23427 23427 23493 23428
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22507 16284 22573 16285
rect 22507 16220 22508 16284
rect 22572 16220 22573 16284
rect 22507 16219 22573 16220
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22139 8396 22205 8397
rect 22139 8332 22140 8396
rect 22204 8332 22205 8396
rect 22139 8331 22205 8332
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 23430 7853 23490 23427
rect 23795 22268 23861 22269
rect 23795 22204 23796 22268
rect 23860 22204 23861 22268
rect 23795 22203 23861 22204
rect 23427 7852 23493 7853
rect 23427 7788 23428 7852
rect 23492 7788 23493 7852
rect 23427 7787 23493 7788
rect 23798 7445 23858 22203
rect 24166 21725 24226 26691
rect 47163 26620 47229 26621
rect 47163 26556 47164 26620
rect 47228 26556 47229 26620
rect 47163 26555 47229 26556
rect 46059 26212 46125 26213
rect 46059 26148 46060 26212
rect 46124 26148 46125 26212
rect 46059 26147 46125 26148
rect 30051 25940 30117 25941
rect 30051 25876 30052 25940
rect 30116 25876 30117 25940
rect 30051 25875 30117 25876
rect 24899 24988 24965 24989
rect 24899 24924 24900 24988
rect 24964 24924 24965 24988
rect 24899 24923 24965 24924
rect 24163 21724 24229 21725
rect 24163 21660 24164 21724
rect 24228 21660 24229 21724
rect 24163 21659 24229 21660
rect 24902 19005 24962 24923
rect 27944 23968 28264 24528
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 27475 23492 27541 23493
rect 27475 23428 27476 23492
rect 27540 23428 27541 23492
rect 27475 23427 27541 23428
rect 27291 22676 27357 22677
rect 27291 22612 27292 22676
rect 27356 22612 27357 22676
rect 27291 22611 27357 22612
rect 26003 22404 26069 22405
rect 26003 22340 26004 22404
rect 26068 22340 26069 22404
rect 26003 22339 26069 22340
rect 24899 19004 24965 19005
rect 24899 18940 24900 19004
rect 24964 18940 24965 19004
rect 24899 18939 24965 18940
rect 24899 18052 24965 18053
rect 24899 17988 24900 18052
rect 24964 17988 24965 18052
rect 24899 17987 24965 17988
rect 24902 13837 24962 17987
rect 24899 13836 24965 13837
rect 24899 13772 24900 13836
rect 24964 13772 24965 13836
rect 24899 13771 24965 13772
rect 24902 7717 24962 13771
rect 26006 10573 26066 22339
rect 26555 21316 26621 21317
rect 26555 21252 26556 21316
rect 26620 21252 26621 21316
rect 26555 21251 26621 21252
rect 26558 18053 26618 21251
rect 27107 18868 27173 18869
rect 27107 18804 27108 18868
rect 27172 18804 27173 18868
rect 27107 18803 27173 18804
rect 26555 18052 26621 18053
rect 26555 17988 26556 18052
rect 26620 17988 26621 18052
rect 26555 17987 26621 17988
rect 26923 17644 26989 17645
rect 26923 17580 26924 17644
rect 26988 17580 26989 17644
rect 26923 17579 26989 17580
rect 26739 14924 26805 14925
rect 26739 14860 26740 14924
rect 26804 14860 26805 14924
rect 26739 14859 26805 14860
rect 26742 12069 26802 14859
rect 26926 12341 26986 17579
rect 27110 17373 27170 18803
rect 27107 17372 27173 17373
rect 27107 17308 27108 17372
rect 27172 17308 27173 17372
rect 27107 17307 27173 17308
rect 26923 12340 26989 12341
rect 26923 12276 26924 12340
rect 26988 12276 26989 12340
rect 26923 12275 26989 12276
rect 26739 12068 26805 12069
rect 26739 12004 26740 12068
rect 26804 12004 26805 12068
rect 26739 12003 26805 12004
rect 27107 12068 27173 12069
rect 27107 12004 27108 12068
rect 27172 12004 27173 12068
rect 27107 12003 27173 12004
rect 26003 10572 26069 10573
rect 26003 10508 26004 10572
rect 26068 10508 26069 10572
rect 26003 10507 26069 10508
rect 24899 7716 24965 7717
rect 24899 7652 24900 7716
rect 24964 7652 24965 7716
rect 24899 7651 24965 7652
rect 23795 7444 23861 7445
rect 23795 7380 23796 7444
rect 23860 7380 23861 7444
rect 23795 7379 23861 7380
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 21219 6356 21285 6357
rect 21219 6292 21220 6356
rect 21284 6292 21285 6356
rect 21219 6291 21285 6292
rect 20667 6220 20733 6221
rect 20667 6156 20668 6220
rect 20732 6156 20733 6220
rect 20667 6155 20733 6156
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17171 5268 17237 5269
rect 17171 5204 17172 5268
rect 17236 5204 17237 5268
rect 17171 5203 17237 5204
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 27110 5677 27170 12003
rect 27294 11525 27354 22611
rect 27478 17917 27538 23427
rect 27944 22880 28264 23904
rect 28763 23492 28829 23493
rect 28763 23428 28764 23492
rect 28828 23428 28829 23492
rect 28763 23427 28829 23428
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27659 19004 27725 19005
rect 27659 18940 27660 19004
rect 27724 18940 27725 19004
rect 27659 18939 27725 18940
rect 27475 17916 27541 17917
rect 27475 17852 27476 17916
rect 27540 17852 27541 17916
rect 27475 17851 27541 17852
rect 27291 11524 27357 11525
rect 27291 11460 27292 11524
rect 27356 11460 27357 11524
rect 27291 11459 27357 11460
rect 27291 11388 27357 11389
rect 27291 11324 27292 11388
rect 27356 11324 27357 11388
rect 27291 11323 27357 11324
rect 27294 9757 27354 11323
rect 27291 9756 27357 9757
rect 27291 9692 27292 9756
rect 27356 9692 27357 9756
rect 27291 9691 27357 9692
rect 27478 5813 27538 17851
rect 27662 16965 27722 18939
rect 27944 18528 28264 19552
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27944 17440 28264 18464
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27659 16964 27725 16965
rect 27659 16900 27660 16964
rect 27724 16900 27725 16964
rect 27659 16899 27725 16900
rect 27944 16352 28264 17376
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27944 14176 28264 15200
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27475 5812 27541 5813
rect 27475 5748 27476 5812
rect 27540 5748 27541 5812
rect 27475 5747 27541 5748
rect 27107 5676 27173 5677
rect 27107 5612 27108 5676
rect 27172 5612 27173 5676
rect 27107 5611 27173 5612
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 27944 5472 28264 6496
rect 28766 6493 28826 23427
rect 30054 23357 30114 25875
rect 44219 25124 44285 25125
rect 44219 25060 44220 25124
rect 44284 25060 44285 25124
rect 44219 25059 44285 25060
rect 34651 24580 34717 24581
rect 32944 24512 33264 24528
rect 34651 24516 34652 24580
rect 34716 24516 34717 24580
rect 34651 24515 34717 24516
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 30235 23492 30301 23493
rect 30235 23428 30236 23492
rect 30300 23428 30301 23492
rect 30235 23427 30301 23428
rect 30971 23492 31037 23493
rect 30971 23428 30972 23492
rect 31036 23428 31037 23492
rect 30971 23427 31037 23428
rect 31523 23492 31589 23493
rect 31523 23428 31524 23492
rect 31588 23428 31589 23492
rect 31523 23427 31589 23428
rect 32443 23492 32509 23493
rect 32443 23428 32444 23492
rect 32508 23428 32509 23492
rect 32443 23427 32509 23428
rect 30051 23356 30117 23357
rect 30051 23292 30052 23356
rect 30116 23292 30117 23356
rect 30051 23291 30117 23292
rect 29315 22268 29381 22269
rect 29315 22204 29316 22268
rect 29380 22204 29381 22268
rect 29315 22203 29381 22204
rect 28947 21996 29013 21997
rect 28947 21932 28948 21996
rect 29012 21932 29013 21996
rect 28947 21931 29013 21932
rect 28950 14109 29010 21931
rect 29318 20093 29378 22203
rect 29315 20092 29381 20093
rect 29315 20028 29316 20092
rect 29380 20028 29381 20092
rect 29315 20027 29381 20028
rect 29499 19412 29565 19413
rect 29499 19348 29500 19412
rect 29564 19348 29565 19412
rect 29499 19347 29565 19348
rect 29502 16557 29562 19347
rect 29499 16556 29565 16557
rect 29499 16492 29500 16556
rect 29564 16492 29565 16556
rect 29499 16491 29565 16492
rect 28947 14108 29013 14109
rect 28947 14044 28948 14108
rect 29012 14044 29013 14108
rect 28947 14043 29013 14044
rect 29502 6901 29562 16491
rect 30238 7309 30298 23427
rect 30974 10981 31034 23427
rect 31339 22132 31405 22133
rect 31339 22068 31340 22132
rect 31404 22068 31405 22132
rect 31339 22067 31405 22068
rect 31155 15196 31221 15197
rect 31155 15132 31156 15196
rect 31220 15132 31221 15196
rect 31155 15131 31221 15132
rect 31158 13837 31218 15131
rect 31155 13836 31221 13837
rect 31155 13772 31156 13836
rect 31220 13772 31221 13836
rect 31155 13771 31221 13772
rect 30971 10980 31037 10981
rect 30971 10916 30972 10980
rect 31036 10916 31037 10980
rect 30971 10915 31037 10916
rect 30235 7308 30301 7309
rect 30235 7244 30236 7308
rect 30300 7244 30301 7308
rect 30235 7243 30301 7244
rect 29499 6900 29565 6901
rect 29499 6836 29500 6900
rect 29564 6836 29565 6900
rect 29499 6835 29565 6836
rect 28763 6492 28829 6493
rect 28763 6428 28764 6492
rect 28828 6428 28829 6492
rect 28763 6427 28829 6428
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 31342 4725 31402 22067
rect 31526 14517 31586 23427
rect 31891 19004 31957 19005
rect 31891 18940 31892 19004
rect 31956 18940 31957 19004
rect 31891 18939 31957 18940
rect 31894 16421 31954 18939
rect 31891 16420 31957 16421
rect 31891 16356 31892 16420
rect 31956 16356 31957 16420
rect 31891 16355 31957 16356
rect 31523 14516 31589 14517
rect 31523 14452 31524 14516
rect 31588 14452 31589 14516
rect 31523 14451 31589 14452
rect 32259 11524 32325 11525
rect 32259 11460 32260 11524
rect 32324 11460 32325 11524
rect 32259 11459 32325 11460
rect 32262 8941 32322 11459
rect 32446 11253 32506 23427
rect 32944 23424 33264 24448
rect 34467 23900 34533 23901
rect 34467 23836 34468 23900
rect 34532 23836 34533 23900
rect 34467 23835 34533 23836
rect 34099 23492 34165 23493
rect 34099 23428 34100 23492
rect 34164 23428 34165 23492
rect 34099 23427 34165 23428
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 32944 19072 33264 20096
rect 33547 19140 33613 19141
rect 33547 19076 33548 19140
rect 33612 19076 33613 19140
rect 33547 19075 33613 19076
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32627 17916 32693 17917
rect 32627 17852 32628 17916
rect 32692 17852 32693 17916
rect 32627 17851 32693 17852
rect 32630 11661 32690 17851
rect 32944 16896 33264 17920
rect 33363 17100 33429 17101
rect 33363 17036 33364 17100
rect 33428 17036 33429 17100
rect 33363 17035 33429 17036
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32811 16148 32877 16149
rect 32811 16084 32812 16148
rect 32876 16084 32877 16148
rect 32811 16083 32877 16084
rect 32627 11660 32693 11661
rect 32627 11596 32628 11660
rect 32692 11596 32693 11660
rect 32627 11595 32693 11596
rect 32814 11389 32874 16083
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32811 11388 32877 11389
rect 32811 11324 32812 11388
rect 32876 11324 32877 11388
rect 32811 11323 32877 11324
rect 32443 11252 32509 11253
rect 32443 11188 32444 11252
rect 32508 11188 32509 11252
rect 32443 11187 32509 11188
rect 32944 10368 33264 11392
rect 33366 11389 33426 17035
rect 33550 13973 33610 19075
rect 33547 13972 33613 13973
rect 33547 13908 33548 13972
rect 33612 13908 33613 13972
rect 33547 13907 33613 13908
rect 33363 11388 33429 11389
rect 33363 11324 33364 11388
rect 33428 11324 33429 11388
rect 33363 11323 33429 11324
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32259 8940 32325 8941
rect 32259 8876 32260 8940
rect 32324 8876 32325 8940
rect 32259 8875 32325 8876
rect 32944 8192 33264 9216
rect 34102 8397 34162 23427
rect 34283 22812 34349 22813
rect 34283 22748 34284 22812
rect 34348 22748 34349 22812
rect 34283 22747 34349 22748
rect 34286 16557 34346 22747
rect 34470 20501 34530 23835
rect 34654 23629 34714 24515
rect 37944 23968 38264 24528
rect 42944 24512 43264 24528
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 40355 24036 40421 24037
rect 40355 23972 40356 24036
rect 40420 23972 40421 24036
rect 40355 23971 40421 23972
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 34651 23628 34717 23629
rect 34651 23564 34652 23628
rect 34716 23564 34717 23628
rect 34651 23563 34717 23564
rect 36491 23628 36557 23629
rect 36491 23564 36492 23628
rect 36556 23564 36557 23628
rect 36491 23563 36557 23564
rect 34467 20500 34533 20501
rect 34467 20436 34468 20500
rect 34532 20436 34533 20500
rect 34467 20435 34533 20436
rect 34654 20365 34714 23563
rect 34835 23220 34901 23221
rect 34835 23156 34836 23220
rect 34900 23156 34901 23220
rect 34835 23155 34901 23156
rect 34651 20364 34717 20365
rect 34651 20300 34652 20364
rect 34716 20300 34717 20364
rect 34651 20299 34717 20300
rect 34467 19276 34533 19277
rect 34467 19212 34468 19276
rect 34532 19212 34533 19276
rect 34467 19211 34533 19212
rect 34470 16965 34530 19211
rect 34467 16964 34533 16965
rect 34467 16900 34468 16964
rect 34532 16900 34533 16964
rect 34467 16899 34533 16900
rect 34283 16556 34349 16557
rect 34283 16492 34284 16556
rect 34348 16492 34349 16556
rect 34283 16491 34349 16492
rect 34283 12068 34349 12069
rect 34283 12004 34284 12068
rect 34348 12004 34349 12068
rect 34283 12003 34349 12004
rect 34286 11117 34346 12003
rect 34467 11252 34533 11253
rect 34467 11188 34468 11252
rect 34532 11188 34533 11252
rect 34467 11187 34533 11188
rect 34283 11116 34349 11117
rect 34283 11052 34284 11116
rect 34348 11052 34349 11116
rect 34283 11051 34349 11052
rect 34286 9621 34346 11051
rect 34470 10165 34530 11187
rect 34467 10164 34533 10165
rect 34467 10100 34468 10164
rect 34532 10100 34533 10164
rect 34467 10099 34533 10100
rect 34283 9620 34349 9621
rect 34283 9556 34284 9620
rect 34348 9556 34349 9620
rect 34283 9555 34349 9556
rect 34838 9349 34898 23155
rect 35939 21996 36005 21997
rect 35939 21932 35940 21996
rect 36004 21932 36005 21996
rect 35939 21931 36005 21932
rect 35755 21588 35821 21589
rect 35755 21524 35756 21588
rect 35820 21524 35821 21588
rect 35755 21523 35821 21524
rect 35203 20500 35269 20501
rect 35203 20436 35204 20500
rect 35268 20436 35269 20500
rect 35203 20435 35269 20436
rect 35019 13292 35085 13293
rect 35019 13228 35020 13292
rect 35084 13228 35085 13292
rect 35019 13227 35085 13228
rect 35022 11525 35082 13227
rect 35206 12341 35266 20435
rect 35387 20364 35453 20365
rect 35387 20300 35388 20364
rect 35452 20300 35453 20364
rect 35387 20299 35453 20300
rect 35203 12340 35269 12341
rect 35203 12276 35204 12340
rect 35268 12276 35269 12340
rect 35203 12275 35269 12276
rect 35019 11524 35085 11525
rect 35019 11460 35020 11524
rect 35084 11460 35085 11524
rect 35019 11459 35085 11460
rect 34835 9348 34901 9349
rect 34835 9284 34836 9348
rect 34900 9284 34901 9348
rect 34835 9283 34901 9284
rect 34099 8396 34165 8397
rect 34099 8332 34100 8396
rect 34164 8332 34165 8396
rect 34099 8331 34165 8332
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 31339 4724 31405 4725
rect 31339 4660 31340 4724
rect 31404 4660 31405 4724
rect 31339 4659 31405 4660
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 3840 33264 4864
rect 35390 4589 35450 20299
rect 35758 16693 35818 21523
rect 35942 17781 36002 21931
rect 35939 17780 36005 17781
rect 35939 17716 35940 17780
rect 36004 17716 36005 17780
rect 35939 17715 36005 17716
rect 35755 16692 35821 16693
rect 35755 16628 35756 16692
rect 35820 16628 35821 16692
rect 35755 16627 35821 16628
rect 36494 4997 36554 23563
rect 36675 23492 36741 23493
rect 36675 23428 36676 23492
rect 36740 23428 36741 23492
rect 36675 23427 36741 23428
rect 36678 5133 36738 23427
rect 37411 23356 37477 23357
rect 37411 23292 37412 23356
rect 37476 23292 37477 23356
rect 37411 23291 37477 23292
rect 36859 18732 36925 18733
rect 36859 18668 36860 18732
rect 36924 18668 36925 18732
rect 36859 18667 36925 18668
rect 36862 16965 36922 18667
rect 37043 18460 37109 18461
rect 37043 18396 37044 18460
rect 37108 18396 37109 18460
rect 37043 18395 37109 18396
rect 36859 16964 36925 16965
rect 36859 16900 36860 16964
rect 36924 16900 36925 16964
rect 36859 16899 36925 16900
rect 37046 10845 37106 18395
rect 37227 12340 37293 12341
rect 37227 12276 37228 12340
rect 37292 12276 37293 12340
rect 37227 12275 37293 12276
rect 37043 10844 37109 10845
rect 37043 10780 37044 10844
rect 37108 10780 37109 10844
rect 37043 10779 37109 10780
rect 37230 5949 37290 12275
rect 37414 9077 37474 23291
rect 37944 22880 38264 23904
rect 38515 23492 38581 23493
rect 38515 23428 38516 23492
rect 38580 23428 38581 23492
rect 38515 23427 38581 23428
rect 39435 23492 39501 23493
rect 39435 23428 39436 23492
rect 39500 23428 39501 23492
rect 39435 23427 39501 23428
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37595 22404 37661 22405
rect 37595 22340 37596 22404
rect 37660 22340 37661 22404
rect 37595 22339 37661 22340
rect 37598 14925 37658 22339
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 38331 18052 38397 18053
rect 38331 17988 38332 18052
rect 38396 17988 38397 18052
rect 38331 17987 38397 17988
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37595 14924 37661 14925
rect 37595 14860 37596 14924
rect 37660 14860 37661 14924
rect 37595 14859 37661 14860
rect 37944 14176 38264 15200
rect 38334 14245 38394 17987
rect 38331 14244 38397 14245
rect 38331 14180 38332 14244
rect 38396 14180 38397 14244
rect 38331 14179 38397 14180
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 38331 12340 38397 12341
rect 38331 12276 38332 12340
rect 38396 12276 38397 12340
rect 38331 12275 38397 12276
rect 38334 12069 38394 12275
rect 38331 12068 38397 12069
rect 38331 12004 38332 12068
rect 38396 12004 38397 12068
rect 38331 12003 38397 12004
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37411 9076 37477 9077
rect 37411 9012 37412 9076
rect 37476 9012 37477 9076
rect 37411 9011 37477 9012
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 38518 7717 38578 23427
rect 39067 21860 39133 21861
rect 39067 21796 39068 21860
rect 39132 21796 39133 21860
rect 39067 21795 39133 21796
rect 38883 19956 38949 19957
rect 38883 19892 38884 19956
rect 38948 19892 38949 19956
rect 38883 19891 38949 19892
rect 38886 19549 38946 19891
rect 38883 19548 38949 19549
rect 38883 19484 38884 19548
rect 38948 19484 38949 19548
rect 38883 19483 38949 19484
rect 38883 18596 38949 18597
rect 38883 18532 38884 18596
rect 38948 18532 38949 18596
rect 38883 18531 38949 18532
rect 38699 16828 38765 16829
rect 38699 16764 38700 16828
rect 38764 16764 38765 16828
rect 38699 16763 38765 16764
rect 38702 11797 38762 16763
rect 38886 15197 38946 18531
rect 38883 15196 38949 15197
rect 38883 15132 38884 15196
rect 38948 15132 38949 15196
rect 38883 15131 38949 15132
rect 38699 11796 38765 11797
rect 38699 11732 38700 11796
rect 38764 11732 38765 11796
rect 38699 11731 38765 11732
rect 39070 11525 39130 21795
rect 39067 11524 39133 11525
rect 39067 11460 39068 11524
rect 39132 11460 39133 11524
rect 39067 11459 39133 11460
rect 39070 9621 39130 11459
rect 39438 11389 39498 23427
rect 39803 22268 39869 22269
rect 39803 22204 39804 22268
rect 39868 22204 39869 22268
rect 39803 22203 39869 22204
rect 39619 20908 39685 20909
rect 39619 20844 39620 20908
rect 39684 20844 39685 20908
rect 39619 20843 39685 20844
rect 39622 11933 39682 20843
rect 39806 20501 39866 22203
rect 39803 20500 39869 20501
rect 39803 20436 39804 20500
rect 39868 20436 39869 20500
rect 39803 20435 39869 20436
rect 40358 20365 40418 23971
rect 40539 23492 40605 23493
rect 40539 23428 40540 23492
rect 40604 23428 40605 23492
rect 40539 23427 40605 23428
rect 42563 23492 42629 23493
rect 42563 23428 42564 23492
rect 42628 23428 42629 23492
rect 42563 23427 42629 23428
rect 40355 20364 40421 20365
rect 40355 20300 40356 20364
rect 40420 20300 40421 20364
rect 40355 20299 40421 20300
rect 39803 18052 39869 18053
rect 39803 17988 39804 18052
rect 39868 17988 39869 18052
rect 39803 17987 39869 17988
rect 39619 11932 39685 11933
rect 39619 11868 39620 11932
rect 39684 11868 39685 11932
rect 39619 11867 39685 11868
rect 39435 11388 39501 11389
rect 39435 11324 39436 11388
rect 39500 11324 39501 11388
rect 39435 11323 39501 11324
rect 39067 9620 39133 9621
rect 39067 9556 39068 9620
rect 39132 9556 39133 9620
rect 39067 9555 39133 9556
rect 38699 8804 38765 8805
rect 38699 8740 38700 8804
rect 38764 8740 38765 8804
rect 38699 8739 38765 8740
rect 38702 7989 38762 8739
rect 38699 7988 38765 7989
rect 38699 7924 38700 7988
rect 38764 7924 38765 7988
rect 38699 7923 38765 7924
rect 38515 7716 38581 7717
rect 38515 7652 38516 7716
rect 38580 7652 38581 7716
rect 38515 7651 38581 7652
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 39806 6629 39866 17987
rect 40355 15332 40421 15333
rect 40355 15268 40356 15332
rect 40420 15268 40421 15332
rect 40355 15267 40421 15268
rect 39987 11116 40053 11117
rect 39987 11052 39988 11116
rect 40052 11052 40053 11116
rect 39987 11051 40053 11052
rect 39990 7445 40050 11051
rect 39987 7444 40053 7445
rect 39987 7380 39988 7444
rect 40052 7380 40053 7444
rect 39987 7379 40053 7380
rect 39803 6628 39869 6629
rect 39803 6564 39804 6628
rect 39868 6564 39869 6628
rect 39803 6563 39869 6564
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37227 5948 37293 5949
rect 37227 5884 37228 5948
rect 37292 5884 37293 5948
rect 37227 5883 37293 5884
rect 37944 5472 38264 6496
rect 40358 6357 40418 15267
rect 40542 8125 40602 23427
rect 41091 22540 41157 22541
rect 41091 22476 41092 22540
rect 41156 22476 41157 22540
rect 41091 22475 41157 22476
rect 40723 20500 40789 20501
rect 40723 20436 40724 20500
rect 40788 20436 40789 20500
rect 40723 20435 40789 20436
rect 40726 14109 40786 20435
rect 41094 20365 41154 22475
rect 41827 20908 41893 20909
rect 41827 20844 41828 20908
rect 41892 20844 41893 20908
rect 41827 20843 41893 20844
rect 41275 20636 41341 20637
rect 41275 20572 41276 20636
rect 41340 20572 41341 20636
rect 41275 20571 41341 20572
rect 41091 20364 41157 20365
rect 41091 20300 41092 20364
rect 41156 20300 41157 20364
rect 41091 20299 41157 20300
rect 40907 14788 40973 14789
rect 40907 14724 40908 14788
rect 40972 14724 40973 14788
rect 40907 14723 40973 14724
rect 40723 14108 40789 14109
rect 40723 14044 40724 14108
rect 40788 14044 40789 14108
rect 40723 14043 40789 14044
rect 40539 8124 40605 8125
rect 40539 8060 40540 8124
rect 40604 8060 40605 8124
rect 40539 8059 40605 8060
rect 40355 6356 40421 6357
rect 40355 6292 40356 6356
rect 40420 6292 40421 6356
rect 40355 6291 40421 6292
rect 40910 6221 40970 14723
rect 41094 13701 41154 20299
rect 41278 15333 41338 20571
rect 41643 19276 41709 19277
rect 41643 19212 41644 19276
rect 41708 19212 41709 19276
rect 41643 19211 41709 19212
rect 41275 15332 41341 15333
rect 41275 15268 41276 15332
rect 41340 15268 41341 15332
rect 41275 15267 41341 15268
rect 41646 15061 41706 19211
rect 41643 15060 41709 15061
rect 41643 14996 41644 15060
rect 41708 14996 41709 15060
rect 41643 14995 41709 14996
rect 41091 13700 41157 13701
rect 41091 13636 41092 13700
rect 41156 13636 41157 13700
rect 41091 13635 41157 13636
rect 41830 11797 41890 20843
rect 42011 20228 42077 20229
rect 42011 20164 42012 20228
rect 42076 20164 42077 20228
rect 42011 20163 42077 20164
rect 41827 11796 41893 11797
rect 41827 11732 41828 11796
rect 41892 11732 41893 11796
rect 41827 11731 41893 11732
rect 41830 10981 41890 11731
rect 41827 10980 41893 10981
rect 41827 10916 41828 10980
rect 41892 10916 41893 10980
rect 41827 10915 41893 10916
rect 42014 7989 42074 20163
rect 42379 20092 42445 20093
rect 42379 20028 42380 20092
rect 42444 20028 42445 20092
rect 42379 20027 42445 20028
rect 42382 19141 42442 20027
rect 42379 19140 42445 19141
rect 42379 19076 42380 19140
rect 42444 19076 42445 19140
rect 42379 19075 42445 19076
rect 42382 10845 42442 19075
rect 42379 10844 42445 10845
rect 42379 10780 42380 10844
rect 42444 10780 42445 10844
rect 42379 10779 42445 10780
rect 42566 8533 42626 23427
rect 42944 23424 43264 24448
rect 43667 24036 43733 24037
rect 43667 23972 43668 24036
rect 43732 23972 43733 24036
rect 43667 23971 43733 23972
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 43670 13565 43730 23971
rect 44035 23084 44101 23085
rect 44035 23020 44036 23084
rect 44100 23020 44101 23084
rect 44035 23019 44101 23020
rect 43667 13564 43733 13565
rect 43667 13500 43668 13564
rect 43732 13500 43733 13564
rect 43667 13499 43733 13500
rect 43667 13428 43733 13429
rect 43667 13364 43668 13428
rect 43732 13364 43733 13428
rect 43667 13363 43733 13364
rect 43483 12612 43549 12613
rect 43483 12548 43484 12612
rect 43548 12548 43549 12612
rect 43483 12547 43549 12548
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 43486 11253 43546 12547
rect 43483 11252 43549 11253
rect 43483 11188 43484 11252
rect 43548 11188 43549 11252
rect 43483 11187 43549 11188
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 43670 9621 43730 13363
rect 43851 11116 43917 11117
rect 43851 11052 43852 11116
rect 43916 11052 43917 11116
rect 43851 11051 43917 11052
rect 43667 9620 43733 9621
rect 43667 9556 43668 9620
rect 43732 9556 43733 9620
rect 43667 9555 43733 9556
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42563 8532 42629 8533
rect 42563 8468 42564 8532
rect 42628 8468 42629 8532
rect 42563 8467 42629 8468
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42011 7988 42077 7989
rect 42011 7924 42012 7988
rect 42076 7924 42077 7988
rect 42011 7923 42077 7924
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 40907 6220 40973 6221
rect 40907 6156 40908 6220
rect 40972 6156 40973 6220
rect 40907 6155 40973 6156
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 36675 5132 36741 5133
rect 36675 5068 36676 5132
rect 36740 5068 36741 5132
rect 36675 5067 36741 5068
rect 36491 4996 36557 4997
rect 36491 4932 36492 4996
rect 36556 4932 36557 4996
rect 36491 4931 36557 4932
rect 35387 4588 35453 4589
rect 35387 4524 35388 4588
rect 35452 4524 35453 4588
rect 35387 4523 35453 4524
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 6016 43264 7040
rect 43854 6901 43914 11051
rect 44038 9621 44098 23019
rect 44222 20229 44282 25059
rect 44955 23492 45021 23493
rect 44955 23428 44956 23492
rect 45020 23428 45021 23492
rect 44955 23427 45021 23428
rect 44219 20228 44285 20229
rect 44219 20164 44220 20228
rect 44284 20164 44285 20228
rect 44219 20163 44285 20164
rect 44771 19140 44837 19141
rect 44771 19076 44772 19140
rect 44836 19076 44837 19140
rect 44771 19075 44837 19076
rect 44219 18868 44285 18869
rect 44219 18804 44220 18868
rect 44284 18804 44285 18868
rect 44219 18803 44285 18804
rect 44222 10165 44282 18803
rect 44403 15876 44469 15877
rect 44403 15812 44404 15876
rect 44468 15812 44469 15876
rect 44403 15811 44469 15812
rect 44406 12205 44466 15811
rect 44774 13837 44834 19075
rect 44771 13836 44837 13837
rect 44771 13772 44772 13836
rect 44836 13772 44837 13836
rect 44771 13771 44837 13772
rect 44403 12204 44469 12205
rect 44403 12140 44404 12204
rect 44468 12140 44469 12204
rect 44403 12139 44469 12140
rect 44771 11932 44837 11933
rect 44771 11868 44772 11932
rect 44836 11868 44837 11932
rect 44771 11867 44837 11868
rect 44219 10164 44285 10165
rect 44219 10100 44220 10164
rect 44284 10100 44285 10164
rect 44219 10099 44285 10100
rect 44035 9620 44101 9621
rect 44035 9556 44036 9620
rect 44100 9556 44101 9620
rect 44035 9555 44101 9556
rect 43851 6900 43917 6901
rect 43851 6836 43852 6900
rect 43916 6836 43917 6900
rect 43851 6835 43917 6836
rect 44774 6493 44834 11867
rect 44958 11797 45018 23427
rect 45323 22404 45389 22405
rect 45323 22340 45324 22404
rect 45388 22340 45389 22404
rect 45323 22339 45389 22340
rect 45139 20908 45205 20909
rect 45139 20844 45140 20908
rect 45204 20844 45205 20908
rect 45139 20843 45205 20844
rect 44955 11796 45021 11797
rect 44955 11732 44956 11796
rect 45020 11732 45021 11796
rect 44955 11731 45021 11732
rect 45142 7445 45202 20843
rect 45326 18053 45386 22339
rect 45323 18052 45389 18053
rect 45323 17988 45324 18052
rect 45388 17988 45389 18052
rect 45323 17987 45389 17988
rect 45323 17508 45389 17509
rect 45323 17444 45324 17508
rect 45388 17444 45389 17508
rect 45323 17443 45389 17444
rect 45326 16421 45386 17443
rect 45323 16420 45389 16421
rect 45323 16356 45324 16420
rect 45388 16356 45389 16420
rect 45323 16355 45389 16356
rect 45507 16420 45573 16421
rect 45507 16356 45508 16420
rect 45572 16356 45573 16420
rect 45507 16355 45573 16356
rect 45139 7444 45205 7445
rect 45139 7380 45140 7444
rect 45204 7380 45205 7444
rect 45139 7379 45205 7380
rect 45510 6765 45570 16355
rect 46062 15333 46122 26147
rect 46979 23900 47045 23901
rect 46979 23836 46980 23900
rect 47044 23836 47045 23900
rect 46979 23835 47045 23836
rect 46243 23492 46309 23493
rect 46243 23428 46244 23492
rect 46308 23428 46309 23492
rect 46243 23427 46309 23428
rect 46795 23492 46861 23493
rect 46795 23428 46796 23492
rect 46860 23428 46861 23492
rect 46795 23427 46861 23428
rect 46059 15332 46125 15333
rect 46059 15268 46060 15332
rect 46124 15268 46125 15332
rect 46059 15267 46125 15268
rect 45691 13564 45757 13565
rect 45691 13500 45692 13564
rect 45756 13500 45757 13564
rect 45691 13499 45757 13500
rect 45694 7037 45754 13499
rect 46246 10165 46306 23427
rect 46427 20228 46493 20229
rect 46427 20164 46428 20228
rect 46492 20164 46493 20228
rect 46427 20163 46493 20164
rect 46430 13293 46490 20163
rect 46798 16421 46858 23427
rect 46982 18869 47042 23835
rect 47166 19141 47226 26555
rect 47944 23968 48264 24528
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 48451 23492 48517 23493
rect 48451 23428 48452 23492
rect 48516 23428 48517 23492
rect 48451 23427 48517 23428
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47163 19140 47229 19141
rect 47163 19076 47164 19140
rect 47228 19076 47229 19140
rect 47163 19075 47229 19076
rect 46979 18868 47045 18869
rect 46979 18804 46980 18868
rect 47044 18804 47045 18868
rect 46979 18803 47045 18804
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47715 18052 47781 18053
rect 47715 17988 47716 18052
rect 47780 17988 47781 18052
rect 47715 17987 47781 17988
rect 46979 17916 47045 17917
rect 46979 17852 46980 17916
rect 47044 17852 47045 17916
rect 46979 17851 47045 17852
rect 46795 16420 46861 16421
rect 46795 16356 46796 16420
rect 46860 16356 46861 16420
rect 46795 16355 46861 16356
rect 46427 13292 46493 13293
rect 46427 13228 46428 13292
rect 46492 13228 46493 13292
rect 46427 13227 46493 13228
rect 46243 10164 46309 10165
rect 46243 10100 46244 10164
rect 46308 10100 46309 10164
rect 46243 10099 46309 10100
rect 45691 7036 45757 7037
rect 45691 6972 45692 7036
rect 45756 6972 45757 7036
rect 45691 6971 45757 6972
rect 45507 6764 45573 6765
rect 45507 6700 45508 6764
rect 45572 6700 45573 6764
rect 45507 6699 45573 6700
rect 44771 6492 44837 6493
rect 44771 6428 44772 6492
rect 44836 6428 44837 6492
rect 44771 6427 44837 6428
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 46798 5677 46858 16355
rect 46982 11933 47042 17851
rect 47347 16692 47413 16693
rect 47347 16628 47348 16692
rect 47412 16628 47413 16692
rect 47347 16627 47413 16628
rect 46979 11932 47045 11933
rect 46979 11868 46980 11932
rect 47044 11868 47045 11932
rect 46979 11867 47045 11868
rect 47350 11389 47410 16627
rect 47718 13429 47778 17987
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47715 13428 47781 13429
rect 47715 13364 47716 13428
rect 47780 13364 47781 13428
rect 47715 13363 47781 13364
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47347 11388 47413 11389
rect 47347 11324 47348 11388
rect 47412 11324 47413 11388
rect 47347 11323 47413 11324
rect 46979 11116 47045 11117
rect 46979 11052 46980 11116
rect 47044 11052 47045 11116
rect 46979 11051 47045 11052
rect 46982 9077 47042 11051
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 46979 9076 47045 9077
rect 46979 9012 46980 9076
rect 47044 9012 47045 9076
rect 46979 9011 47045 9012
rect 46982 6765 47042 9011
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 48454 8261 48514 23427
rect 48635 20772 48701 20773
rect 48635 20708 48636 20772
rect 48700 20708 48701 20772
rect 48635 20707 48701 20708
rect 48638 13565 48698 20707
rect 49187 19412 49253 19413
rect 49187 19348 49188 19412
rect 49252 19348 49253 19412
rect 49187 19347 49253 19348
rect 48819 19140 48885 19141
rect 48819 19076 48820 19140
rect 48884 19076 48885 19140
rect 48819 19075 48885 19076
rect 48635 13564 48701 13565
rect 48635 13500 48636 13564
rect 48700 13500 48701 13564
rect 48635 13499 48701 13500
rect 48822 9077 48882 19075
rect 49190 14109 49250 19347
rect 49923 18868 49989 18869
rect 49923 18804 49924 18868
rect 49988 18804 49989 18868
rect 49923 18803 49989 18804
rect 49926 14789 49986 18803
rect 49923 14788 49989 14789
rect 49923 14724 49924 14788
rect 49988 14724 49989 14788
rect 49923 14723 49989 14724
rect 49187 14108 49253 14109
rect 49187 14044 49188 14108
rect 49252 14044 49253 14108
rect 49187 14043 49253 14044
rect 48819 9076 48885 9077
rect 48819 9012 48820 9076
rect 48884 9012 48885 9076
rect 48819 9011 48885 9012
rect 48451 8260 48517 8261
rect 48451 8196 48452 8260
rect 48516 8196 48517 8260
rect 48451 8195 48517 8196
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 46979 6764 47045 6765
rect 46979 6700 46980 6764
rect 47044 6700 47045 6764
rect 46979 6699 47045 6700
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 46795 5676 46861 5677
rect 46795 5612 46796 5676
rect 46860 5612 46861 5676
rect 46795 5611 46861 5612
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_2  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1679235063
transform 1 0 11684 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1679235063
transform 1 0 7544 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _107_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1679235063
transform 1 0 3588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1679235063
transform 1 0 16836 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1679235063
transform 1 0 13432 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1679235063
transform 1 0 5704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1679235063
transform 1 0 9292 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1679235063
transform 1 0 10764 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1679235063
transform 1 0 6716 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1679235063
transform 1 0 3588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1679235063
transform 1 0 11684 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1679235063
transform 1 0 16008 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1679235063
transform 1 0 11224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1679235063
transform 1 0 6808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1679235063
transform 1 0 3588 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1679235063
transform 1 0 6072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1679235063
transform 1 0 11776 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1679235063
transform 1 0 7176 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1679235063
transform 1 0 3496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1679235063
transform 1 0 19412 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1679235063
transform 1 0 21988 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1679235063
transform 1 0 4968 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _128_
timestamp 1679235063
transform 1 0 4232 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1679235063
transform 1 0 24564 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1679235063
transform 1 0 6072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1679235063
transform 1 0 2392 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1679235063
transform 1 0 5704 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1679235063
transform 1 0 6440 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1679235063
transform 1 0 37444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1679235063
transform 1 0 37260 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1679235063
transform 1 0 37996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1679235063
transform 1 0 43608 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1679235063
transform 1 0 39192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1679235063
transform 1 0 38456 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1679235063
transform 1 0 38088 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1679235063
transform 1 0 44068 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1679235063
transform 1 0 38364 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1679235063
transform 1 0 37812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1679235063
transform 1 0 38548 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1679235063
transform 1 0 44804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1679235063
transform 1 0 40020 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1679235063
transform 1 0 40940 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1679235063
transform 1 0 40020 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1679235063
transform 1 0 44068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1679235063
transform 1 0 41860 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1679235063
transform 1 0 39008 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1679235063
transform 1 0 40480 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1679235063
transform 1 0 44252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1679235063
transform 1 0 41124 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1679235063
transform 1 0 39652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1679235063
transform 1 0 42228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1679235063
transform 1 0 44344 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1679235063
transform 1 0 45080 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1679235063
transform 1 0 42596 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1679235063
transform 1 0 45540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1679235063
transform 1 0 46460 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1679235063
transform 1 0 45908 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1679235063
transform 1 0 45172 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1679235063
transform 1 0 3128 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _165_
timestamp 1679235063
transform 1 0 2392 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1679235063
transform 1 0 5428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _167_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 4140 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _168_
timestamp 1679235063
transform 1 0 7820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _169_
timestamp 1679235063
transform 1 0 7728 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _170_
timestamp 1679235063
transform 1 0 3956 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _171_
timestamp 1679235063
transform 1 0 6532 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _172_
timestamp 1679235063
transform 1 0 5888 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _173_
timestamp 1679235063
transform 1 0 9108 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1679235063
transform 1 0 14260 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _175_
timestamp 1679235063
transform 1 0 23644 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _176_
timestamp 1679235063
transform 1 0 3128 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1679235063
transform 1 0 19412 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1679235063
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _179_
timestamp 1679235063
transform 1 0 18492 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _180_
timestamp 1679235063
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _181_
timestamp 1679235063
transform 1 0 18400 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _182_
timestamp 1679235063
transform 1 0 11040 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _183_
timestamp 1679235063
transform 1 0 13708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 1679235063
transform 1 0 14628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1679235063
transform 1 0 28612 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1679235063
transform 1 0 28796 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _187_
timestamp 1679235063
transform 1 0 31464 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 1679235063
transform 1 0 17112 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1679235063
transform 1 0 27324 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _190_
timestamp 1679235063
transform 1 0 24564 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1679235063
transform 1 0 27140 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _192_
timestamp 1679235063
transform 1 0 31464 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _193_
timestamp 1679235063
transform 1 0 16836 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _194_
timestamp 1679235063
transform 1 0 16100 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1679235063
transform 1 0 16928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1679235063
transform 1 0 18676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1679235063
transform 1 0 20240 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 44252 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1679235063
transform 1 0 36892 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1679235063
transform 1 0 44252 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1679235063
transform 1 0 34960 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1679235063
transform 1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1679235063
transform 1 0 12236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1679235063
transform 1 0 2668 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1679235063
transform 1 0 10212 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1679235063
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1679235063
transform 1 0 10212 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1679235063
transform 1 0 12788 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1679235063
transform 1 0 35788 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1679235063
transform 1 0 46828 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1679235063
transform 1 0 35972 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1679235063
transform 1 0 48300 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1679235063
transform 1 0 47656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1679235063
transform 1 0 45448 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1679235063
transform 1 0 47196 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1679235063
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1679235063
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1679235063
transform 1 0 9200 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1679235063
transform 1 0 28244 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1679235063
transform 1 0 36892 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1679235063
transform 1 0 38916 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1679235063
transform 1 0 46368 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1679235063
transform 1 0 47288 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1679235063
transform 1 0 47564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1679235063
transform 1 0 47564 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1679235063
transform 1 0 48668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1679235063
transform 1 0 6532 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1679235063
transform 1 0 44804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1679235063
transform 1 0 10672 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1679235063
transform 1 0 14812 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1679235063
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1679235063
transform 1 0 5704 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1679235063
transform 1 0 6440 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1679235063
transform 1 0 3864 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1679235063
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1679235063
transform 1 0 6716 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1679235063
transform 1 0 3312 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1679235063
transform 1 0 3220 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1679235063
transform 1 0 3312 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1679235063
transform 1 0 3220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1679235063
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1679235063
transform 1 0 8280 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1679235063
transform 1 0 1656 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1679235063
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1679235063
transform 1 0 2760 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1679235063
transform 1 0 6440 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1679235063
transform 1 0 3312 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1679235063
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1679235063
transform 1 0 17940 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1679235063
transform 1 0 22540 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1679235063
transform 1 0 5520 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1679235063
transform 1 0 25116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1679235063
transform 1 0 37996 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1679235063
transform 1 0 36892 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A
timestamp 1679235063
transform 1 0 38548 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A
timestamp 1679235063
transform 1 0 39744 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1679235063
transform 1 0 38088 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1679235063
transform 1 0 38640 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1679235063
transform 1 0 37996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1679235063
transform 1 0 37628 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1679235063
transform 1 0 39008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1679235063
transform 1 0 40204 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1679235063
transform 1 0 40756 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1679235063
transform 1 0 41492 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1679235063
transform 1 0 43884 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1679235063
transform 1 0 39560 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1679235063
transform 1 0 40572 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1679235063
transform 1 0 41768 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1679235063
transform 1 0 38640 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1679235063
transform 1 0 41952 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1679235063
transform 1 0 42136 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A
timestamp 1679235063
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__A
timestamp 1679235063
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A
timestamp 1679235063
transform 1 0 1472 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1679235063
transform 1 0 3312 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1679235063
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A
timestamp 1679235063
transform 1 0 29072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A
timestamp 1679235063
transform 1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1679235063
transform 1 0 18584 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 9016 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 6532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 9016 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 16192 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 13616 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 11592 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 19412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 17480 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 17940 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 11592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__S
timestamp 1679235063
transform 1 0 18124 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 3864 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 18216 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 16468 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 17572 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 13984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 18216 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 18768 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 15272 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 12604 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 12420 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 13984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 11592 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 6532 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 8832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 14352 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 9292 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 9108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 11776 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 14168 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 23000 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20608 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 23276 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1679235063
transform 1 0 30084 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1679235063
transform 1 0 13984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1679235063
transform 1 0 14168 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1679235063
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1679235063
transform 1 0 20056 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1679235063
transform 1 0 14168 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1679235063
transform 1 0 9292 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1679235063
transform 1 0 22724 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1679235063
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1679235063
transform 1 0 32752 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1679235063
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1679235063
transform 1 0 35052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1679235063
transform 1 0 37628 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1679235063
transform 1 0 33672 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1679235063
transform 1 0 34316 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1679235063
transform 1 0 47196 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1679235063
transform 1 0 44344 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout203_A
timestamp 1679235063
transform 1 0 23552 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout204_A
timestamp 1679235063
transform 1 0 14168 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout205_A
timestamp 1679235063
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout206_A
timestamp 1679235063
transform 1 0 14260 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout207_A
timestamp 1679235063
transform 1 0 9016 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout208_A
timestamp 1679235063
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout209_A
timestamp 1679235063
transform 1 0 31740 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout210_A
timestamp 1679235063
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout211_A
timestamp 1679235063
transform 1 0 44528 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout212_A
timestamp 1679235063
transform 1 0 46828 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout213_A
timestamp 1679235063
transform 1 0 44712 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout214_A
timestamp 1679235063
transform 1 0 43332 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout215_A
timestamp 1679235063
transform 1 0 45080 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold10_A
timestamp 1679235063
transform 1 0 44620 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold58_A
timestamp 1679235063
transform 1 0 39468 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold157_A
timestamp 1679235063
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold168_A
timestamp 1679235063
transform 1 0 5060 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold211_A
timestamp 1679235063
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold240_A
timestamp 1679235063
transform 1 0 47196 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold253_A
timestamp 1679235063
transform 1 0 48300 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold281_A
timestamp 1679235063
transform 1 0 44436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold282_A
timestamp 1679235063
transform 1 0 3036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold307_A
timestamp 1679235063
transform 1 0 3312 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold313_A
timestamp 1679235063
transform 1 0 9200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold319_A
timestamp 1679235063
transform 1 0 34500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold320_A
timestamp 1679235063
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold323_A
timestamp 1679235063
transform 1 0 41952 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold329_A
timestamp 1679235063
transform 1 0 3312 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold334_A
timestamp 1679235063
transform 1 0 47564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold340_A
timestamp 1679235063
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold342_A
timestamp 1679235063
transform 1 0 48300 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold349_A
timestamp 1679235063
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold351_A
timestamp 1679235063
transform 1 0 46736 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold354_A
timestamp 1679235063
transform 1 0 16836 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold358_A
timestamp 1679235063
transform 1 0 42136 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold360_A
timestamp 1679235063
transform 1 0 6716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold363_A
timestamp 1679235063
transform 1 0 44988 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold364_A
timestamp 1679235063
transform 1 0 5152 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold370_A
timestamp 1679235063
transform 1 0 44804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold371_A
timestamp 1679235063
transform 1 0 44620 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold372_A
timestamp 1679235063
transform 1 0 42320 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold373_A
timestamp 1679235063
transform 1 0 39560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold374_A
timestamp 1679235063
transform 1 0 45816 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold377_A
timestamp 1679235063
transform 1 0 3220 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold378_A
timestamp 1679235063
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold380_A
timestamp 1679235063
transform 1 0 43700 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold381_A
timestamp 1679235063
transform 1 0 47288 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold386_A
timestamp 1679235063
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1679235063
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1679235063
transform 1 0 3036 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1679235063
transform 1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1679235063
transform 1 0 2760 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1679235063
transform 1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1679235063
transform 1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1679235063
transform 1 0 2300 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1679235063
transform 1 0 3036 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1679235063
transform 1 0 3404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1679235063
transform 1 0 3220 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1679235063
transform 1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1679235063
transform 1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1679235063
transform 1 0 2668 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1679235063
transform 1 0 2392 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1679235063
transform 1 0 2852 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1679235063
transform 1 0 3312 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1679235063
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1679235063
transform 1 0 4508 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1679235063
transform 1 0 2852 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1679235063
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1679235063
transform 1 0 2668 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1679235063
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1679235063
transform 1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1679235063
transform 1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1679235063
transform 1 0 2116 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1679235063
transform 1 0 2852 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1679235063
transform 1 0 3036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1679235063
transform 1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1679235063
transform 1 0 2116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1679235063
transform 1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1679235063
transform 1 0 44620 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1679235063
transform 1 0 44252 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1679235063
transform 1 0 47564 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1679235063
transform 1 0 44804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1679235063
transform 1 0 47288 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1679235063
transform 1 0 47564 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1679235063
transform 1 0 47564 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1679235063
transform 1 0 43148 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1679235063
transform 1 0 46920 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1679235063
transform 1 0 46644 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1679235063
transform 1 0 44528 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1679235063
transform 1 0 44988 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1679235063
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1679235063
transform 1 0 47564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1679235063
transform 1 0 42044 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1679235063
transform 1 0 45172 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1679235063
transform 1 0 44068 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1679235063
transform 1 0 46276 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1679235063
transform 1 0 45448 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1679235063
transform 1 0 46000 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1679235063
transform 1 0 42964 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1679235063
transform 1 0 43516 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1679235063
transform 1 0 47564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1679235063
transform 1 0 46644 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1679235063
transform 1 0 45816 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1679235063
transform 1 0 47564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1679235063
transform 1 0 42780 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1679235063
transform 1 0 45448 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1679235063
transform 1 0 43884 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1679235063
transform 1 0 41860 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1679235063
transform 1 0 12236 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1679235063
transform 1 0 47288 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1679235063
transform 1 0 44988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1679235063
transform 1 0 38456 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1679235063
transform 1 0 39284 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1679235063
transform 1 0 41860 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1679235063
transform 1 0 42136 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1679235063
transform 1 0 43056 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1679235063
transform 1 0 43792 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1679235063
transform 1 0 45172 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1679235063
transform 1 0 44988 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1679235063
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1679235063
transform 1 0 47564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1679235063
transform 1 0 44988 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1679235063
transform 1 0 47104 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1679235063
transform 1 0 47104 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1679235063
transform 1 0 47564 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1679235063
transform 1 0 44528 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1679235063
transform 1 0 46920 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1679235063
transform 1 0 43700 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1679235063
transform 1 0 46276 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1679235063
transform 1 0 47564 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1679235063
transform 1 0 9384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1679235063
transform 1 0 20332 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1679235063
transform 1 0 13984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1679235063
transform 1 0 42044 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1679235063
transform 1 0 46828 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1679235063
transform 1 0 5704 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1679235063
transform 1 0 3312 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1679235063
transform 1 0 44988 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1679235063
transform 1 0 29164 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1679235063
transform 1 0 31280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1679235063
transform 1 0 33396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1679235063
transform 1 0 35512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1679235063
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1679235063
transform 1 0 44620 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1679235063
transform 1 0 47472 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1679235063
transform 1 0 46000 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1679235063
transform 1 0 45632 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1679235063
transform 1 0 46460 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1679235063
transform 1 0 45264 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1679235063
transform 1 0 44988 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1679235063
transform 1 0 16744 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1679235063
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output123_A
timestamp 1679235063
transform 1 0 5336 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output126_A
timestamp 1679235063
transform 1 0 3312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output171_A
timestamp 1679235063
transform 1 0 9016 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output190_A
timestamp 1679235063
transform 1 0 11960 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 25024 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21344 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 16744 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20424 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19320 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23368 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__D
timestamp 1679235063
transform 1 0 10120 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 9384 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 9384 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2__D
timestamp 1679235063
transform 1 0 11592 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 11776 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 18860 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 16744 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21896 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 39284 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 37444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 36800 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 39376 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__D
timestamp 1679235063
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 44620 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 47564 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 46092 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 47012 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 41860 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 44712 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 44804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 42044 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 39284 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24472 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 25576 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 21344 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 24012 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 18584 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 19412 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19872 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 9108 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 7544 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 6716 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 7544 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 7544 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 9016 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 9200 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 3864 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 41124 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 41860 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 35328 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 29072 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 27140 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 23828 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 22908 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 26220 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 26404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 22080 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 23736 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23000 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 16560 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 18124 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l2_in_1__S
timestamp 1679235063
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 27048 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 26864 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 26312 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 25576 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 24564 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 28888 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 28520 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 24564 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 24472 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 18768 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 18400 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 18584 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 29164 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 29440 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 26496 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 24932 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 25116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 19688 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 19596 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 19320 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 28888 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 26496 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 20700 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 21896 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 21344 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 12788 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 31740 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 17112 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 20608 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 21344 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l2_in_1__A0
timestamp 1679235063
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l2_in_1__S
timestamp 1679235063
transform 1 0 15640 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l3_in_0__S
timestamp 1679235063
transform 1 0 10856 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 5428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 35604 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 35512 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 29256 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 25208 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 23920 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 23736 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 23184 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_37.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 42044 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_37.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 44344 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_37.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 30544 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_37.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 29164 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_37.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 24288 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_45.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 44620 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_45.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 44712 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_45.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 42136 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_45.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 34224 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 44620 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 27140 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 20516 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_1__S
timestamp 1679235063
transform 1 0 19228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 29716 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 34316 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 29900 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 34316 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 34132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 34132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 26404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 26588 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 27968 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 44528 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 41308 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 40296 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 33856 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 34040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 29716 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 29900 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 46828 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 47012 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 36064 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 35880 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 33856 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 34040 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 47196 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 46828 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 47196 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 34868 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 34316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 37076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 36892 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 35512 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 36984 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 41768 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 41952 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 42044 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 34500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 39560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 35604 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 30636 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 31832 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 41952 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 42136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 41768 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 31648 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 27784 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 27968 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 28244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 34132 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 34500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 31464 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 28060 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 30728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 26404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 26588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 30176 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 30912 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 25484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 25484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 32292 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 34500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 30360 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 30636 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31556 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 31740 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 29532 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 30912 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 30728 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 47104 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 44436 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 44712 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 41032 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 41216 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 41676 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 22816 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 28152 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 34316 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 26496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l2_in_1__S
timestamp 1679235063
transform 1 0 33304 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 26312 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 41400 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 41584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 35236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 39560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 37444 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 47196 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 47012 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 47288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 47748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 45356 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 44620 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 34776 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3312 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 49036 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 45172 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 41860 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 35880 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 37628 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l2_in_1__A0
timestamp 1679235063
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l3_in_0__S
timestamp 1679235063
transform 1 0 35420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 47196 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 45172 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 49128 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 44712 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 47564 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 49312 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 41860 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 39468 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 44804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l2_in_1__S
timestamp 1679235063
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 47012 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 46828 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 49220 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 47380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 39468 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 47196 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 44528 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 44620 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 39468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 42136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 44344 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 33212 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 29716 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 27140 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 24472 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26956 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 26588 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 28520 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 24012 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 29164 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 30728 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 25760 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_28.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25944 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 23092 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_30.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 22632 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 22816 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3220 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_32.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16836 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18308 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_34.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18216 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 4692 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 29164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 19136 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_40.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14168 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_40.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14168 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_42.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_42.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16652 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_46.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 9016 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_48.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 12696 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_50.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 9108 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_50.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_50.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_58.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_58.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13616 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_58.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 11776 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_58.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 6532 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_58.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 9200 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 2208 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17940 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16100 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16192 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 16284 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 13248 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 14260 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13156 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10396 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 10304 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 10764 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11684 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11592 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 10120 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 8464 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14260 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15456 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 15548 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 19044 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_
timestamp 1679235063
transform 1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13984 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 17204 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_
timestamp 1679235063
transform 1 0 17296 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_
timestamp 1679235063
transform 1 0 16928 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__259 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16468 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 14536 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_
timestamp 1679235063
transform 1 0 18492 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_
timestamp 1679235063
transform 1 0 17572 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18676 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12052 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_
timestamp 1679235063
transform 1 0 17848 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_
timestamp 1679235063
transform 1 0 15456 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_
timestamp 1679235063
transform 1 0 17940 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12696 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12788 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_
timestamp 1679235063
transform 1 0 12972 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_
timestamp 1679235063
transform 1 0 16928 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__260
timestamp 1679235063
transform 1 0 15824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_
timestamp 1679235063
transform 1 0 15456 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_
timestamp 1679235063
transform 1 0 14996 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17756 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 7544 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 7728 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 17204 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_
timestamp 1679235063
transform 1 0 14260 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_
timestamp 1679235063
transform 1 0 15732 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9108 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_
timestamp 1679235063
transform 1 0 12972 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_
timestamp 1679235063
transform 1 0 11684 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__261
timestamp 1679235063
transform 1 0 10672 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_
timestamp 1679235063
transform 1 0 11960 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_
timestamp 1679235063
transform 1 0 11776 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14996 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12604 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 13156 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14352 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_
timestamp 1679235063
transform 1 0 17940 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_
timestamp 1679235063
transform 1 0 12972 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11960 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_
timestamp 1679235063
transform 1 0 14260 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_
timestamp 1679235063
transform 1 0 12972 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_
timestamp 1679235063
transform 1 0 15180 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__262
timestamp 1679235063
transform 1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 11408 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_
timestamp 1679235063
transform 1 0 11868 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 27140 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 22264 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 22172 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14536 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 25208 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 24012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 23092 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 20976 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20976 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 24104 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 22264 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 24840 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 19320 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24564 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 23644 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 21620 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 27508 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 18124 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 28796 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 27140 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16560 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1679235063
transform 1 0 14720 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1679235063
transform 1 0 22264 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1679235063
transform 1 0 20884 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1679235063
transform 1 0 16468 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1679235063
transform 1 0 15640 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1679235063
transform 1 0 21344 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1679235063
transform 1 0 20516 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1679235063
transform 1 0 33028 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1679235063
transform 1 0 30636 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1679235063
transform 1 0 35236 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1679235063
transform 1 0 35972 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1679235063
transform 1 0 31372 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1679235063
transform 1 0 31556 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1679235063
transform 1 0 37352 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1679235063
transform 1 0 35972 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout203
timestamp 1679235063
transform 1 0 21988 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout204
timestamp 1679235063
transform 1 0 17940 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout205
timestamp 1679235063
transform 1 0 27140 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout206 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23276 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  fanout207
timestamp 1679235063
transform 1 0 19412 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout208 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16928 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout209
timestamp 1679235063
transform 1 0 30544 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  fanout210 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 36616 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout211
timestamp 1679235063
transform 1 0 34868 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout212 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 32384 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout213
timestamp 1679235063
transform 1 0 43700 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout214
timestamp 1679235063
transform 1 0 48576 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout215
timestamp 1679235063
transform 1 0 48852 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17
timestamp 1679235063
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24
timestamp 1679235063
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1679235063
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1679235063
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp 1679235063
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 7820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1679235063
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1679235063
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95
timestamp 1679235063
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1679235063
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1679235063
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp 1679235063
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1679235063
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_159
timestamp 1679235063
transform 1 0 15732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1679235063
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1679235063
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1679235063
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1679235063
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1679235063
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_205
timestamp 1679235063
transform 1 0 19964 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_211
timestamp 1679235063
transform 1 0 20516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1679235063
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1679235063
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1679235063
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_255
timestamp 1679235063
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1679235063
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1679235063
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1679235063
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_293 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_299
timestamp 1679235063
transform 1 0 28612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_303
timestamp 1679235063
transform 1 0 28980 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1679235063
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1679235063
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_321
timestamp 1679235063
transform 1 0 30636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_326
timestamp 1679235063
transform 1 0 31096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1679235063
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_337
timestamp 1679235063
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_345
timestamp 1679235063
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_349
timestamp 1679235063
transform 1 0 33212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_353
timestamp 1679235063
transform 1 0 33580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1679235063
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_365
timestamp 1679235063
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_372
timestamp 1679235063
transform 1 0 35328 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_376
timestamp 1679235063
transform 1 0 35696 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_388
timestamp 1679235063
transform 1 0 36800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1679235063
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1679235063
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1679235063
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_421
timestamp 1679235063
transform 1 0 39836 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_429
timestamp 1679235063
transform 1 0 40572 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1679235063
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1679235063
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1679235063
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1679235063
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_477
timestamp 1679235063
transform 1 0 44988 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_485
timestamp 1679235063
transform 1 0 45724 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1679235063
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_505
timestamp 1679235063
transform 1 0 47564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1679235063
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1679235063
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_9
timestamp 1679235063
transform 1 0 1932 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_19
timestamp 1679235063
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_31
timestamp 1679235063
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_43
timestamp 1679235063
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1679235063
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1679235063
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_69
timestamp 1679235063
transform 1 0 7452 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_77
timestamp 1679235063
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_86
timestamp 1679235063
transform 1 0 9016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_98
timestamp 1679235063
transform 1 0 10120 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1679235063
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1679235063
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1679235063
transform 1 0 12236 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_130
timestamp 1679235063
transform 1 0 13064 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_142
timestamp 1679235063
transform 1 0 14168 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1679235063
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1679235063
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1679235063
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_194
timestamp 1679235063
transform 1 0 18952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1679235063
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1679235063
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1679235063
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_229
timestamp 1679235063
transform 1 0 22172 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1679235063
transform 1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_243
timestamp 1679235063
transform 1 0 23460 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_266
timestamp 1679235063
transform 1 0 25576 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1679235063
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_281
timestamp 1679235063
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_294
timestamp 1679235063
transform 1 0 28152 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_300
timestamp 1679235063
transform 1 0 28704 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_322
timestamp 1679235063
transform 1 0 30728 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1679235063
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1679235063
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1679235063
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1679235063
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1679235063
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1679235063
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1679235063
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1679235063
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1679235063
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1679235063
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1679235063
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1679235063
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1679235063
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1679235063
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_461
timestamp 1679235063
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_465
timestamp 1679235063
transform 1 0 43884 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_482
timestamp 1679235063
transform 1 0 45448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1679235063
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_505
timestamp 1679235063
transform 1 0 47564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1679235063
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1679235063
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1679235063
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1679235063
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1679235063
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1679235063
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1679235063
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1679235063
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_77
timestamp 1679235063
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_81
timestamp 1679235063
transform 1 0 8556 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1679235063
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp 1679235063
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_93
timestamp 1679235063
transform 1 0 9660 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_105
timestamp 1679235063
transform 1 0 10764 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_117
timestamp 1679235063
transform 1 0 11868 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_129
timestamp 1679235063
transform 1 0 12972 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1679235063
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1679235063
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_153
timestamp 1679235063
transform 1 0 15180 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_161
timestamp 1679235063
transform 1 0 15916 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1679235063
transform 1 0 16468 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_171
timestamp 1679235063
transform 1 0 16836 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_175
timestamp 1679235063
transform 1 0 17204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1679235063
transform 1 0 18308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1679235063
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1679235063
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_207
timestamp 1679235063
transform 1 0 20148 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_215
timestamp 1679235063
transform 1 0 20884 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_237
timestamp 1679235063
transform 1 0 22908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_241
timestamp 1679235063
transform 1 0 23276 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1679235063
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1679235063
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_275
timestamp 1679235063
transform 1 0 26404 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_291
timestamp 1679235063
transform 1 0 27876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_303
timestamp 1679235063
transform 1 0 28980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1679235063
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1679235063
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_319
timestamp 1679235063
transform 1 0 30452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_331
timestamp 1679235063
transform 1 0 31556 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_343
timestamp 1679235063
transform 1 0 32660 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_355
timestamp 1679235063
transform 1 0 33764 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1679235063
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1679235063
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1679235063
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1679235063
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1679235063
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1679235063
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1679235063
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1679235063
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1679235063
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1679235063
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1679235063
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1679235063
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1679235063
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1679235063
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_505
timestamp 1679235063
transform 1 0 47564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1679235063
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1679235063
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_9
timestamp 1679235063
transform 1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_17
timestamp 1679235063
transform 1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_23
timestamp 1679235063
transform 1 0 3220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_35
timestamp 1679235063
transform 1 0 4324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1679235063
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1679235063
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1679235063
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1679235063
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1679235063
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_101
timestamp 1679235063
transform 1 0 10396 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 1679235063
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1679235063
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1679235063
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1679235063
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1679235063
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1679235063
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1679235063
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1679235063
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1679235063
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_206
timestamp 1679235063
transform 1 0 20056 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp 1679235063
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1679235063
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_235
timestamp 1679235063
transform 1 0 22724 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_246
timestamp 1679235063
transform 1 0 23736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_271
timestamp 1679235063
transform 1 0 26036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1679235063
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1679235063
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_304
timestamp 1679235063
transform 1 0 29072 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_316
timestamp 1679235063
transform 1 0 30176 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_328
timestamp 1679235063
transform 1 0 31280 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1679235063
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1679235063
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1679235063
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1679235063
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1679235063
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1679235063
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1679235063
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_399
timestamp 1679235063
transform 1 0 37812 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_403
timestamp 1679235063
transform 1 0 38180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_415
timestamp 1679235063
transform 1 0 39284 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_427
timestamp 1679235063
transform 1 0 40388 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_439
timestamp 1679235063
transform 1 0 41492 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1679235063
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1679235063
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1679235063
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1679235063
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_485
timestamp 1679235063
transform 1 0 45724 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1679235063
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_507
timestamp 1679235063
transform 1 0 47748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1679235063
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1679235063
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_9
timestamp 1679235063
transform 1 0 1932 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1679235063
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1679235063
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1679235063
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1679235063
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1679235063
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1679235063
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1679235063
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1679235063
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1679235063
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1679235063
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1679235063
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1679235063
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1679235063
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1679235063
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1679235063
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1679235063
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1679235063
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1679235063
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_189
timestamp 1679235063
transform 1 0 18492 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1679235063
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1679235063
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_208
timestamp 1679235063
transform 1 0 20240 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_214
timestamp 1679235063
transform 1 0 20792 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_236
timestamp 1679235063
transform 1 0 22816 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_240
timestamp 1679235063
transform 1 0 23184 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1679235063
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1679235063
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_258
timestamp 1679235063
transform 1 0 24840 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_283
timestamp 1679235063
transform 1 0 27140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_295
timestamp 1679235063
transform 1 0 28244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1679235063
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1679235063
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1679235063
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1679235063
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1679235063
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1679235063
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1679235063
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1679235063
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1679235063
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_391
timestamp 1679235063
transform 1 0 37076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_397
timestamp 1679235063
transform 1 0 37628 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1679235063
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_409
timestamp 1679235063
transform 1 0 38732 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_417
timestamp 1679235063
transform 1 0 39468 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1679235063
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1679235063
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1679235063
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1679235063
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1679235063
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1679235063
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_477
timestamp 1679235063
transform 1 0 44988 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_485
timestamp 1679235063
transform 1 0 45724 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_490
timestamp 1679235063
transform 1 0 46184 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_497
timestamp 1679235063
transform 1 0 46828 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_502
timestamp 1679235063
transform 1 0 47288 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_507
timestamp 1679235063
transform 1 0 47748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1679235063
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1679235063
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1679235063
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1679235063
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1679235063
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1679235063
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1679235063
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1679235063
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1679235063
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1679235063
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1679235063
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1679235063
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1679235063
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1679235063
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1679235063
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1679235063
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1679235063
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1679235063
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1679235063
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1679235063
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1679235063
transform 1 0 17204 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1679235063
transform 1 0 17572 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_184
timestamp 1679235063
transform 1 0 18032 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_196
timestamp 1679235063
transform 1 0 19136 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_208
timestamp 1679235063
transform 1 0 20240 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1679235063
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_225
timestamp 1679235063
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_229
timestamp 1679235063
transform 1 0 22172 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_233
timestamp 1679235063
transform 1 0 22540 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_245
timestamp 1679235063
transform 1 0 23644 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_252
timestamp 1679235063
transform 1 0 24288 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_264
timestamp 1679235063
transform 1 0 25392 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1679235063
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1679235063
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1679235063
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1679235063
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1679235063
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1679235063
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1679235063
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1679235063
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_342
timestamp 1679235063
transform 1 0 32568 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_354
timestamp 1679235063
transform 1 0 33672 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_366
timestamp 1679235063
transform 1 0 34776 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_378
timestamp 1679235063
transform 1 0 35880 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_390
timestamp 1679235063
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_393
timestamp 1679235063
transform 1 0 37260 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_401
timestamp 1679235063
transform 1 0 37996 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_404
timestamp 1679235063
transform 1 0 38272 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_410
timestamp 1679235063
transform 1 0 38824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_418
timestamp 1679235063
transform 1 0 39560 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_422
timestamp 1679235063
transform 1 0 39928 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_434
timestamp 1679235063
transform 1 0 41032 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_446
timestamp 1679235063
transform 1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1679235063
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1679235063
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_473
timestamp 1679235063
transform 1 0 44620 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_481
timestamp 1679235063
transform 1 0 45356 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_484
timestamp 1679235063
transform 1 0 45632 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1679235063
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_507
timestamp 1679235063
transform 1 0 47748 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1679235063
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1679235063
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1679235063
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_17
timestamp 1679235063
transform 1 0 2668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1679235063
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1679235063
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1679235063
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1679235063
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1679235063
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1679235063
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1679235063
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1679235063
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1679235063
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1679235063
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1679235063
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1679235063
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1679235063
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1679235063
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1679235063
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_153
timestamp 1679235063
transform 1 0 15180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_159
timestamp 1679235063
transform 1 0 15732 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_163
timestamp 1679235063
transform 1 0 16100 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_170
timestamp 1679235063
transform 1 0 16744 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_182
timestamp 1679235063
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1679235063
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1679235063
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_202
timestamp 1679235063
transform 1 0 19688 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_208
timestamp 1679235063
transform 1 0 20240 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_217
timestamp 1679235063
transform 1 0 21068 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_226
timestamp 1679235063
transform 1 0 21896 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_238
timestamp 1679235063
transform 1 0 23000 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1679235063
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1679235063
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_263
timestamp 1679235063
transform 1 0 25300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_275
timestamp 1679235063
transform 1 0 26404 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_287
timestamp 1679235063
transform 1 0 27508 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_299
timestamp 1679235063
transform 1 0 28612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1679235063
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1679235063
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_319
timestamp 1679235063
transform 1 0 30452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_331
timestamp 1679235063
transform 1 0 31556 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_335
timestamp 1679235063
transform 1 0 31924 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_347
timestamp 1679235063
transform 1 0 33028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_359
timestamp 1679235063
transform 1 0 34132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1679235063
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1679235063
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1679235063
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1679235063
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1679235063
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1679235063
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1679235063
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1679235063
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1679235063
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1679235063
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_457
timestamp 1679235063
transform 1 0 43148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_461
timestamp 1679235063
transform 1 0 43516 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_466
timestamp 1679235063
transform 1 0 43976 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_477
timestamp 1679235063
transform 1 0 44988 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_490
timestamp 1679235063
transform 1 0 46184 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_495
timestamp 1679235063
transform 1 0 46644 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_500
timestamp 1679235063
transform 1 0 47104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_505
timestamp 1679235063
transform 1 0 47564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1679235063
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1679235063
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_9
timestamp 1679235063
transform 1 0 1932 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1679235063
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1679235063
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1679235063
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1679235063
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1679235063
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1679235063
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1679235063
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1679235063
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1679235063
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1679235063
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1679235063
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1679235063
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_119
timestamp 1679235063
transform 1 0 12052 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_123
timestamp 1679235063
transform 1 0 12420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_138
timestamp 1679235063
transform 1 0 13800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_142
timestamp 1679235063
transform 1 0 14168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_146
timestamp 1679235063
transform 1 0 14536 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_150
timestamp 1679235063
transform 1 0 14904 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_154
timestamp 1679235063
transform 1 0 15272 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1679235063
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1679235063
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 1679235063
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_186
timestamp 1679235063
transform 1 0 18216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_198
timestamp 1679235063
transform 1 0 19320 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_210
timestamp 1679235063
transform 1 0 20424 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1679235063
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1679235063
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_235
timestamp 1679235063
transform 1 0 22724 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_243
timestamp 1679235063
transform 1 0 23460 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_252
timestamp 1679235063
transform 1 0 24288 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_264
timestamp 1679235063
transform 1 0 25392 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1679235063
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1679235063
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1679235063
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_307
timestamp 1679235063
transform 1 0 29348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_311
timestamp 1679235063
transform 1 0 29716 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_320
timestamp 1679235063
transform 1 0 30544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1679235063
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1679235063
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_347
timestamp 1679235063
transform 1 0 33028 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_354
timestamp 1679235063
transform 1 0 33672 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_366
timestamp 1679235063
transform 1 0 34776 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_378
timestamp 1679235063
transform 1 0 35880 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_390
timestamp 1679235063
transform 1 0 36984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_393
timestamp 1679235063
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_401
timestamp 1679235063
transform 1 0 37996 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_406
timestamp 1679235063
transform 1 0 38456 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_410
timestamp 1679235063
transform 1 0 38824 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_422
timestamp 1679235063
transform 1 0 39928 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_434
timestamp 1679235063
transform 1 0 41032 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_446
timestamp 1679235063
transform 1 0 42136 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1679235063
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_461
timestamp 1679235063
transform 1 0 43516 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_479
timestamp 1679235063
transform 1 0 45172 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_484
timestamp 1679235063
transform 1 0 45632 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_491
timestamp 1679235063
transform 1 0 46276 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_498
timestamp 1679235063
transform 1 0 46920 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_507
timestamp 1679235063
transform 1 0 47748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1679235063
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1679235063
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_9
timestamp 1679235063
transform 1 0 1932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_16
timestamp 1679235063
transform 1 0 2576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1679235063
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1679235063
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1679235063
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1679235063
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1679235063
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1679235063
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1679235063
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 1679235063
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_89
timestamp 1679235063
transform 1 0 9292 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_92
timestamp 1679235063
transform 1 0 9568 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_104
timestamp 1679235063
transform 1 0 10672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_118
timestamp 1679235063
transform 1 0 11960 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_125
timestamp 1679235063
transform 1 0 12604 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_129
timestamp 1679235063
transform 1 0 12972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_133
timestamp 1679235063
transform 1 0 13340 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1679235063
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1679235063
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_146
timestamp 1679235063
transform 1 0 14536 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_162
timestamp 1679235063
transform 1 0 16008 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_166
timestamp 1679235063
transform 1 0 16376 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_175
timestamp 1679235063
transform 1 0 17204 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_188
timestamp 1679235063
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1679235063
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_202
timestamp 1679235063
transform 1 0 19688 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_216
timestamp 1679235063
transform 1 0 20976 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_228
timestamp 1679235063
transform 1 0 22080 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_240
timestamp 1679235063
transform 1 0 23184 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1679235063
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_253
timestamp 1679235063
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_261
timestamp 1679235063
transform 1 0 25116 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_270
timestamp 1679235063
transform 1 0 25944 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_282
timestamp 1679235063
transform 1 0 27048 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_298
timestamp 1679235063
transform 1 0 28520 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1679235063
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1679235063
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_319
timestamp 1679235063
transform 1 0 30452 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_331
timestamp 1679235063
transform 1 0 31556 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_347
timestamp 1679235063
transform 1 0 33028 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_359
timestamp 1679235063
transform 1 0 34132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1679235063
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1679235063
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_375
timestamp 1679235063
transform 1 0 35604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_387
timestamp 1679235063
transform 1 0 36708 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_399
timestamp 1679235063
transform 1 0 37812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_411
timestamp 1679235063
transform 1 0 38916 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1679235063
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1679235063
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1679235063
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1679235063
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_457
timestamp 1679235063
transform 1 0 43148 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_465
timestamp 1679235063
transform 1 0 43884 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_471
timestamp 1679235063
transform 1 0 44436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1679235063
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_479
timestamp 1679235063
transform 1 0 45172 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_485
timestamp 1679235063
transform 1 0 45724 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_505
timestamp 1679235063
transform 1 0 47564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1679235063
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1679235063
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_9
timestamp 1679235063
transform 1 0 1932 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_13
timestamp 1679235063
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_25
timestamp 1679235063
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_37
timestamp 1679235063
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1679235063
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1679235063
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1679235063
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1679235063
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_81
timestamp 1679235063
transform 1 0 8556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_85
timestamp 1679235063
transform 1 0 8924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_90
timestamp 1679235063
transform 1 0 9384 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_97
timestamp 1679235063
transform 1 0 10028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_104
timestamp 1679235063
transform 1 0 10672 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp 1679235063
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_119
timestamp 1679235063
transform 1 0 12052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_126
timestamp 1679235063
transform 1 0 12696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_138
timestamp 1679235063
transform 1 0 13800 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_142
timestamp 1679235063
transform 1 0 14168 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_154
timestamp 1679235063
transform 1 0 15272 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1679235063
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_173
timestamp 1679235063
transform 1 0 17020 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_185
timestamp 1679235063
transform 1 0 18124 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_198
timestamp 1679235063
transform 1 0 19320 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_210
timestamp 1679235063
transform 1 0 20424 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1679235063
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_227
timestamp 1679235063
transform 1 0 21988 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_243
timestamp 1679235063
transform 1 0 23460 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_255
timestamp 1679235063
transform 1 0 24564 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_267
timestamp 1679235063
transform 1 0 25668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1679235063
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_281
timestamp 1679235063
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_295
timestamp 1679235063
transform 1 0 28244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_299
timestamp 1679235063
transform 1 0 28612 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_308
timestamp 1679235063
transform 1 0 29440 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_320
timestamp 1679235063
transform 1 0 30544 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_332
timestamp 1679235063
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_337
timestamp 1679235063
transform 1 0 32108 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_349
timestamp 1679235063
transform 1 0 33212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_361
timestamp 1679235063
transform 1 0 34316 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_365
timestamp 1679235063
transform 1 0 34684 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_375
timestamp 1679235063
transform 1 0 35604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_387
timestamp 1679235063
transform 1 0 36708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1679235063
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_393
timestamp 1679235063
transform 1 0 37260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_399
timestamp 1679235063
transform 1 0 37812 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_403
timestamp 1679235063
transform 1 0 38180 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_409
timestamp 1679235063
transform 1 0 38732 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_416
timestamp 1679235063
transform 1 0 39376 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_423
timestamp 1679235063
transform 1 0 40020 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_427
timestamp 1679235063
transform 1 0 40388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_439
timestamp 1679235063
transform 1 0 41492 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1679235063
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_449
timestamp 1679235063
transform 1 0 42412 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_459
timestamp 1679235063
transform 1 0 43332 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_464
timestamp 1679235063
transform 1 0 43792 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_471
timestamp 1679235063
transform 1 0 44436 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_479
timestamp 1679235063
transform 1 0 45172 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_486
timestamp 1679235063
transform 1 0 45816 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_494
timestamp 1679235063
transform 1 0 46552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_502
timestamp 1679235063
transform 1 0 47288 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_507
timestamp 1679235063
transform 1 0 47748 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1679235063
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1679235063
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_9
timestamp 1679235063
transform 1 0 1932 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1679235063
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1679235063
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1679235063
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1679235063
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1679235063
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1679235063
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_77
timestamp 1679235063
transform 1 0 8188 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1679235063
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp 1679235063
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_93
timestamp 1679235063
transform 1 0 9660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_100
timestamp 1679235063
transform 1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_107
timestamp 1679235063
transform 1 0 10948 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_114
timestamp 1679235063
transform 1 0 11592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_126
timestamp 1679235063
transform 1 0 12696 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1679235063
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp 1679235063
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_144
timestamp 1679235063
transform 1 0 14352 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1679235063
transform 1 0 14812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_161
timestamp 1679235063
transform 1 0 15916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_185
timestamp 1679235063
transform 1 0 18124 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_192
timestamp 1679235063
transform 1 0 18768 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp 1679235063
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_208
timestamp 1679235063
transform 1 0 20240 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_220
timestamp 1679235063
transform 1 0 21344 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_232
timestamp 1679235063
transform 1 0 22448 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_238
timestamp 1679235063
transform 1 0 23000 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1679235063
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_255
timestamp 1679235063
transform 1 0 24564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_259
timestamp 1679235063
transform 1 0 24932 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_268
timestamp 1679235063
transform 1 0 25760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_280
timestamp 1679235063
transform 1 0 26864 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_294
timestamp 1679235063
transform 1 0 28152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1679235063
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1679235063
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_319
timestamp 1679235063
transform 1 0 30452 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_331
timestamp 1679235063
transform 1 0 31556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_336
timestamp 1679235063
transform 1 0 32016 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_347
timestamp 1679235063
transform 1 0 33028 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_351
timestamp 1679235063
transform 1 0 33396 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_361
timestamp 1679235063
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_365
timestamp 1679235063
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_375
timestamp 1679235063
transform 1 0 35604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_387
timestamp 1679235063
transform 1 0 36708 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_391
timestamp 1679235063
transform 1 0 37076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_395
timestamp 1679235063
transform 1 0 37444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_403
timestamp 1679235063
transform 1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_411
timestamp 1679235063
transform 1 0 38916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_418
timestamp 1679235063
transform 1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_421
timestamp 1679235063
transform 1 0 39836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_427
timestamp 1679235063
transform 1 0 40388 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_433
timestamp 1679235063
transform 1 0 40940 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_442
timestamp 1679235063
transform 1 0 41768 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_445
timestamp 1679235063
transform 1 0 42044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_450
timestamp 1679235063
transform 1 0 42504 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_455
timestamp 1679235063
transform 1 0 42964 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_462
timestamp 1679235063
transform 1 0 43608 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_469
timestamp 1679235063
transform 1 0 44252 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_481
timestamp 1679235063
transform 1 0 45356 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_486
timestamp 1679235063
transform 1 0 45816 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_494
timestamp 1679235063
transform 1 0 46552 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_502
timestamp 1679235063
transform 1 0 47288 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_506
timestamp 1679235063
transform 1 0 47656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1679235063
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1679235063
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_15
timestamp 1679235063
transform 1 0 2484 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1679235063
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1679235063
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_51
timestamp 1679235063
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1679235063
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_72
timestamp 1679235063
transform 1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_79
timestamp 1679235063
transform 1 0 8372 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_97
timestamp 1679235063
transform 1 0 10028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_101
timestamp 1679235063
transform 1 0 10396 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1679235063
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1679235063
transform 1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_125
timestamp 1679235063
transform 1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_138
timestamp 1679235063
transform 1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_144
timestamp 1679235063
transform 1 0 14352 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_154
timestamp 1679235063
transform 1 0 15272 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1679235063
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp 1679235063
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1679235063
transform 1 0 17756 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_189
timestamp 1679235063
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_192
timestamp 1679235063
transform 1 0 18768 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_214
timestamp 1679235063
transform 1 0 20792 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1679235063
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1679235063
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_247
timestamp 1679235063
transform 1 0 23828 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_251
timestamp 1679235063
transform 1 0 24196 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_262
timestamp 1679235063
transform 1 0 25208 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1679235063
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_281
timestamp 1679235063
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_293
timestamp 1679235063
transform 1 0 28060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_317
timestamp 1679235063
transform 1 0 30268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_323
timestamp 1679235063
transform 1 0 30820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1679235063
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_337
timestamp 1679235063
transform 1 0 32108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_349
timestamp 1679235063
transform 1 0 33212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_362
timestamp 1679235063
transform 1 0 34408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_366
timestamp 1679235063
transform 1 0 34776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_376
timestamp 1679235063
transform 1 0 35696 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_388
timestamp 1679235063
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1679235063
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_403
timestamp 1679235063
transform 1 0 38180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_410
timestamp 1679235063
transform 1 0 38824 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_414
timestamp 1679235063
transform 1 0 39192 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_417
timestamp 1679235063
transform 1 0 39468 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_429
timestamp 1679235063
transform 1 0 40572 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_437
timestamp 1679235063
transform 1 0 41308 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1679235063
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_449
timestamp 1679235063
transform 1 0 42412 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_454
timestamp 1679235063
transform 1 0 42872 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_458
timestamp 1679235063
transform 1 0 43240 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_463
timestamp 1679235063
transform 1 0 43700 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_471
timestamp 1679235063
transform 1 0 44436 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_475
timestamp 1679235063
transform 1 0 44804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_482
timestamp 1679235063
transform 1 0 45448 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_502
timestamp 1679235063
transform 1 0 47288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_507
timestamp 1679235063
transform 1 0 47748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1679235063
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1679235063
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_9
timestamp 1679235063
transform 1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_17
timestamp 1679235063
transform 1 0 2668 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_24
timestamp 1679235063
transform 1 0 3312 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_31
timestamp 1679235063
transform 1 0 3956 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_43
timestamp 1679235063
transform 1 0 5060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_49
timestamp 1679235063
transform 1 0 5612 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_62
timestamp 1679235063
transform 1 0 6808 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_70
timestamp 1679235063
transform 1 0 7544 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1679235063
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1679235063
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_101
timestamp 1679235063
transform 1 0 10396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_113
timestamp 1679235063
transform 1 0 11500 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_125
timestamp 1679235063
transform 1 0 12604 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1679235063
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1679235063
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_147
timestamp 1679235063
transform 1 0 14628 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_160
timestamp 1679235063
transform 1 0 15824 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_184
timestamp 1679235063
transform 1 0 18032 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_188
timestamp 1679235063
transform 1 0 18400 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1679235063
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_203
timestamp 1679235063
transform 1 0 19780 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_225
timestamp 1679235063
transform 1 0 21804 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_249
timestamp 1679235063
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1679235063
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_263
timestamp 1679235063
transform 1 0 25300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_267
timestamp 1679235063
transform 1 0 25668 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_278
timestamp 1679235063
transform 1 0 26680 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_290
timestamp 1679235063
transform 1 0 27784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_294
timestamp 1679235063
transform 1 0 28152 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1679235063
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1679235063
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_331
timestamp 1679235063
transform 1 0 31556 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_355
timestamp 1679235063
transform 1 0 33764 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1679235063
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1679235063
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_376
timestamp 1679235063
transform 1 0 35696 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_388
timestamp 1679235063
transform 1 0 36800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_392
timestamp 1679235063
transform 1 0 37168 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_403
timestamp 1679235063
transform 1 0 38180 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_410
timestamp 1679235063
transform 1 0 38824 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_416
timestamp 1679235063
transform 1 0 39376 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_421
timestamp 1679235063
transform 1 0 39836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_427
timestamp 1679235063
transform 1 0 40388 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_441
timestamp 1679235063
transform 1 0 41676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_455
timestamp 1679235063
transform 1 0 42964 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_462
timestamp 1679235063
transform 1 0 43608 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_466
timestamp 1679235063
transform 1 0 43976 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_473
timestamp 1679235063
transform 1 0 44620 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_481
timestamp 1679235063
transform 1 0 45356 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_493
timestamp 1679235063
transform 1 0 46460 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_499
timestamp 1679235063
transform 1 0 47012 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_505
timestamp 1679235063
transform 1 0 47564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1679235063
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1679235063
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_9
timestamp 1679235063
transform 1 0 1932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_16
timestamp 1679235063
transform 1 0 2576 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_21
timestamp 1679235063
transform 1 0 3036 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_28
timestamp 1679235063
transform 1 0 3680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_35
timestamp 1679235063
transform 1 0 4324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_41
timestamp 1679235063
transform 1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_47
timestamp 1679235063
transform 1 0 5428 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1679235063
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1679235063
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 1679235063
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_77
timestamp 1679235063
transform 1 0 8188 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_86
timestamp 1679235063
transform 1 0 9016 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_98
timestamp 1679235063
transform 1 0 10120 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1679235063
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1679235063
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1679235063
transform 1 0 11960 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_128
timestamp 1679235063
transform 1 0 12880 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_152
timestamp 1679235063
transform 1 0 15088 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1679235063
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1679235063
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1679235063
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_218
timestamp 1679235063
transform 1 0 21160 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1679235063
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_236
timestamp 1679235063
transform 1 0 22816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_241
timestamp 1679235063
transform 1 0 23276 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_263
timestamp 1679235063
transform 1 0 25300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_267
timestamp 1679235063
transform 1 0 25668 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1679235063
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_281
timestamp 1679235063
transform 1 0 26956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_287
timestamp 1679235063
transform 1 0 27508 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_311
timestamp 1679235063
transform 1 0 29716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_318
timestamp 1679235063
transform 1 0 30360 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_323
timestamp 1679235063
transform 1 0 30820 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1679235063
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1679235063
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_359
timestamp 1679235063
transform 1 0 34132 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_372
timestamp 1679235063
transform 1 0 35328 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_376
timestamp 1679235063
transform 1 0 35696 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_388
timestamp 1679235063
transform 1 0 36800 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1679235063
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_403
timestamp 1679235063
transform 1 0 38180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_415
timestamp 1679235063
transform 1 0 39284 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_423
timestamp 1679235063
transform 1 0 40020 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_427
timestamp 1679235063
transform 1 0 40388 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_432
timestamp 1679235063
transform 1 0 40848 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_446
timestamp 1679235063
transform 1 0 42136 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_449
timestamp 1679235063
transform 1 0 42412 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_461
timestamp 1679235063
transform 1 0 43516 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_475
timestamp 1679235063
transform 1 0 44804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_489
timestamp 1679235063
transform 1 0 46092 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_493
timestamp 1679235063
transform 1 0 46460 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_500
timestamp 1679235063
transform 1 0 47104 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_507
timestamp 1679235063
transform 1 0 47748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1679235063
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1679235063
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_15
timestamp 1679235063
transform 1 0 2484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_22
timestamp 1679235063
transform 1 0 3128 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1679235063
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1679235063
transform 1 0 4876 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_45
timestamp 1679235063
transform 1 0 5244 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_49
timestamp 1679235063
transform 1 0 5612 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_54
timestamp 1679235063
transform 1 0 6072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_62
timestamp 1679235063
transform 1 0 6808 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_70
timestamp 1679235063
transform 1 0 7544 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1679235063
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1679235063
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1679235063
transform 1 0 9384 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_100
timestamp 1679235063
transform 1 0 10304 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_112
timestamp 1679235063
transform 1 0 11408 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_125
timestamp 1679235063
transform 1 0 12604 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1679235063
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1679235063
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_163
timestamp 1679235063
transform 1 0 16100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1679235063
transform 1 0 16744 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_181
timestamp 1679235063
transform 1 0 17756 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1679235063
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1679235063
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_219
timestamp 1679235063
transform 1 0 21252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_223
timestamp 1679235063
transform 1 0 21620 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_233
timestamp 1679235063
transform 1 0 22540 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_246
timestamp 1679235063
transform 1 0 23736 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1679235063
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1679235063
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_264
timestamp 1679235063
transform 1 0 25392 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_272
timestamp 1679235063
transform 1 0 26128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_278
timestamp 1679235063
transform 1 0 26680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_299
timestamp 1679235063
transform 1 0 28612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1679235063
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1679235063
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_320
timestamp 1679235063
transform 1 0 30544 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_326
timestamp 1679235063
transform 1 0 31096 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_336
timestamp 1679235063
transform 1 0 32016 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_351
timestamp 1679235063
transform 1 0 33396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1679235063
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1679235063
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_387
timestamp 1679235063
transform 1 0 36708 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_393
timestamp 1679235063
transform 1 0 37260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_404
timestamp 1679235063
transform 1 0 38272 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_416
timestamp 1679235063
transform 1 0 39376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_421
timestamp 1679235063
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_431
timestamp 1679235063
transform 1 0 40756 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_439
timestamp 1679235063
transform 1 0 41492 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_447
timestamp 1679235063
transform 1 0 42228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_461
timestamp 1679235063
transform 1 0 43516 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_467
timestamp 1679235063
transform 1 0 44068 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_474
timestamp 1679235063
transform 1 0 44712 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_479
timestamp 1679235063
transform 1 0 45172 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_485
timestamp 1679235063
transform 1 0 45724 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_505
timestamp 1679235063
transform 1 0 47564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1679235063
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1679235063
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_9
timestamp 1679235063
transform 1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_17
timestamp 1679235063
transform 1 0 2668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_23
timestamp 1679235063
transform 1 0 3220 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_29
timestamp 1679235063
transform 1 0 3772 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_43
timestamp 1679235063
transform 1 0 5060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_51
timestamp 1679235063
transform 1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1679235063
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_60
timestamp 1679235063
transform 1 0 6624 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_66
timestamp 1679235063
transform 1 0 7176 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_74
timestamp 1679235063
transform 1 0 7912 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_86
timestamp 1679235063
transform 1 0 9016 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_98
timestamp 1679235063
transform 1 0 10120 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1679235063
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1679235063
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_116
timestamp 1679235063
transform 1 0 11776 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_127
timestamp 1679235063
transform 1 0 12788 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_154
timestamp 1679235063
transform 1 0 15272 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1679235063
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_169
timestamp 1679235063
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1679235063
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_194
timestamp 1679235063
transform 1 0 18952 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1679235063
transform 1 0 19504 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1679235063
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 1679235063
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp 1679235063
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_244
timestamp 1679235063
transform 1 0 23552 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_249
timestamp 1679235063
transform 1 0 24012 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_271
timestamp 1679235063
transform 1 0 26036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_277
timestamp 1679235063
transform 1 0 26588 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_281
timestamp 1679235063
transform 1 0 26956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_293
timestamp 1679235063
transform 1 0 28060 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_297
timestamp 1679235063
transform 1 0 28428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_307
timestamp 1679235063
transform 1 0 29348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_311
timestamp 1679235063
transform 1 0 29716 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_333
timestamp 1679235063
transform 1 0 31740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_337
timestamp 1679235063
transform 1 0 32108 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_341
timestamp 1679235063
transform 1 0 32476 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_351
timestamp 1679235063
transform 1 0 33396 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_375
timestamp 1679235063
transform 1 0 35604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_388
timestamp 1679235063
transform 1 0 36800 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1679235063
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_404
timestamp 1679235063
transform 1 0 38272 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_416
timestamp 1679235063
transform 1 0 39376 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_428
timestamp 1679235063
transform 1 0 40480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_440
timestamp 1679235063
transform 1 0 41584 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_449
timestamp 1679235063
transform 1 0 42412 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_454
timestamp 1679235063
transform 1 0 42872 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_468
timestamp 1679235063
transform 1 0 44160 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_482
timestamp 1679235063
transform 1 0 45448 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_496
timestamp 1679235063
transform 1 0 46736 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_507
timestamp 1679235063
transform 1 0 47748 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1679235063
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1679235063
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_9
timestamp 1679235063
transform 1 0 1932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_13
timestamp 1679235063
transform 1 0 2300 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_18
timestamp 1679235063
transform 1 0 2760 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1679235063
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_31
timestamp 1679235063
transform 1 0 3956 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_38
timestamp 1679235063
transform 1 0 4600 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_46
timestamp 1679235063
transform 1 0 5336 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_52
timestamp 1679235063
transform 1 0 5888 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_58
timestamp 1679235063
transform 1 0 6440 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_70
timestamp 1679235063
transform 1 0 7544 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1679235063
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_91
timestamp 1679235063
transform 1 0 9476 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_101
timestamp 1679235063
transform 1 0 10396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_125
timestamp 1679235063
transform 1 0 12604 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1679235063
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1679235063
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_144
timestamp 1679235063
transform 1 0 14352 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_155
timestamp 1679235063
transform 1 0 15364 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_168
timestamp 1679235063
transform 1 0 16560 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_181
timestamp 1679235063
transform 1 0 17756 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1679235063
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1679235063
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_202
timestamp 1679235063
transform 1 0 19688 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_208
timestamp 1679235063
transform 1 0 20240 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1679235063
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_243
timestamp 1679235063
transform 1 0 23460 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1679235063
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1679235063
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_275
timestamp 1679235063
transform 1 0 26404 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_279
timestamp 1679235063
transform 1 0 26772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_300
timestamp 1679235063
transform 1 0 28704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1679235063
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_319
timestamp 1679235063
transform 1 0 30452 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_343
timestamp 1679235063
transform 1 0 32660 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_356
timestamp 1679235063
transform 1 0 33856 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_360
timestamp 1679235063
transform 1 0 34224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_365
timestamp 1679235063
transform 1 0 34684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_377
timestamp 1679235063
transform 1 0 35788 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_402
timestamp 1679235063
transform 1 0 38088 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_414
timestamp 1679235063
transform 1 0 39192 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_421
timestamp 1679235063
transform 1 0 39836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_431
timestamp 1679235063
transform 1 0 40756 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_443
timestamp 1679235063
transform 1 0 41860 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_451
timestamp 1679235063
transform 1 0 42596 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_458
timestamp 1679235063
transform 1 0 43240 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_472
timestamp 1679235063
transform 1 0 44528 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_481
timestamp 1679235063
transform 1 0 45356 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_494
timestamp 1679235063
transform 1 0 46552 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_498
timestamp 1679235063
transform 1 0 46920 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_505
timestamp 1679235063
transform 1 0 47564 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1679235063
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1679235063
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1679235063
transform 1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_13
timestamp 1679235063
transform 1 0 2300 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_18
timestamp 1679235063
transform 1 0 2760 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_26
timestamp 1679235063
transform 1 0 3496 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_32
timestamp 1679235063
transform 1 0 4048 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_42
timestamp 1679235063
transform 1 0 4968 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_48
timestamp 1679235063
transform 1 0 5520 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1679235063
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1679235063
transform 1 0 6808 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_74
timestamp 1679235063
transform 1 0 7912 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_86
timestamp 1679235063
transform 1 0 9016 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_98
timestamp 1679235063
transform 1 0 10120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1679235063
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1679235063
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_138
timestamp 1679235063
transform 1 0 13800 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_142
timestamp 1679235063
transform 1 0 14168 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1679235063
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1679235063
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_171
timestamp 1679235063
transform 1 0 16836 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_176
timestamp 1679235063
transform 1 0 17296 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1679235063
transform 1 0 19504 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_204
timestamp 1679235063
transform 1 0 19872 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1679235063
transform 1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1679235063
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1679235063
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_247
timestamp 1679235063
transform 1 0 23828 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_260
timestamp 1679235063
transform 1 0 25024 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_273
timestamp 1679235063
transform 1 0 26220 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1679235063
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1679235063
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_292
timestamp 1679235063
transform 1 0 27968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_317
timestamp 1679235063
transform 1 0 30268 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_332
timestamp 1679235063
transform 1 0 31648 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1679235063
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_348
timestamp 1679235063
transform 1 0 33120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_373
timestamp 1679235063
transform 1 0 35420 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_386
timestamp 1679235063
transform 1 0 36616 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1679235063
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_415
timestamp 1679235063
transform 1 0 39284 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_427
timestamp 1679235063
transform 1 0 40388 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_439
timestamp 1679235063
transform 1 0 41492 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_446
timestamp 1679235063
transform 1 0 42136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_449
timestamp 1679235063
transform 1 0 42412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_455
timestamp 1679235063
transform 1 0 42964 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_459
timestamp 1679235063
transform 1 0 43332 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_464
timestamp 1679235063
transform 1 0 43792 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_472
timestamp 1679235063
transform 1 0 44528 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_480
timestamp 1679235063
transform 1 0 45264 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_494
timestamp 1679235063
transform 1 0 46552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_502
timestamp 1679235063
transform 1 0 47288 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_507
timestamp 1679235063
transform 1 0 47748 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1679235063
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1679235063
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_14
timestamp 1679235063
transform 1 0 2392 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_19
timestamp 1679235063
transform 1 0 2852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1679235063
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1679235063
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_34
timestamp 1679235063
transform 1 0 4232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_46
timestamp 1679235063
transform 1 0 5336 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_58
timestamp 1679235063
transform 1 0 6440 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_70
timestamp 1679235063
transform 1 0 7544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1679235063
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1679235063
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_96
timestamp 1679235063
transform 1 0 9936 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_120
timestamp 1679235063
transform 1 0 12144 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_127
timestamp 1679235063
transform 1 0 12788 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1679235063
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1679235063
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_164
timestamp 1679235063
transform 1 0 16192 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1679235063
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_192
timestamp 1679235063
transform 1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_199
timestamp 1679235063
transform 1 0 19412 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1679235063
transform 1 0 20424 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_214
timestamp 1679235063
transform 1 0 20792 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_226
timestamp 1679235063
transform 1 0 21896 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_241
timestamp 1679235063
transform 1 0 23276 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_248
timestamp 1679235063
transform 1 0 23920 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1679235063
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_275
timestamp 1679235063
transform 1 0 26404 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_288
timestamp 1679235063
transform 1 0 27600 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_294
timestamp 1679235063
transform 1 0 28152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1679235063
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1679235063
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_314
timestamp 1679235063
transform 1 0 29992 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_318
timestamp 1679235063
transform 1 0 30360 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_341
timestamp 1679235063
transform 1 0 32476 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_354
timestamp 1679235063
transform 1 0 33672 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_358
timestamp 1679235063
transform 1 0 34040 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1679235063
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1679235063
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_387
timestamp 1679235063
transform 1 0 36708 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_400
timestamp 1679235063
transform 1 0 37904 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_413
timestamp 1679235063
transform 1 0 39100 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1679235063
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1679235063
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_431
timestamp 1679235063
transform 1 0 40756 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_443
timestamp 1679235063
transform 1 0 41860 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_455
timestamp 1679235063
transform 1 0 42964 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_467
timestamp 1679235063
transform 1 0 44068 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_474
timestamp 1679235063
transform 1 0 44712 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_477
timestamp 1679235063
transform 1 0 44988 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_489
timestamp 1679235063
transform 1 0 46092 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_503
timestamp 1679235063
transform 1 0 47380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_507
timestamp 1679235063
transform 1 0 47748 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1679235063
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1679235063
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_15
timestamp 1679235063
transform 1 0 2484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_20
timestamp 1679235063
transform 1 0 2944 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_30
timestamp 1679235063
transform 1 0 3864 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_42
timestamp 1679235063
transform 1 0 4968 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1679235063
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1679235063
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1679235063
transform 1 0 6624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_63
timestamp 1679235063
transform 1 0 6900 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_73
timestamp 1679235063
transform 1 0 7820 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_85
timestamp 1679235063
transform 1 0 8924 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_97
timestamp 1679235063
transform 1 0 10028 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1679235063
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1679235063
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_124
timestamp 1679235063
transform 1 0 12512 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_128
timestamp 1679235063
transform 1 0 12880 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_138
timestamp 1679235063
transform 1 0 13800 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_144
timestamp 1679235063
transform 1 0 14352 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1679235063
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_171
timestamp 1679235063
transform 1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_177
timestamp 1679235063
transform 1 0 17388 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1679235063
transform 1 0 17756 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_194
timestamp 1679235063
transform 1 0 18952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_207
timestamp 1679235063
transform 1 0 20148 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_211
timestamp 1679235063
transform 1 0 20516 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1679235063
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_227
timestamp 1679235063
transform 1 0 21988 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_232
timestamp 1679235063
transform 1 0 22448 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_245
timestamp 1679235063
transform 1 0 23644 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_269
timestamp 1679235063
transform 1 0 25852 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_276
timestamp 1679235063
transform 1 0 26496 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1679235063
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_291
timestamp 1679235063
transform 1 0 27876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_295
timestamp 1679235063
transform 1 0 28244 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_316
timestamp 1679235063
transform 1 0 30176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_331
timestamp 1679235063
transform 1 0 31556 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1679235063
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1679235063
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_359
timestamp 1679235063
transform 1 0 34132 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_366
timestamp 1679235063
transform 1 0 34776 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_370
timestamp 1679235063
transform 1 0 35144 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_382
timestamp 1679235063
transform 1 0 36248 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_390
timestamp 1679235063
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1679235063
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_418
timestamp 1679235063
transform 1 0 39560 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_430
timestamp 1679235063
transform 1 0 40664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_442
timestamp 1679235063
transform 1 0 41768 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_449
timestamp 1679235063
transform 1 0 42412 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_459
timestamp 1679235063
transform 1 0 43332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_471
timestamp 1679235063
transform 1 0 44436 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_477
timestamp 1679235063
transform 1 0 44988 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_483
timestamp 1679235063
transform 1 0 45540 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_490
timestamp 1679235063
transform 1 0 46184 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_502
timestamp 1679235063
transform 1 0 47288 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_507
timestamp 1679235063
transform 1 0 47748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1679235063
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1679235063
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_21
timestamp 1679235063
transform 1 0 3036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1679235063
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_34
timestamp 1679235063
transform 1 0 4232 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_46
timestamp 1679235063
transform 1 0 5336 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_58
timestamp 1679235063
transform 1 0 6440 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_70
timestamp 1679235063
transform 1 0 7544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1679235063
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_87
timestamp 1679235063
transform 1 0 9108 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1679235063
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_122
timestamp 1679235063
transform 1 0 12328 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_135
timestamp 1679235063
transform 1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_141
timestamp 1679235063
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_146
timestamp 1679235063
transform 1 0 14536 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_159
timestamp 1679235063
transform 1 0 15732 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_184
timestamp 1679235063
transform 1 0 18032 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_197
timestamp 1679235063
transform 1 0 19228 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_200
timestamp 1679235063
transform 1 0 19504 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_211
timestamp 1679235063
transform 1 0 20516 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_235
timestamp 1679235063
transform 1 0 22724 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_239
timestamp 1679235063
transform 1 0 23092 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1679235063
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1679235063
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_275
timestamp 1679235063
transform 1 0 26404 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_279
timestamp 1679235063
transform 1 0 26772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_303
timestamp 1679235063
transform 1 0 28980 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1679235063
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_317
timestamp 1679235063
transform 1 0 30268 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_320
timestamp 1679235063
transform 1 0 30544 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_343
timestamp 1679235063
transform 1 0 32660 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_358
timestamp 1679235063
transform 1 0 34040 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1679235063
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_369
timestamp 1679235063
transform 1 0 35052 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_380
timestamp 1679235063
transform 1 0 36064 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_404
timestamp 1679235063
transform 1 0 38272 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_416
timestamp 1679235063
transform 1 0 39376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_421
timestamp 1679235063
transform 1 0 39836 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_431
timestamp 1679235063
transform 1 0 40756 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_443
timestamp 1679235063
transform 1 0 41860 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_455
timestamp 1679235063
transform 1 0 42964 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_467
timestamp 1679235063
transform 1 0 44068 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_474
timestamp 1679235063
transform 1 0 44712 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_483
timestamp 1679235063
transform 1 0 45540 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_493
timestamp 1679235063
transform 1 0 46460 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_505
timestamp 1679235063
transform 1 0 47564 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1679235063
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1679235063
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_21
timestamp 1679235063
transform 1 0 3036 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_25
timestamp 1679235063
transform 1 0 3404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_30
timestamp 1679235063
transform 1 0 3864 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_42
timestamp 1679235063
transform 1 0 4968 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1679235063
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1679235063
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1679235063
transform 1 0 6808 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_74
timestamp 1679235063
transform 1 0 7912 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_86
timestamp 1679235063
transform 1 0 9016 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_98
timestamp 1679235063
transform 1 0 10120 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1679235063
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1679235063
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_123
timestamp 1679235063
transform 1 0 12420 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_136
timestamp 1679235063
transform 1 0 13616 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_149
timestamp 1679235063
transform 1 0 14812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_162
timestamp 1679235063
transform 1 0 16008 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_173
timestamp 1679235063
transform 1 0 17020 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1679235063
transform 1 0 18032 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_188
timestamp 1679235063
transform 1 0 18400 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1679235063
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1679235063
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1679235063
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_236
timestamp 1679235063
transform 1 0 22816 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_240
timestamp 1679235063
transform 1 0 23184 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_250
timestamp 1679235063
transform 1 0 24104 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_256
timestamp 1679235063
transform 1 0 24656 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1679235063
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1679235063
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_303
timestamp 1679235063
transform 1 0 28980 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_327
timestamp 1679235063
transform 1 0 31188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1679235063
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1679235063
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_342
timestamp 1679235063
transform 1 0 32568 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_346
timestamp 1679235063
transform 1 0 32936 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_368
timestamp 1679235063
transform 1 0 34960 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_375
timestamp 1679235063
transform 1 0 35604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1679235063
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1679235063
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_404
timestamp 1679235063
transform 1 0 38272 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_417
timestamp 1679235063
transform 1 0 39468 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_429
timestamp 1679235063
transform 1 0 40572 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_441
timestamp 1679235063
transform 1 0 41676 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1679235063
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_449
timestamp 1679235063
transform 1 0 42412 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_459
timestamp 1679235063
transform 1 0 43332 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_471
timestamp 1679235063
transform 1 0 44436 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_477
timestamp 1679235063
transform 1 0 44988 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_487
timestamp 1679235063
transform 1 0 45908 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_499
timestamp 1679235063
transform 1 0 47012 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1679235063
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_505
timestamp 1679235063
transform 1 0 47564 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_511
timestamp 1679235063
transform 1 0 48116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_515
timestamp 1679235063
transform 1 0 48484 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1679235063
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1679235063
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_21
timestamp 1679235063
transform 1 0 3036 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1679235063
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_34
timestamp 1679235063
transform 1 0 4232 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_46
timestamp 1679235063
transform 1 0 5336 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_58
timestamp 1679235063
transform 1 0 6440 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_70
timestamp 1679235063
transform 1 0 7544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1679235063
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1679235063
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1679235063
transform 1 0 9200 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_98
timestamp 1679235063
transform 1 0 10120 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_110
timestamp 1679235063
transform 1 0 11224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_135
timestamp 1679235063
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1679235063
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_152
timestamp 1679235063
transform 1 0 15088 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_165
timestamp 1679235063
transform 1 0 16284 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_171
timestamp 1679235063
transform 1 0 16836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_181
timestamp 1679235063
transform 1 0 17756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1679235063
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_199
timestamp 1679235063
transform 1 0 19412 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1679235063
transform 1 0 20424 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_237
timestamp 1679235063
transform 1 0 22908 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1679235063
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_253
timestamp 1679235063
transform 1 0 24380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_256
timestamp 1679235063
transform 1 0 24656 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_266
timestamp 1679235063
transform 1 0 25576 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_290
timestamp 1679235063
transform 1 0 27784 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_294
timestamp 1679235063
transform 1 0 28152 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1679235063
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1679235063
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_331
timestamp 1679235063
transform 1 0 31556 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_344
timestamp 1679235063
transform 1 0 32752 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_357
timestamp 1679235063
transform 1 0 33948 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_361
timestamp 1679235063
transform 1 0 34316 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1679235063
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_387
timestamp 1679235063
transform 1 0 36708 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_411
timestamp 1679235063
transform 1 0 38916 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1679235063
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_421
timestamp 1679235063
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_431
timestamp 1679235063
transform 1 0 40756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_443
timestamp 1679235063
transform 1 0 41860 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_455
timestamp 1679235063
transform 1 0 42964 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_467
timestamp 1679235063
transform 1 0 44068 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_474
timestamp 1679235063
transform 1 0 44712 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_477
timestamp 1679235063
transform 1 0 44988 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_487
timestamp 1679235063
transform 1 0 45908 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_499
timestamp 1679235063
transform 1 0 47012 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_511
timestamp 1679235063
transform 1 0 48116 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_515
timestamp 1679235063
transform 1 0 48484 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1679235063
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1679235063
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_21
timestamp 1679235063
transform 1 0 3036 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_25
timestamp 1679235063
transform 1 0 3404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_30
timestamp 1679235063
transform 1 0 3864 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_42
timestamp 1679235063
transform 1 0 4968 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1679235063
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_61
timestamp 1679235063
transform 1 0 6716 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_71
timestamp 1679235063
transform 1 0 7636 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_83
timestamp 1679235063
transform 1 0 8740 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_96
timestamp 1679235063
transform 1 0 9936 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_100
timestamp 1679235063
transform 1 0 10304 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1679235063
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_115
timestamp 1679235063
transform 1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_126
timestamp 1679235063
transform 1 0 12696 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_139
timestamp 1679235063
transform 1 0 13892 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_163
timestamp 1679235063
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1679235063
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_175
timestamp 1679235063
transform 1 0 17204 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_180
timestamp 1679235063
transform 1 0 17664 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_191
timestamp 1679235063
transform 1 0 18676 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_204
timestamp 1679235063
transform 1 0 19872 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_217
timestamp 1679235063
transform 1 0 21068 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1679235063
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_238
timestamp 1679235063
transform 1 0 23000 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_248
timestamp 1679235063
transform 1 0 23920 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_259
timestamp 1679235063
transform 1 0 24932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_263
timestamp 1679235063
transform 1 0 25300 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_273
timestamp 1679235063
transform 1 0 26220 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1679235063
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1679235063
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_292
timestamp 1679235063
transform 1 0 27968 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_305
timestamp 1679235063
transform 1 0 29164 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_318
timestamp 1679235063
transform 1 0 30360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_322
timestamp 1679235063
transform 1 0 30728 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_332
timestamp 1679235063
transform 1 0 31648 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1679235063
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_348
timestamp 1679235063
transform 1 0 33120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_361
timestamp 1679235063
transform 1 0 34316 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_365
timestamp 1679235063
transform 1 0 34684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_376
timestamp 1679235063
transform 1 0 35696 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_389
timestamp 1679235063
transform 1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_399
timestamp 1679235063
transform 1 0 37812 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_421
timestamp 1679235063
transform 1 0 39836 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_434
timestamp 1679235063
transform 1 0 41032 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 1679235063
transform 1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_449
timestamp 1679235063
transform 1 0 42412 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_459
timestamp 1679235063
transform 1 0 43332 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_471
timestamp 1679235063
transform 1 0 44436 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_477
timestamp 1679235063
transform 1 0 44988 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_487
timestamp 1679235063
transform 1 0 45908 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_491
timestamp 1679235063
transform 1 0 46276 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_505
timestamp 1679235063
transform 1 0 47564 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_511
timestamp 1679235063
transform 1 0 48116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_515
timestamp 1679235063
transform 1 0 48484 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_524
timestamp 1679235063
transform 1 0 49312 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1679235063
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_21
timestamp 1679235063
transform 1 0 3036 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1679235063
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_34
timestamp 1679235063
transform 1 0 4232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_46
timestamp 1679235063
transform 1 0 5336 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_58
timestamp 1679235063
transform 1 0 6440 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_70
timestamp 1679235063
transform 1 0 7544 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1679235063
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1679235063
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_88
timestamp 1679235063
transform 1 0 9200 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_94
timestamp 1679235063
transform 1 0 9752 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_118
timestamp 1679235063
transform 1 0 11960 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_131
timestamp 1679235063
transform 1 0 13156 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1679235063
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1679235063
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_152
timestamp 1679235063
transform 1 0 15088 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_165
timestamp 1679235063
transform 1 0 16284 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_169
timestamp 1679235063
transform 1 0 16652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_179
timestamp 1679235063
transform 1 0 17572 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_192
timestamp 1679235063
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_201
timestamp 1679235063
transform 1 0 19596 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_211
timestamp 1679235063
transform 1 0 20516 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_224
timestamp 1679235063
transform 1 0 21712 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_228
timestamp 1679235063
transform 1 0 22080 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_233
timestamp 1679235063
transform 1 0 22540 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_246
timestamp 1679235063
transform 1 0 23736 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_253
timestamp 1679235063
transform 1 0 24380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_256
timestamp 1679235063
transform 1 0 24656 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_266
timestamp 1679235063
transform 1 0 25576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_278
timestamp 1679235063
transform 1 0 26680 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_291
timestamp 1679235063
transform 1 0 27876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_303
timestamp 1679235063
transform 1 0 28980 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1679235063
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1679235063
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_320
timestamp 1679235063
transform 1 0 30544 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_324
timestamp 1679235063
transform 1 0 30912 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_329
timestamp 1679235063
transform 1 0 31372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_342
timestamp 1679235063
transform 1 0 32568 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_355
timestamp 1679235063
transform 1 0 33764 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1679235063
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_367
timestamp 1679235063
transform 1 0 34868 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_379
timestamp 1679235063
transform 1 0 35972 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_391
timestamp 1679235063
transform 1 0 37076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_415
timestamp 1679235063
transform 1 0 39284 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1679235063
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_421
timestamp 1679235063
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_443
timestamp 1679235063
transform 1 0 41860 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_455
timestamp 1679235063
transform 1 0 42964 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_467
timestamp 1679235063
transform 1 0 44068 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_474
timestamp 1679235063
transform 1 0 44712 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_477
timestamp 1679235063
transform 1 0 44988 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_489
timestamp 1679235063
transform 1 0 46092 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_496
timestamp 1679235063
transform 1 0 46736 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_508
timestamp 1679235063
transform 1 0 47840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_520
timestamp 1679235063
transform 1 0 48944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_526
timestamp 1679235063
transform 1 0 49496 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1679235063
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 1679235063
transform 1 0 3036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_25
timestamp 1679235063
transform 1 0 3404 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_30
timestamp 1679235063
transform 1 0 3864 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_42
timestamp 1679235063
transform 1 0 4968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1679235063
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1679235063
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_68
timestamp 1679235063
transform 1 0 7360 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_81
timestamp 1679235063
transform 1 0 8556 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_88
timestamp 1679235063
transform 1 0 9200 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_98
timestamp 1679235063
transform 1 0 10120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1679235063
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1679235063
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_116
timestamp 1679235063
transform 1 0 11776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_127
timestamp 1679235063
transform 1 0 12788 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_140
timestamp 1679235063
transform 1 0 13984 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1679235063
transform 1 0 15180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1679235063
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_173
timestamp 1679235063
transform 1 0 17020 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_184
timestamp 1679235063
transform 1 0 18032 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_192
timestamp 1679235063
transform 1 0 18768 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_217
timestamp 1679235063
transform 1 0 21068 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1679235063
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_236
timestamp 1679235063
transform 1 0 22816 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_249
timestamp 1679235063
transform 1 0 24012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_262
timestamp 1679235063
transform 1 0 25208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_275
timestamp 1679235063
transform 1 0 26404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1679235063
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1679235063
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_292
timestamp 1679235063
transform 1 0 27968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_304
timestamp 1679235063
transform 1 0 29072 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_308
timestamp 1679235063
transform 1 0 29440 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_318
timestamp 1679235063
transform 1 0 30360 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_322
timestamp 1679235063
transform 1 0 30728 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_332
timestamp 1679235063
transform 1 0 31648 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1679235063
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_348
timestamp 1679235063
transform 1 0 33120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_361
timestamp 1679235063
transform 1 0 34316 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_365
timestamp 1679235063
transform 1 0 34684 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_389
timestamp 1679235063
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_393
timestamp 1679235063
transform 1 0 37260 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_400
timestamp 1679235063
transform 1 0 37904 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_424
timestamp 1679235063
transform 1 0 40112 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_428
timestamp 1679235063
transform 1 0 40480 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_440
timestamp 1679235063
transform 1 0 41584 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_449
timestamp 1679235063
transform 1 0 42412 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_459
timestamp 1679235063
transform 1 0 43332 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_471
timestamp 1679235063
transform 1 0 44436 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_483
timestamp 1679235063
transform 1 0 45540 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_495
timestamp 1679235063
transform 1 0 46644 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_502
timestamp 1679235063
transform 1 0 47288 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_509
timestamp 1679235063
transform 1 0 47932 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_519
timestamp 1679235063
transform 1 0 48852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1679235063
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_21
timestamp 1679235063
transform 1 0 3036 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_29
timestamp 1679235063
transform 1 0 3772 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_32
timestamp 1679235063
transform 1 0 4048 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_42
timestamp 1679235063
transform 1 0 4968 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_54
timestamp 1679235063
transform 1 0 6072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_66
timestamp 1679235063
transform 1 0 7176 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_79
timestamp 1679235063
transform 1 0 8372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_85
timestamp 1679235063
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_96
timestamp 1679235063
transform 1 0 9936 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_108
timestamp 1679235063
transform 1 0 11040 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_121
timestamp 1679235063
transform 1 0 12236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_134
timestamp 1679235063
transform 1 0 13432 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1679235063
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_152
timestamp 1679235063
transform 1 0 15088 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_156
timestamp 1679235063
transform 1 0 15456 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_166
timestamp 1679235063
transform 1 0 16376 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_178
timestamp 1679235063
transform 1 0 17480 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_191
timestamp 1679235063
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1679235063
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_208
timestamp 1679235063
transform 1 0 20240 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_214
timestamp 1679235063
transform 1 0 20792 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_236
timestamp 1679235063
transform 1 0 22816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_240
timestamp 1679235063
transform 1 0 23184 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1679235063
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_257
timestamp 1679235063
transform 1 0 24748 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_279
timestamp 1679235063
transform 1 0 26772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_285
timestamp 1679235063
transform 1 0 27324 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_296
timestamp 1679235063
transform 1 0 28336 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_300
timestamp 1679235063
transform 1 0 28704 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1679235063
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_313
timestamp 1679235063
transform 1 0 29900 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_335
timestamp 1679235063
transform 1 0 31924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_348
timestamp 1679235063
transform 1 0 33120 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_361
timestamp 1679235063
transform 1 0 34316 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1679235063
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_387
timestamp 1679235063
transform 1 0 36708 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_400
timestamp 1679235063
transform 1 0 37904 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_413
timestamp 1679235063
transform 1 0 39100 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1679235063
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_421
timestamp 1679235063
transform 1 0 39836 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_432
timestamp 1679235063
transform 1 0 40848 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_444
timestamp 1679235063
transform 1 0 41952 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_456
timestamp 1679235063
transform 1 0 43056 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_468
timestamp 1679235063
transform 1 0 44160 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_477
timestamp 1679235063
transform 1 0 44988 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_487
timestamp 1679235063
transform 1 0 45908 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_499
timestamp 1679235063
transform 1 0 47012 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_511
timestamp 1679235063
transform 1 0 48116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_523
timestamp 1679235063
transform 1 0 49220 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1679235063
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_21
timestamp 1679235063
transform 1 0 3036 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_25
timestamp 1679235063
transform 1 0 3404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_30
timestamp 1679235063
transform 1 0 3864 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_42
timestamp 1679235063
transform 1 0 4968 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1679235063
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_63
timestamp 1679235063
transform 1 0 6900 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_73
timestamp 1679235063
transform 1 0 7820 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_85
timestamp 1679235063
transform 1 0 8924 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_97
timestamp 1679235063
transform 1 0 10028 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1679235063
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_117
timestamp 1679235063
transform 1 0 11868 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_128
timestamp 1679235063
transform 1 0 12880 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_132
timestamp 1679235063
transform 1 0 13248 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_141
timestamp 1679235063
transform 1 0 14076 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_153
timestamp 1679235063
transform 1 0 15180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1679235063
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_169
timestamp 1679235063
transform 1 0 16652 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_172
timestamp 1679235063
transform 1 0 16928 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_194
timestamp 1679235063
transform 1 0 18952 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_218
timestamp 1679235063
transform 1 0 21160 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1679235063
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_235
timestamp 1679235063
transform 1 0 22724 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_259
timestamp 1679235063
transform 1 0 24932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_272
timestamp 1679235063
transform 1 0 26128 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1679235063
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_291
timestamp 1679235063
transform 1 0 27876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_315
timestamp 1679235063
transform 1 0 30084 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_328
timestamp 1679235063
transform 1 0 31280 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_339
timestamp 1679235063
transform 1 0 32292 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_362
timestamp 1679235063
transform 1 0 34408 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_375
timestamp 1679235063
transform 1 0 35604 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_388
timestamp 1679235063
transform 1 0 36800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1679235063
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_403
timestamp 1679235063
transform 1 0 38180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_427
timestamp 1679235063
transform 1 0 40388 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_431
timestamp 1679235063
transform 1 0 40756 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_441
timestamp 1679235063
transform 1 0 41676 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1679235063
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_449
timestamp 1679235063
transform 1 0 42412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_459
timestamp 1679235063
transform 1 0 43332 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_471
timestamp 1679235063
transform 1 0 44436 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_483
timestamp 1679235063
transform 1 0 45540 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_495
timestamp 1679235063
transform 1 0 46644 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_502
timestamp 1679235063
transform 1 0 47288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_505
timestamp 1679235063
transform 1 0 47564 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_515
timestamp 1679235063
transform 1 0 48484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_523
timestamp 1679235063
transform 1 0 49220 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1679235063
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_21
timestamp 1679235063
transform 1 0 3036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1679235063
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_34
timestamp 1679235063
transform 1 0 4232 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_46
timestamp 1679235063
transform 1 0 5336 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_58
timestamp 1679235063
transform 1 0 6440 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_70
timestamp 1679235063
transform 1 0 7544 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1679235063
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_87
timestamp 1679235063
transform 1 0 9108 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_93
timestamp 1679235063
transform 1 0 9660 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_105
timestamp 1679235063
transform 1 0 10764 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_129
timestamp 1679235063
transform 1 0 12972 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_133
timestamp 1679235063
transform 1 0 13340 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1679235063
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1679235063
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_163
timestamp 1679235063
transform 1 0 16100 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_171
timestamp 1679235063
transform 1 0 16836 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_175
timestamp 1679235063
transform 1 0 17204 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_185
timestamp 1679235063
transform 1 0 18124 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1679235063
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1679235063
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_203
timestamp 1679235063
transform 1 0 19780 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_207
timestamp 1679235063
transform 1 0 20148 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_228
timestamp 1679235063
transform 1 0 22080 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_241
timestamp 1679235063
transform 1 0 23276 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1679235063
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1679235063
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_258
timestamp 1679235063
transform 1 0 24840 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_262
timestamp 1679235063
transform 1 0 25208 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_284
timestamp 1679235063
transform 1 0 27232 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_291
timestamp 1679235063
transform 1 0 27876 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_295
timestamp 1679235063
transform 1 0 28244 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1679235063
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1679235063
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_320
timestamp 1679235063
transform 1 0 30544 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_326
timestamp 1679235063
transform 1 0 31096 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_349
timestamp 1679235063
transform 1 0 33212 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1679235063
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1679235063
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_376
timestamp 1679235063
transform 1 0 35696 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_382
timestamp 1679235063
transform 1 0 36248 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_404
timestamp 1679235063
transform 1 0 38272 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_417
timestamp 1679235063
transform 1 0 39468 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_421
timestamp 1679235063
transform 1 0 39836 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_443
timestamp 1679235063
transform 1 0 41860 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_455
timestamp 1679235063
transform 1 0 42964 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_467
timestamp 1679235063
transform 1 0 44068 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_474
timestamp 1679235063
transform 1 0 44712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_477
timestamp 1679235063
transform 1 0 44988 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_487
timestamp 1679235063
transform 1 0 45908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_499
timestamp 1679235063
transform 1 0 47012 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_511
timestamp 1679235063
transform 1 0 48116 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_523
timestamp 1679235063
transform 1 0 49220 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1679235063
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_21
timestamp 1679235063
transform 1 0 3036 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_25
timestamp 1679235063
transform 1 0 3404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_30
timestamp 1679235063
transform 1 0 3864 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_42
timestamp 1679235063
transform 1 0 4968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1679235063
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1679235063
transform 1 0 6532 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_64
timestamp 1679235063
transform 1 0 6992 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_76
timestamp 1679235063
transform 1 0 8096 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_101
timestamp 1679235063
transform 1 0 10396 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1679235063
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1679235063
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_119
timestamp 1679235063
transform 1 0 12052 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_123
timestamp 1679235063
transform 1 0 12420 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_145
timestamp 1679235063
transform 1 0 14444 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_158
timestamp 1679235063
transform 1 0 15640 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1679235063
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1679235063
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_180
timestamp 1679235063
transform 1 0 17664 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_187
timestamp 1679235063
transform 1 0 18308 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_197
timestamp 1679235063
transform 1 0 19228 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1679235063
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1679235063
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_231
timestamp 1679235063
transform 1 0 22356 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_235
timestamp 1679235063
transform 1 0 22724 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_256
timestamp 1679235063
transform 1 0 24656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_263
timestamp 1679235063
transform 1 0 25300 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_274
timestamp 1679235063
transform 1 0 26312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1679235063
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_303
timestamp 1679235063
transform 1 0 28980 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_315
timestamp 1679235063
transform 1 0 30084 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_319
timestamp 1679235063
transform 1 0 30452 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_329
timestamp 1679235063
transform 1 0 31372 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1679235063
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_341
timestamp 1679235063
transform 1 0 32476 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_352
timestamp 1679235063
transform 1 0 33488 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_360
timestamp 1679235063
transform 1 0 34224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_382
timestamp 1679235063
transform 1 0 36248 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1679235063
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1679235063
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_403
timestamp 1679235063
transform 1 0 38180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_427
timestamp 1679235063
transform 1 0 40388 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_431
timestamp 1679235063
transform 1 0 40756 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_441
timestamp 1679235063
transform 1 0 41676 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1679235063
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_449
timestamp 1679235063
transform 1 0 42412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_459
timestamp 1679235063
transform 1 0 43332 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_471
timestamp 1679235063
transform 1 0 44436 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_483
timestamp 1679235063
transform 1 0 45540 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_495
timestamp 1679235063
transform 1 0 46644 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1679235063
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_517
timestamp 1679235063
transform 1 0 48668 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1679235063
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1679235063
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_21
timestamp 1679235063
transform 1 0 3036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1679235063
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_47
timestamp 1679235063
transform 1 0 5428 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_52
timestamp 1679235063
transform 1 0 5888 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_58
timestamp 1679235063
transform 1 0 6440 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_70
timestamp 1679235063
transform 1 0 7544 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1679235063
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_89
timestamp 1679235063
transform 1 0 9292 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_99
timestamp 1679235063
transform 1 0 10212 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_123
timestamp 1679235063
transform 1 0 12420 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_128
timestamp 1679235063
transform 1 0 12880 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1679235063
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1679235063
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_163
timestamp 1679235063
transform 1 0 16100 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_178
timestamp 1679235063
transform 1 0 17480 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_191
timestamp 1679235063
transform 1 0 18676 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1679235063
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_203
timestamp 1679235063
transform 1 0 19780 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_216
timestamp 1679235063
transform 1 0 20976 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_231
timestamp 1679235063
transform 1 0 22356 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_237
timestamp 1679235063
transform 1 0 22908 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_248
timestamp 1679235063
transform 1 0 23920 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1679235063
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_259
timestamp 1679235063
transform 1 0 24932 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_263
timestamp 1679235063
transform 1 0 25300 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_274
timestamp 1679235063
transform 1 0 26312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_287
timestamp 1679235063
transform 1 0 27508 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_300
timestamp 1679235063
transform 1 0 28704 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1679235063
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_320
timestamp 1679235063
transform 1 0 30544 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_326
timestamp 1679235063
transform 1 0 31096 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_340
timestamp 1679235063
transform 1 0 32384 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_353
timestamp 1679235063
transform 1 0 33580 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_357
timestamp 1679235063
transform 1 0 33948 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1679235063
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_365
timestamp 1679235063
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_376
timestamp 1679235063
transform 1 0 35696 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_380
timestamp 1679235063
transform 1 0 36064 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_402
timestamp 1679235063
transform 1 0 38088 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_415
timestamp 1679235063
transform 1 0 39284 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1679235063
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_421
timestamp 1679235063
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_443
timestamp 1679235063
transform 1 0 41860 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_455
timestamp 1679235063
transform 1 0 42964 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_467
timestamp 1679235063
transform 1 0 44068 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_474
timestamp 1679235063
transform 1 0 44712 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_477
timestamp 1679235063
transform 1 0 44988 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_487
timestamp 1679235063
transform 1 0 45908 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_499
timestamp 1679235063
transform 1 0 47012 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_505
timestamp 1679235063
transform 1 0 47564 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_515
timestamp 1679235063
transform 1 0 48484 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_523
timestamp 1679235063
transform 1 0 49220 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1679235063
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1679235063
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1679235063
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_45
timestamp 1679235063
transform 1 0 5244 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1679235063
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_63
timestamp 1679235063
transform 1 0 6900 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_73
timestamp 1679235063
transform 1 0 7820 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_85
timestamp 1679235063
transform 1 0 8924 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_97
timestamp 1679235063
transform 1 0 10028 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1679235063
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_119
timestamp 1679235063
transform 1 0 12052 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_132
timestamp 1679235063
transform 1 0 13248 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_136
timestamp 1679235063
transform 1 0 13616 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_141
timestamp 1679235063
transform 1 0 14076 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_153
timestamp 1679235063
transform 1 0 15180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1679235063
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1679235063
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1679235063
transform 1 0 17572 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_206
timestamp 1679235063
transform 1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_210
timestamp 1679235063
transform 1 0 20424 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1679235063
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1679235063
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_236
timestamp 1679235063
transform 1 0 22816 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_240
timestamp 1679235063
transform 1 0 23184 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_251
timestamp 1679235063
transform 1 0 24196 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_264
timestamp 1679235063
transform 1 0 25392 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_268
timestamp 1679235063
transform 1 0 25760 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1679235063
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_285
timestamp 1679235063
transform 1 0 27324 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_296
timestamp 1679235063
transform 1 0 28336 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_300
timestamp 1679235063
transform 1 0 28704 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_311
timestamp 1679235063
transform 1 0 29716 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_318
timestamp 1679235063
transform 1 0 30360 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_322
timestamp 1679235063
transform 1 0 30728 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1679235063
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_339
timestamp 1679235063
transform 1 0 32292 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_351
timestamp 1679235063
transform 1 0 33396 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_364
timestamp 1679235063
transform 1 0 34592 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_368
timestamp 1679235063
transform 1 0 34960 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_375
timestamp 1679235063
transform 1 0 35604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_390
timestamp 1679235063
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1679235063
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_403
timestamp 1679235063
transform 1 0 38180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_427
timestamp 1679235063
transform 1 0 40388 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_440
timestamp 1679235063
transform 1 0 41584 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_449
timestamp 1679235063
transform 1 0 42412 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_459
timestamp 1679235063
transform 1 0 43332 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_471
timestamp 1679235063
transform 1 0 44436 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_483
timestamp 1679235063
transform 1 0 45540 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_495
timestamp 1679235063
transform 1 0 46644 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1679235063
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_519
timestamp 1679235063
transform 1 0 48852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1679235063
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1679235063
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_21
timestamp 1679235063
transform 1 0 3036 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1679235063
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_47
timestamp 1679235063
transform 1 0 5428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_67
timestamp 1679235063
transform 1 0 7268 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_72
timestamp 1679235063
transform 1 0 7728 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1679235063
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1679235063
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_90
timestamp 1679235063
transform 1 0 9384 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_102
timestamp 1679235063
transform 1 0 10488 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1679235063
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1679235063
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_141
timestamp 1679235063
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_144
timestamp 1679235063
transform 1 0 14352 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_154
timestamp 1679235063
transform 1 0 15272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_169
timestamp 1679235063
transform 1 0 16652 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1679235063
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1679235063
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1679235063
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_234
timestamp 1679235063
transform 1 0 22632 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_238
timestamp 1679235063
transform 1 0 23000 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1679235063
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_257
timestamp 1679235063
transform 1 0 24748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_279
timestamp 1679235063
transform 1 0 26772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_303
timestamp 1679235063
transform 1 0 28980 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1679235063
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1679235063
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_320
timestamp 1679235063
transform 1 0 30544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_327
timestamp 1679235063
transform 1 0 31188 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_342
timestamp 1679235063
transform 1 0 32568 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_355
timestamp 1679235063
transform 1 0 33764 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1679235063
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1679235063
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_376
timestamp 1679235063
transform 1 0 35696 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_389
timestamp 1679235063
transform 1 0 36892 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_393
timestamp 1679235063
transform 1 0 37260 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_405
timestamp 1679235063
transform 1 0 38364 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_418
timestamp 1679235063
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1679235063
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_432
timestamp 1679235063
transform 1 0 40848 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_444
timestamp 1679235063
transform 1 0 41952 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_456
timestamp 1679235063
transform 1 0 43056 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_468
timestamp 1679235063
transform 1 0 44160 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_477
timestamp 1679235063
transform 1 0 44988 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_487
timestamp 1679235063
transform 1 0 45908 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_499
timestamp 1679235063
transform 1 0 47012 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_511
timestamp 1679235063
transform 1 0 48116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_523
timestamp 1679235063
transform 1 0 49220 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1679235063
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_21
timestamp 1679235063
transform 1 0 3036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_41
timestamp 1679235063
transform 1 0 4876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_45
timestamp 1679235063
transform 1 0 5244 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1679235063
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1679235063
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_75
timestamp 1679235063
transform 1 0 8004 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_80
timestamp 1679235063
transform 1 0 8464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_86
timestamp 1679235063
transform 1 0 9016 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_98
timestamp 1679235063
transform 1 0 10120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1679235063
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_113
timestamp 1679235063
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_120
timestamp 1679235063
transform 1 0 12144 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_132
timestamp 1679235063
transform 1 0 13248 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_156
timestamp 1679235063
transform 1 0 15456 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_160
timestamp 1679235063
transform 1 0 15824 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1679235063
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_169
timestamp 1679235063
transform 1 0 16652 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_172
timestamp 1679235063
transform 1 0 16928 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_194
timestamp 1679235063
transform 1 0 18952 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_199
timestamp 1679235063
transform 1 0 19412 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1679235063
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1679235063
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_236
timestamp 1679235063
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_260
timestamp 1679235063
transform 1 0 25024 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_266
timestamp 1679235063
transform 1 0 25576 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1679235063
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1679235063
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_292
timestamp 1679235063
transform 1 0 27968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_304
timestamp 1679235063
transform 1 0 29072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_310
timestamp 1679235063
transform 1 0 29624 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_322
timestamp 1679235063
transform 1 0 30728 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1679235063
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1679235063
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_359
timestamp 1679235063
transform 1 0 34132 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_365
timestamp 1679235063
transform 1 0 34684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_376
timestamp 1679235063
transform 1 0 35696 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1679235063
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_399
timestamp 1679235063
transform 1 0 37812 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_421
timestamp 1679235063
transform 1 0 39836 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_434
timestamp 1679235063
transform 1 0 41032 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_446
timestamp 1679235063
transform 1 0 42136 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_449
timestamp 1679235063
transform 1 0 42412 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_459
timestamp 1679235063
transform 1 0 43332 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_471
timestamp 1679235063
transform 1 0 44436 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_483
timestamp 1679235063
transform 1 0 45540 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_495
timestamp 1679235063
transform 1 0 46644 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1679235063
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_505
timestamp 1679235063
transform 1 0 47564 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_517
timestamp 1679235063
transform 1 0 48668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1679235063
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1679235063
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_21
timestamp 1679235063
transform 1 0 3036 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1679235063
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1679235063
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_67
timestamp 1679235063
transform 1 0 7268 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_72
timestamp 1679235063
transform 1 0 7728 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1679235063
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_91
timestamp 1679235063
transform 1 0 9476 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_101
timestamp 1679235063
transform 1 0 10396 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_113
timestamp 1679235063
transform 1 0 11500 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_125
timestamp 1679235063
transform 1 0 12604 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1679235063
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_143
timestamp 1679235063
transform 1 0 14260 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_165
timestamp 1679235063
transform 1 0 16284 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_170
timestamp 1679235063
transform 1 0 16744 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_181
timestamp 1679235063
transform 1 0 17756 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1679235063
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_197
timestamp 1679235063
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_209
timestamp 1679235063
transform 1 0 20332 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_215
timestamp 1679235063
transform 1 0 20884 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_237
timestamp 1679235063
transform 1 0 22908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1679235063
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_253
timestamp 1679235063
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_265
timestamp 1679235063
transform 1 0 25484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_278
timestamp 1679235063
transform 1 0 26680 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_284
timestamp 1679235063
transform 1 0 27232 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_295
timestamp 1679235063
transform 1 0 28244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_303
timestamp 1679235063
transform 1 0 28980 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1679235063
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1679235063
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_320
timestamp 1679235063
transform 1 0 30544 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_333
timestamp 1679235063
transform 1 0 31740 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_346
timestamp 1679235063
transform 1 0 32936 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_359
timestamp 1679235063
transform 1 0 34132 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1679235063
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1679235063
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_387
timestamp 1679235063
transform 1 0 36708 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_394
timestamp 1679235063
transform 1 0 37352 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_418
timestamp 1679235063
transform 1 0 39560 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_421
timestamp 1679235063
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_432
timestamp 1679235063
transform 1 0 40848 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_444
timestamp 1679235063
transform 1 0 41952 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_456
timestamp 1679235063
transform 1 0 43056 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_468
timestamp 1679235063
transform 1 0 44160 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_477
timestamp 1679235063
transform 1 0 44988 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_487
timestamp 1679235063
transform 1 0 45908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_499
timestamp 1679235063
transform 1 0 47012 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_511
timestamp 1679235063
transform 1 0 48116 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_523
timestamp 1679235063
transform 1 0 49220 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1679235063
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1679235063
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_41
timestamp 1679235063
transform 1 0 4876 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_45
timestamp 1679235063
transform 1 0 5244 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1679235063
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1679235063
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_75
timestamp 1679235063
transform 1 0 8004 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_95
timestamp 1679235063
transform 1 0 9844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_100
timestamp 1679235063
transform 1 0 10304 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1679235063
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_113
timestamp 1679235063
transform 1 0 11500 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1679235063
transform 1 0 11960 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_128
timestamp 1679235063
transform 1 0 12880 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_140
timestamp 1679235063
transform 1 0 13984 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_153
timestamp 1679235063
transform 1 0 15180 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1679235063
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_169
timestamp 1679235063
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_178
timestamp 1679235063
transform 1 0 17480 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_202
timestamp 1679235063
transform 1 0 19688 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_215
timestamp 1679235063
transform 1 0 20884 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1679235063
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1679235063
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_248
timestamp 1679235063
transform 1 0 23920 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_272
timestamp 1679235063
transform 1 0 26128 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1679235063
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_292
timestamp 1679235063
transform 1 0 27968 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_296
timestamp 1679235063
transform 1 0 28336 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_307
timestamp 1679235063
transform 1 0 29348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_320
timestamp 1679235063
transform 1 0 30544 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_333
timestamp 1679235063
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1679235063
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_348
timestamp 1679235063
transform 1 0 33120 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_352
timestamp 1679235063
transform 1 0 33488 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_376
timestamp 1679235063
transform 1 0 35696 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_389
timestamp 1679235063
transform 1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_393
timestamp 1679235063
transform 1 0 37260 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_400
timestamp 1679235063
transform 1 0 37904 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_424
timestamp 1679235063
transform 1 0 40112 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_437
timestamp 1679235063
transform 1 0 41308 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_441
timestamp 1679235063
transform 1 0 41676 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1679235063
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_449
timestamp 1679235063
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_459
timestamp 1679235063
transform 1 0 43332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_471
timestamp 1679235063
transform 1 0 44436 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_483
timestamp 1679235063
transform 1 0 45540 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_495
timestamp 1679235063
transform 1 0 46644 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_502
timestamp 1679235063
transform 1 0 47288 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_505
timestamp 1679235063
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_515
timestamp 1679235063
transform 1 0 48484 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1679235063
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1679235063
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_21
timestamp 1679235063
transform 1 0 3036 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1679235063
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_47
timestamp 1679235063
transform 1 0 5428 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_67
timestamp 1679235063
transform 1 0 7268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_72
timestamp 1679235063
transform 1 0 7728 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1679235063
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1679235063
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_103
timestamp 1679235063
transform 1 0 10580 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_108
timestamp 1679235063
transform 1 0 11040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_114
timestamp 1679235063
transform 1 0 11592 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_134
timestamp 1679235063
transform 1 0 13432 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1679235063
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_147
timestamp 1679235063
transform 1 0 14628 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_171
timestamp 1679235063
transform 1 0 16836 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_176
timestamp 1679235063
transform 1 0 17296 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1679235063
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_199
timestamp 1679235063
transform 1 0 19412 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_210
timestamp 1679235063
transform 1 0 20424 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_223
timestamp 1679235063
transform 1 0 21620 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_236
timestamp 1679235063
transform 1 0 22816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_240
timestamp 1679235063
transform 1 0 23184 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1679235063
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_255
timestamp 1679235063
transform 1 0 24564 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_266
timestamp 1679235063
transform 1 0 25576 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_279
timestamp 1679235063
transform 1 0 26772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_294
timestamp 1679235063
transform 1 0 28152 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1679235063
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1679235063
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_319
timestamp 1679235063
transform 1 0 30452 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_344
timestamp 1679235063
transform 1 0 32752 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_357
timestamp 1679235063
transform 1 0 33948 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1679235063
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1679235063
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_376
timestamp 1679235063
transform 1 0 35696 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_390
timestamp 1679235063
transform 1 0 36984 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_403
timestamp 1679235063
transform 1 0 38180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_416
timestamp 1679235063
transform 1 0 39376 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_421
timestamp 1679235063
transform 1 0 39836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_432
timestamp 1679235063
transform 1 0 40848 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_445
timestamp 1679235063
transform 1 0 42044 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_457
timestamp 1679235063
transform 1 0 43148 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_469
timestamp 1679235063
transform 1 0 44252 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1679235063
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_477
timestamp 1679235063
transform 1 0 44988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_487
timestamp 1679235063
transform 1 0 45908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_499
timestamp 1679235063
transform 1 0 47012 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_511
timestamp 1679235063
transform 1 0 48116 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_523
timestamp 1679235063
transform 1 0 49220 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1679235063
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_21
timestamp 1679235063
transform 1 0 3036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_25
timestamp 1679235063
transform 1 0 3404 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1679235063
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1679235063
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_65
timestamp 1679235063
transform 1 0 7084 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_85
timestamp 1679235063
transform 1 0 8924 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_92
timestamp 1679235063
transform 1 0 9568 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1679235063
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1679235063
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_125
timestamp 1679235063
transform 1 0 12604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_129
timestamp 1679235063
transform 1 0 12972 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_146
timestamp 1679235063
transform 1 0 14536 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1679235063
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1679235063
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_191
timestamp 1679235063
transform 1 0 18676 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_195
timestamp 1679235063
transform 1 0 19044 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_220
timestamp 1679235063
transform 1 0 21344 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_225
timestamp 1679235063
transform 1 0 21804 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_230
timestamp 1679235063
transform 1 0 22264 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_241
timestamp 1679235063
transform 1 0 23276 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_254
timestamp 1679235063
transform 1 0 24472 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1679235063
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_283
timestamp 1679235063
transform 1 0 27140 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_289
timestamp 1679235063
transform 1 0 27692 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_313
timestamp 1679235063
transform 1 0 29900 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_326
timestamp 1679235063
transform 1 0 31096 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1679235063
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1679235063
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_348
timestamp 1679235063
transform 1 0 33120 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_352
timestamp 1679235063
transform 1 0 33488 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_373
timestamp 1679235063
transform 1 0 35420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_377
timestamp 1679235063
transform 1 0 35788 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_389
timestamp 1679235063
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1679235063
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_415
timestamp 1679235063
transform 1 0 39284 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_428
timestamp 1679235063
transform 1 0 40480 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_441
timestamp 1679235063
transform 1 0 41676 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1679235063
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1679235063
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_459
timestamp 1679235063
transform 1 0 43332 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_474
timestamp 1679235063
transform 1 0 44712 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_486
timestamp 1679235063
transform 1 0 45816 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_498
timestamp 1679235063
transform 1 0 46920 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_505
timestamp 1679235063
transform 1 0 47564 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_515
timestamp 1679235063
transform 1 0 48484 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1679235063
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1679235063
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_21
timestamp 1679235063
transform 1 0 3036 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_29
timestamp 1679235063
transform 1 0 3772 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_32
timestamp 1679235063
transform 1 0 4048 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1679235063
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1679235063
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1679235063
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_85
timestamp 1679235063
transform 1 0 8924 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_88
timestamp 1679235063
transform 1 0 9200 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_98
timestamp 1679235063
transform 1 0 10120 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_118
timestamp 1679235063
transform 1 0 11960 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1679235063
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_145
timestamp 1679235063
transform 1 0 14444 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_150
timestamp 1679235063
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1679235063
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1679235063
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1679235063
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_210
timestamp 1679235063
transform 1 0 20424 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_237
timestamp 1679235063
transform 1 0 22908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1679235063
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1679235063
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_259
timestamp 1679235063
transform 1 0 24932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_263
timestamp 1679235063
transform 1 0 25300 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_284
timestamp 1679235063
transform 1 0 27232 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_297
timestamp 1679235063
transform 1 0 28428 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_305
timestamp 1679235063
transform 1 0 29164 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_311
timestamp 1679235063
transform 1 0 29716 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_333
timestamp 1679235063
transform 1 0 31740 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_358
timestamp 1679235063
transform 1 0 34040 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1679235063
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_387
timestamp 1679235063
transform 1 0 36708 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_413
timestamp 1679235063
transform 1 0 39100 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_418
timestamp 1679235063
transform 1 0 39560 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1679235063
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_433
timestamp 1679235063
transform 1 0 40940 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_439
timestamp 1679235063
transform 1 0 41492 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_464
timestamp 1679235063
transform 1 0 43792 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_472
timestamp 1679235063
transform 1 0 44528 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_477
timestamp 1679235063
transform 1 0 44988 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_487
timestamp 1679235063
transform 1 0 45908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_499
timestamp 1679235063
transform 1 0 47012 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_511
timestamp 1679235063
transform 1 0 48116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_523
timestamp 1679235063
transform 1 0 49220 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_3
timestamp 1679235063
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1679235063
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1679235063
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1679235063
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_69
timestamp 1679235063
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_73
timestamp 1679235063
transform 1 0 7820 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1679235063
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1679235063
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1679235063
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_126
timestamp 1679235063
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1679235063
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1679235063
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_169
timestamp 1679235063
transform 1 0 16652 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_172
timestamp 1679235063
transform 1 0 16928 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_177
timestamp 1679235063
transform 1 0 17388 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_197
timestamp 1679235063
transform 1 0 19228 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1679235063
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1679235063
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_243
timestamp 1679235063
transform 1 0 23460 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_248
timestamp 1679235063
transform 1 0 23920 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_254
timestamp 1679235063
transform 1 0 24472 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1679235063
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_285
timestamp 1679235063
transform 1 0 27324 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_297
timestamp 1679235063
transform 1 0 28428 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_309
timestamp 1679235063
transform 1 0 29532 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_315
timestamp 1679235063
transform 1 0 30084 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_326
timestamp 1679235063
transform 1 0 31096 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1679235063
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_337
timestamp 1679235063
transform 1 0 32108 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_346
timestamp 1679235063
transform 1 0 32936 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_370
timestamp 1679235063
transform 1 0 35144 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_376
timestamp 1679235063
transform 1 0 35696 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_388
timestamp 1679235063
transform 1 0 36800 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1679235063
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_418
timestamp 1679235063
transform 1 0 39560 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_422
timestamp 1679235063
transform 1 0 39928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_432
timestamp 1679235063
transform 1 0 40848 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_444
timestamp 1679235063
transform 1 0 41952 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_449
timestamp 1679235063
transform 1 0 42412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_459
timestamp 1679235063
transform 1 0 43332 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_471
timestamp 1679235063
transform 1 0 44436 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_481
timestamp 1679235063
transform 1 0 45356 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_495
timestamp 1679235063
transform 1 0 46644 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1679235063
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_505
timestamp 1679235063
transform 1 0 47564 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_512
timestamp 1679235063
transform 1 0 48208 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_525
timestamp 1679235063
transform 1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_3
timestamp 1679235063
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_8
timestamp 1679235063
transform 1 0 1840 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1679235063
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1679235063
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1679235063
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1679235063
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1679235063
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1679235063
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1679235063
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_85
timestamp 1679235063
transform 1 0 8924 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_92
timestamp 1679235063
transform 1 0 9568 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1679235063
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_113
timestamp 1679235063
transform 1 0 11500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_120
timestamp 1679235063
transform 1 0 12144 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1679235063
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1679235063
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1679235063
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1679235063
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1679235063
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_174
timestamp 1679235063
transform 1 0 17112 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1679235063
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1679235063
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_219
timestamp 1679235063
transform 1 0 21252 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_225
timestamp 1679235063
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_243
timestamp 1679235063
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1679235063
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_255
timestamp 1679235063
transform 1 0 24564 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_266
timestamp 1679235063
transform 1 0 25576 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_278
timestamp 1679235063
transform 1 0 26680 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_281
timestamp 1679235063
transform 1 0 26956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_287
timestamp 1679235063
transform 1 0 27508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_300
timestamp 1679235063
transform 1 0 28704 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1679235063
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_319
timestamp 1679235063
transform 1 0 30452 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_331
timestamp 1679235063
transform 1 0 31556 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_335
timestamp 1679235063
transform 1 0 31924 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1679235063
transform 1 0 32108 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_348
timestamp 1679235063
transform 1 0 33120 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_360
timestamp 1679235063
transform 1 0 34224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1679235063
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_376
timestamp 1679235063
transform 1 0 35696 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_389
timestamp 1679235063
transform 1 0 36892 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_393
timestamp 1679235063
transform 1 0 37260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_404
timestamp 1679235063
transform 1 0 38272 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_417
timestamp 1679235063
transform 1 0 39468 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1679235063
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_432
timestamp 1679235063
transform 1 0 40848 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_444
timestamp 1679235063
transform 1 0 41952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_449
timestamp 1679235063
transform 1 0 42412 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_459
timestamp 1679235063
transform 1 0 43332 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_471
timestamp 1679235063
transform 1 0 44436 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1679235063
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1679235063
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_487
timestamp 1679235063
transform 1 0 45908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_499
timestamp 1679235063
transform 1 0 47012 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_503
timestamp 1679235063
transform 1 0 47380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_505
timestamp 1679235063
transform 1 0 47564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_511
timestamp 1679235063
transform 1 0 48116 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_525
timestamp 1679235063
transform 1 0 49404 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 48208 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1679235063
transform 1 0 47748 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1679235063
transform 1 0 8280 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1679235063
transform 1 0 12328 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold5 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6900 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1679235063
transform 1 0 18400 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1679235063
transform 1 0 19412 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1679235063
transform 1 0 12144 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1679235063
transform 1 0 19504 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold10
timestamp 1679235063
transform 1 0 44160 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1679235063
transform 1 0 42596 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1679235063
transform 1 0 30912 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1679235063
transform 1 0 28244 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1679235063
transform 1 0 42596 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1679235063
transform 1 0 41124 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1679235063
transform 1 0 9660 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1679235063
transform 1 0 7912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1679235063
transform 1 0 41216 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1679235063
transform 1 0 7084 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1679235063
transform 1 0 46276 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1679235063
transform 1 0 9200 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold22
timestamp 1679235063
transform 1 0 24472 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold23
timestamp 1679235063
transform 1 0 25944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1679235063
transform 1 0 42228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1679235063
transform 1 0 23368 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1679235063
transform 1 0 37444 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1679235063
transform 1 0 42596 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 12144 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1679235063
transform 1 0 47748 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1679235063
transform 1 0 4232 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1679235063
transform 1 0 19688 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1679235063
transform 1 0 42320 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1679235063
transform 1 0 43424 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1679235063
transform 1 0 43332 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1679235063
transform 1 0 10488 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1679235063
transform 1 0 9200 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1679235063
transform 1 0 5704 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1679235063
transform 1 0 3496 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1679235063
transform 1 0 45172 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1679235063
transform 1 0 5336 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold41
timestamp 1679235063
transform 1 0 36064 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1679235063
transform 1 0 13064 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1679235063
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold44
timestamp 1679235063
transform 1 0 34868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold45
timestamp 1679235063
transform 1 0 44804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold46
timestamp 1679235063
transform 1 0 40020 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1679235063
transform 1 0 16836 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold48
timestamp 1679235063
transform 1 0 7176 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold49
timestamp 1679235063
transform 1 0 46276 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold50
timestamp 1679235063
transform 1 0 29716 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold51
timestamp 1679235063
transform 1 0 26312 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold52
timestamp 1679235063
transform 1 0 8280 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold53
timestamp 1679235063
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold54
timestamp 1679235063
transform 1 0 45172 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold55
timestamp 1679235063
transform 1 0 47380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold56
timestamp 1679235063
transform 1 0 7084 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold57
timestamp 1679235063
transform 1 0 21988 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold58
timestamp 1679235063
transform 1 0 34040 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold59
timestamp 1679235063
transform 1 0 43700 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold60
timestamp 1679235063
transform 1 0 9660 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold61
timestamp 1679235063
transform 1 0 9384 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold62
timestamp 1679235063
transform 1 0 47748 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold63
timestamp 1679235063
transform 1 0 18216 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold64
timestamp 1679235063
transform 1 0 44804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold65
timestamp 1679235063
transform 1 0 38548 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold66
timestamp 1679235063
transform 1 0 5336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold67
timestamp 1679235063
transform 1 0 28704 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold68
timestamp 1679235063
transform 1 0 4232 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold69
timestamp 1679235063
transform 1 0 9384 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold70
timestamp 1679235063
transform 1 0 27140 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold71
timestamp 1679235063
transform 1 0 20792 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold72
timestamp 1679235063
transform 1 0 43424 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold73
timestamp 1679235063
transform 1 0 30820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold74
timestamp 1679235063
transform 1 0 45172 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold75
timestamp 1679235063
transform 1 0 7176 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold76
timestamp 1679235063
transform 1 0 25944 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold77
timestamp 1679235063
transform 1 0 40020 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold78
timestamp 1679235063
transform 1 0 9292 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold79
timestamp 1679235063
transform 1 0 24656 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold80
timestamp 1679235063
transform 1 0 9568 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold81
timestamp 1679235063
transform 1 0 19780 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold82
timestamp 1679235063
transform 1 0 26128 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold83
timestamp 1679235063
transform 1 0 6808 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold84
timestamp 1679235063
transform 1 0 41124 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold85
timestamp 1679235063
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold86
timestamp 1679235063
transform 1 0 13248 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold87
timestamp 1679235063
transform 1 0 30912 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold88
timestamp 1679235063
transform 1 0 10488 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold89
timestamp 1679235063
transform 1 0 5336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold90
timestamp 1679235063
transform 1 0 22908 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold91
timestamp 1679235063
transform 1 0 10488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold92
timestamp 1679235063
transform 1 0 39836 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold93
timestamp 1679235063
transform 1 0 25208 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold94
timestamp 1679235063
transform 1 0 43700 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold95
timestamp 1679235063
transform 1 0 14536 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold96
timestamp 1679235063
transform 1 0 43700 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold97
timestamp 1679235063
transform 1 0 10488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold98
timestamp 1679235063
transform 1 0 41216 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold99
timestamp 1679235063
transform 1 0 39744 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold100
timestamp 1679235063
transform 1 0 38640 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold101
timestamp 1679235063
transform 1 0 20608 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold102
timestamp 1679235063
transform 1 0 46552 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold103
timestamp 1679235063
transform 1 0 28244 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold104
timestamp 1679235063
transform 1 0 41400 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold105
timestamp 1679235063
transform 1 0 15640 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold106
timestamp 1679235063
transform 1 0 48484 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold107
timestamp 1679235063
transform 1 0 21712 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold108
timestamp 1679235063
transform 1 0 33580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold109
timestamp 1679235063
transform 1 0 28612 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold110
timestamp 1679235063
transform 1 0 42228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold111
timestamp 1679235063
transform 1 0 47380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold112
timestamp 1679235063
transform 1 0 7084 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold113
timestamp 1679235063
transform 1 0 14444 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold114
timestamp 1679235063
transform 1 0 38456 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold115
timestamp 1679235063
transform 1 0 45724 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold116
timestamp 1679235063
transform 1 0 13064 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold117
timestamp 1679235063
transform 1 0 45172 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold118
timestamp 1679235063
transform 1 0 45172 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold119
timestamp 1679235063
transform 1 0 45908 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold120
timestamp 1679235063
transform 1 0 39652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold121
timestamp 1679235063
transform 1 0 16744 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold122
timestamp 1679235063
transform 1 0 41400 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold123
timestamp 1679235063
transform 1 0 38640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold124
timestamp 1679235063
transform 1 0 9384 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold125
timestamp 1679235063
transform 1 0 10764 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold126
timestamp 1679235063
transform 1 0 28796 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold127
timestamp 1679235063
transform 1 0 32292 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold128
timestamp 1679235063
transform 1 0 45172 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold129
timestamp 1679235063
transform 1 0 43700 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold130
timestamp 1679235063
transform 1 0 23368 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold131
timestamp 1679235063
transform 1 0 29716 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold132
timestamp 1679235063
transform 1 0 27508 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold133
timestamp 1679235063
transform 1 0 42228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold134
timestamp 1679235063
transform 1 0 27416 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold135
timestamp 1679235063
transform 1 0 3128 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold136
timestamp 1679235063
transform 1 0 10764 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold137
timestamp 1679235063
transform 1 0 31096 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold138
timestamp 1679235063
transform 1 0 5704 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold139
timestamp 1679235063
transform 1 0 36064 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold140
timestamp 1679235063
transform 1 0 42596 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold141
timestamp 1679235063
transform 1 0 5704 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold142
timestamp 1679235063
transform 1 0 46276 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold143
timestamp 1679235063
transform 1 0 48484 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold144
timestamp 1679235063
transform 1 0 45908 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold145
timestamp 1679235063
transform 1 0 9384 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold146
timestamp 1679235063
transform 1 0 7912 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold147
timestamp 1679235063
transform 1 0 9660 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold148
timestamp 1679235063
transform 1 0 25944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold149
timestamp 1679235063
transform 1 0 47104 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold150
timestamp 1679235063
transform 1 0 48116 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold151
timestamp 1679235063
transform 1 0 48484 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold152
timestamp 1679235063
transform 1 0 47380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold153
timestamp 1679235063
transform 1 0 9660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold154
timestamp 1679235063
transform 1 0 10028 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold155
timestamp 1679235063
transform 1 0 11132 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold156
timestamp 1679235063
transform 1 0 13432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold157
timestamp 1679235063
transform 1 0 7912 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold158
timestamp 1679235063
transform 1 0 4232 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold159
timestamp 1679235063
transform 1 0 17112 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold160
timestamp 1679235063
transform 1 0 16468 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold161
timestamp 1679235063
transform 1 0 19504 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold162
timestamp 1679235063
transform 1 0 14536 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold163
timestamp 1679235063
transform 1 0 41216 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold164
timestamp 1679235063
transform 1 0 42320 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold165
timestamp 1679235063
transform 1 0 17572 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold166
timestamp 1679235063
transform 1 0 20424 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold167
timestamp 1679235063
transform 1 0 11776 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold168
timestamp 1679235063
transform 1 0 4232 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold169
timestamp 1679235063
transform 1 0 42320 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold170
timestamp 1679235063
transform 1 0 43700 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold171
timestamp 1679235063
transform 1 0 27140 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold172
timestamp 1679235063
transform 1 0 29716 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold173
timestamp 1679235063
transform 1 0 21344 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold174
timestamp 1679235063
transform 1 0 20240 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold175
timestamp 1679235063
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold176
timestamp 1679235063
transform 1 0 9384 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold177
timestamp 1679235063
transform 1 0 30820 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold178
timestamp 1679235063
transform 1 0 32292 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold179
timestamp 1679235063
transform 1 0 40940 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold180
timestamp 1679235063
transform 1 0 40020 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold181
timestamp 1679235063
transform 1 0 9292 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold182
timestamp 1679235063
transform 1 0 9476 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold183
timestamp 1679235063
transform 1 0 8188 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold184
timestamp 1679235063
transform 1 0 10304 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold185
timestamp 1679235063
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold186
timestamp 1679235063
transform 1 0 7360 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold187
timestamp 1679235063
transform 1 0 41216 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold188
timestamp 1679235063
transform 1 0 42412 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold189
timestamp 1679235063
transform 1 0 44804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold190
timestamp 1679235063
transform 1 0 45908 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold191
timestamp 1679235063
transform 1 0 24564 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold192
timestamp 1679235063
transform 1 0 18584 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold193
timestamp 1679235063
transform 1 0 23368 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold194
timestamp 1679235063
transform 1 0 24656 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold195
timestamp 1679235063
transform 1 0 41216 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold196
timestamp 1679235063
transform 1 0 42596 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold197
timestamp 1679235063
transform 1 0 5336 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold198
timestamp 1679235063
transform 1 0 4600 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold199
timestamp 1679235063
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold200
timestamp 1679235063
transform 1 0 11684 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold201
timestamp 1679235063
transform 1 0 25944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold202
timestamp 1679235063
transform 1 0 29716 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold203
timestamp 1679235063
transform 1 0 43700 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold204
timestamp 1679235063
transform 1 0 43700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold205
timestamp 1679235063
transform 1 0 42596 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold206
timestamp 1679235063
transform 1 0 43700 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold207
timestamp 1679235063
transform 1 0 15640 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold208
timestamp 1679235063
transform 1 0 18492 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold209
timestamp 1679235063
transform 1 0 43332 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold210
timestamp 1679235063
transform 1 0 43700 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold211
timestamp 1679235063
transform 1 0 4600 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold212
timestamp 1679235063
transform 1 0 6808 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold213
timestamp 1679235063
transform 1 0 43700 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold214
timestamp 1679235063
transform 1 0 42228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold215
timestamp 1679235063
transform 1 0 15640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold216
timestamp 1679235063
transform 1 0 19688 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold217
timestamp 1679235063
transform 1 0 4600 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold218
timestamp 1679235063
transform 1 0 11960 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold219
timestamp 1679235063
transform 1 0 11868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold220
timestamp 1679235063
transform 1 0 10672 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold221
timestamp 1679235063
transform 1 0 43332 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold222
timestamp 1679235063
transform 1 0 44804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold223
timestamp 1679235063
transform 1 0 37444 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold224
timestamp 1679235063
transform 1 0 37444 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold225
timestamp 1679235063
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold226
timestamp 1679235063
transform 1 0 4232 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold227
timestamp 1679235063
transform 1 0 8004 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold228
timestamp 1679235063
transform 1 0 6808 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold229
timestamp 1679235063
transform 1 0 46276 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold230
timestamp 1679235063
transform 1 0 46276 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold231
timestamp 1679235063
transform 1 0 44804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold232
timestamp 1679235063
transform 1 0 46828 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold233
timestamp 1679235063
transform 1 0 4232 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold234
timestamp 1679235063
transform 1 0 4600 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold235
timestamp 1679235063
transform 1 0 45172 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold236
timestamp 1679235063
transform 1 0 43516 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold237
timestamp 1679235063
transform 1 0 45172 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold238
timestamp 1679235063
transform 1 0 45172 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold239
timestamp 1679235063
transform 1 0 10488 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold240
timestamp 1679235063
transform 1 0 33488 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold241
timestamp 1679235063
transform 1 0 4232 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold242
timestamp 1679235063
transform 1 0 5336 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold243
timestamp 1679235063
transform 1 0 42596 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold244
timestamp 1679235063
transform 1 0 42228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold245
timestamp 1679235063
transform 1 0 6624 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold246
timestamp 1679235063
transform 1 0 5704 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold247
timestamp 1679235063
transform 1 0 20792 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold248
timestamp 1679235063
transform 1 0 23552 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold249
timestamp 1679235063
transform 1 0 43332 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold250
timestamp 1679235063
transform 1 0 41124 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold251
timestamp 1679235063
transform 1 0 37444 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold252
timestamp 1679235063
transform 1 0 34868 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold253
timestamp 1679235063
transform 1 0 46276 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold254
timestamp 1679235063
transform 1 0 47380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold255
timestamp 1679235063
transform 1 0 28520 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold256
timestamp 1679235063
transform 1 0 25944 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold257
timestamp 1679235063
transform 1 0 10488 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold258
timestamp 1679235063
transform 1 0 9292 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold259
timestamp 1679235063
transform 1 0 19504 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold260
timestamp 1679235063
transform 1 0 18584 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold261
timestamp 1679235063
transform 1 0 45172 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold262
timestamp 1679235063
transform 1 0 46276 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold263
timestamp 1679235063
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold264
timestamp 1679235063
transform 1 0 1656 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold265
timestamp 1679235063
transform 1 0 6808 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold266
timestamp 1679235063
transform 1 0 6808 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold267
timestamp 1679235063
transform 1 0 20332 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold268
timestamp 1679235063
transform 1 0 21988 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold269
timestamp 1679235063
transform 1 0 20792 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold270
timestamp 1679235063
transform 1 0 24564 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold271
timestamp 1679235063
transform 1 0 42596 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold272
timestamp 1679235063
transform 1 0 45172 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold273
timestamp 1679235063
transform 1 0 47748 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold274
timestamp 1679235063
transform 1 0 45908 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold275
timestamp 1679235063
transform 1 0 33396 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold276
timestamp 1679235063
transform 1 0 32292 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold277
timestamp 1679235063
transform 1 0 29808 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold278
timestamp 1679235063
transform 1 0 28520 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold279
timestamp 1679235063
transform 1 0 40848 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold280
timestamp 1679235063
transform 1 0 38640 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold281
timestamp 1679235063
transform 1 0 47380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold282
timestamp 1679235063
transform 1 0 1656 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold283
timestamp 1679235063
transform 1 0 43424 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold284
timestamp 1679235063
transform 1 0 45908 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold285
timestamp 1679235063
transform 1 0 8280 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold286
timestamp 1679235063
transform 1 0 9384 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold287
timestamp 1679235063
transform 1 0 24840 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold288
timestamp 1679235063
transform 1 0 28336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold289
timestamp 1679235063
transform 1 0 10488 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold290
timestamp 1679235063
transform 1 0 6808 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold291
timestamp 1679235063
transform 1 0 6440 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold292
timestamp 1679235063
transform 1 0 4600 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold293
timestamp 1679235063
transform 1 0 29716 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold294
timestamp 1679235063
transform 1 0 29808 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold295
timestamp 1679235063
transform 1 0 7912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold296
timestamp 1679235063
transform 1 0 9752 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold297
timestamp 1679235063
transform 1 0 25024 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold298
timestamp 1679235063
transform 1 0 27048 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold299
timestamp 1679235063
transform 1 0 23828 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold300
timestamp 1679235063
transform 1 0 23368 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold301
timestamp 1679235063
transform 1 0 11868 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold302
timestamp 1679235063
transform 1 0 24840 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold303
timestamp 1679235063
transform 1 0 17480 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold304
timestamp 1679235063
transform 1 0 15180 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold305
timestamp 1679235063
transform 1 0 21988 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold306
timestamp 1679235063
transform 1 0 28336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold307
timestamp 1679235063
transform 1 0 7912 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold308
timestamp 1679235063
transform 1 0 12512 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold309
timestamp 1679235063
transform 1 0 41032 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold310
timestamp 1679235063
transform 1 0 39928 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold311
timestamp 1679235063
transform 1 0 5704 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold312
timestamp 1679235063
transform 1 0 4232 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold313
timestamp 1679235063
transform 1 0 9384 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold314
timestamp 1679235063
transform 1 0 29348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold315
timestamp 1679235063
transform 1 0 22264 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold316
timestamp 1679235063
transform 1 0 23368 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold317
timestamp 1679235063
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold318
timestamp 1679235063
transform 1 0 34868 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold319
timestamp 1679235063
transform 1 0 33580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold320
timestamp 1679235063
transform 1 0 5336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold321
timestamp 1679235063
transform 1 0 5336 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold322
timestamp 1679235063
transform 1 0 10028 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold323
timestamp 1679235063
transform 1 0 40020 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold324
timestamp 1679235063
transform 1 0 24932 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold325
timestamp 1679235063
transform 1 0 15272 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold326
timestamp 1679235063
transform 1 0 42596 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold327
timestamp 1679235063
transform 1 0 9292 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold328
timestamp 1679235063
transform 1 0 47380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold329
timestamp 1679235063
transform 1 0 10856 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold330
timestamp 1679235063
transform 1 0 44804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold331
timestamp 1679235063
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold332
timestamp 1679235063
transform 1 0 45908 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold333
timestamp 1679235063
transform 1 0 37444 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold334
timestamp 1679235063
transform 1 0 45724 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold335
timestamp 1679235063
transform 1 0 29716 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold336
timestamp 1679235063
transform 1 0 24840 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold337
timestamp 1679235063
transform 1 0 11868 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold338
timestamp 1679235063
transform 1 0 40756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold339
timestamp 1679235063
transform 1 0 42596 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold340
timestamp 1679235063
transform 1 0 14444 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold341
timestamp 1679235063
transform 1 0 32476 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold342
timestamp 1679235063
transform 1 0 46276 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold343
timestamp 1679235063
transform 1 0 14536 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold344
timestamp 1679235063
transform 1 0 37444 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold345
timestamp 1679235063
transform 1 0 46276 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold346
timestamp 1679235063
transform 1 0 36340 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold347
timestamp 1679235063
transform 1 0 43332 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold348
timestamp 1679235063
transform 1 0 13340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold349
timestamp 1679235063
transform 1 0 8188 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold350
timestamp 1679235063
transform 1 0 29716 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold351
timestamp 1679235063
transform 1 0 46552 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold352
timestamp 1679235063
transform 1 0 43700 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold353
timestamp 1679235063
transform 1 0 32292 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold354
timestamp 1679235063
transform 1 0 17020 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold355
timestamp 1679235063
transform 1 0 42596 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold356
timestamp 1679235063
transform 1 0 22724 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold357
timestamp 1679235063
transform 1 0 43332 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold358
timestamp 1679235063
transform 1 0 41124 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold359
timestamp 1679235063
transform 1 0 46276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold360
timestamp 1679235063
transform 1 0 7912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold361
timestamp 1679235063
transform 1 0 28612 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold362
timestamp 1679235063
transform 1 0 27784 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold363
timestamp 1679235063
transform 1 0 45080 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold364
timestamp 1679235063
transform 1 0 4232 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold365
timestamp 1679235063
transform 1 0 9384 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold366
timestamp 1679235063
transform 1 0 42596 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold367
timestamp 1679235063
transform 1 0 27324 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold368
timestamp 1679235063
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold369
timestamp 1679235063
transform 1 0 6808 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold370
timestamp 1679235063
transform 1 0 42228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold371
timestamp 1679235063
transform 1 0 30820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold372
timestamp 1679235063
transform 1 0 46184 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold373
timestamp 1679235063
transform 1 0 40020 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold374
timestamp 1679235063
transform 1 0 48484 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold375
timestamp 1679235063
transform 1 0 8280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold376
timestamp 1679235063
transform 1 0 8188 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold377
timestamp 1679235063
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold378
timestamp 1679235063
transform 1 0 27140 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold379
timestamp 1679235063
transform 1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold380
timestamp 1679235063
transform 1 0 48484 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold381
timestamp 1679235063
transform 1 0 48668 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold382
timestamp 1679235063
transform 1 0 48668 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold383
timestamp 1679235063
transform 1 0 48576 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold384
timestamp 1679235063
transform 1 0 48484 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold385
timestamp 1679235063
transform 1 0 47380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold386
timestamp 1679235063
transform 1 0 7912 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold387
timestamp 1679235063
transform 1 0 9108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold388
timestamp 1679235063
transform 1 0 10212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold389
timestamp 1679235063
transform 1 0 9384 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold390
timestamp 1679235063
transform 1 0 10488 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1679235063
transform 1 0 9384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1679235063
transform 1 0 47012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1679235063
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1679235063
transform 1 0 1564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1679235063
transform 1 0 1564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1679235063
transform 1 0 2300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1679235063
transform 1 0 1564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1679235063
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1679235063
transform 1 0 1564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1679235063
transform 1 0 1564 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1679235063
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1679235063
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1679235063
transform 1 0 1564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1679235063
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1679235063
transform 1 0 1564 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1679235063
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1679235063
transform 1 0 1564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1679235063
transform 1 0 1564 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1679235063
transform 1 0 3036 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1679235063
transform 1 0 4048 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1679235063
transform 1 0 1564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1679235063
transform 1 0 3404 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1679235063
transform 1 0 1564 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1679235063
transform 1 0 3128 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1679235063
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1679235063
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1679235063
transform 1 0 1564 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input28
timestamp 1679235063
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1679235063
transform 1 0 1564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1679235063
transform 1 0 1564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1679235063
transform 1 0 1564 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1679235063
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1679235063
transform 1 0 43332 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input34
timestamp 1679235063
transform 1 0 48852 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1679235063
transform 1 0 47748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1679235063
transform 1 0 45448 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1679235063
transform 1 0 48852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1679235063
transform 1 0 41768 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1679235063
transform 1 0 47196 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1679235063
transform 1 0 43516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1679235063
transform 1 0 46920 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1679235063
transform 1 0 47196 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1679235063
transform 1 0 46920 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1679235063
transform 1 0 49036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1679235063
transform 1 0 45356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1679235063
transform 1 0 47748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1679235063
transform 1 0 36616 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1679235063
transform 1 0 44160 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1679235063
transform 1 0 45540 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1679235063
transform 1 0 46000 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1679235063
transform 1 0 46920 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1679235063
transform 1 0 46368 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1679235063
transform 1 0 42688 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1679235063
transform 1 0 48484 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1679235063
transform 1 0 48852 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1679235063
transform 1 0 49036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1679235063
transform 1 0 47288 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1679235063
transform 1 0 49036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1679235063
transform 1 0 47840 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1679235063
transform 1 0 47748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1679235063
transform 1 0 46644 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1679235063
transform 1 0 35236 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1679235063
transform 1 0 11684 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1679235063
transform 1 0 47748 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1679235063
transform 1 0 45172 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1679235063
transform 1 0 39652 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1679235063
transform 1 0 40756 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1679235063
transform 1 0 42044 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1679235063
transform 1 0 42596 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input70
timestamp 1679235063
transform 1 0 42596 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1679235063
transform 1 0 42596 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input72
timestamp 1679235063
transform 1 0 45172 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1679235063
transform 1 0 43884 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1679235063
transform 1 0 21252 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1679235063
transform 1 0 45816 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1679235063
transform 1 0 45172 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1679235063
transform 1 0 47748 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input78
timestamp 1679235063
transform 1 0 45632 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input79
timestamp 1679235063
transform 1 0 46460 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input80
timestamp 1679235063
transform 1 0 45540 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input81
timestamp 1679235063
transform 1 0 43608 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input82
timestamp 1679235063
transform 1 0 43240 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input83
timestamp 1679235063
transform 1 0 44528 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input84
timestamp 1679235063
transform 1 0 45632 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1679235063
transform 1 0 9016 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1679235063
transform 1 0 23644 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1679235063
transform 1 0 13432 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input88
timestamp 1679235063
transform 1 0 41216 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input89
timestamp 1679235063
transform 1 0 47748 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1679235063
transform 1 0 6716 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input91
timestamp 1679235063
transform 1 0 11684 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input92
timestamp 1679235063
transform 1 0 44988 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1679235063
transform 1 0 28704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1679235063
transform 1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1679235063
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1679235063
transform 1 0 35052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input97
timestamp 1679235063
transform 1 0 37444 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1679235063
transform 1 0 44160 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input99
timestamp 1679235063
transform 1 0 44896 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input100
timestamp 1679235063
transform 1 0 45356 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input101
timestamp 1679235063
transform 1 0 46736 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input102
timestamp 1679235063
transform 1 0 46184 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1679235063
transform 1 0 46184 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input104
timestamp 1679235063
transform 1 0 43424 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input105
timestamp 1679235063
transform 1 0 24104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1679235063
transform 1 0 37536 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output107 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 40664 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1679235063
transform 1 0 3404 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1679235063
transform 1 0 1564 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1679235063
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1679235063
transform 1 0 1564 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1679235063
transform 1 0 1564 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1679235063
transform 1 0 1564 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1679235063
transform 1 0 1564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1679235063
transform 1 0 1564 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1679235063
transform 1 0 3404 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1679235063
transform 1 0 1564 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1679235063
transform 1 0 1564 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1679235063
transform 1 0 1564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1679235063
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1679235063
transform 1 0 3956 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1679235063
transform 1 0 3956 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1679235063
transform 1 0 5796 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1679235063
transform 1 0 5796 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1679235063
transform 1 0 6532 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1679235063
transform 1 0 3956 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1679235063
transform 1 0 5796 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1679235063
transform 1 0 6532 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1679235063
transform 1 0 8372 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1679235063
transform 1 0 9108 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1679235063
transform 1 0 1564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1679235063
transform 1 0 1564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1679235063
transform 1 0 1564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1679235063
transform 1 0 1564 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1679235063
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1679235063
transform 1 0 1564 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1679235063
transform 1 0 1564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1679235063
transform 1 0 1564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1679235063
transform 1 0 45816 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1679235063
transform 1 0 47932 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1679235063
transform 1 0 47932 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1679235063
transform 1 0 46092 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1679235063
transform 1 0 47932 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1679235063
transform 1 0 47932 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1679235063
transform 1 0 47932 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1679235063
transform 1 0 45816 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1679235063
transform 1 0 47932 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1679235063
transform 1 0 47932 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1679235063
transform 1 0 47932 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1679235063
transform 1 0 43976 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1679235063
transform 1 0 46092 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1679235063
transform 1 0 47932 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1679235063
transform 1 0 47932 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1679235063
transform 1 0 47932 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1679235063
transform 1 0 47932 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1679235063
transform 1 0 47932 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1679235063
transform 1 0 47932 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1679235063
transform 1 0 47932 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1679235063
transform 1 0 47932 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1679235063
transform 1 0 47932 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1679235063
transform 1 0 45816 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1679235063
transform 1 0 45816 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1679235063
transform 1 0 46092 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1679235063
transform 1 0 47932 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1679235063
transform 1 0 47932 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1679235063
transform 1 0 47932 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1679235063
transform 1 0 45816 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1679235063
transform 1 0 47932 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1679235063
transform 1 0 3956 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1679235063
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1679235063
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1679235063
transform 1 0 9752 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1679235063
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1679235063
transform 1 0 10488 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1679235063
transform 1 0 11960 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1679235063
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1679235063
transform 1 0 12328 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1679235063
transform 1 0 13064 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1679235063
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1679235063
transform 1 0 3404 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1679235063
transform 1 0 13064 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1679235063
transform 1 0 14904 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1679235063
transform 1 0 15272 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1679235063
transform 1 0 14904 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1679235063
transform 1 0 17480 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1679235063
transform 1 0 14904 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1679235063
transform 1 0 17756 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1679235063
transform 1 0 17480 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1679235063
transform 1 0 21988 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1679235063
transform 1 0 21988 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1679235063
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1679235063
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1679235063
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1679235063
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1679235063
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1679235063
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1679235063
transform 1 0 7452 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1679235063
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1679235063
transform 1 0 11776 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1679235063
transform 1 0 14260 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1679235063
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output202
timestamp 1679235063
transform 1 0 17480 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1679235063
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1679235063
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1679235063
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1679235063
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1679235063
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1679235063
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1679235063
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1679235063
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1679235063
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1679235063
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1679235063
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1679235063
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1679235063
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1679235063
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1679235063
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1679235063
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1679235063
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1679235063
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1679235063
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1679235063
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1679235063
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1679235063
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1679235063
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1679235063
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1679235063
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1679235063
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1679235063
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1679235063
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1679235063
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1679235063
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1679235063
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1679235063
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1679235063
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1679235063
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1679235063
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1679235063
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1679235063
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1679235063
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1679235063
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1679235063
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1679235063
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1679235063
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1679235063
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1679235063
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1679235063
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1679235063
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1679235063
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1679235063
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1679235063
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1679235063
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1679235063
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1679235063
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1679235063
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1679235063
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1679235063
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1679235063
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1679235063
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1679235063
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1679235063
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1679235063
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1679235063
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1679235063
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1679235063
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1679235063
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1679235063
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1679235063
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1679235063
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1679235063
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1679235063
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1679235063
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1679235063
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1679235063
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1679235063
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1679235063
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1679235063
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1679235063
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1679235063
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1679235063
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1679235063
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1679235063
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1679235063
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1679235063
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 26864 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24932 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 23092 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22816 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20700 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 17112 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17020 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20240 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 17112 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19136 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20884 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 19688 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20792 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20976 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 19320 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19596 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19596 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 17848 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19228 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19596 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 19412 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20792 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24288 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 23184 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24932 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 27140 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 25392 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 27140 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 28060 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 24840 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24840 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 25392 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 21068 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 28244 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 30084 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 31280 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 32568 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 34868 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 34960 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 34868 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 36432 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 37444 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 34868 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 37444 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 35972 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 33764 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 34868 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 33488 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 30636 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 32292 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 30728 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 29348 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 28336 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 28336 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 26772 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 28428 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 29900 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 30820 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 32292 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 31924 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 29716 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 27876 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 26864 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 41676 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 30820 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 29900 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 32108 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 33580 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 33304 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 34868 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 34868 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 32292 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 33764 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 37444 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 37076 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 37444 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 38272 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 37720 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 37996 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 36432 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 34408 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 36248 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 38548 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 38548 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 40020 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 40020 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 38272 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 38548 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 40020 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 37996 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 37444 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 37076 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 33120 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 29716 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 25944 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24840 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24564 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24012 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24564 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24564 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24196 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23460 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22172 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19964 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18952 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19320 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21620 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17664 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14536 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14260 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14260 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12604 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11132 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10580 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11960 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13616 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14444 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14996 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30912 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 27508 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_2_
timestamp 1679235063
transform 1 0 22816 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_1.mux_l1_in_3__263
timestamp 1679235063
transform 1 0 26220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_3_
timestamp 1679235063
transform 1 0 22080 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 25484 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l2_in_1_
timestamp 1679235063
transform 1 0 24104 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 22448 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16008 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24748 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 23368 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_3.mux_l2_in_1__216
timestamp 1679235063
transform 1 0 9108 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l2_in_1_
timestamp 1679235063
transform 1 0 17848 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 17848 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25760 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24564 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_5.mux_l2_in_1__219
timestamp 1679235063
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l2_in_1_
timestamp 1679235063
transform 1 0 18124 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l3_in_0_
timestamp 1679235063
transform 1 0 17296 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_0_
timestamp 1679235063
transform 1 0 26680 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24380 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_2_
timestamp 1679235063
transform 1 0 19596 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22908 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l2_in_1_
timestamp 1679235063
transform 1 0 19688 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_7.mux_l2_in_1__221
timestamp 1679235063
transform 1 0 21160 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19596 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16468 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27416 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_1_
timestamp 1679235063
transform 1 0 25484 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_2_
timestamp 1679235063
transform 1 0 20700 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_11.mux_l1_in_3__264
timestamp 1679235063
transform 1 0 17020 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_3_
timestamp 1679235063
transform 1 0 20424 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23092 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l2_in_1_
timestamp 1679235063
transform 1 0 20240 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6532 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27140 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_1_
timestamp 1679235063
transform 1 0 23276 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_2_
timestamp 1679235063
transform 1 0 20884 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20792 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_13.mux_l2_in_1__265
timestamp 1679235063
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l2_in_1_
timestamp 1679235063
transform 1 0 19504 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l3_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 12420 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27600 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_1_
timestamp 1679235063
transform 1 0 23276 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_2_
timestamp 1679235063
transform 1 0 21988 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22448 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l2_in_1_
timestamp 1679235063
transform 1 0 20056 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_21.mux_l2_in_1__266
timestamp 1679235063
transform 1 0 3956 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l3_in_0_
timestamp 1679235063
transform 1 0 16928 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_0_
timestamp 1679235063
transform 1 0 29716 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_1_
timestamp 1679235063
transform 1 0 27140 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_2_
timestamp 1679235063
transform 1 0 23184 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l2_in_0_
timestamp 1679235063
transform 1 0 25852 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l2_in_1_
timestamp 1679235063
transform 1 0 23184 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_29.mux_l2_in_1__267
timestamp 1679235063
transform 1 0 30084 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l3_in_0_
timestamp 1679235063
transform 1 0 20148 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6532 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l1_in_0_
timestamp 1679235063
transform 1 0 32292 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l1_in_1_
timestamp 1679235063
transform 1 0 28888 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l2_in_0_
timestamp 1679235063
transform 1 0 27876 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_37.mux_l2_in_1__217
timestamp 1679235063
transform 1 0 22264 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l2_in_1_
timestamp 1679235063
transform 1 0 23276 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l3_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17112 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l1_in_0_
timestamp 1679235063
transform 1 0 32292 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l2_in_0_
timestamp 1679235063
transform 1 0 27876 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l2_in_1_
timestamp 1679235063
transform 1 0 27600 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_45.mux_l2_in_1__218
timestamp 1679235063
transform 1 0 37076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l3_in_0_
timestamp 1679235063
transform 1 0 23644 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30268 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l2_in_0_
timestamp 1679235063
transform 1 0 25944 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l2_in_1_
timestamp 1679235063
transform 1 0 21988 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_53.mux_l2_in_1__220
timestamp 1679235063
transform 1 0 24564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19504 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 29716 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 33120 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 27140 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 32292 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_0.mux_l2_in_1__222
timestamp 1679235063
transform 1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 29532 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 33488 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 41860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 33304 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 33580 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 28428 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 33764 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 33488 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_2.mux_l2_in_1__225
timestamp 1679235063
transform 1 0 34132 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 35972 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 44436 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 34868 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 32660 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_2_
timestamp 1679235063
transform 1 0 32844 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 34776 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l2_in_1_
timestamp 1679235063
transform 1 0 35788 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_4.mux_l2_in_1__229
timestamp 1679235063
transform 1 0 39284 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l3_in_0_
timestamp 1679235063
transform 1 0 38640 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 42964 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 36064 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 33488 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_2_
timestamp 1679235063
transform 1 0 35972 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_3_
timestamp 1679235063
transform 1 0 34868 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_6.mux_l1_in_3__232
timestamp 1679235063
transform 1 0 33396 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 34868 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 37444 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 38272 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 43332 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 34868 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 32936 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_2_
timestamp 1679235063
transform 1 0 37444 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_3_
timestamp 1679235063
transform 1 0 31004 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_10.mux_l1_in_3__223
timestamp 1679235063
transform 1 0 31648 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 35236 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l2_in_1_
timestamp 1679235063
transform 1 0 34868 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l3_in_0_
timestamp 1679235063
transform 1 0 35972 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 43976 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 32936 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_1_
timestamp 1679235063
transform 1 0 30820 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_2_
timestamp 1679235063
transform 1 0 27140 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 31740 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_12.mux_l2_in_1__224
timestamp 1679235063
transform 1 0 31556 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l2_in_1_
timestamp 1679235063
transform 1 0 32568 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l3_in_0_
timestamp 1679235063
transform 1 0 37444 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 44436 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 29900 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_1_
timestamp 1679235063
transform 1 0 29716 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_2_
timestamp 1679235063
transform 1 0 26772 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 29716 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l2_in_1_
timestamp 1679235063
transform 1 0 28428 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_20.mux_l2_in_1__226
timestamp 1679235063
transform 1 0 30084 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l3_in_0_
timestamp 1679235063
transform 1 0 32568 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 42596 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 29716 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_1_
timestamp 1679235063
transform 1 0 29532 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_2_
timestamp 1679235063
transform 1 0 25852 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 31924 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_28.mux_l2_in_1__227
timestamp 1679235063
transform 1 0 27232 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l2_in_1_
timestamp 1679235063
transform 1 0 28244 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l3_in_0_
timestamp 1679235063
transform 1 0 34500 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 39100 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30544 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l1_in_1_
timestamp 1679235063
transform 1 0 30820 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l2_in_0_
timestamp 1679235063
transform 1 0 33028 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l2_in_1_
timestamp 1679235063
transform 1 0 31004 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_36.mux_l2_in_1__228
timestamp 1679235063
transform 1 0 32292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l3_in_0_
timestamp 1679235063
transform 1 0 33580 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 39744 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30452 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l1_in_1_
timestamp 1679235063
transform 1 0 29716 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_44.mux_l1_in_1__230
timestamp 1679235063
transform 1 0 34132 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 31188 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 37168 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l1_in_0_
timestamp 1679235063
transform 1 0 28428 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l1_in_1_
timestamp 1679235063
transform 1 0 27232 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_52.mux_l1_in_1__231
timestamp 1679235063
transform 1 0 28980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l2_in_0_
timestamp 1679235063
transform 1 0 32292 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 38548 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 33120 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 40020 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 24656 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_0.mux_l1_in_3__233
timestamp 1679235063
transform 1 0 34132 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 29716 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 36064 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 28520 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 30268 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 37536 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 34868 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 40020 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 30912 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 38640 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 34868 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_2.mux_l2_in_1__239
timestamp 1679235063
transform 1 0 47012 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 32292 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 44436 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 36064 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 40020 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 36064 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l2_in_1_
timestamp 1679235063
transform 1 0 30912 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_4.mux_l2_in_1__249
timestamp 1679235063
transform 1 0 32292 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l3_in_0_
timestamp 1679235063
transform 1 0 32108 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 38548 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 40848 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_2_
timestamp 1679235063
transform 1 0 32568 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 39652 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 35972 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_6.mux_l2_in_1__257
timestamp 1679235063
transform 1 0 43424 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 37444 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 30912 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1679235063
transform 1 0 40020 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_1_
timestamp 1679235063
transform 1 0 41216 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_2_
timestamp 1679235063
transform 1 0 34868 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 40480 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l2_in_1_
timestamp 1679235063
transform 1 0 36156 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_8.mux_l2_in_1__258
timestamp 1679235063
transform 1 0 47012 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l3_in_0_
timestamp 1679235063
transform 1 0 37352 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 47012 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 36064 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 40204 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 38732 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l2_in_1_
timestamp 1679235063
transform 1 0 32292 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_10.mux_l2_in_1__234
timestamp 1679235063
transform 1 0 31096 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l3_in_0_
timestamp 1679235063
transform 1 0 32752 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 40020 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 40020 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 40848 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_12.mux_l2_in_1__235
timestamp 1679235063
transform 1 0 44436 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l2_in_1_
timestamp 1679235063
transform 1 0 37076 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l3_in_0_
timestamp 1679235063
transform 1 0 38456 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 39284 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 40756 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 40848 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l2_in_1_
timestamp 1679235063
transform 1 0 35144 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_14.mux_l2_in_1__236
timestamp 1679235063
transform 1 0 44436 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l3_in_0_
timestamp 1679235063
transform 1 0 38640 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 35328 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1679235063
transform 1 0 40020 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 40756 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_16.mux_l2_in_1__237
timestamp 1679235063
transform 1 0 44436 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l2_in_1_
timestamp 1679235063
transform 1 0 37076 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l3_in_0_
timestamp 1679235063
transform 1 0 36064 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 39284 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 38272 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 40204 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_18.mux_l2_in_1__238
timestamp 1679235063
transform 1 0 34500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l2_in_1_
timestamp 1679235063
transform 1 0 32384 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l3_in_0_
timestamp 1679235063
transform 1 0 32292 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 27600 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27508 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l1_in_1_
timestamp 1679235063
transform 1 0 25392 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_20.mux_l1_in_1__240
timestamp 1679235063
transform 1 0 29716 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 25300 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25576 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_22.mux_l1_in_1__241
timestamp 1679235063
transform 1 0 22172 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l1_in_1_
timestamp 1679235063
transform 1 0 25392 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27140 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24196 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_24.mux_l1_in_1__242
timestamp 1679235063
transform 1 0 20056 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14536 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27048 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_26.mux_l1_in_1__243
timestamp 1679235063
transform 1 0 23828 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l1_in_1_
timestamp 1679235063
transform 1 0 24564 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22908 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_28.mux_l2_in_0__244
timestamp 1679235063
transform 1 0 19412 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6532 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18124 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_30.mux_l2_in_0__245
timestamp 1679235063
transform 1 0 19412 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3956 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16928 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16928 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_32.mux_l2_in_0__246
timestamp 1679235063
transform 1 0 14352 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14260 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19320 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_34.mux_l2_in_0__247
timestamp 1679235063
transform 1 0 18492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l1_in_0_
timestamp 1679235063
transform 1 0 28336 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_36.mux_l1_in_1__248
timestamp 1679235063
transform 1 0 23276 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l1_in_1_
timestamp 1679235063
transform 1 0 21712 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_40.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14352 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_40.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13064 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_40.mux_l2_in_0__250
timestamp 1679235063
transform 1 0 13524 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8096 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_42.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16744 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_42.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14812 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_42.mux_l2_in_0__251
timestamp 1679235063
transform 1 0 3956 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12420 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_44.mux_l2_in_0__252
timestamp 1679235063
transform 1 0 8740 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9752 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12328 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_46.mux_l2_in_0__253
timestamp 1679235063
transform 1 0 2852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_48.mux_l2_in_0__254
timestamp 1679235063
transform 1 0 10396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14352 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_50.mux_l2_in_0__255
timestamp 1679235063
transform 1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3496 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_58.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19596 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_58.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_58.mux_l2_in_0__256
timestamp 1679235063
transform 1 0 12328 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 2760 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1679235063
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1679235063
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1679235063
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1679235063
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1679235063
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1679235063
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1679235063
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1679235063
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1679235063
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1679235063
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1679235063
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1679235063
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1679235063
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1679235063
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1679235063
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1679235063
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1679235063
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1679235063
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1679235063
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1679235063
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1679235063
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1679235063
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1679235063
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1679235063
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1679235063
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1679235063
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1679235063
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1679235063
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1679235063
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1679235063
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1679235063
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1679235063
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1679235063
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1679235063
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1679235063
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1679235063
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1679235063
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1679235063
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1679235063
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1679235063
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1679235063
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1679235063
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1679235063
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1679235063
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1679235063
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1679235063
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1679235063
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1679235063
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1679235063
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1679235063
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1679235063
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1679235063
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1679235063
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1679235063
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1679235063
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1679235063
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1679235063
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1679235063
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1679235063
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1679235063
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1679235063
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1679235063
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1679235063
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1679235063
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1679235063
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1679235063
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1679235063
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1679235063
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1679235063
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1679235063
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1679235063
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1679235063
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1679235063
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1679235063
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1679235063
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1679235063
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1679235063
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1679235063
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1679235063
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1679235063
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1679235063
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1679235063
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1679235063
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1679235063
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1679235063
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1679235063
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1679235063
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1679235063
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1679235063
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1679235063
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1679235063
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1679235063
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1679235063
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1679235063
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1679235063
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1679235063
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1679235063
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1679235063
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1679235063
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1679235063
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1679235063
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1679235063
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1679235063
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1679235063
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1679235063
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1679235063
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1679235063
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1679235063
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1679235063
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1679235063
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1679235063
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1679235063
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1679235063
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1679235063
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1679235063
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1679235063
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1679235063
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1679235063
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1679235063
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1679235063
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1679235063
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1679235063
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1679235063
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1679235063
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1679235063
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1679235063
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1679235063
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1679235063
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1679235063
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1679235063
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1679235063
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1679235063
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1679235063
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1679235063
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1679235063
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1679235063
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1679235063
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1679235063
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1679235063
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1679235063
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1679235063
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1679235063
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1679235063
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1679235063
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1679235063
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1679235063
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1679235063
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1679235063
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1679235063
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1679235063
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1679235063
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1679235063
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1679235063
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1679235063
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1679235063
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1679235063
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1679235063
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1679235063
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1679235063
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1679235063
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1679235063
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1679235063
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1679235063
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1679235063
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1679235063
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1679235063
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1679235063
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1679235063
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1679235063
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1679235063
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1679235063
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1679235063
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1679235063
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1679235063
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1679235063
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1679235063
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1679235063
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1679235063
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1679235063
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1679235063
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1679235063
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1679235063
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1679235063
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1679235063
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1679235063
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1679235063
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1679235063
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1679235063
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1679235063
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1679235063
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1679235063
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1679235063
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1679235063
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1679235063
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1679235063
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1679235063
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1679235063
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1679235063
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1679235063
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1679235063
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1679235063
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1679235063
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1679235063
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1679235063
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1679235063
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1679235063
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1679235063
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1679235063
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1679235063
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1679235063
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1679235063
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1679235063
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1679235063
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1679235063
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1679235063
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1679235063
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1679235063
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1679235063
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1679235063
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1679235063
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1679235063
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1679235063
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1679235063
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1679235063
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1679235063
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1679235063
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1679235063
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1679235063
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1679235063
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1679235063
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1679235063
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1679235063
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1679235063
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1679235063
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1679235063
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1679235063
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1679235063
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1679235063
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1679235063
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1679235063
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1679235063
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1679235063
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1679235063
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1679235063
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1679235063
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1679235063
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1679235063
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1679235063
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1679235063
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1679235063
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1679235063
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1679235063
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1679235063
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1679235063
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1679235063
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1679235063
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1679235063
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1679235063
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1679235063
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1679235063
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1679235063
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1679235063
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1679235063
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1679235063
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1679235063
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1679235063
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1679235063
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1679235063
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1679235063
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1679235063
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1679235063
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1679235063
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1679235063
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1679235063
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1679235063
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1679235063
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1679235063
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1679235063
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1679235063
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1679235063
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1679235063
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1679235063
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1679235063
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1679235063
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1679235063
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1679235063
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1679235063
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1679235063
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1679235063
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1679235063
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1679235063
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1679235063
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1679235063
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1679235063
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1679235063
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1679235063
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1679235063
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1679235063
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1679235063
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1679235063
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1679235063
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1679235063
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1679235063
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1679235063
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1679235063
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1679235063
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1679235063
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1679235063
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1679235063
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1679235063
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1679235063
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1679235063
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1679235063
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1679235063
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1679235063
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1679235063
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1679235063
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1679235063
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1679235063
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1679235063
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1679235063
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1679235063
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1679235063
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1679235063
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1679235063
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1679235063
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1679235063
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1679235063
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1679235063
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1679235063
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1679235063
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1679235063
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1679235063
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1679235063
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1679235063
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1679235063
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1679235063
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1679235063
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1679235063
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1679235063
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1679235063
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1679235063
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1679235063
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1679235063
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1679235063
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1679235063
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1679235063
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1679235063
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1679235063
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1679235063
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1679235063
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1679235063
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1679235063
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1679235063
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1679235063
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1679235063
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1679235063
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1679235063
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1679235063
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1679235063
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1679235063
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1679235063
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1679235063
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1679235063
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1679235063
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1679235063
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1679235063
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1679235063
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1679235063
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1679235063
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1679235063
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1679235063
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1679235063
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1679235063
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1679235063
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1679235063
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1679235063
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1679235063
transform 1 0 26864 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1679235063
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1679235063
transform 1 0 32016 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1679235063
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1679235063
transform 1 0 37168 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1679235063
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1679235063
transform 1 0 42320 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1679235063
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1679235063
transform 1 0 47472 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 49238 26200 49294 27000 0 FreeSans 224 90 0 0 ccff_head_1
port 3 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1582 26200 1638 27000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[20]
port 18 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[21]
port 19 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[22]
port 20 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[23]
port 21 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[24]
port 22 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[25]
port 23 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[26]
port 24 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[27]
port 25 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[28]
port 26 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[29]
port 27 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 28 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 29 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 30 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 31 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 32 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 33 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 34 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 35 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 36 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 37 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 38 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 39 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 40 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 41 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 42 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 43 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 44 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 45 nsew signal tristate
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 46 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 47 nsew signal tristate
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 chanx_left_out[20]
port 48 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 chanx_left_out[21]
port 49 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 chanx_left_out[22]
port 50 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_out[23]
port 51 nsew signal tristate
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 chanx_left_out[24]
port 52 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 chanx_left_out[25]
port 53 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 chanx_left_out[26]
port 54 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 chanx_left_out[27]
port 55 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_out[28]
port 56 nsew signal tristate
flabel metal3 s 0 25576 800 25696 0 FreeSans 480 0 0 0 chanx_left_out[29]
port 57 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal3 s 50200 13608 51000 13728 0 FreeSans 480 0 0 0 chanx_right_in_0[0]
port 66 nsew signal input
flabel metal3 s 50200 17688 51000 17808 0 FreeSans 480 0 0 0 chanx_right_in_0[10]
port 67 nsew signal input
flabel metal3 s 50200 18096 51000 18216 0 FreeSans 480 0 0 0 chanx_right_in_0[11]
port 68 nsew signal input
flabel metal3 s 50200 18504 51000 18624 0 FreeSans 480 0 0 0 chanx_right_in_0[12]
port 69 nsew signal input
flabel metal3 s 50200 18912 51000 19032 0 FreeSans 480 0 0 0 chanx_right_in_0[13]
port 70 nsew signal input
flabel metal3 s 50200 19320 51000 19440 0 FreeSans 480 0 0 0 chanx_right_in_0[14]
port 71 nsew signal input
flabel metal3 s 50200 19728 51000 19848 0 FreeSans 480 0 0 0 chanx_right_in_0[15]
port 72 nsew signal input
flabel metal3 s 50200 20136 51000 20256 0 FreeSans 480 0 0 0 chanx_right_in_0[16]
port 73 nsew signal input
flabel metal3 s 50200 20544 51000 20664 0 FreeSans 480 0 0 0 chanx_right_in_0[17]
port 74 nsew signal input
flabel metal3 s 50200 20952 51000 21072 0 FreeSans 480 0 0 0 chanx_right_in_0[18]
port 75 nsew signal input
flabel metal3 s 50200 21360 51000 21480 0 FreeSans 480 0 0 0 chanx_right_in_0[19]
port 76 nsew signal input
flabel metal3 s 50200 14016 51000 14136 0 FreeSans 480 0 0 0 chanx_right_in_0[1]
port 77 nsew signal input
flabel metal3 s 50200 21768 51000 21888 0 FreeSans 480 0 0 0 chanx_right_in_0[20]
port 78 nsew signal input
flabel metal3 s 50200 22176 51000 22296 0 FreeSans 480 0 0 0 chanx_right_in_0[21]
port 79 nsew signal input
flabel metal3 s 50200 22584 51000 22704 0 FreeSans 480 0 0 0 chanx_right_in_0[22]
port 80 nsew signal input
flabel metal3 s 50200 22992 51000 23112 0 FreeSans 480 0 0 0 chanx_right_in_0[23]
port 81 nsew signal input
flabel metal3 s 50200 23400 51000 23520 0 FreeSans 480 0 0 0 chanx_right_in_0[24]
port 82 nsew signal input
flabel metal3 s 50200 23808 51000 23928 0 FreeSans 480 0 0 0 chanx_right_in_0[25]
port 83 nsew signal input
flabel metal3 s 50200 24216 51000 24336 0 FreeSans 480 0 0 0 chanx_right_in_0[26]
port 84 nsew signal input
flabel metal3 s 50200 24624 51000 24744 0 FreeSans 480 0 0 0 chanx_right_in_0[27]
port 85 nsew signal input
flabel metal3 s 50200 25032 51000 25152 0 FreeSans 480 0 0 0 chanx_right_in_0[28]
port 86 nsew signal input
flabel metal3 s 50200 25440 51000 25560 0 FreeSans 480 0 0 0 chanx_right_in_0[29]
port 87 nsew signal input
flabel metal3 s 50200 14424 51000 14544 0 FreeSans 480 0 0 0 chanx_right_in_0[2]
port 88 nsew signal input
flabel metal3 s 50200 14832 51000 14952 0 FreeSans 480 0 0 0 chanx_right_in_0[3]
port 89 nsew signal input
flabel metal3 s 50200 15240 51000 15360 0 FreeSans 480 0 0 0 chanx_right_in_0[4]
port 90 nsew signal input
flabel metal3 s 50200 15648 51000 15768 0 FreeSans 480 0 0 0 chanx_right_in_0[5]
port 91 nsew signal input
flabel metal3 s 50200 16056 51000 16176 0 FreeSans 480 0 0 0 chanx_right_in_0[6]
port 92 nsew signal input
flabel metal3 s 50200 16464 51000 16584 0 FreeSans 480 0 0 0 chanx_right_in_0[7]
port 93 nsew signal input
flabel metal3 s 50200 16872 51000 16992 0 FreeSans 480 0 0 0 chanx_right_in_0[8]
port 94 nsew signal input
flabel metal3 s 50200 17280 51000 17400 0 FreeSans 480 0 0 0 chanx_right_in_0[9]
port 95 nsew signal input
flabel metal3 s 50200 1368 51000 1488 0 FreeSans 480 0 0 0 chanx_right_out_0[0]
port 96 nsew signal tristate
flabel metal3 s 50200 5448 51000 5568 0 FreeSans 480 0 0 0 chanx_right_out_0[10]
port 97 nsew signal tristate
flabel metal3 s 50200 5856 51000 5976 0 FreeSans 480 0 0 0 chanx_right_out_0[11]
port 98 nsew signal tristate
flabel metal3 s 50200 6264 51000 6384 0 FreeSans 480 0 0 0 chanx_right_out_0[12]
port 99 nsew signal tristate
flabel metal3 s 50200 6672 51000 6792 0 FreeSans 480 0 0 0 chanx_right_out_0[13]
port 100 nsew signal tristate
flabel metal3 s 50200 7080 51000 7200 0 FreeSans 480 0 0 0 chanx_right_out_0[14]
port 101 nsew signal tristate
flabel metal3 s 50200 7488 51000 7608 0 FreeSans 480 0 0 0 chanx_right_out_0[15]
port 102 nsew signal tristate
flabel metal3 s 50200 7896 51000 8016 0 FreeSans 480 0 0 0 chanx_right_out_0[16]
port 103 nsew signal tristate
flabel metal3 s 50200 8304 51000 8424 0 FreeSans 480 0 0 0 chanx_right_out_0[17]
port 104 nsew signal tristate
flabel metal3 s 50200 8712 51000 8832 0 FreeSans 480 0 0 0 chanx_right_out_0[18]
port 105 nsew signal tristate
flabel metal3 s 50200 9120 51000 9240 0 FreeSans 480 0 0 0 chanx_right_out_0[19]
port 106 nsew signal tristate
flabel metal3 s 50200 1776 51000 1896 0 FreeSans 480 0 0 0 chanx_right_out_0[1]
port 107 nsew signal tristate
flabel metal3 s 50200 9528 51000 9648 0 FreeSans 480 0 0 0 chanx_right_out_0[20]
port 108 nsew signal tristate
flabel metal3 s 50200 9936 51000 10056 0 FreeSans 480 0 0 0 chanx_right_out_0[21]
port 109 nsew signal tristate
flabel metal3 s 50200 10344 51000 10464 0 FreeSans 480 0 0 0 chanx_right_out_0[22]
port 110 nsew signal tristate
flabel metal3 s 50200 10752 51000 10872 0 FreeSans 480 0 0 0 chanx_right_out_0[23]
port 111 nsew signal tristate
flabel metal3 s 50200 11160 51000 11280 0 FreeSans 480 0 0 0 chanx_right_out_0[24]
port 112 nsew signal tristate
flabel metal3 s 50200 11568 51000 11688 0 FreeSans 480 0 0 0 chanx_right_out_0[25]
port 113 nsew signal tristate
flabel metal3 s 50200 11976 51000 12096 0 FreeSans 480 0 0 0 chanx_right_out_0[26]
port 114 nsew signal tristate
flabel metal3 s 50200 12384 51000 12504 0 FreeSans 480 0 0 0 chanx_right_out_0[27]
port 115 nsew signal tristate
flabel metal3 s 50200 12792 51000 12912 0 FreeSans 480 0 0 0 chanx_right_out_0[28]
port 116 nsew signal tristate
flabel metal3 s 50200 13200 51000 13320 0 FreeSans 480 0 0 0 chanx_right_out_0[29]
port 117 nsew signal tristate
flabel metal3 s 50200 2184 51000 2304 0 FreeSans 480 0 0 0 chanx_right_out_0[2]
port 118 nsew signal tristate
flabel metal3 s 50200 2592 51000 2712 0 FreeSans 480 0 0 0 chanx_right_out_0[3]
port 119 nsew signal tristate
flabel metal3 s 50200 3000 51000 3120 0 FreeSans 480 0 0 0 chanx_right_out_0[4]
port 120 nsew signal tristate
flabel metal3 s 50200 3408 51000 3528 0 FreeSans 480 0 0 0 chanx_right_out_0[5]
port 121 nsew signal tristate
flabel metal3 s 50200 3816 51000 3936 0 FreeSans 480 0 0 0 chanx_right_out_0[6]
port 122 nsew signal tristate
flabel metal3 s 50200 4224 51000 4344 0 FreeSans 480 0 0 0 chanx_right_out_0[7]
port 123 nsew signal tristate
flabel metal3 s 50200 4632 51000 4752 0 FreeSans 480 0 0 0 chanx_right_out_0[8]
port 124 nsew signal tristate
flabel metal3 s 50200 5040 51000 5160 0 FreeSans 480 0 0 0 chanx_right_out_0[9]
port 125 nsew signal tristate
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 126 nsew signal input
flabel metal2 s 27986 26200 28042 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 127 nsew signal input
flabel metal2 s 28630 26200 28686 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 128 nsew signal input
flabel metal2 s 29274 26200 29330 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 129 nsew signal input
flabel metal2 s 29918 26200 29974 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 130 nsew signal input
flabel metal2 s 30562 26200 30618 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 131 nsew signal input
flabel metal2 s 31206 26200 31262 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 132 nsew signal input
flabel metal2 s 31850 26200 31906 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 133 nsew signal input
flabel metal2 s 32494 26200 32550 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 134 nsew signal input
flabel metal2 s 33138 26200 33194 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 135 nsew signal input
flabel metal2 s 33782 26200 33838 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 136 nsew signal input
flabel metal2 s 22190 26200 22246 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 137 nsew signal input
flabel metal2 s 34426 26200 34482 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 138 nsew signal input
flabel metal2 s 35070 26200 35126 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 139 nsew signal input
flabel metal2 s 35714 26200 35770 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 140 nsew signal input
flabel metal2 s 36358 26200 36414 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 141 nsew signal input
flabel metal2 s 37002 26200 37058 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 142 nsew signal input
flabel metal2 s 37646 26200 37702 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 143 nsew signal input
flabel metal2 s 38290 26200 38346 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 144 nsew signal input
flabel metal2 s 38934 26200 38990 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 145 nsew signal input
flabel metal2 s 39578 26200 39634 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 146 nsew signal input
flabel metal2 s 40222 26200 40278 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 147 nsew signal input
flabel metal2 s 22834 26200 22890 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 148 nsew signal input
flabel metal2 s 23478 26200 23534 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 149 nsew signal input
flabel metal2 s 24122 26200 24178 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 150 nsew signal input
flabel metal2 s 24766 26200 24822 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 151 nsew signal input
flabel metal2 s 25410 26200 25466 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 152 nsew signal input
flabel metal2 s 26054 26200 26110 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 153 nsew signal input
flabel metal2 s 26698 26200 26754 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 154 nsew signal input
flabel metal2 s 27342 26200 27398 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 155 nsew signal input
flabel metal2 s 2226 26200 2282 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 156 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 157 nsew signal tristate
flabel metal2 s 9310 26200 9366 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 158 nsew signal tristate
flabel metal2 s 9954 26200 10010 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 159 nsew signal tristate
flabel metal2 s 10598 26200 10654 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 160 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 161 nsew signal tristate
flabel metal2 s 11886 26200 11942 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 162 nsew signal tristate
flabel metal2 s 12530 26200 12586 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 163 nsew signal tristate
flabel metal2 s 13174 26200 13230 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 164 nsew signal tristate
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 165 nsew signal tristate
flabel metal2 s 14462 26200 14518 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 166 nsew signal tristate
flabel metal2 s 2870 26200 2926 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 167 nsew signal tristate
flabel metal2 s 15106 26200 15162 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 168 nsew signal tristate
flabel metal2 s 15750 26200 15806 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 169 nsew signal tristate
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 170 nsew signal tristate
flabel metal2 s 17038 26200 17094 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 171 nsew signal tristate
flabel metal2 s 17682 26200 17738 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 172 nsew signal tristate
flabel metal2 s 18326 26200 18382 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 173 nsew signal tristate
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 174 nsew signal tristate
flabel metal2 s 19614 26200 19670 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 175 nsew signal tristate
flabel metal2 s 20258 26200 20314 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 176 nsew signal tristate
flabel metal2 s 20902 26200 20958 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 177 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 178 nsew signal tristate
flabel metal2 s 4158 26200 4214 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 179 nsew signal tristate
flabel metal2 s 4802 26200 4858 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 180 nsew signal tristate
flabel metal2 s 5446 26200 5502 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 181 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 182 nsew signal tristate
flabel metal2 s 6734 26200 6790 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 183 nsew signal tristate
flabel metal2 s 7378 26200 7434 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 184 nsew signal tristate
flabel metal2 s 8022 26200 8078 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 185 nsew signal tristate
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 42154 26200 42210 27000 0 FreeSans 224 90 0 0 prog_reset
port 200 nsew signal input
flabel metal2 s 42798 26200 42854 27000 0 FreeSans 224 90 0 0 reset
port 201 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 202 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 203 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 204 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 205 nsew signal input
flabel metal2 s 43442 26200 43498 27000 0 FreeSans 224 90 0 0 test_enable
port 206 nsew signal input
flabel metal2 s 45374 26200 45430 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 207 nsew signal input
flabel metal2 s 46018 26200 46074 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 208 nsew signal input
flabel metal2 s 46662 26200 46718 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 209 nsew signal input
flabel metal2 s 47306 26200 47362 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 210 nsew signal input
flabel metal2 s 47950 26200 48006 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 211 nsew signal input
flabel metal2 s 48594 26200 48650 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 212 nsew signal input
flabel metal2 s 44086 26200 44142 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 213 nsew signal input
flabel metal2 s 44730 26200 44786 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 214 nsew signal input
flabel metal2 s 1122 0 1178 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_inpad_0_
port 215 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_1__pin_inpad_0_
port 216 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_2__pin_inpad_0_
port 217 nsew signal tristate
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_3__pin_inpad_0_
port 218 nsew signal tristate
rlabel metal1 25484 23936 25484 23936 0 VGND
rlabel metal1 25484 24480 25484 24480 0 VPWR
rlabel metal1 21574 2482 21574 2482 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 20286 3502 20286 3502 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 19504 2958 19504 2958 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 17986 4114 17986 4114 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 20562 20978 20562 20978 0 cbx_1__0_.cbx_8__0_.ccff_head
rlabel metal1 18032 6834 18032 6834 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
rlabel metal1 19458 15674 19458 15674 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
rlabel metal1 14582 13804 14582 13804 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
rlabel metal1 18262 8806 18262 8806 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
rlabel metal2 15594 8806 15594 8806 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
rlabel metal1 18722 9486 18722 9486 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
rlabel metal1 13708 8398 13708 8398 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
rlabel metal1 15180 9350 15180 9350 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
rlabel metal1 12374 10064 12374 10064 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
rlabel metal2 8326 10166 8326 10166 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
rlabel metal1 7774 12274 7774 12274 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
rlabel metal1 9614 11152 9614 11152 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
rlabel metal1 8234 12750 8234 12750 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
rlabel metal1 6762 14348 6762 14348 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
rlabel metal1 12466 14960 12466 14960 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
rlabel metal2 14490 15232 14490 15232 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18262 6766 18262 6766 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 18860 4590 18860 4590 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 14812 13906 14812 13906 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17020 13974 17020 13974 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18354 14042 18354 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17296 7310 17296 7310 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 14858 11186 14858 11186 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16836 14042 16836 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 18170 7514 18170 7514 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 18216 7446 18216 7446 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 16376 6630 16376 6630 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel via2 13202 13379 13202 13379 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15410 9146 15410 9146 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 17802 5202 17802 5202 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 12098 15130 12098 15130 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13432 13906 13432 13906 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14352 13974 14352 13974 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13110 8398 13110 8398 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13110 11186 13110 11186 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 13110 11118 13110 11118 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 13294 8602 13294 8602 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 16698 8602 16698 8602 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 15226 9010 15226 9010 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 9384 15062 9384 15062 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12190 10234 12190 10234 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 13478 6732 13478 6732 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 8648 15130 8648 15130 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17342 15334 17342 15334 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14122 14246 14122 14246 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 13478 9350 13478 9350 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10350 12954 10350 12954 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12512 12410 12512 12410 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 12650 9146 12650 9146 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 12052 10778 12052 10778 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 11362 10098 11362 10098 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 12466 16320 12466 16320 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11362 15130 11362 15130 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 14490 6358 14490 6358 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 12926 16218 12926 16218 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14766 15708 14766 15708 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16330 15402 16330 15402 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 13478 11356 13478 11356 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11960 16218 11960 16218 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 11822 16014 11822 16014 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 12558 10166 12558 10166 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 14904 14042 14904 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 10902 15742 10902 15742 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 17618 3162 17618 3162 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 22540 2482 22540 2482 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 27278 4182 27278 4182 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 23000 3910 23000 3910 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 20056 3434 20056 3434 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 25116 4658 25116 4658 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 25760 2618 25760 2618 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 22632 2550 22632 2550 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 24334 4590 24334 4590 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 17296 4046 17296 4046 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal2 23874 4352 23874 4352 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 9200 1734 9200 1734 0 ccff_head
rlabel metal1 48944 13906 48944 13906 0 ccff_head_1
rlabel metal2 41354 1622 41354 1622 0 ccff_tail
rlabel metal2 1610 24354 1610 24354 0 ccff_tail_0
rlabel metal2 3266 1989 3266 1989 0 chanx_left_in[0]
rlabel metal1 1472 5678 1472 5678 0 chanx_left_in[10]
rlabel metal1 1472 6290 1472 6290 0 chanx_left_in[11]
rlabel metal1 2162 6766 2162 6766 0 chanx_left_in[12]
rlabel metal1 1426 6766 1426 6766 0 chanx_left_in[13]
rlabel metal1 1472 7378 1472 7378 0 chanx_left_in[14]
rlabel metal1 1472 7854 1472 7854 0 chanx_left_in[15]
rlabel metal2 1610 8245 1610 8245 0 chanx_left_in[16]
rlabel metal1 2346 8908 2346 8908 0 chanx_left_in[17]
rlabel metal1 1472 8942 1472 8942 0 chanx_left_in[18]
rlabel metal1 1886 9554 1886 9554 0 chanx_left_in[19]
rlabel metal1 2346 2380 2346 2380 0 chanx_left_in[1]
rlabel metal2 2806 8415 2806 8415 0 chanx_left_in[20]
rlabel metal1 2346 10608 2346 10608 0 chanx_left_in[21]
rlabel metal1 1610 10676 1610 10676 0 chanx_left_in[22]
rlabel metal2 1610 10676 1610 10676 0 chanx_left_in[23]
rlabel metal3 1717 11356 1717 11356 0 chanx_left_in[24]
rlabel metal1 4232 9554 4232 9554 0 chanx_left_in[25]
rlabel metal1 1472 11730 1472 11730 0 chanx_left_in[26]
rlabel metal3 2484 12648 2484 12648 0 chanx_left_in[27]
rlabel metal1 1472 12818 1472 12818 0 chanx_left_in[28]
rlabel metal3 1786 13396 1786 13396 0 chanx_left_in[29]
rlabel metal1 1610 2448 1610 2448 0 chanx_left_in[2]
rlabel metal1 1472 3026 1472 3026 0 chanx_left_in[3]
rlabel metal1 1472 3502 1472 3502 0 chanx_left_in[4]
rlabel metal1 2346 4080 2346 4080 0 chanx_left_in[5]
rlabel metal1 1472 4114 1472 4114 0 chanx_left_in[6]
rlabel metal1 1518 4522 1518 4522 0 chanx_left_in[7]
rlabel metal1 1472 5134 1472 5134 0 chanx_left_in[8]
rlabel metal2 2806 5457 2806 5457 0 chanx_left_in[9]
rlabel metal2 2806 13583 2806 13583 0 chanx_left_out[0]
rlabel metal2 2806 18275 2806 18275 0 chanx_left_out[10]
rlabel metal3 1372 18292 1372 18292 0 chanx_left_out[11]
rlabel metal2 2898 19227 2898 19227 0 chanx_left_out[12]
rlabel metal2 2806 19737 2806 19737 0 chanx_left_out[13]
rlabel metal2 2990 19720 2990 19720 0 chanx_left_out[14]
rlabel metal2 3358 20689 3358 20689 0 chanx_left_out[15]
rlabel via2 3910 20349 3910 20349 0 chanx_left_out[16]
rlabel metal3 1004 20740 1004 20740 0 chanx_left_out[17]
rlabel metal2 2852 21148 2852 21148 0 chanx_left_out[18]
rlabel metal3 1694 21556 1694 21556 0 chanx_left_out[19]
rlabel metal3 820 14212 820 14212 0 chanx_left_out[1]
rlabel metal2 3266 22015 3266 22015 0 chanx_left_out[20]
rlabel metal3 1579 22372 1579 22372 0 chanx_left_out[21]
rlabel metal2 3726 22457 3726 22457 0 chanx_left_out[22]
rlabel metal2 3266 23103 3266 23103 0 chanx_left_out[23]
rlabel metal1 6348 21454 6348 21454 0 chanx_left_out[24]
rlabel metal2 3404 21556 3404 21556 0 chanx_left_out[25]
rlabel metal1 6256 19890 6256 19890 0 chanx_left_out[26]
rlabel metal1 6670 20502 6670 20502 0 chanx_left_out[27]
rlabel via2 4094 25211 4094 25211 0 chanx_left_out[28]
rlabel via1 9798 22073 9798 22073 0 chanx_left_out[29]
rlabel metal3 1004 14620 1004 14620 0 chanx_left_out[2]
rlabel metal3 1004 15028 1004 15028 0 chanx_left_out[3]
rlabel metal3 1004 15436 1004 15436 0 chanx_left_out[4]
rlabel metal3 1004 15844 1004 15844 0 chanx_left_out[5]
rlabel metal3 1004 16252 1004 16252 0 chanx_left_out[6]
rlabel metal3 1004 16660 1004 16660 0 chanx_left_out[7]
rlabel metal3 958 17068 958 17068 0 chanx_left_out[8]
rlabel metal3 1372 17476 1372 17476 0 chanx_left_out[9]
rlabel metal3 47572 13668 47572 13668 0 chanx_right_in_0[0]
rlabel metal3 48308 17748 48308 17748 0 chanx_right_in_0[10]
rlabel metal1 47840 14994 47840 14994 0 chanx_right_in_0[11]
rlabel metal2 49864 15436 49864 15436 0 chanx_right_in_0[12]
rlabel metal1 48852 17238 48852 17238 0 chanx_right_in_0[13]
rlabel metal3 49849 19380 49849 19380 0 chanx_right_in_0[14]
rlabel metal3 49872 19788 49872 19788 0 chanx_right_in_0[15]
rlabel metal3 44275 13260 44275 13260 0 chanx_right_in_0[16]
rlabel metal1 50462 19346 50462 19346 0 chanx_right_in_0[17]
rlabel metal2 46782 16762 46782 16762 0 chanx_right_in_0[18]
rlabel metal3 48262 21420 48262 21420 0 chanx_right_in_0[19]
rlabel metal3 49757 14076 49757 14076 0 chanx_right_in_0[1]
rlabel metal1 50186 20706 50186 20706 0 chanx_right_in_0[20]
rlabel metal1 47104 13906 47104 13906 0 chanx_right_in_0[21]
rlabel metal2 36754 17935 36754 17935 0 chanx_right_in_0[22]
rlabel metal1 50370 17374 50370 17374 0 chanx_right_in_0[23]
rlabel metal1 45862 7378 45862 7378 0 chanx_right_in_0[24]
rlabel metal1 46276 6290 46276 6290 0 chanx_right_in_0[25]
rlabel metal2 49956 17238 49956 17238 0 chanx_right_in_0[26]
rlabel metal2 46598 5746 46598 5746 0 chanx_right_in_0[27]
rlabel metal2 41354 22593 41354 22593 0 chanx_right_in_0[28]
rlabel metal3 44712 13532 44712 13532 0 chanx_right_in_0[29]
rlabel metal3 50010 14484 50010 14484 0 chanx_right_in_0[2]
rlabel metal3 48124 14892 48124 14892 0 chanx_right_in_0[3]
rlabel metal2 45816 13804 45816 13804 0 chanx_right_in_0[4]
rlabel metal3 49964 15708 49964 15708 0 chanx_right_in_0[5]
rlabel metal3 48837 16116 48837 16116 0 chanx_right_in_0[6]
rlabel metal3 49021 16524 49021 16524 0 chanx_right_in_0[7]
rlabel metal3 48170 16932 48170 16932 0 chanx_right_in_0[8]
rlabel metal3 48484 17476 48484 17476 0 chanx_right_in_0[9]
rlabel metal3 48492 1428 48492 1428 0 chanx_right_out_0[0]
rlabel metal1 49312 4658 49312 4658 0 chanx_right_out_0[10]
rlabel metal2 49174 5593 49174 5593 0 chanx_right_out_0[11]
rlabel metal3 49504 6324 49504 6324 0 chanx_right_out_0[12]
rlabel metal1 49266 5746 49266 5746 0 chanx_right_out_0[13]
rlabel metal1 49220 6358 49220 6358 0 chanx_right_out_0[14]
rlabel metal2 49174 7191 49174 7191 0 chanx_right_out_0[15]
rlabel metal2 46874 8177 46874 8177 0 chanx_right_out_0[16]
rlabel metal1 49266 7446 49266 7446 0 chanx_right_out_0[17]
rlabel metal1 49220 7922 49220 7922 0 chanx_right_out_0[18]
rlabel metal2 49174 8857 49174 8857 0 chanx_right_out_0[19]
rlabel metal3 48538 1836 48538 1836 0 chanx_right_out_0[1]
rlabel metal3 48584 9588 48584 9588 0 chanx_right_out_0[20]
rlabel metal1 49220 9010 49220 9010 0 chanx_right_out_0[21]
rlabel metal1 49312 9622 49312 9622 0 chanx_right_out_0[22]
rlabel metal2 49174 10455 49174 10455 0 chanx_right_out_0[23]
rlabel metal1 49266 10710 49266 10710 0 chanx_right_out_0[24]
rlabel metal2 49174 11407 49174 11407 0 chanx_right_out_0[25]
rlabel metal2 49174 11917 49174 11917 0 chanx_right_out_0[26]
rlabel metal3 49734 12444 49734 12444 0 chanx_right_out_0[27]
rlabel via2 49174 12835 49174 12835 0 chanx_right_out_0[28]
rlabel metal3 49734 13260 49734 13260 0 chanx_right_out_0[29]
rlabel metal3 49412 2244 49412 2244 0 chanx_right_out_0[2]
rlabel metal3 48584 2652 48584 2652 0 chanx_right_out_0[3]
rlabel metal3 49504 3060 49504 3060 0 chanx_right_out_0[4]
rlabel metal3 49734 3468 49734 3468 0 chanx_right_out_0[5]
rlabel metal1 49220 3094 49220 3094 0 chanx_right_out_0[6]
rlabel metal2 49174 3927 49174 3927 0 chanx_right_out_0[7]
rlabel metal1 47610 5134 47610 5134 0 chanx_right_out_0[8]
rlabel metal1 49220 4114 49220 4114 0 chanx_right_out_0[9]
rlabel metal3 21137 23460 21137 23460 0 chany_top_in[0]
rlabel metal1 32200 22134 32200 22134 0 chany_top_in[10]
rlabel metal2 35650 6647 35650 6647 0 chany_top_in[11]
rlabel metal2 26128 12420 26128 12420 0 chany_top_in[12]
rlabel metal1 39238 8398 39238 8398 0 chany_top_in[13]
rlabel metal1 33074 13872 33074 13872 0 chany_top_in[14]
rlabel metal2 36754 9928 36754 9928 0 chany_top_in[15]
rlabel metal2 31878 22236 31878 22236 0 chany_top_in[16]
rlabel metal3 33488 11220 33488 11220 0 chany_top_in[17]
rlabel metal3 34109 23188 34109 23188 0 chany_top_in[18]
rlabel metal3 33971 23460 33971 23460 0 chany_top_in[19]
rlabel metal1 21298 21522 21298 21522 0 chany_top_in[1]
rlabel metal2 33902 24548 33902 24548 0 chany_top_in[20]
rlabel metal2 35512 19108 35512 19108 0 chany_top_in[21]
rlabel metal2 35834 26231 35834 26231 0 chany_top_in[22]
rlabel metal3 37099 23324 37099 23324 0 chany_top_in[23]
rlabel metal2 41354 8024 41354 8024 0 chany_top_in[24]
rlabel metal3 38111 23460 38111 23460 0 chany_top_in[25]
rlabel metal2 38318 26173 38318 26173 0 chany_top_in[26]
rlabel metal3 39215 23460 39215 23460 0 chany_top_in[27]
rlabel metal2 39192 17204 39192 17204 0 chany_top_in[28]
rlabel metal3 40779 20604 40779 20604 0 chany_top_in[29]
rlabel metal2 20746 7820 20746 7820 0 chany_top_in[2]
rlabel metal2 23789 26316 23789 26316 0 chany_top_in[3]
rlabel metal2 14122 7667 14122 7667 0 chany_top_in[4]
rlabel via2 40066 8517 40066 8517 0 chany_top_in[5]
rlabel metal1 48484 19142 48484 19142 0 chany_top_in[6]
rlabel via3 5773 11764 5773 11764 0 chany_top_in[7]
rlabel metal1 4922 21046 4922 21046 0 chany_top_in[8]
rlabel metal4 35972 19856 35972 19856 0 chany_top_in[9]
rlabel metal2 2254 24252 2254 24252 0 chany_top_out[0]
rlabel metal1 8464 24242 8464 24242 0 chany_top_out[10]
rlabel metal2 9154 25041 9154 25041 0 chany_top_out[11]
rlabel metal2 10258 24429 10258 24429 0 chany_top_out[12]
rlabel metal2 10718 25041 10718 25041 0 chany_top_out[13]
rlabel metal2 11270 24728 11270 24728 0 chany_top_out[14]
rlabel metal1 12466 22100 12466 22100 0 chany_top_out[15]
rlabel metal2 12466 25279 12466 25279 0 chany_top_out[16]
rlabel metal2 13386 24735 13386 24735 0 chany_top_out[17]
rlabel metal2 13846 24422 13846 24422 0 chany_top_out[18]
rlabel metal1 14030 24242 14030 24242 0 chany_top_out[19]
rlabel metal2 4370 21835 4370 21835 0 chany_top_out[1]
rlabel metal1 14720 23766 14720 23766 0 chany_top_out[20]
rlabel metal2 15870 24497 15870 24497 0 chany_top_out[21]
rlabel metal2 16422 24728 16422 24728 0 chany_top_out[22]
rlabel metal1 16606 23766 16606 23766 0 chany_top_out[23]
rlabel metal1 17848 22066 17848 22066 0 chany_top_out[24]
rlabel metal1 17250 24106 17250 24106 0 chany_top_out[25]
rlabel metal2 18998 25034 18998 25034 0 chany_top_out[26]
rlabel metal1 18998 24242 18998 24242 0 chany_top_out[27]
rlabel metal2 20286 24796 20286 24796 0 chany_top_out[28]
rlabel metal2 21298 25279 21298 25279 0 chany_top_out[29]
rlabel metal1 3404 24242 3404 24242 0 chany_top_out[2]
rlabel metal1 4094 23766 4094 23766 0 chany_top_out[3]
rlabel metal2 5106 24429 5106 24429 0 chany_top_out[4]
rlabel metal2 5474 24966 5474 24966 0 chany_top_out[5]
rlabel metal2 6118 24728 6118 24728 0 chany_top_out[6]
rlabel metal1 5842 24276 5842 24276 0 chany_top_out[7]
rlabel metal1 7682 22542 7682 22542 0 chany_top_out[8]
rlabel metal2 7866 24735 7866 24735 0 chany_top_out[9]
rlabel metal1 16100 19754 16100 19754 0 clknet_0_prog_clk
rlabel metal2 16330 5508 16330 5508 0 clknet_4_0_0_prog_clk
rlabel metal1 35880 12750 35880 12750 0 clknet_4_10_0_prog_clk
rlabel metal1 34500 14382 34500 14382 0 clknet_4_11_0_prog_clk
rlabel metal1 32292 18802 32292 18802 0 clknet_4_12_0_prog_clk
rlabel metal1 24610 22542 24610 22542 0 clknet_4_13_0_prog_clk
rlabel metal2 34914 16320 34914 16320 0 clknet_4_14_0_prog_clk
rlabel metal2 37490 22882 37490 22882 0 clknet_4_15_0_prog_clk
rlabel metal1 10626 13362 10626 13362 0 clknet_4_1_0_prog_clk
rlabel metal2 21850 5916 21850 5916 0 clknet_4_2_0_prog_clk
rlabel metal1 21252 13362 21252 13362 0 clknet_4_3_0_prog_clk
rlabel metal2 8510 18462 8510 18462 0 clknet_4_4_0_prog_clk
rlabel metal1 15801 22066 15801 22066 0 clknet_4_5_0_prog_clk
rlabel metal2 20746 20230 20746 20230 0 clknet_4_6_0_prog_clk
rlabel metal2 17894 20400 17894 20400 0 clknet_4_7_0_prog_clk
rlabel metal2 32338 13056 32338 13056 0 clknet_4_8_0_prog_clk
rlabel metal1 29946 14450 29946 14450 0 clknet_4_9_0_prog_clk
rlabel metal2 11730 1622 11730 1622 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 13846 1622 13846 1622 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 15962 823 15962 823 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 18078 823 18078 823 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 28796 2414 28796 2414 0 gfpga_pad_io_soc_in[0]
rlabel metal1 30912 2414 30912 2414 0 gfpga_pad_io_soc_in[1]
rlabel metal2 33166 1989 33166 1989 0 gfpga_pad_io_soc_in[2]
rlabel metal1 35144 2414 35144 2414 0 gfpga_pad_io_soc_in[3]
rlabel metal1 20102 4046 20102 4046 0 gfpga_pad_io_soc_out[0]
rlabel metal1 21643 2958 21643 2958 0 gfpga_pad_io_soc_out[1]
rlabel metal1 23644 3434 23644 3434 0 gfpga_pad_io_soc_out[2]
rlabel metal2 26542 1554 26542 1554 0 gfpga_pad_io_soc_out[3]
rlabel metal2 37122 1520 37122 1520 0 isol_n
rlabel metal2 10534 3196 10534 3196 0 net1
rlabel metal1 16790 18258 16790 18258 0 net10
rlabel metal1 17250 15572 17250 15572 0 net100
rlabel via2 16054 17085 16054 17085 0 net101
rlabel via2 12834 15555 12834 15555 0 net102
rlabel metal2 17342 18275 17342 18275 0 net103
rlabel metal2 16054 19023 16054 19023 0 net104
rlabel metal1 33718 21862 33718 21862 0 net105
rlabel metal2 14398 21539 14398 21539 0 net106
rlabel metal1 39514 2414 39514 2414 0 net107
rlabel metal2 10258 18802 10258 18802 0 net108
rlabel metal1 1794 13260 1794 13260 0 net109
rlabel via2 19550 14909 19550 14909 0 net11
rlabel metal1 5336 18122 5336 18122 0 net110
rlabel metal2 1794 18326 1794 18326 0 net111
rlabel metal1 1794 19856 1794 19856 0 net112
rlabel metal1 1794 20468 1794 20468 0 net113
rlabel metal1 1794 20944 1794 20944 0 net114
rlabel metal1 1794 21454 1794 21454 0 net115
rlabel metal2 3634 19414 3634 19414 0 net116
rlabel metal1 1794 21964 1794 21964 0 net117
rlabel metal1 1794 22644 1794 22644 0 net118
rlabel metal2 1794 22457 1794 22457 0 net119
rlabel metal2 1794 8857 1794 8857 0 net12
rlabel metal2 11270 16252 11270 16252 0 net120
rlabel metal1 3910 16150 3910 16150 0 net121
rlabel metal1 16169 24854 16169 24854 0 net122
rlabel via2 15134 18955 15134 18955 0 net123
rlabel metal1 5520 20910 5520 20910 0 net124
rlabel metal1 5520 21590 5520 21590 0 net125
rlabel metal1 4002 18700 4002 18700 0 net126
rlabel metal1 6026 19788 6026 19788 0 net127
rlabel metal2 2714 15776 2714 15776 0 net128
rlabel metal2 5796 12716 5796 12716 0 net129
rlabel via2 1794 9435 1794 9435 0 net13
rlabel metal1 6026 12614 6026 12614 0 net130
rlabel metal1 1886 14382 1886 14382 0 net131
rlabel metal1 2277 14994 2277 14994 0 net132
rlabel metal2 3634 14756 3634 14756 0 net133
rlabel metal2 1794 15691 1794 15691 0 net134
rlabel metal2 12834 17323 12834 17323 0 net135
rlabel metal1 1840 17170 1840 17170 0 net136
rlabel metal1 1794 17612 1794 17612 0 net137
rlabel metal1 2277 18258 2277 18258 0 net138
rlabel metal1 41814 4114 41814 4114 0 net139
rlabel metal2 16054 2655 16054 2655 0 net14
rlabel metal2 40250 6256 40250 6256 0 net140
rlabel metal1 47932 5202 47932 5202 0 net141
rlabel metal2 42642 7344 42642 7344 0 net142
rlabel metal2 42550 7276 42550 7276 0 net143
rlabel metal2 40342 7752 40342 7752 0 net144
rlabel metal1 47886 6766 47886 6766 0 net145
rlabel metal1 45862 8398 45862 8398 0 net146
rlabel metal2 39330 7922 39330 7922 0 net147
rlabel metal2 47150 8602 47150 8602 0 net148
rlabel metal1 47932 8466 47932 8466 0 net149
rlabel metal1 15134 16218 15134 16218 0 net15
rlabel metal2 39422 3740 39422 3740 0 net150
rlabel metal1 43792 10166 43792 10166 0 net151
rlabel metal2 39882 9214 39882 9214 0 net152
rlabel metal1 47426 9554 47426 9554 0 net153
rlabel metal1 47978 9996 47978 9996 0 net154
rlabel metal2 45402 9520 45402 9520 0 net155
rlabel metal1 47978 11152 47978 11152 0 net156
rlabel metal1 46322 8058 46322 8058 0 net157
rlabel metal1 46690 15334 46690 15334 0 net158
rlabel metal1 46644 12682 46644 12682 0 net159
rlabel metal1 17756 16150 17756 16150 0 net16
rlabel metal1 46184 12954 46184 12954 0 net160
rlabel metal1 44344 2414 44344 2414 0 net161
rlabel metal1 45816 3026 45816 3026 0 net162
rlabel metal2 40434 4318 40434 4318 0 net163
rlabel metal1 47978 2448 47978 2448 0 net164
rlabel metal2 38410 5984 38410 5984 0 net165
rlabel metal1 47564 3502 47564 3502 0 net166
rlabel metal2 40158 6256 40158 6256 0 net167
rlabel metal2 39238 5882 39238 5882 0 net168
rlabel metal1 3680 19822 3680 19822 0 net169
rlabel via2 1794 10523 1794 10523 0 net17
rlabel metal1 7406 24140 7406 24140 0 net170
rlabel metal2 17250 17612 17250 17612 0 net171
rlabel via2 3450 12291 3450 12291 0 net172
rlabel metal2 16652 20332 16652 20332 0 net173
rlabel metal2 10534 23732 10534 23732 0 net174
rlabel metal2 17986 17663 17986 17663 0 net175
rlabel metal1 9384 24242 9384 24242 0 net176
rlabel metal3 17894 19108 17894 19108 0 net177
rlabel metal2 12742 22355 12742 22355 0 net178
rlabel metal1 13294 24174 13294 24174 0 net179
rlabel metal3 32844 22440 32844 22440 0 net18
rlabel metal2 2622 16694 2622 16694 0 net180
rlabel metal2 14674 23494 14674 23494 0 net181
rlabel metal2 15226 21546 15226 21546 0 net182
rlabel metal1 16054 23086 16054 23086 0 net183
rlabel metal2 15042 24378 15042 24378 0 net184
rlabel metal1 17342 23494 17342 23494 0 net185
rlabel metal1 15180 24174 15180 24174 0 net186
rlabel metal1 18400 23698 18400 23698 0 net187
rlabel metal1 18538 24174 18538 24174 0 net188
rlabel metal1 31832 22610 31832 22610 0 net189
rlabel metal2 5934 12852 5934 12852 0 net19
rlabel metal2 17158 5185 17158 5185 0 net190
rlabel metal2 2162 18802 2162 18802 0 net191
rlabel metal1 4140 10642 4140 10642 0 net192
rlabel metal1 2116 14518 2116 14518 0 net193
rlabel via3 7659 9588 7659 9588 0 net194
rlabel metal2 4324 22610 4324 22610 0 net195
rlabel metal2 2438 20367 2438 20367 0 net196
rlabel metal1 7590 19890 7590 19890 0 net197
rlabel metal3 7935 18700 7935 18700 0 net198
rlabel metal1 14398 3366 14398 3366 0 net199
rlabel metal1 47334 16558 47334 16558 0 net2
rlabel metal3 6394 12444 6394 12444 0 net20
rlabel metal1 15456 2414 15456 2414 0 net200
rlabel metal1 17894 3026 17894 3026 0 net201
rlabel metal1 17710 2346 17710 2346 0 net202
rlabel metal2 20746 11220 20746 11220 0 net203
rlabel metal2 17066 5474 17066 5474 0 net204
rlabel metal2 18584 21590 18584 21590 0 net205
rlabel metal2 17986 17102 17986 17102 0 net206
rlabel metal1 7498 14790 7498 14790 0 net207
rlabel metal1 17848 12818 17848 12818 0 net208
rlabel metal2 33350 9282 33350 9282 0 net209
rlabel metal2 1794 12563 1794 12563 0 net21
rlabel metal1 36708 12614 36708 12614 0 net210
rlabel metal1 34960 19754 34960 19754 0 net211
rlabel metal1 27147 23018 27147 23018 0 net212
rlabel metal1 43247 23018 43247 23018 0 net213
rlabel metal1 44712 8058 44712 8058 0 net214
rlabel metal2 16974 21471 16974 21471 0 net215
rlabel via2 9154 19669 9154 19669 0 net216
rlabel metal1 23184 13906 23184 13906 0 net217
rlabel metal2 37122 20672 37122 20672 0 net218
rlabel metal1 18124 14314 18124 14314 0 net219
rlabel metal1 3266 13906 3266 13906 0 net22
rlabel metal1 24610 17748 24610 17748 0 net220
rlabel metal1 20516 13226 20516 13226 0 net221
rlabel metal1 29440 16218 29440 16218 0 net222
rlabel metal1 31556 5746 31556 5746 0 net223
rlabel metal1 31648 13838 31648 13838 0 net224
rlabel metal2 34178 15810 34178 15810 0 net225
rlabel metal1 29900 9622 29900 9622 0 net226
rlabel metal1 27968 8874 27968 8874 0 net227
rlabel metal2 31510 6987 31510 6987 0 net228
rlabel metal1 38548 7922 38548 7922 0 net229
rlabel metal1 1978 12818 1978 12818 0 net23
rlabel metal2 34178 9452 34178 9452 0 net230
rlabel metal1 28566 9894 28566 9894 0 net231
rlabel metal1 33488 6426 33488 6426 0 net232
rlabel metal1 32959 19822 32959 19822 0 net233
rlabel metal1 32430 15368 32430 15368 0 net234
rlabel metal1 37628 16490 37628 16490 0 net235
rlabel metal1 43746 14450 43746 14450 0 net236
rlabel metal1 38180 12206 38180 12206 0 net237
rlabel metal1 34408 12750 34408 12750 0 net238
rlabel metal2 37490 16184 37490 16184 0 net239
rlabel metal1 23644 19958 23644 19958 0 net24
rlabel metal1 25852 15062 25852 15062 0 net240
rlabel metal2 25760 12580 25760 12580 0 net241
rlabel metal1 21091 11798 21091 11798 0 net242
rlabel metal2 24978 10506 24978 10506 0 net243
rlabel metal1 19320 6834 19320 6834 0 net244
rlabel metal1 19228 5746 19228 5746 0 net245
rlabel metal1 14766 8942 14766 8942 0 net246
rlabel metal1 19642 12818 19642 12818 0 net247
rlabel metal1 22724 10030 22724 10030 0 net248
rlabel metal2 31326 16660 31326 16660 0 net249
rlabel metal1 37398 4488 37398 4488 0 net25
rlabel metal1 13018 14994 13018 14994 0 net250
rlabel metal4 15180 13532 15180 13532 0 net251
rlabel metal1 11822 19142 11822 19142 0 net252
rlabel metal1 10534 19346 10534 19346 0 net253
rlabel metal2 11546 17884 11546 17884 0 net254
rlabel metal2 14766 21471 14766 21471 0 net255
rlabel metal3 12788 18972 12788 18972 0 net256
rlabel metal2 36386 23647 36386 23647 0 net257
rlabel metal1 36754 21862 36754 21862 0 net258
rlabel metal1 16928 5746 16928 5746 0 net259
rlabel metal1 17204 7446 17204 7446 0 net26
rlabel metal2 15870 7106 15870 7106 0 net260
rlabel metal1 10948 7922 10948 7922 0 net261
rlabel metal1 16422 6290 16422 6290 0 net262
rlabel metal1 23414 10710 23414 10710 0 net263
rlabel metal2 18262 11424 18262 11424 0 net264
rlabel metal1 19734 19822 19734 19822 0 net265
rlabel metal1 19734 21420 19734 21420 0 net266
rlabel metal1 27232 19414 27232 19414 0 net267
rlabel metal2 48622 15164 48622 15164 0 net268
rlabel metal2 48438 17476 48438 17476 0 net269
rlabel metal1 1886 3638 1886 3638 0 net27
rlabel metal1 9614 2822 9614 2822 0 net270
rlabel metal1 13248 3026 13248 3026 0 net271
rlabel metal1 7314 15130 7314 15130 0 net272
rlabel metal1 18400 5270 18400 5270 0 net273
rlabel metal2 20102 3910 20102 3910 0 net274
rlabel metal2 14582 8908 14582 8908 0 net275
rlabel metal2 20286 7242 20286 7242 0 net276
rlabel via2 5198 10251 5198 10251 0 net277
rlabel metal1 43516 20570 43516 20570 0 net278
rlabel metal2 31602 7684 31602 7684 0 net279
rlabel metal1 18032 7378 18032 7378 0 net28
rlabel metal1 29348 3502 29348 3502 0 net280
rlabel metal2 43286 19652 43286 19652 0 net281
rlabel metal1 40066 14416 40066 14416 0 net282
rlabel metal2 10350 9350 10350 9350 0 net283
rlabel metal1 9062 17850 9062 17850 0 net284
rlabel metal2 41906 21556 41906 21556 0 net285
rlabel metal1 7590 17306 7590 17306 0 net286
rlabel metal2 45954 16252 45954 16252 0 net287
rlabel metal1 10120 16558 10120 16558 0 net288
rlabel metal2 18446 9061 18446 9061 0 net289
rlabel via1 2438 4029 2438 4029 0 net29
rlabel metal1 27830 8602 27830 8602 0 net290
rlabel metal2 42642 17340 42642 17340 0 net291
rlabel metal1 24380 4794 24380 4794 0 net292
rlabel metal1 37858 17306 37858 17306 0 net293
rlabel metal2 43746 23868 43746 23868 0 net294
rlabel metal2 12788 23324 12788 23324 0 net295
rlabel metal3 48553 20740 48553 20740 0 net296
rlabel metal2 4922 14212 4922 14212 0 net297
rlabel metal1 20056 6426 20056 6426 0 net298
rlabel metal1 43378 16762 43378 16762 0 net299
rlabel metal2 14260 7718 14260 7718 0 net3
rlabel metal2 19734 5304 19734 5304 0 net30
rlabel metal2 42274 15946 42274 15946 0 net300
rlabel metal2 43746 12988 43746 12988 0 net301
rlabel metal2 11730 14076 11730 14076 0 net302
rlabel metal1 9614 13294 9614 13294 0 net303
rlabel metal1 5842 14518 5842 14518 0 net304
rlabel metal1 1702 23664 1702 23664 0 net305
rlabel metal1 46092 18938 46092 18938 0 net306
rlabel metal2 6854 15946 6854 15946 0 net307
rlabel metal1 34408 5678 34408 5678 0 net308
rlabel metal2 10718 8670 10718 8670 0 net309
rlabel metal1 9062 11186 9062 11186 0 net31
rlabel metal2 6854 18496 6854 18496 0 net310
rlabel metal2 34914 6970 34914 6970 0 net311
rlabel metal1 45126 17034 45126 17034 0 net312
rlabel metal1 40940 10234 40940 10234 0 net313
rlabel metal1 18216 18258 18216 18258 0 net314
rlabel metal1 7360 14042 7360 14042 0 net315
rlabel metal1 43608 21998 43608 21998 0 net316
rlabel metal1 30452 22066 30452 22066 0 net317
rlabel metal1 23598 6324 23598 6324 0 net318
rlabel metal1 7360 13294 7360 13294 0 net319
rlabel metal1 14168 8602 14168 8602 0 net32
rlabel metal2 12006 8092 12006 8092 0 net320
rlabel metal1 45356 15130 45356 15130 0 net321
rlabel metal1 46506 18258 46506 18258 0 net322
rlabel metal1 6210 12886 6210 12886 0 net323
rlabel metal1 23184 4046 23184 4046 0 net324
rlabel metal1 1702 12138 1702 12138 0 net325
rlabel metal1 42274 13328 42274 13328 0 net326
rlabel metal1 21436 20978 21436 20978 0 net327
rlabel metal2 10074 14212 10074 14212 0 net328
rlabel metal2 47426 21114 47426 21114 0 net329
rlabel metal1 40710 15062 40710 15062 0 net33
rlabel metal2 18906 6086 18906 6086 0 net330
rlabel metal2 45494 20740 45494 20740 0 net331
rlabel metal1 38962 9690 38962 9690 0 net332
rlabel metal1 5336 17306 5336 17306 0 net333
rlabel metal2 29394 7684 29394 7684 0 net334
rlabel metal2 5750 17850 5750 17850 0 net335
rlabel metal2 9798 20026 9798 20026 0 net336
rlabel metal2 28382 16524 28382 16524 0 net337
rlabel metal1 21758 6290 21758 6290 0 net338
rlabel metal2 45954 20094 45954 20094 0 net339
rlabel via2 16146 11067 16146 11067 0 net34
rlabel metal1 30176 6290 30176 6290 0 net340
rlabel metal1 45264 13906 45264 13906 0 net341
rlabel metal2 7866 11934 7866 11934 0 net342
rlabel metal1 25990 17714 25990 17714 0 net343
rlabel metal1 38916 12410 38916 12410 0 net344
rlabel metal1 12489 20434 12489 20434 0 net345
rlabel metal1 25162 6426 25162 6426 0 net346
rlabel metal1 8832 12614 8832 12614 0 net347
rlabel metal1 20608 15538 20608 15538 0 net348
rlabel metal1 26956 8058 26956 8058 0 net349
rlabel metal1 18584 13498 18584 13498 0 net35
rlabel metal1 9292 11050 9292 11050 0 net350
rlabel metal2 39974 12988 39974 12988 0 net351
rlabel metal1 15778 7514 15778 7514 0 net352
rlabel metal1 14076 21658 14076 21658 0 net353
rlabel metal1 31234 6426 31234 6426 0 net354
rlabel metal1 13754 15946 13754 15946 0 net355
rlabel metal1 5980 18054 5980 18054 0 net356
rlabel metal2 23598 5508 23598 5508 0 net357
rlabel metal1 15870 8874 15870 8874 0 net358
rlabel metal2 32890 13583 32890 13583 0 net359
rlabel via2 45494 6613 45494 6613 0 net36
rlabel metal2 25898 8704 25898 8704 0 net360
rlabel metal1 39468 18190 39468 18190 0 net361
rlabel metal1 15042 7310 15042 7310 0 net362
rlabel metal2 38502 18785 38502 18785 0 net363
rlabel metal1 18722 20468 18722 20468 0 net364
rlabel metal2 25162 24072 25162 24072 0 net365
rlabel metal2 40434 10302 40434 10302 0 net366
rlabel via2 32246 12835 32246 12835 0 net367
rlabel metal2 21436 13260 21436 13260 0 net368
rlabel metal1 37207 23290 37207 23290 0 net369
rlabel metal3 21252 22984 21252 22984 0 net37
rlabel metal1 24886 13192 24886 13192 0 net370
rlabel metal2 42090 14688 42090 14688 0 net371
rlabel metal1 16468 6426 16468 6426 0 net372
rlabel metal1 38410 20978 38410 20978 0 net373
rlabel metal2 21206 10608 21206 10608 0 net374
rlabel metal1 33442 7514 33442 7514 0 net375
rlabel metal1 27508 14450 27508 14450 0 net376
rlabel metal2 37766 11968 37766 11968 0 net377
rlabel metal3 37697 22372 37697 22372 0 net378
rlabel metal1 13754 20264 13754 20264 0 net379
rlabel via2 16146 20451 16146 20451 0 net38
rlabel metal2 19642 17544 19642 17544 0 net380
rlabel via2 39146 11339 39146 11339 0 net381
rlabel via2 19734 24123 19734 24123 0 net382
rlabel metal1 14812 18598 14812 18598 0 net383
rlabel metal2 38318 14773 38318 14773 0 net384
rlabel metal1 35696 20978 35696 20978 0 net385
rlabel metal2 38594 16422 38594 16422 0 net386
rlabel metal1 39790 13226 39790 13226 0 net387
rlabel metal1 20332 16490 20332 16490 0 net388
rlabel metal2 32292 21862 32292 21862 0 net389
rlabel metal2 1794 24480 1794 24480 0 net39
rlabel metal1 37582 10506 37582 10506 0 net390
rlabel metal2 11270 10030 11270 10030 0 net391
rlabel metal1 11500 21114 11500 21114 0 net392
rlabel metal1 27508 18190 27508 18190 0 net393
rlabel metal2 30682 7939 30682 7939 0 net394
rlabel metal4 30084 24616 30084 24616 0 net395
rlabel via2 34730 18309 34730 18309 0 net396
rlabel metal2 24058 8007 24058 8007 0 net397
rlabel metal1 30360 6630 30360 6630 0 net398
rlabel metal1 27968 7514 27968 7514 0 net399
rlabel metal1 1794 5576 1794 5576 0 net4
rlabel metal2 42826 13872 42826 13872 0 net40
rlabel metal2 38962 13957 38962 13957 0 net400
rlabel metal1 27968 8058 27968 8058 0 net401
rlabel metal1 3864 12954 3864 12954 0 net402
rlabel metal1 11040 9146 11040 9146 0 net403
rlabel metal2 30130 19669 30130 19669 0 net404
rlabel metal1 10028 15402 10028 15402 0 net405
rlabel metal1 36524 8466 36524 8466 0 net406
rlabel via2 32890 17221 32890 17221 0 net407
rlabel metal2 6440 12852 6440 12852 0 net408
rlabel metal2 46966 24021 46966 24021 0 net409
rlabel metal2 19366 21777 19366 21777 0 net41
rlabel via2 38594 21573 38594 21573 0 net410
rlabel metal2 32062 24344 32062 24344 0 net411
rlabel metal1 14214 13294 14214 13294 0 net412
rlabel metal1 10258 13498 10258 13498 0 net413
rlabel metal2 14030 11730 14030 11730 0 net414
rlabel metal2 26634 16218 26634 16218 0 net415
rlabel metal1 48254 14382 48254 14382 0 net416
rlabel metal2 48806 16388 48806 16388 0 net417
rlabel metal1 47794 17204 47794 17204 0 net418
rlabel metal2 42688 21046 42688 21046 0 net419
rlabel metal1 19550 15130 19550 15130 0 net42
rlabel metal1 9430 2414 9430 2414 0 net420
rlabel metal1 9430 3060 9430 3060 0 net421
rlabel metal2 12374 3196 12374 3196 0 net422
rlabel metal1 14490 2958 14490 2958 0 net423
rlabel metal1 8280 14586 8280 14586 0 net424
rlabel metal1 4876 17238 4876 17238 0 net425
rlabel metal2 18446 5372 18446 5372 0 net426
rlabel metal2 17158 8160 17158 8160 0 net427
rlabel metal2 12190 7446 12190 7446 0 net428
rlabel metal1 16790 8534 16790 8534 0 net429
rlabel metal2 34730 17391 34730 17391 0 net43
rlabel metal2 42642 19414 42642 19414 0 net430
rlabel metal1 38134 20332 38134 20332 0 net431
rlabel metal1 18860 3502 18860 3502 0 net432
rlabel metal1 21206 4250 21206 4250 0 net433
rlabel metal2 12098 24616 12098 24616 0 net434
rlabel metal2 18906 22457 18906 22457 0 net435
rlabel metal1 42826 20434 42826 20434 0 net436
rlabel metal1 43470 21658 43470 21658 0 net437
rlabel metal1 28060 3502 28060 3502 0 net438
rlabel metal2 29118 3230 29118 3230 0 net439
rlabel metal3 18492 15368 18492 15368 0 net44
rlabel metal2 22034 7310 22034 7310 0 net440
rlabel metal1 20010 6698 20010 6698 0 net441
rlabel metal2 9706 9452 9706 9452 0 net442
rlabel metal1 11040 9486 11040 9486 0 net443
rlabel metal2 30958 7548 30958 7548 0 net444
rlabel metal2 28382 9928 28382 9928 0 net445
rlabel metal1 41584 14042 41584 14042 0 net446
rlabel via2 40158 14331 40158 14331 0 net447
rlabel metal2 9982 17442 9982 17442 0 net448
rlabel metal2 14214 18496 14214 18496 0 net449
rlabel metal1 41722 21930 41722 21930 0 net45
rlabel metal2 9246 16660 9246 16660 0 net450
rlabel metal2 17986 16014 17986 16014 0 net451
rlabel metal1 8556 15606 8556 15606 0 net452
rlabel metal1 12834 17578 12834 17578 0 net453
rlabel metal1 41216 20910 41216 20910 0 net454
rlabel metal1 43240 22066 43240 22066 0 net455
rlabel metal1 46322 16524 46322 16524 0 net456
rlabel metal1 44022 15572 44022 15572 0 net457
rlabel metal2 24518 8636 24518 8636 0 net458
rlabel metal2 19274 13294 19274 13294 0 net459
rlabel metal2 19918 15980 19918 15980 0 net46
rlabel metal2 24058 4046 24058 4046 0 net460
rlabel metal2 24886 4284 24886 4284 0 net461
rlabel metal1 42090 16762 42090 16762 0 net462
rlabel metal1 32982 17544 32982 17544 0 net463
rlabel metal2 6026 13396 6026 13396 0 net464
rlabel metal2 15042 20927 15042 20927 0 net465
rlabel metal1 10856 14042 10856 14042 0 net466
rlabel metal2 13754 14195 13754 14195 0 net467
rlabel metal2 25990 8636 25990 8636 0 net468
rlabel metal1 29992 11322 29992 11322 0 net469
rlabel metal2 19182 17918 19182 17918 0 net47
rlabel metal1 42642 24140 42642 24140 0 net470
rlabel metal2 27278 24276 27278 24276 0 net471
rlabel metal2 43286 13124 43286 13124 0 net472
rlabel metal1 39422 12716 39422 12716 0 net473
rlabel metal1 16468 16558 16468 16558 0 net474
rlabel metal1 20631 18394 20631 18394 0 net475
rlabel metal1 42872 16558 42872 16558 0 net476
rlabel metal1 39882 17000 39882 17000 0 net477
rlabel metal1 5704 13158 5704 13158 0 net478
rlabel metal1 16514 22610 16514 22610 0 net479
rlabel metal1 18584 15130 18584 15130 0 net48
rlabel metal2 44390 16388 44390 16388 0 net480
rlabel metal1 39882 16184 39882 16184 0 net481
rlabel metal1 19734 6324 19734 6324 0 net482
rlabel metal1 20194 7514 20194 7514 0 net483
rlabel metal1 10534 8534 10534 8534 0 net484
rlabel metal3 12167 15028 12167 15028 0 net485
rlabel metal1 12972 7378 12972 7378 0 net486
rlabel metal2 12834 10404 12834 10404 0 net487
rlabel metal1 44620 14994 44620 14994 0 net488
rlabel metal2 45494 15776 45494 15776 0 net489
rlabel metal1 45448 7514 45448 7514 0 net49
rlabel metal2 37490 17612 37490 17612 0 net490
rlabel metal1 30544 16490 30544 16490 0 net491
rlabel metal2 6026 14212 6026 14212 0 net492
rlabel metal2 10810 16337 10810 16337 0 net493
rlabel metal1 8280 15062 8280 15062 0 net494
rlabel metal1 7728 15674 7728 15674 0 net495
rlabel metal1 45218 18768 45218 18768 0 net496
rlabel metal1 43654 19924 43654 19924 0 net497
rlabel metal1 46644 21386 46644 21386 0 net498
rlabel metal1 33327 2550 33327 2550 0 net499
rlabel metal1 14168 10778 14168 10778 0 net5
rlabel metal1 41032 20774 41032 20774 0 net50
rlabel metal2 7130 13838 7130 13838 0 net500
rlabel metal2 13938 19941 13938 19941 0 net501
rlabel metal1 46092 23290 46092 23290 0 net502
rlabel metal2 32798 24548 32798 24548 0 net503
rlabel metal1 45678 16558 45678 16558 0 net504
rlabel metal1 40135 17102 40135 17102 0 net505
rlabel via1 12282 21539 12282 21539 0 net506
rlabel metal2 34178 24514 34178 24514 0 net507
rlabel metal1 7222 13940 7222 13940 0 net508
rlabel metal1 14766 21998 14766 21998 0 net509
rlabel metal1 33350 6188 33350 6188 0 net51
rlabel metal1 43516 14994 43516 14994 0 net510
rlabel metal2 37398 13923 37398 13923 0 net511
rlabel metal1 7222 16150 7222 16150 0 net512
rlabel metal2 18170 22593 18170 22593 0 net513
rlabel metal1 26358 6732 26358 6732 0 net514
rlabel metal2 24242 7616 24242 7616 0 net515
rlabel metal2 40710 10234 40710 10234 0 net516
rlabel metal1 39054 11186 39054 11186 0 net517
rlabel metal1 35236 7378 35236 7378 0 net518
rlabel metal1 33902 6834 33902 6834 0 net519
rlabel metal3 40503 23460 40503 23460 0 net52
rlabel metal1 47242 14586 47242 14586 0 net520
rlabel metal1 46184 21046 46184 21046 0 net521
rlabel metal1 29486 21998 29486 21998 0 net522
rlabel metal1 27048 24174 27048 24174 0 net523
rlabel metal1 11086 11798 11086 11798 0 net524
rlabel metal1 13984 12886 13984 12886 0 net525
rlabel metal2 20194 5236 20194 5236 0 net526
rlabel metal1 19320 6426 19320 6426 0 net527
rlabel metal2 45862 20230 45862 20230 0 net528
rlabel metal1 38318 20536 38318 20536 0 net529
rlabel metal2 41078 7922 41078 7922 0 net53
rlabel metal1 4784 20570 4784 20570 0 net530
rlabel metal2 2346 24106 2346 24106 0 net531
rlabel metal1 7268 18938 7268 18938 0 net532
rlabel via2 15226 19805 15226 19805 0 net533
rlabel metal2 21022 6086 21022 6086 0 net534
rlabel metal2 21942 8738 21942 8738 0 net535
rlabel metal2 22034 4556 22034 4556 0 net536
rlabel metal2 20562 7310 20562 7310 0 net537
rlabel metal1 44252 22406 44252 22406 0 net538
rlabel metal2 39974 8874 39974 8874 0 net539
rlabel metal1 20056 21862 20056 21862 0 net54
rlabel metal2 48438 19380 48438 19380 0 net540
rlabel metal2 44022 17918 44022 17918 0 net541
rlabel metal1 35098 6698 35098 6698 0 net542
rlabel metal2 30774 7446 30774 7446 0 net543
rlabel metal1 28750 7344 28750 7344 0 net544
rlabel metal1 27324 13226 27324 13226 0 net545
rlabel metal2 38594 10030 38594 10030 0 net546
rlabel metal1 38134 10064 38134 10064 0 net547
rlabel metal2 39606 19941 39606 19941 0 net548
rlabel metal2 2346 15810 2346 15810 0 net549
rlabel metal4 18676 16592 18676 16592 0 net55
rlabel metal1 43792 20026 43792 20026 0 net550
rlabel metal1 38870 19448 38870 19448 0 net551
rlabel metal1 9200 13906 9200 13906 0 net552
rlabel metal1 11960 14586 11960 14586 0 net553
rlabel metal1 25898 15674 25898 15674 0 net554
rlabel metal1 25845 13702 25845 13702 0 net555
rlabel metal2 7222 10574 7222 10574 0 net556
rlabel metal1 8418 18870 8418 18870 0 net557
rlabel metal1 6854 16558 6854 16558 0 net558
rlabel metal2 10994 17833 10994 17833 0 net559
rlabel metal1 21390 15572 21390 15572 0 net56
rlabel metal2 30406 6324 30406 6324 0 net560
rlabel metal1 30544 6426 30544 6426 0 net561
rlabel metal2 9430 21148 9430 21148 0 net562
rlabel metal2 13754 19550 13754 19550 0 net563
rlabel metal1 25944 7854 25944 7854 0 net564
rlabel metal1 26450 9146 26450 9146 0 net565
rlabel metal2 24702 6732 24702 6732 0 net566
rlabel metal1 23920 8058 23920 8058 0 net567
rlabel metal2 12558 21318 12558 21318 0 net568
rlabel metal1 25392 24038 25392 24038 0 net569
rlabel metal3 40779 15300 40779 15300 0 net57
rlabel metal1 17894 6426 17894 6426 0 net570
rlabel metal1 16928 8058 16928 8058 0 net571
rlabel metal2 22218 16218 22218 16218 0 net572
rlabel metal1 24472 17102 24472 17102 0 net573
rlabel metal1 8970 19346 8970 19346 0 net574
rlabel metal1 20138 17850 20138 17850 0 net575
rlabel metal2 41722 13124 41722 13124 0 net576
rlabel metal2 40618 13107 40618 13107 0 net577
rlabel metal1 7452 13158 7452 13158 0 net578
rlabel metal1 4968 12954 4968 12954 0 net579
rlabel metal1 17756 8466 17756 8466 0 net58
rlabel metal1 9890 22950 9890 22950 0 net580
rlabel metal1 28658 18394 28658 18394 0 net581
rlabel metal2 22954 5372 22954 5372 0 net582
rlabel metal1 23782 5882 23782 5882 0 net583
rlabel metal1 6854 11152 6854 11152 0 net584
rlabel metal2 32890 7072 32890 7072 0 net585
rlabel metal1 35098 8058 35098 8058 0 net586
rlabel metal2 6026 17238 6026 17238 0 net587
rlabel metal2 6026 23171 6026 23171 0 net588
rlabel metal2 10534 16796 10534 16796 0 net589
rlabel metal1 35834 24820 35834 24820 0 net59
rlabel metal1 40296 13498 40296 13498 0 net590
rlabel metal2 25254 6970 25254 6970 0 net591
rlabel metal1 15778 6834 15778 6834 0 net592
rlabel metal1 41262 23732 41262 23732 0 net593
rlabel metal1 10258 10642 10258 10642 0 net594
rlabel metal1 46598 15028 46598 15028 0 net595
rlabel metal2 11546 20196 11546 20196 0 net596
rlabel viali 43740 19346 43740 19346 0 net597
rlabel metal1 20148 7854 20148 7854 0 net598
rlabel metal1 43746 20468 43746 20468 0 net599
rlabel metal1 2346 6664 2346 6664 0 net6
rlabel metal2 13570 17731 13570 17731 0 net60
rlabel metal1 38226 8602 38226 8602 0 net600
rlabel metal1 47426 13498 47426 13498 0 net601
rlabel metal1 38824 13294 38824 13294 0 net602
rlabel metal1 26634 14586 26634 14586 0 net603
rlabel metal1 15686 6256 15686 6256 0 net604
rlabel metal2 41446 12036 41446 12036 0 net605
rlabel metal1 41446 15028 41446 15028 0 net606
rlabel metal3 14973 16660 14973 16660 0 net607
rlabel metal2 38364 10676 38364 10676 0 net608
rlabel metal1 46368 14042 46368 14042 0 net609
rlabel metal3 41101 14756 41101 14756 0 net61
rlabel metal1 13110 18768 13110 18768 0 net610
rlabel metal1 33626 7344 33626 7344 0 net611
rlabel metal1 47380 14382 47380 14382 0 net612
rlabel metal2 37030 15113 37030 15113 0 net613
rlabel metal1 39974 11730 39974 11730 0 net614
rlabel metal1 14260 17306 14260 17306 0 net615
rlabel metal1 7130 19380 7130 19380 0 net616
rlabel metal1 29624 23698 29624 23698 0 net617
rlabel metal1 47012 12886 47012 12886 0 net618
rlabel metal2 44390 14212 44390 14212 0 net619
rlabel metal1 13432 12818 13432 12818 0 net62
rlabel metal1 32660 6426 32660 6426 0 net620
rlabel metal1 17250 14450 17250 14450 0 net621
rlabel metal1 41768 20434 41768 20434 0 net622
rlabel metal2 23414 6970 23414 6970 0 net623
rlabel metal2 43746 18428 43746 18428 0 net624
rlabel viali 38686 10644 38686 10644 0 net625
rlabel metal2 45954 17340 45954 17340 0 net626
rlabel metal1 10810 20944 10810 20944 0 net627
rlabel metal2 29302 6596 29302 6596 0 net628
rlabel metal1 28428 6834 28428 6834 0 net629
rlabel metal2 14950 6222 14950 6222 0 net63
rlabel metal1 45724 22746 45724 22746 0 net630
rlabel metal1 4002 12750 4002 12750 0 net631
rlabel metal2 9430 11084 9430 11084 0 net632
rlabel metal2 43286 14212 43286 14212 0 net633
rlabel metal1 27738 7854 27738 7854 0 net634
rlabel metal1 10810 8976 10810 8976 0 net635
rlabel metal1 6624 14586 6624 14586 0 net636
rlabel metal2 42642 18428 42642 18428 0 net637
rlabel metal1 31326 24038 31326 24038 0 net638
rlabel metal2 46874 22916 46874 22916 0 net639
rlabel metal1 31188 18054 31188 18054 0 net64
rlabel metal1 36110 8432 36110 8432 0 net640
rlabel metal2 48530 20298 48530 20298 0 net641
rlabel metal1 8924 10778 8924 10778 0 net642
rlabel metal2 8878 13124 8878 13124 0 net643
rlabel metal1 9016 16082 9016 16082 0 net644
rlabel metal1 27002 12954 27002 12954 0 net645
rlabel metal1 11546 7990 11546 7990 0 net646
rlabel metal1 45954 21556 45954 21556 0 net647
rlabel metal1 48852 14042 48852 14042 0 net648
rlabel metal2 49358 15028 49358 15028 0 net649
rlabel metal1 28520 20842 28520 20842 0 net65
rlabel metal2 49266 15606 49266 15606 0 net650
rlabel metal1 49082 16422 49082 16422 0 net651
rlabel metal1 48300 16422 48300 16422 0 net652
rlabel metal1 9246 2482 9246 2482 0 net653
rlabel metal1 9062 2958 9062 2958 0 net654
rlabel metal1 10488 2618 10488 2618 0 net655
rlabel metal1 9844 3162 9844 3162 0 net656
rlabel metal2 11178 3332 11178 3332 0 net657
rlabel metal2 38686 8449 38686 8449 0 net66
rlabel metal1 34132 9554 34132 9554 0 net67
rlabel metal1 41630 9010 41630 9010 0 net68
rlabel metal2 35282 18819 35282 18819 0 net69
rlabel metal2 1794 6256 1794 6256 0 net7
rlabel metal1 36754 20434 36754 20434 0 net70
rlabel metal1 35190 20434 35190 20434 0 net71
rlabel metal3 39974 21964 39974 21964 0 net72
rlabel metal3 34086 20876 34086 20876 0 net73
rlabel metal1 23598 20774 23598 20774 0 net74
rlabel metal1 30912 17510 30912 17510 0 net75
rlabel via2 45494 15555 45494 15555 0 net76
rlabel metal2 32246 19040 32246 19040 0 net77
rlabel metal2 44206 11407 44206 11407 0 net78
rlabel metal1 37260 20230 37260 20230 0 net79
rlabel metal2 1794 7072 1794 7072 0 net8
rlabel metal2 35144 20842 35144 20842 0 net80
rlabel metal1 35420 18666 35420 18666 0 net81
rlabel via2 36570 20485 36570 20485 0 net82
rlabel via2 35374 20349 35374 20349 0 net83
rlabel metal1 42412 22066 42412 22066 0 net84
rlabel metal1 17342 21862 17342 21862 0 net85
rlabel metal1 30820 16014 30820 16014 0 net86
rlabel metal2 33442 16031 33442 16031 0 net87
rlabel metal2 34914 14246 34914 14246 0 net88
rlabel metal2 36018 18819 36018 18819 0 net89
rlabel metal2 20194 9044 20194 9044 0 net9
rlabel metal1 17204 18054 17204 18054 0 net90
rlabel metal1 14950 22610 14950 22610 0 net91
rlabel metal1 29900 17646 29900 17646 0 net92
rlabel metal1 26864 2550 26864 2550 0 net93
rlabel metal2 30866 3264 30866 3264 0 net94
rlabel metal1 32936 2618 32936 2618 0 net95
rlabel metal1 34776 2618 34776 2618 0 net96
rlabel metal1 37306 2482 37306 2482 0 net97
rlabel metal1 44344 7174 44344 7174 0 net98
rlabel metal2 40526 16711 40526 16711 0 net99
rlabel metal2 39238 2098 39238 2098 0 prog_clk
rlabel metal2 44390 7939 44390 7939 0 prog_reset
rlabel metal2 33948 9452 33948 9452 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 40434 14251 40434 14251 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 42412 3570 42412 3570 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 34454 14790 34454 14790 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 32890 11628 32890 11628 0 sb_1__0_.mem_left_track_1.ccff_head
rlabel metal2 20930 16626 20930 16626 0 sb_1__0_.mem_left_track_1.ccff_tail
rlabel metal1 27600 19346 27600 19346 0 sb_1__0_.mem_left_track_1.mem_out\[0\]
rlabel metal2 24702 14977 24702 14977 0 sb_1__0_.mem_left_track_1.mem_out\[1\]
rlabel metal1 20194 14484 20194 14484 0 sb_1__0_.mem_left_track_11.ccff_head
rlabel metal1 9430 17102 9430 17102 0 sb_1__0_.mem_left_track_11.ccff_tail
rlabel metal1 17020 13838 17020 13838 0 sb_1__0_.mem_left_track_11.mem_out\[0\]
rlabel metal1 20838 14892 20838 14892 0 sb_1__0_.mem_left_track_11.mem_out\[1\]
rlabel metal1 19228 21454 19228 21454 0 sb_1__0_.mem_left_track_13.ccff_tail
rlabel metal1 21436 19142 21436 19142 0 sb_1__0_.mem_left_track_13.mem_out\[0\]
rlabel metal2 20194 19567 20194 19567 0 sb_1__0_.mem_left_track_13.mem_out\[1\]
rlabel metal1 17526 20910 17526 20910 0 sb_1__0_.mem_left_track_21.ccff_tail
rlabel metal1 21252 16082 21252 16082 0 sb_1__0_.mem_left_track_21.mem_out\[0\]
rlabel metal2 17250 21216 17250 21216 0 sb_1__0_.mem_left_track_21.mem_out\[1\]
rlabel metal3 18492 19652 18492 19652 0 sb_1__0_.mem_left_track_29.ccff_tail
rlabel metal2 12742 21488 12742 21488 0 sb_1__0_.mem_left_track_29.mem_out\[0\]
rlabel metal2 17250 21760 17250 21760 0 sb_1__0_.mem_left_track_29.mem_out\[1\]
rlabel metal2 7866 18972 7866 18972 0 sb_1__0_.mem_left_track_3.ccff_tail
rlabel metal2 14582 19873 14582 19873 0 sb_1__0_.mem_left_track_3.mem_out\[0\]
rlabel metal2 16698 20604 16698 20604 0 sb_1__0_.mem_left_track_3.mem_out\[1\]
rlabel metal1 28520 21998 28520 21998 0 sb_1__0_.mem_left_track_37.ccff_tail
rlabel metal1 27853 19686 27853 19686 0 sb_1__0_.mem_left_track_37.mem_out\[0\]
rlabel metal1 27462 18054 27462 18054 0 sb_1__0_.mem_left_track_37.mem_out\[1\]
rlabel metal2 11822 24208 11822 24208 0 sb_1__0_.mem_left_track_45.ccff_tail
rlabel metal2 39974 24361 39974 24361 0 sb_1__0_.mem_left_track_45.mem_out\[0\]
rlabel metal1 33258 22440 33258 22440 0 sb_1__0_.mem_left_track_45.mem_out\[1\]
rlabel metal1 8234 17238 8234 17238 0 sb_1__0_.mem_left_track_5.ccff_tail
rlabel metal1 17986 19890 17986 19890 0 sb_1__0_.mem_left_track_5.mem_out\[0\]
rlabel metal1 21712 17510 21712 17510 0 sb_1__0_.mem_left_track_5.mem_out\[1\]
rlabel metal2 42734 24225 42734 24225 0 sb_1__0_.mem_left_track_53.mem_out\[0\]
rlabel via2 19366 20315 19366 20315 0 sb_1__0_.mem_left_track_53.mem_out\[1\]
rlabel metal1 26956 18394 26956 18394 0 sb_1__0_.mem_left_track_7.mem_out\[0\]
rlabel metal1 20286 13328 20286 13328 0 sb_1__0_.mem_left_track_7.mem_out\[1\]
rlabel metal1 15778 21454 15778 21454 0 sb_1__0_.mem_right_track_0.ccff_head
rlabel metal1 34270 16626 34270 16626 0 sb_1__0_.mem_right_track_0.ccff_tail
rlabel metal1 30314 21012 30314 21012 0 sb_1__0_.mem_right_track_0.mem_out\[0\]
rlabel metal1 33166 16626 33166 16626 0 sb_1__0_.mem_right_track_0.mem_out\[1\]
rlabel metal2 39238 12070 39238 12070 0 sb_1__0_.mem_right_track_10.ccff_head
rlabel metal1 40894 10676 40894 10676 0 sb_1__0_.mem_right_track_10.ccff_tail
rlabel metal2 31786 8160 31786 8160 0 sb_1__0_.mem_right_track_10.mem_out\[0\]
rlabel metal1 35742 13362 35742 13362 0 sb_1__0_.mem_right_track_10.mem_out\[1\]
rlabel metal1 38134 13804 38134 13804 0 sb_1__0_.mem_right_track_12.ccff_tail
rlabel metal1 34086 7854 34086 7854 0 sb_1__0_.mem_right_track_12.mem_out\[0\]
rlabel metal1 32522 15538 32522 15538 0 sb_1__0_.mem_right_track_12.mem_out\[1\]
rlabel metal2 36662 16218 36662 16218 0 sb_1__0_.mem_right_track_2.ccff_tail
rlabel metal2 39146 18445 39146 18445 0 sb_1__0_.mem_right_track_2.mem_out\[0\]
rlabel metal1 39238 17680 39238 17680 0 sb_1__0_.mem_right_track_2.mem_out\[1\]
rlabel metal1 32430 10166 32430 10166 0 sb_1__0_.mem_right_track_20.ccff_tail
rlabel metal1 32430 20264 32430 20264 0 sb_1__0_.mem_right_track_20.mem_out\[0\]
rlabel metal1 30682 13838 30682 13838 0 sb_1__0_.mem_right_track_20.mem_out\[1\]
rlabel metal2 34914 8058 34914 8058 0 sb_1__0_.mem_right_track_28.ccff_tail
rlabel metal1 26588 9486 26588 9486 0 sb_1__0_.mem_right_track_28.mem_out\[0\]
rlabel metal2 32614 13974 32614 13974 0 sb_1__0_.mem_right_track_28.mem_out\[1\]
rlabel metal2 34270 8636 34270 8636 0 sb_1__0_.mem_right_track_36.ccff_tail
rlabel metal1 32200 6290 32200 6290 0 sb_1__0_.mem_right_track_36.mem_out\[0\]
rlabel metal1 37398 9554 37398 9554 0 sb_1__0_.mem_right_track_36.mem_out\[1\]
rlabel metal1 39330 13804 39330 13804 0 sb_1__0_.mem_right_track_4.ccff_tail
rlabel metal1 36800 15946 36800 15946 0 sb_1__0_.mem_right_track_4.mem_out\[0\]
rlabel metal2 39882 14654 39882 14654 0 sb_1__0_.mem_right_track_4.mem_out\[1\]
rlabel metal1 31418 9078 31418 9078 0 sb_1__0_.mem_right_track_44.ccff_tail
rlabel metal1 33580 6766 33580 6766 0 sb_1__0_.mem_right_track_44.mem_out\[0\]
rlabel metal1 28842 17714 28842 17714 0 sb_1__0_.mem_right_track_52.mem_out\[0\]
rlabel metal1 36800 9146 36800 9146 0 sb_1__0_.mem_right_track_6.mem_out\[0\]
rlabel metal2 35558 13673 35558 13673 0 sb_1__0_.mem_right_track_6.mem_out\[1\]
rlabel metal2 36846 23443 36846 23443 0 sb_1__0_.mem_top_track_0.ccff_tail
rlabel via2 40710 23205 40710 23205 0 sb_1__0_.mem_top_track_0.mem_out\[0\]
rlabel metal2 27646 20791 27646 20791 0 sb_1__0_.mem_top_track_0.mem_out\[1\]
rlabel metal1 39100 20774 39100 20774 0 sb_1__0_.mem_top_track_10.ccff_head
rlabel metal2 36202 18564 36202 18564 0 sb_1__0_.mem_top_track_10.ccff_tail
rlabel metal1 40894 20332 40894 20332 0 sb_1__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 38364 17510 38364 17510 0 sb_1__0_.mem_top_track_10.mem_out\[1\]
rlabel metal1 41262 18122 41262 18122 0 sb_1__0_.mem_top_track_12.ccff_tail
rlabel metal2 38594 19448 38594 19448 0 sb_1__0_.mem_top_track_12.mem_out\[0\]
rlabel metal3 39514 16252 39514 16252 0 sb_1__0_.mem_top_track_12.mem_out\[1\]
rlabel metal1 39974 15878 39974 15878 0 sb_1__0_.mem_top_track_14.ccff_tail
rlabel metal1 47794 18700 47794 18700 0 sb_1__0_.mem_top_track_14.mem_out\[0\]
rlabel metal2 35834 15147 35834 15147 0 sb_1__0_.mem_top_track_14.mem_out\[1\]
rlabel metal1 38962 14790 38962 14790 0 sb_1__0_.mem_top_track_16.ccff_tail
rlabel metal1 41170 16626 41170 16626 0 sb_1__0_.mem_top_track_16.mem_out\[0\]
rlabel metal2 40618 13821 40618 13821 0 sb_1__0_.mem_top_track_16.mem_out\[1\]
rlabel metal1 40986 13940 40986 13940 0 sb_1__0_.mem_top_track_18.ccff_tail
rlabel metal1 39284 15334 39284 15334 0 sb_1__0_.mem_top_track_18.mem_out\[0\]
rlabel metal1 39054 14518 39054 14518 0 sb_1__0_.mem_top_track_18.mem_out\[1\]
rlabel metal1 39146 23664 39146 23664 0 sb_1__0_.mem_top_track_2.ccff_tail
rlabel metal1 35742 8942 35742 8942 0 sb_1__0_.mem_top_track_2.mem_out\[0\]
rlabel metal1 35512 22066 35512 22066 0 sb_1__0_.mem_top_track_2.mem_out\[1\]
rlabel metal1 24932 15470 24932 15470 0 sb_1__0_.mem_top_track_20.ccff_tail
rlabel via2 28566 14773 28566 14773 0 sb_1__0_.mem_top_track_20.mem_out\[0\]
rlabel metal1 25484 13498 25484 13498 0 sb_1__0_.mem_top_track_22.ccff_tail
rlabel metal1 26588 14042 26588 14042 0 sb_1__0_.mem_top_track_22.mem_out\[0\]
rlabel metal1 24150 13362 24150 13362 0 sb_1__0_.mem_top_track_24.ccff_tail
rlabel metal1 26358 12682 26358 12682 0 sb_1__0_.mem_top_track_24.mem_out\[0\]
rlabel metal2 21390 12954 21390 12954 0 sb_1__0_.mem_top_track_26.ccff_tail
rlabel metal1 25116 7378 25116 7378 0 sb_1__0_.mem_top_track_26.mem_out\[0\]
rlabel metal1 19044 10098 19044 10098 0 sb_1__0_.mem_top_track_28.ccff_tail
rlabel metal1 23506 10030 23506 10030 0 sb_1__0_.mem_top_track_28.mem_out\[0\]
rlabel metal2 18722 10336 18722 10336 0 sb_1__0_.mem_top_track_30.ccff_tail
rlabel metal2 20838 6766 20838 6766 0 sb_1__0_.mem_top_track_30.mem_out\[0\]
rlabel metal1 19964 5202 19964 5202 0 sb_1__0_.mem_top_track_32.ccff_tail
rlabel metal1 20608 8398 20608 8398 0 sb_1__0_.mem_top_track_32.mem_out\[0\]
rlabel metal1 20286 12750 20286 12750 0 sb_1__0_.mem_top_track_34.ccff_tail
rlabel metal1 20424 9350 20424 9350 0 sb_1__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 22586 13804 22586 13804 0 sb_1__0_.mem_top_track_36.ccff_tail
rlabel metal2 22816 9010 22816 9010 0 sb_1__0_.mem_top_track_36.mem_out\[0\]
rlabel metal2 34086 20740 34086 20740 0 sb_1__0_.mem_top_track_4.ccff_tail
rlabel metal1 36662 21522 36662 21522 0 sb_1__0_.mem_top_track_4.mem_out\[0\]
rlabel metal2 36662 20553 36662 20553 0 sb_1__0_.mem_top_track_4.mem_out\[1\]
rlabel metal1 13754 14892 13754 14892 0 sb_1__0_.mem_top_track_40.ccff_tail
rlabel metal1 15042 11696 15042 11696 0 sb_1__0_.mem_top_track_40.mem_out\[0\]
rlabel metal1 16008 17510 16008 17510 0 sb_1__0_.mem_top_track_42.ccff_tail
rlabel metal1 16238 15130 16238 15130 0 sb_1__0_.mem_top_track_42.mem_out\[0\]
rlabel metal1 12880 19278 12880 19278 0 sb_1__0_.mem_top_track_44.ccff_tail
rlabel metal2 16146 16898 16146 16898 0 sb_1__0_.mem_top_track_44.mem_out\[0\]
rlabel metal2 9614 18513 9614 18513 0 sb_1__0_.mem_top_track_46.ccff_tail
rlabel metal2 13018 15419 13018 15419 0 sb_1__0_.mem_top_track_46.mem_out\[0\]
rlabel metal2 5750 18972 5750 18972 0 sb_1__0_.mem_top_track_48.ccff_tail
rlabel metal1 13708 19686 13708 19686 0 sb_1__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 14950 21420 14950 21420 0 sb_1__0_.mem_top_track_50.ccff_tail
rlabel metal1 15686 19278 15686 19278 0 sb_1__0_.mem_top_track_50.mem_out\[0\]
rlabel metal2 18630 22304 18630 22304 0 sb_1__0_.mem_top_track_58.mem_out\[0\]
rlabel metal2 39606 14552 39606 14552 0 sb_1__0_.mem_top_track_6.ccff_tail
rlabel metal2 35558 20638 35558 20638 0 sb_1__0_.mem_top_track_6.mem_out\[0\]
rlabel metal2 37214 23018 37214 23018 0 sb_1__0_.mem_top_track_6.mem_out\[1\]
rlabel metal2 39514 17068 39514 17068 0 sb_1__0_.mem_top_track_8.mem_out\[0\]
rlabel metal1 38410 21352 38410 21352 0 sb_1__0_.mem_top_track_8.mem_out\[1\]
rlabel metal1 7866 10030 7866 10030 0 sb_1__0_.mux_left_track_1.out
rlabel metal1 26772 18666 26772 18666 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 26220 18734 26220 18734 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23322 12682 23322 12682 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24288 14994 24288 14994 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23322 17578 23322 17578 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23966 15130 23966 15130 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 20930 17952 20930 17952 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7774 15538 7774 15538 0 sb_1__0_.mux_left_track_11.out
rlabel metal1 24564 18734 24564 18734 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24518 18394 24518 18394 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20884 11594 20884 11594 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20562 11322 20562 11322 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20286 16558 20286 16558 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 20056 15130 20056 15130 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 17342 13158 17342 13158 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 12512 7514 12512 7514 0 sb_1__0_.mux_left_track_13.out
rlabel metal2 21666 21760 21666 21760 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22034 21267 22034 21267 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20700 15674 20700 15674 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20838 21386 20838 21386 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19412 19958 19412 19958 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 19136 15980 19136 15980 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 5382 9350 5382 9350 0 sb_1__0_.mux_left_track_21.out
rlabel metal1 24012 22678 24012 22678 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 23322 22406 23322 22406 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21344 15946 21344 15946 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18538 22134 18538 22134 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 17342 21114 17342 21114 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel via3 16997 20740 16997 20740 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12972 12342 12972 12342 0 sb_1__0_.mux_left_track_29.out
rlabel metal1 26358 21012 26358 21012 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 26726 20570 26726 20570 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23414 15946 23414 15946 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 25622 20774 25622 20774 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22218 20026 22218 20026 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 20194 19023 20194 19023 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9982 12750 9982 12750 0 sb_1__0_.mux_left_track_3.out
rlabel metal2 22494 21879 22494 21879 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 23506 19363 23506 19363 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22034 21726 22034 21726 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 17894 17323 17894 17323 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17434 18598 17434 18598 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 14398 13498 14398 13498 0 sb_1__0_.mux_left_track_37.out
rlabel metal1 32108 21658 32108 21658 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 28612 18734 28612 18734 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24150 16422 24150 16422 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23506 14042 23506 14042 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 21206 15215 21206 15215 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11822 7480 11822 7480 0 sb_1__0_.mux_left_track_45.out
rlabel metal2 30498 23426 30498 23426 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24288 22610 24288 22610 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 25852 22746 25852 22746 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 12006 7395 12006 7395 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 2530 11152 2530 11152 0 sb_1__0_.mux_left_track_5.out
rlabel metal1 23322 19414 23322 19414 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23506 19482 23506 19482 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21666 19482 21666 19482 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17940 14586 17940 14586 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel via3 17365 16660 17365 16660 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 6762 14790 6762 14790 0 sb_1__0_.mux_left_track_53.out
rlabel metal1 26450 22100 26450 22100 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20010 21046 20010 21046 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21436 20570 21436 20570 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel via3 19435 20740 19435 20740 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 6624 12750 6624 12750 0 sb_1__0_.mux_left_track_7.out
rlabel metal1 24104 15470 24104 15470 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 23322 15674 23322 15674 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19918 12410 19918 12410 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22586 14790 22586 14790 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19872 13498 19872 13498 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18262 14552 18262 14552 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 43608 12750 43608 12750 0 sb_1__0_.mux_right_track_0.out
rlabel metal1 29670 20774 29670 20774 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33258 14586 33258 14586 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 27232 15130 27232 15130 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33994 16660 33994 16660 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 33718 16286 33718 16286 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 33580 16422 33580 16422 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 44022 8262 44022 8262 0 sb_1__0_.mux_right_track_10.out
rlabel metal1 35466 13294 35466 13294 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 35558 13226 35558 13226 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 35374 9520 35374 9520 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33511 8534 33511 8534 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel via1 36478 9641 36478 9641 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 35650 8602 35650 8602 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 36018 8704 36018 8704 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 44482 12682 44482 12682 0 sb_1__0_.mux_right_track_12.out
rlabel metal1 32522 15470 32522 15470 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 30866 15674 30866 15674 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 31510 10744 31510 10744 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37950 13804 37950 13804 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32982 10438 32982 10438 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 37996 14042 37996 14042 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 45770 12818 45770 12818 0 sb_1__0_.mux_right_track_2.out
rlabel metal1 33810 19482 33810 19482 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33902 17850 33902 17850 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32890 14552 32890 14552 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 36478 17068 36478 17068 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 34132 16218 34132 16218 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 37306 17034 37306 17034 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 44252 8942 44252 8942 0 sb_1__0_.mux_right_track_20.out
rlabel metal1 30222 15504 30222 15504 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 29946 15470 29946 15470 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 27876 12138 27876 12138 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 32430 9826 32430 9826 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32660 10030 32660 10030 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 33580 10166 33580 10166 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 43286 7208 43286 7208 0 sb_1__0_.mux_right_track_28.out
rlabel metal1 32430 14484 32430 14484 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 32338 14416 32338 14416 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 28750 9180 28750 9180 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 34132 14314 34132 14314 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 34914 9350 34914 9350 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 38962 7378 38962 7378 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 44942 7480 44942 7480 0 sb_1__0_.mux_right_track_36.out
rlabel metal1 32154 16048 32154 16048 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 32798 14960 32798 14960 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 34086 9928 34086 9928 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 33994 8976 33994 8976 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 39974 7412 39974 7412 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 45080 15402 45080 15402 0 sb_1__0_.mux_right_track_4.out
rlabel metal1 35098 17306 35098 17306 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34684 17238 34684 17238 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34592 11866 34592 11866 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 38318 13821 38318 13821 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 39790 12716 39790 12716 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 40043 14042 40043 14042 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 37214 7208 37214 7208 0 sb_1__0_.mux_right_track_44.out
rlabel metal1 30866 16966 30866 16966 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 30682 9962 30682 9962 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35098 7922 35098 7922 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 41032 5678 41032 5678 0 sb_1__0_.mux_right_track_52.out
rlabel metal2 31970 15232 31970 15232 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 32706 11152 32706 11152 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33994 11526 33994 11526 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 45770 7820 45770 7820 0 sb_1__0_.mux_right_track_6.out
rlabel metal2 35374 17680 35374 17680 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34408 15130 34408 15130 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37444 10098 37444 10098 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 34960 8806 34960 8806 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 36524 13838 36524 13838 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 38088 10234 38088 10234 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 38502 10744 38502 10744 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 17250 5202 17250 5202 0 sb_1__0_.mux_top_track_0.out
rlabel metal1 34132 21998 34132 21998 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 37950 23783 37950 23783 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 26266 21114 26266 21114 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 29762 20774 29762 20774 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 31464 22678 31464 22678 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 29624 21658 29624 21658 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal3 31855 18972 31855 18972 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 17342 24480 17342 24480 0 sb_1__0_.mux_top_track_10.out
rlabel metal1 39054 19890 39054 19890 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39698 19822 39698 19822 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33258 18836 33258 18836 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32384 16218 32384 16218 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32706 18870 32706 18870 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel via2 39330 14501 39330 14501 0 sb_1__0_.mux_top_track_12.out
rlabel metal1 41446 18258 41446 18258 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40526 18054 40526 18054 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37628 16762 37628 16762 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 38778 18581 38778 18581 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel via2 35374 14059 35374 14059 0 sb_1__0_.mux_top_track_14.out
rlabel metal1 41262 17238 41262 17238 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40020 17306 40020 17306 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36294 15674 36294 15674 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 35880 13906 35880 13906 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 38962 23001 38962 23001 0 sb_1__0_.mux_top_track_16.out
rlabel metal1 40664 16218 40664 16218 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39606 15912 39606 15912 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37122 12138 37122 12138 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 36202 14790 36202 14790 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal3 16698 20060 16698 20060 0 sb_1__0_.mux_top_track_18.out
rlabel metal1 39560 14926 39560 14926 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39008 15130 39008 15130 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32614 14994 32614 14994 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 27830 16320 27830 16320 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 38686 22831 38686 22831 0 sb_1__0_.mux_top_track_2.out
rlabel metal1 39146 24276 39146 24276 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39560 24106 39560 24106 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32062 21352 32062 21352 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 38686 24072 38686 24072 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 34638 21862 34638 21862 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 32338 23885 32338 23885 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 14352 19414 14352 19414 0 sb_1__0_.mux_top_track_20.out
rlabel metal1 27554 16456 27554 16456 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 25438 16150 25438 16150 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 25392 17306 25392 17306 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13386 6800 13386 6800 0 sb_1__0_.mux_top_track_22.out
rlabel metal1 24150 14382 24150 14382 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24472 14314 24472 14314 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19688 11118 19688 11118 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14674 8058 14674 8058 0 sb_1__0_.mux_top_track_24.out
rlabel metal1 23782 13396 23782 13396 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23966 11594 23966 11594 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14766 7888 14766 7888 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 18722 9061 18722 9061 0 sb_1__0_.mux_top_track_26.out
rlabel metal1 21206 12682 21206 12682 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23460 10166 23460 10166 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20792 12614 20792 12614 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 6394 13991 6394 13991 0 sb_1__0_.mux_top_track_28.out
rlabel metal1 18630 10132 18630 10132 0 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 18170 9945 18170 9945 0 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4048 15674 4048 15674 0 sb_1__0_.mux_top_track_30.out
rlabel metal1 21712 9690 21712 9690 0 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17986 10778 17986 10778 0 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel via3 19573 18020 19573 18020 0 sb_1__0_.mux_top_track_32.out
rlabel metal2 16974 10608 16974 10608 0 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14490 6798 14490 6798 0 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3496 12206 3496 12206 0 sb_1__0_.mux_top_track_34.out
rlabel metal1 18354 11322 18354 11322 0 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 19366 12699 19366 12699 0 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 4002 14501 4002 14501 0 sb_1__0_.mux_top_track_36.out
rlabel metal1 22678 14042 22678 14042 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22172 13770 22172 13770 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22034 13923 22034 13923 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21206 24072 21206 24072 0 sb_1__0_.mux_top_track_4.out
rlabel metal1 36340 21658 36340 21658 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40112 21114 40112 21114 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32614 21862 32614 21862 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 32522 20128 32522 20128 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17112 24174 17112 24174 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 9154 8364 9154 8364 0 sb_1__0_.mux_top_track_40.out
rlabel metal1 14306 11594 14306 11594 0 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12650 13617 12650 13617 0 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 8418 8466 8418 8466 0 sb_1__0_.mux_top_track_42.out
rlabel metal1 16054 15674 16054 15674 0 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 14927 18020 14927 18020 0 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9522 7514 9522 7514 0 sb_1__0_.mux_top_track_44.out
rlabel metal1 15548 17306 15548 17306 0 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12466 18513 12466 18513 0 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6578 8602 6578 8602 0 sb_1__0_.mux_top_track_46.out
rlabel metal1 12052 15674 12052 15674 0 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10304 19482 10304 19482 0 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 7774 9180 7774 9180 0 sb_1__0_.mux_top_track_48.out
rlabel metal1 15778 18394 15778 18394 0 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 12811 20876 12811 20876 0 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6854 9622 6854 9622 0 sb_1__0_.mux_top_track_50.out
rlabel metal2 15594 20502 15594 20502 0 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 13823 13668 13823 13668 0 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 2806 10234 2806 10234 0 sb_1__0_.mux_top_track_58.out
rlabel metal2 19642 21760 19642 21760 0 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_0_X
rlabel via3 15709 20740 15709 20740 0 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28658 19856 28658 19856 0 sb_1__0_.mux_top_track_6.out
rlabel metal1 38548 22202 38548 22202 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40480 22746 40480 22746 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32614 19448 32614 19448 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 39698 23460 39698 23460 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 36294 23834 36294 23834 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 37490 24480 37490 24480 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel via2 29210 24157 29210 24157 0 sb_1__0_.mux_top_track_8.out
rlabel metal2 40066 21726 40066 21726 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 41262 21760 41262 21760 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34960 17850 34960 17850 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 39192 21658 39192 21658 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 36202 21896 36202 21896 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 37628 22134 37628 22134 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 44942 9860 44942 9860 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
rlabel metal1 45494 10030 45494 10030 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
rlabel metal1 46276 9554 46276 9554 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
rlabel metal3 45793 20876 45793 20876 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
rlabel metal1 48944 17170 48944 17170 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
rlabel metal2 48576 16252 48576 16252 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
rlabel via2 16882 23715 16882 23715 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
rlabel metal2 37674 21471 37674 21471 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
rlabel metal2 1150 1095 1150 1095 0 top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 21758 16048 21758 16048 0 top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 19596 13362 19596 13362 0 top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 21850 10880 21850 10880 0 top_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 27000
<< end >>
