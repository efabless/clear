magic
tech sky130A
magscale 1 2
timestamp 1625786074
<< locali >>
rect 15393 14943 15427 15113
rect 18981 13991 19015 14977
rect 6285 11543 6319 11645
rect 6193 10591 6227 10693
rect 8861 9367 8895 9673
rect 8769 8891 8803 9061
rect 13093 8823 13127 9129
rect 3341 8279 3375 8585
rect 8953 6647 8987 6817
rect 16405 6239 16439 6409
rect 2697 5627 2731 5865
rect 13185 5559 13219 5865
rect 12449 5083 12483 5253
rect 10241 3587 10275 3689
<< viali >>
rect 15393 15113 15427 15147
rect 15393 14909 15427 14943
rect 18981 14977 19015 15011
rect 1593 14569 1627 14603
rect 1961 14569 1995 14603
rect 2697 14569 2731 14603
rect 4629 14569 4663 14603
rect 8953 14569 8987 14603
rect 10149 14569 10183 14603
rect 11437 14569 11471 14603
rect 13277 14569 13311 14603
rect 13553 14569 13587 14603
rect 14933 14569 14967 14603
rect 17233 14569 17267 14603
rect 1869 14501 1903 14535
rect 2237 14501 2271 14535
rect 3249 14501 3283 14535
rect 3893 14501 3927 14535
rect 4261 14501 4295 14535
rect 4813 14501 4847 14535
rect 4997 14501 5031 14535
rect 5457 14501 5491 14535
rect 6745 14501 6779 14535
rect 7573 14501 7607 14535
rect 7757 14501 7791 14535
rect 13461 14501 13495 14535
rect 14013 14501 14047 14535
rect 14565 14501 14599 14535
rect 15117 14501 15151 14535
rect 15761 14501 15795 14535
rect 16773 14501 16807 14535
rect 16957 14501 16991 14535
rect 17693 14501 17727 14535
rect 18061 14501 18095 14535
rect 1501 14433 1535 14467
rect 2605 14433 2639 14467
rect 3065 14433 3099 14467
rect 3433 14433 3467 14467
rect 3617 14433 3651 14467
rect 4077 14433 4111 14467
rect 4445 14433 4479 14467
rect 5641 14433 5675 14467
rect 6009 14433 6043 14467
rect 6377 14433 6411 14467
rect 6561 14433 6595 14467
rect 6929 14433 6963 14467
rect 8861 14433 8895 14467
rect 9321 14433 9355 14467
rect 9597 14433 9631 14467
rect 9965 14433 9999 14467
rect 10241 14433 10275 14467
rect 10609 14433 10643 14467
rect 10885 14433 10919 14467
rect 11253 14433 11287 14467
rect 11529 14433 11563 14467
rect 11897 14433 11931 14467
rect 12173 14433 12207 14467
rect 12541 14433 12575 14467
rect 12817 14433 12851 14467
rect 13093 14433 13127 14467
rect 13829 14433 13863 14467
rect 14197 14433 14231 14467
rect 14749 14433 14783 14467
rect 15301 14433 15335 14467
rect 15485 14433 15519 14467
rect 15945 14433 15979 14467
rect 16589 14433 16623 14467
rect 17417 14433 17451 14467
rect 18429 14433 18463 14467
rect 16313 14365 16347 14399
rect 2421 14297 2455 14331
rect 9505 14297 9539 14331
rect 12081 14297 12115 14331
rect 14381 14297 14415 14331
rect 17877 14297 17911 14331
rect 18245 14297 18279 14331
rect 2973 14229 3007 14263
rect 5917 14229 5951 14263
rect 6193 14229 6227 14263
rect 7481 14229 7515 14263
rect 8677 14229 8711 14263
rect 10793 14229 10827 14263
rect 12725 14229 12759 14263
rect 15669 14229 15703 14263
rect 16497 14229 16531 14263
rect 17601 14229 17635 14263
rect 1961 14025 1995 14059
rect 4077 14025 4111 14059
rect 4721 14025 4755 14059
rect 6653 14025 6687 14059
rect 13737 14025 13771 14059
rect 15117 14025 15151 14059
rect 15577 14025 15611 14059
rect 16589 14025 16623 14059
rect 16773 14025 16807 14059
rect 17693 14025 17727 14059
rect 2237 13957 2271 13991
rect 2605 13957 2639 13991
rect 2881 13957 2915 13991
rect 3249 13957 3283 13991
rect 3525 13957 3559 13991
rect 3985 13957 4019 13991
rect 6193 13957 6227 13991
rect 13277 13957 13311 13991
rect 13461 13957 13495 13991
rect 14381 13957 14415 13991
rect 17877 13957 17911 13991
rect 18245 13957 18279 13991
rect 18981 13957 19015 13991
rect 17049 13889 17083 13923
rect 1409 13821 1443 13855
rect 1593 13821 1627 13855
rect 1777 13821 1811 13855
rect 2421 13821 2455 13855
rect 2789 13821 2823 13855
rect 3065 13821 3099 13855
rect 3433 13821 3467 13855
rect 3709 13821 3743 13855
rect 3801 13821 3835 13855
rect 4261 13821 4295 13855
rect 4537 13821 4571 13855
rect 6009 13821 6043 13855
rect 6469 13821 6503 13855
rect 13645 13821 13679 13855
rect 14565 13821 14599 13855
rect 15301 13821 15335 13855
rect 15761 13821 15795 13855
rect 16405 13821 16439 13855
rect 17233 13821 17267 13855
rect 17417 13821 17451 13855
rect 18429 13821 18463 13855
rect 2053 13753 2087 13787
rect 17601 13753 17635 13787
rect 18061 13753 18095 13787
rect 13921 13685 13955 13719
rect 3341 13481 3375 13515
rect 17049 13481 17083 13515
rect 17233 13481 17267 13515
rect 17601 13481 17635 13515
rect 1869 13413 1903 13447
rect 2973 13413 3007 13447
rect 3525 13413 3559 13447
rect 17417 13413 17451 13447
rect 18153 13413 18187 13447
rect 1501 13345 1535 13379
rect 2145 13345 2179 13379
rect 2605 13345 2639 13379
rect 2706 13345 2740 13379
rect 3157 13345 3191 13379
rect 16865 13345 16899 13379
rect 17969 13345 18003 13379
rect 18429 13345 18463 13379
rect 3893 13277 3927 13311
rect 17785 13277 17819 13311
rect 1685 13209 1719 13243
rect 2329 13209 2363 13243
rect 2881 13209 2915 13243
rect 4353 13209 4387 13243
rect 18245 13209 18279 13243
rect 1961 13141 1995 13175
rect 2421 13141 2455 13175
rect 4169 13141 4203 13175
rect 2973 12937 3007 12971
rect 17509 12937 17543 12971
rect 3525 12869 3559 12903
rect 2697 12801 2731 12835
rect 18245 12801 18279 12835
rect 1501 12733 1535 12767
rect 1685 12733 1719 12767
rect 3341 12733 3375 12767
rect 17785 12733 17819 12767
rect 18429 12733 18463 12767
rect 1869 12665 1903 12699
rect 2513 12665 2547 12699
rect 17417 12665 17451 12699
rect 18061 12665 18095 12699
rect 1961 12597 1995 12631
rect 2145 12597 2179 12631
rect 2605 12597 2639 12631
rect 3249 12597 3283 12631
rect 3801 12597 3835 12631
rect 17969 12597 18003 12631
rect 3065 12393 3099 12427
rect 2697 12325 2731 12359
rect 4169 12325 4203 12359
rect 1501 12257 1535 12291
rect 1869 12257 1903 12291
rect 2605 12257 2639 12291
rect 4793 12257 4827 12291
rect 17601 12257 17635 12291
rect 18061 12257 18095 12291
rect 18429 12257 18463 12291
rect 2789 12189 2823 12223
rect 3525 12189 3559 12223
rect 4537 12189 4571 12223
rect 17785 12189 17819 12223
rect 1685 12121 1719 12155
rect 17877 12121 17911 12155
rect 1961 12053 1995 12087
rect 2237 12053 2271 12087
rect 3341 12053 3375 12087
rect 3893 12053 3927 12087
rect 5917 12053 5951 12087
rect 18337 12053 18371 12087
rect 5733 11849 5767 11883
rect 2329 11713 2363 11747
rect 2513 11713 2547 11747
rect 1501 11645 1535 11679
rect 2237 11645 2271 11679
rect 2789 11645 2823 11679
rect 4261 11645 4295 11679
rect 6285 11645 6319 11679
rect 6469 11645 6503 11679
rect 6725 11645 6759 11679
rect 7941 11645 7975 11679
rect 9045 11645 9079 11679
rect 17877 11645 17911 11679
rect 3034 11577 3068 11611
rect 4506 11577 4540 11611
rect 8769 11577 8803 11611
rect 17785 11577 17819 11611
rect 18429 11577 18463 11611
rect 1593 11509 1627 11543
rect 1869 11509 1903 11543
rect 4169 11509 4203 11543
rect 5641 11509 5675 11543
rect 6285 11509 6319 11543
rect 7849 11509 7883 11543
rect 17509 11509 17543 11543
rect 18061 11509 18095 11543
rect 18337 11509 18371 11543
rect 3157 11305 3191 11339
rect 3985 11305 4019 11339
rect 5273 11305 5307 11339
rect 5825 11305 5859 11339
rect 18061 11305 18095 11339
rect 7950 11237 7984 11271
rect 11560 11237 11594 11271
rect 17049 11237 17083 11271
rect 17325 11237 17359 11271
rect 1501 11169 1535 11203
rect 2237 11169 2271 11203
rect 3065 11169 3099 11203
rect 4905 11169 4939 11203
rect 5365 11169 5399 11203
rect 6193 11169 6227 11203
rect 6745 11169 6779 11203
rect 8217 11169 8251 11203
rect 11805 11169 11839 11203
rect 13562 11169 13596 11203
rect 17877 11169 17911 11203
rect 18429 11169 18463 11203
rect 2329 11101 2363 11135
rect 2513 11101 2547 11135
rect 3341 11101 3375 11135
rect 5181 11101 5215 11135
rect 6285 11101 6319 11135
rect 6469 11101 6503 11135
rect 13829 11101 13863 11135
rect 17601 11101 17635 11135
rect 1685 11033 1719 11067
rect 3525 11033 3559 11067
rect 4169 11033 4203 11067
rect 12449 11033 12483 11067
rect 17785 11033 17819 11067
rect 18245 11033 18279 11067
rect 1869 10965 1903 10999
rect 2697 10965 2731 10999
rect 5733 10965 5767 10999
rect 6837 10965 6871 10999
rect 10425 10965 10459 10999
rect 11897 10965 11931 10999
rect 16957 10965 16991 10999
rect 2513 10761 2547 10795
rect 4169 10761 4203 10795
rect 13553 10761 13587 10795
rect 6193 10693 6227 10727
rect 1869 10625 1903 10659
rect 2053 10625 2087 10659
rect 5733 10625 5767 10659
rect 7021 10625 7055 10659
rect 11345 10625 11379 10659
rect 12357 10625 12391 10659
rect 13277 10625 13311 10659
rect 14933 10625 14967 10659
rect 17509 10625 17543 10659
rect 2145 10557 2179 10591
rect 3718 10557 3752 10591
rect 3985 10557 4019 10591
rect 5549 10557 5583 10591
rect 6101 10557 6135 10591
rect 6193 10557 6227 10591
rect 6837 10557 6871 10591
rect 6929 10557 6963 10591
rect 7389 10557 7423 10591
rect 7645 10557 7679 10591
rect 10234 10557 10268 10591
rect 10425 10557 10459 10591
rect 16589 10557 16623 10591
rect 16773 10557 16807 10591
rect 1501 10489 1535 10523
rect 9974 10489 10008 10523
rect 11161 10489 11195 10523
rect 12173 10489 12207 10523
rect 13001 10489 13035 10523
rect 14666 10489 14700 10523
rect 17325 10489 17359 10523
rect 17877 10489 17911 10523
rect 18061 10489 18095 10523
rect 18429 10489 18463 10523
rect 1593 10421 1627 10455
rect 2605 10421 2639 10455
rect 5089 10421 5123 10455
rect 5457 10421 5491 10455
rect 5917 10421 5951 10455
rect 6469 10421 6503 10455
rect 8769 10421 8803 10455
rect 8861 10421 8895 10455
rect 10793 10421 10827 10455
rect 11253 10421 11287 10455
rect 11805 10421 11839 10455
rect 12265 10421 12299 10455
rect 12633 10421 12667 10455
rect 13093 10421 13127 10455
rect 16957 10421 16991 10455
rect 17417 10421 17451 10455
rect 18337 10421 18371 10455
rect 1869 10217 1903 10251
rect 1961 10217 1995 10251
rect 2421 10217 2455 10251
rect 2881 10217 2915 10251
rect 3433 10217 3467 10251
rect 3709 10217 3743 10251
rect 4905 10217 4939 10251
rect 5273 10217 5307 10251
rect 5641 10217 5675 10251
rect 6101 10217 6135 10251
rect 6561 10217 6595 10251
rect 9873 10217 9907 10251
rect 10425 10217 10459 10251
rect 10885 10217 10919 10251
rect 11253 10217 11287 10251
rect 11713 10217 11747 10251
rect 12357 10217 12391 10251
rect 12909 10217 12943 10251
rect 13737 10217 13771 10251
rect 16589 10217 16623 10251
rect 17233 10217 17267 10251
rect 17601 10217 17635 10251
rect 17693 10217 17727 10251
rect 18061 10217 18095 10251
rect 4813 10149 4847 10183
rect 5733 10149 5767 10183
rect 7818 10149 7852 10183
rect 9965 10149 9999 10183
rect 2789 10081 2823 10115
rect 3985 10081 4019 10115
rect 6469 10081 6503 10115
rect 6929 10081 6963 10115
rect 7573 10081 7607 10115
rect 10793 10081 10827 10115
rect 11621 10081 11655 10115
rect 12817 10081 12851 10115
rect 15209 10081 15243 10115
rect 15476 10081 15510 10115
rect 18153 10081 18187 10115
rect 1777 10013 1811 10047
rect 2973 10013 3007 10047
rect 5089 10013 5123 10047
rect 5917 10013 5951 10047
rect 6653 10013 6687 10047
rect 9781 10013 9815 10047
rect 11069 10013 11103 10047
rect 11805 10013 11839 10047
rect 13093 10013 13127 10047
rect 16957 10013 16991 10047
rect 17141 10013 17175 10047
rect 18245 10013 18279 10047
rect 2329 9945 2363 9979
rect 13369 9945 13403 9979
rect 1409 9877 1443 9911
rect 3249 9877 3283 9911
rect 4445 9877 4479 9911
rect 7297 9877 7331 9911
rect 8953 9877 8987 9911
rect 10333 9877 10367 9911
rect 12081 9877 12115 9911
rect 12449 9877 12483 9911
rect 13553 9877 13587 9911
rect 16773 9877 16807 9911
rect 5457 9673 5491 9707
rect 8861 9673 8895 9707
rect 8953 9673 8987 9707
rect 9137 9673 9171 9707
rect 7389 9605 7423 9639
rect 3433 9537 3467 9571
rect 4261 9537 4295 9571
rect 6101 9537 6135 9571
rect 7021 9537 7055 9571
rect 1777 9469 1811 9503
rect 2321 9469 2355 9503
rect 2421 9469 2455 9503
rect 4077 9469 4111 9503
rect 4721 9469 4755 9503
rect 1501 9401 1535 9435
rect 2697 9401 2731 9435
rect 3249 9401 3283 9435
rect 5825 9401 5859 9435
rect 6837 9401 6871 9435
rect 7481 9401 7515 9435
rect 15669 9605 15703 9639
rect 15853 9605 15887 9639
rect 9689 9537 9723 9571
rect 10425 9537 10459 9571
rect 10517 9537 10551 9571
rect 11069 9537 11103 9571
rect 12081 9537 12115 9571
rect 12357 9537 12391 9571
rect 13093 9537 13127 9571
rect 16497 9537 16531 9571
rect 17601 9537 17635 9571
rect 9505 9469 9539 9503
rect 10333 9469 10367 9503
rect 12909 9469 12943 9503
rect 15137 9469 15171 9503
rect 15393 9469 15427 9503
rect 13277 9401 13311 9435
rect 13553 9401 13587 9435
rect 16313 9401 16347 9435
rect 17325 9401 17359 9435
rect 17877 9401 17911 9435
rect 18061 9401 18095 9435
rect 18245 9401 18279 9435
rect 18429 9401 18463 9435
rect 1593 9333 1627 9367
rect 1961 9333 1995 9367
rect 2145 9333 2179 9367
rect 2605 9333 2639 9367
rect 2881 9333 2915 9367
rect 3341 9333 3375 9367
rect 3709 9333 3743 9367
rect 4169 9333 4203 9367
rect 4537 9333 4571 9367
rect 4905 9333 4939 9367
rect 5917 9333 5951 9367
rect 6469 9333 6503 9367
rect 6929 9333 6963 9367
rect 8861 9333 8895 9367
rect 9597 9333 9631 9367
rect 9965 9333 9999 9367
rect 11161 9333 11195 9367
rect 12449 9333 12483 9367
rect 12817 9333 12851 9367
rect 14013 9333 14047 9367
rect 15945 9333 15979 9367
rect 16405 9333 16439 9367
rect 16957 9333 16991 9367
rect 17417 9333 17451 9367
rect 3249 9129 3283 9163
rect 3617 9129 3651 9163
rect 5825 9129 5859 9163
rect 10057 9129 10091 9163
rect 10977 9129 11011 9163
rect 11989 9129 12023 9163
rect 12449 9129 12483 9163
rect 13001 9129 13035 9163
rect 13093 9129 13127 9163
rect 15577 9129 15611 9163
rect 16221 9129 16255 9163
rect 16589 9129 16623 9163
rect 17049 9129 17083 9163
rect 17417 9129 17451 9163
rect 5641 9061 5675 9095
rect 6285 9061 6319 9095
rect 6653 9061 6687 9095
rect 7564 9061 7598 9095
rect 8769 9061 8803 9095
rect 12357 9061 12391 9095
rect 1409 8993 1443 9027
rect 2125 8993 2159 9027
rect 6193 8993 6227 9027
rect 7297 8993 7331 9027
rect 1869 8925 1903 8959
rect 3433 8925 3467 8959
rect 6469 8925 6503 8959
rect 9597 8993 9631 9027
rect 10425 8993 10459 9027
rect 10517 8993 10551 9027
rect 12817 8993 12851 9027
rect 8953 8925 8987 8959
rect 9689 8925 9723 8959
rect 9873 8925 9907 8959
rect 10609 8925 10643 8959
rect 12541 8925 12575 8959
rect 3985 8857 4019 8891
rect 8769 8857 8803 8891
rect 13645 9061 13679 9095
rect 16129 9061 16163 9095
rect 13553 8993 13587 9027
rect 15485 8993 15519 9027
rect 17877 8993 17911 9027
rect 18429 8993 18463 9027
rect 13737 8925 13771 8959
rect 15669 8925 15703 8959
rect 16681 8925 16715 8959
rect 16865 8925 16899 8959
rect 17509 8925 17543 8959
rect 17601 8925 17635 8959
rect 18245 8925 18279 8959
rect 13185 8857 13219 8891
rect 14105 8857 14139 8891
rect 15025 8857 15059 8891
rect 1593 8789 1627 8823
rect 8677 8789 8711 8823
rect 9229 8789 9263 8823
rect 11069 8789 11103 8823
rect 13093 8789 13127 8823
rect 15117 8789 15151 8823
rect 18061 8789 18095 8823
rect 3341 8585 3375 8619
rect 3525 8585 3559 8619
rect 16037 8585 16071 8619
rect 16589 8585 16623 8619
rect 17049 8585 17083 8619
rect 2973 8517 3007 8551
rect 2881 8381 2915 8415
rect 2636 8313 2670 8347
rect 3157 8313 3191 8347
rect 6101 8517 6135 8551
rect 6469 8517 6503 8551
rect 8033 8517 8067 8551
rect 9965 8517 9999 8551
rect 11529 8517 11563 8551
rect 16313 8517 16347 8551
rect 5825 8449 5859 8483
rect 7849 8449 7883 8483
rect 9045 8449 9079 8483
rect 9137 8449 9171 8483
rect 13737 8449 13771 8483
rect 14657 8449 14691 8483
rect 16129 8449 16163 8483
rect 17601 8449 17635 8483
rect 4741 8381 4775 8415
rect 4997 8381 5031 8415
rect 6285 8381 6319 8415
rect 8953 8381 8987 8415
rect 10149 8381 10183 8415
rect 11713 8381 11747 8415
rect 11969 8381 12003 8415
rect 17417 8381 17451 8415
rect 17877 8381 17911 8415
rect 18337 8381 18371 8415
rect 5549 8313 5583 8347
rect 7582 8313 7616 8347
rect 10394 8313 10428 8347
rect 13645 8313 13679 8347
rect 14013 8313 14047 8347
rect 14924 8313 14958 8347
rect 16773 8313 16807 8347
rect 17509 8313 17543 8347
rect 18521 8313 18555 8347
rect 1501 8245 1535 8279
rect 3341 8245 3375 8279
rect 3617 8245 3651 8279
rect 5181 8245 5215 8279
rect 5641 8245 5675 8279
rect 8585 8245 8619 8279
rect 13093 8245 13127 8279
rect 13185 8245 13219 8279
rect 13553 8245 13587 8279
rect 18061 8245 18095 8279
rect 1869 8041 1903 8075
rect 2513 8041 2547 8075
rect 2973 8041 3007 8075
rect 3433 8041 3467 8075
rect 4261 8041 4295 8075
rect 5181 8041 5215 8075
rect 5733 8041 5767 8075
rect 6561 8041 6595 8075
rect 6929 8041 6963 8075
rect 7757 8041 7791 8075
rect 8217 8041 8251 8075
rect 8677 8041 8711 8075
rect 16313 8041 16347 8075
rect 16773 8041 16807 8075
rect 16957 8041 16991 8075
rect 17141 8041 17175 8075
rect 17509 8041 17543 8075
rect 1593 7973 1627 8007
rect 6193 7973 6227 8007
rect 7021 7973 7055 8007
rect 7849 7973 7883 8007
rect 12112 7973 12146 8007
rect 13001 7973 13035 8007
rect 14013 7973 14047 8007
rect 14841 7973 14875 8007
rect 18337 7973 18371 8007
rect 1961 7905 1995 7939
rect 3341 7905 3375 7939
rect 4353 7905 4387 7939
rect 6101 7905 6135 7939
rect 8585 7905 8619 7939
rect 9137 7905 9171 7939
rect 13461 7905 13495 7939
rect 14933 7905 14967 7939
rect 15200 7905 15234 7939
rect 17601 7905 17635 7939
rect 18153 7905 18187 7939
rect 2605 7837 2639 7871
rect 2697 7837 2731 7871
rect 3617 7837 3651 7871
rect 4537 7837 4571 7871
rect 5273 7837 5307 7871
rect 5457 7837 5491 7871
rect 6285 7837 6319 7871
rect 7113 7837 7147 7871
rect 8033 7837 8067 7871
rect 8769 7837 8803 7871
rect 12357 7837 12391 7871
rect 13277 7837 13311 7871
rect 13369 7837 13403 7871
rect 17693 7837 17727 7871
rect 3893 7769 3927 7803
rect 10425 7769 10459 7803
rect 12817 7769 12851 7803
rect 18521 7769 18555 7803
rect 1501 7701 1535 7735
rect 2145 7701 2179 7735
rect 4813 7701 4847 7735
rect 7389 7701 7423 7735
rect 10977 7701 11011 7735
rect 13829 7701 13863 7735
rect 16497 7701 16531 7735
rect 16681 7701 16715 7735
rect 17969 7701 18003 7735
rect 3157 7497 3191 7531
rect 3985 7497 4019 7531
rect 5089 7497 5123 7531
rect 6469 7497 6503 7531
rect 11897 7497 11931 7531
rect 2881 7429 2915 7463
rect 3893 7429 3927 7463
rect 5641 7429 5675 7463
rect 6285 7429 6319 7463
rect 10057 7429 10091 7463
rect 10149 7429 10183 7463
rect 12173 7429 12207 7463
rect 15853 7429 15887 7463
rect 17509 7429 17543 7463
rect 2145 7361 2179 7395
rect 3525 7361 3559 7395
rect 4813 7361 4847 7395
rect 5365 7361 5399 7395
rect 7113 7361 7147 7395
rect 8401 7361 8435 7395
rect 12817 7361 12851 7395
rect 13553 7361 13587 7395
rect 13645 7361 13679 7395
rect 16405 7361 16439 7395
rect 18153 7361 18187 7395
rect 1409 7293 1443 7327
rect 1961 7293 1995 7327
rect 2421 7293 2455 7327
rect 3065 7293 3099 7327
rect 3341 7293 3375 7327
rect 4629 7293 4663 7327
rect 4721 7293 4755 7327
rect 6009 7293 6043 7327
rect 7573 7293 7607 7327
rect 8677 7293 8711 7327
rect 11529 7293 11563 7327
rect 11713 7293 11747 7327
rect 12633 7293 12667 7327
rect 12725 7293 12759 7327
rect 14289 7293 14323 7327
rect 16681 7293 16715 7327
rect 17325 7293 17359 7327
rect 17601 7293 17635 7327
rect 17969 7293 18003 7327
rect 1593 7225 1627 7259
rect 2329 7225 2363 7259
rect 6837 7225 6871 7259
rect 8922 7225 8956 7259
rect 11262 7225 11296 7259
rect 13461 7225 13495 7259
rect 14556 7225 14590 7259
rect 16221 7225 16255 7259
rect 18337 7225 18371 7259
rect 18521 7225 18555 7259
rect 1777 7157 1811 7191
rect 2789 7157 2823 7191
rect 4261 7157 4295 7191
rect 6929 7157 6963 7191
rect 7389 7157 7423 7191
rect 7757 7157 7791 7191
rect 8125 7157 8159 7191
rect 8217 7157 8251 7191
rect 12265 7157 12299 7191
rect 13093 7157 13127 7191
rect 13921 7157 13955 7191
rect 15669 7157 15703 7191
rect 16313 7157 16347 7191
rect 17141 7157 17175 7191
rect 17785 7157 17819 7191
rect 3525 6953 3559 6987
rect 5733 6953 5767 6987
rect 7757 6953 7791 6987
rect 8125 6953 8159 6987
rect 11989 6953 12023 6987
rect 12817 6953 12851 6987
rect 13645 6953 13679 6987
rect 15761 6953 15795 6987
rect 16405 6953 16439 6987
rect 16865 6953 16899 6987
rect 17601 6953 17635 6987
rect 3341 6885 3375 6919
rect 7665 6885 7699 6919
rect 8493 6885 8527 6919
rect 11161 6885 11195 6919
rect 12909 6885 12943 6919
rect 16037 6885 16071 6919
rect 1593 6817 1627 6851
rect 1777 6817 1811 6851
rect 1961 6817 1995 6851
rect 2329 6817 2363 6851
rect 2605 6817 2639 6851
rect 2881 6817 2915 6851
rect 4609 6817 4643 6851
rect 7205 6817 7239 6851
rect 8585 6817 8619 6851
rect 8953 6817 8987 6851
rect 13737 6817 13771 6851
rect 14197 6817 14231 6851
rect 14648 6817 14682 6851
rect 15853 6817 15887 6851
rect 16773 6817 16807 6851
rect 18337 6817 18371 6851
rect 4353 6749 4387 6783
rect 6377 6749 6411 6783
rect 7941 6749 7975 6783
rect 8769 6749 8803 6783
rect 2145 6681 2179 6715
rect 2973 6681 3007 6715
rect 9137 6749 9171 6783
rect 10977 6749 11011 6783
rect 11069 6749 11103 6783
rect 12081 6749 12115 6783
rect 12173 6749 12207 6783
rect 13001 6749 13035 6783
rect 13829 6749 13863 6783
rect 14381 6749 14415 6783
rect 17049 6749 17083 6783
rect 17693 6749 17727 6783
rect 17785 6749 17819 6783
rect 12449 6681 12483 6715
rect 13277 6681 13311 6715
rect 17233 6681 17267 6715
rect 18521 6681 18555 6715
rect 1501 6613 1535 6647
rect 2421 6613 2455 6647
rect 2697 6613 2731 6647
rect 3249 6613 3283 6647
rect 7297 6613 7331 6647
rect 8953 6613 8987 6647
rect 9505 6613 9539 6647
rect 11529 6613 11563 6647
rect 11621 6613 11655 6647
rect 16313 6613 16347 6647
rect 18061 6613 18095 6647
rect 3525 6409 3559 6443
rect 8033 6409 8067 6443
rect 14749 6409 14783 6443
rect 16405 6409 16439 6443
rect 17141 6409 17175 6443
rect 17509 6409 17543 6443
rect 5273 6341 5307 6375
rect 9229 6341 9263 6375
rect 10701 6341 10735 6375
rect 3433 6273 3467 6307
rect 6101 6273 6135 6307
rect 7021 6273 7055 6307
rect 8677 6273 8711 6307
rect 15393 6273 15427 6307
rect 16129 6273 16163 6307
rect 16957 6341 16991 6375
rect 16681 6273 16715 6307
rect 1961 6205 1995 6239
rect 3177 6205 3211 6239
rect 4898 6205 4932 6239
rect 5825 6205 5859 6239
rect 6837 6205 6871 6239
rect 6929 6205 6963 6239
rect 7297 6205 7331 6239
rect 8401 6205 8435 6239
rect 10342 6205 10376 6239
rect 10609 6205 10643 6239
rect 10885 6205 10919 6239
rect 11713 6205 11747 6239
rect 13185 6205 13219 6239
rect 15117 6205 15151 6239
rect 16405 6205 16439 6239
rect 17325 6205 17359 6239
rect 17601 6205 17635 6239
rect 17877 6205 17911 6239
rect 1593 6137 1627 6171
rect 4638 6137 4672 6171
rect 11958 6137 11992 6171
rect 13430 6137 13464 6171
rect 18337 6137 18371 6171
rect 18521 6137 18555 6171
rect 1501 6069 1535 6103
rect 1777 6069 1811 6103
rect 2053 6069 2087 6103
rect 5457 6069 5491 6103
rect 5917 6069 5951 6103
rect 6469 6069 6503 6103
rect 8493 6069 8527 6103
rect 8861 6069 8895 6103
rect 13093 6069 13127 6103
rect 14565 6069 14599 6103
rect 15209 6069 15243 6103
rect 15577 6069 15611 6103
rect 15945 6069 15979 6103
rect 16037 6069 16071 6103
rect 16497 6069 16531 6103
rect 17785 6069 17819 6103
rect 18061 6069 18095 6103
rect 1777 5865 1811 5899
rect 2513 5865 2547 5899
rect 2697 5865 2731 5899
rect 3341 5865 3375 5899
rect 3893 5865 3927 5899
rect 4261 5865 4295 5899
rect 5181 5865 5215 5899
rect 6377 5865 6411 5899
rect 11897 5865 11931 5899
rect 13185 5865 13219 5899
rect 15853 5865 15887 5899
rect 18061 5865 18095 5899
rect 1593 5797 1627 5831
rect 2421 5797 2455 5831
rect 1961 5729 1995 5763
rect 2237 5729 2271 5763
rect 2789 5797 2823 5831
rect 5089 5797 5123 5831
rect 4353 5729 4387 5763
rect 6009 5729 6043 5763
rect 7389 5729 7423 5763
rect 9137 5729 9171 5763
rect 12357 5729 12391 5763
rect 3433 5661 3467 5695
rect 3525 5661 3559 5695
rect 4537 5661 4571 5695
rect 5273 5661 5307 5695
rect 11989 5661 12023 5695
rect 12173 5661 12207 5695
rect 2697 5593 2731 5627
rect 6929 5593 6963 5627
rect 12541 5593 12575 5627
rect 17141 5797 17175 5831
rect 18337 5797 18371 5831
rect 13277 5729 13311 5763
rect 14105 5729 14139 5763
rect 14648 5729 14682 5763
rect 16221 5729 16255 5763
rect 16313 5729 16347 5763
rect 17049 5729 17083 5763
rect 17601 5729 17635 5763
rect 17877 5729 17911 5763
rect 14381 5661 14415 5695
rect 16405 5661 16439 5695
rect 17233 5661 17267 5695
rect 15761 5593 15795 5627
rect 18521 5593 18555 5627
rect 1501 5525 1535 5559
rect 2053 5525 2087 5559
rect 2973 5525 3007 5559
rect 4721 5525 4755 5559
rect 6193 5525 6227 5559
rect 7297 5525 7331 5559
rect 9321 5525 9355 5559
rect 9597 5525 9631 5559
rect 11529 5525 11563 5559
rect 13185 5525 13219 5559
rect 16681 5525 16715 5559
rect 17785 5525 17819 5559
rect 2881 5321 2915 5355
rect 3709 5321 3743 5355
rect 4905 5321 4939 5355
rect 9413 5321 9447 5355
rect 10885 5321 10919 5355
rect 11253 5321 11287 5355
rect 14565 5321 14599 5355
rect 14841 5321 14875 5355
rect 15025 5321 15059 5355
rect 15669 5321 15703 5355
rect 16037 5321 16071 5355
rect 2421 5253 2455 5287
rect 2789 5253 2823 5287
rect 12449 5253 12483 5287
rect 15301 5253 15335 5287
rect 3341 5185 3375 5219
rect 3525 5185 3559 5219
rect 4353 5185 4387 5219
rect 1409 5117 1443 5151
rect 1593 5117 1627 5151
rect 2329 5117 2363 5151
rect 2605 5117 2639 5151
rect 3249 5117 3283 5151
rect 6285 5117 6319 5151
rect 7593 5117 7627 5151
rect 7849 5117 7883 5151
rect 8033 5117 8067 5151
rect 9505 5117 9539 5151
rect 9761 5117 9795 5151
rect 10977 5117 11011 5151
rect 14013 5185 14047 5219
rect 15945 5185 15979 5219
rect 16589 5185 16623 5219
rect 17509 5185 17543 5219
rect 18521 5185 18555 5219
rect 12668 5117 12702 5151
rect 13829 5117 13863 5151
rect 14473 5117 14507 5151
rect 16405 5117 16439 5151
rect 17417 5117 17451 5151
rect 17877 5117 17911 5151
rect 18337 5117 18371 5151
rect 1961 5049 1995 5083
rect 4077 5049 4111 5083
rect 6018 5049 6052 5083
rect 8300 5049 8334 5083
rect 12449 5049 12483 5083
rect 15485 5049 15519 5083
rect 17325 5049 17359 5083
rect 1869 4981 1903 5015
rect 2145 4981 2179 5015
rect 4169 4981 4203 5015
rect 6469 4981 6503 5015
rect 11437 4981 11471 5015
rect 12771 4981 12805 5015
rect 14105 4981 14139 5015
rect 15117 4981 15151 5015
rect 16497 4981 16531 5015
rect 16957 4981 16991 5015
rect 18061 4981 18095 5015
rect 2329 4777 2363 4811
rect 2881 4777 2915 4811
rect 3985 4777 4019 4811
rect 4169 4777 4203 4811
rect 4537 4777 4571 4811
rect 4997 4777 5031 4811
rect 5365 4777 5399 4811
rect 6653 4777 6687 4811
rect 6929 4777 6963 4811
rect 16681 4777 16715 4811
rect 17049 4777 17083 4811
rect 1593 4709 1627 4743
rect 3065 4709 3099 4743
rect 11446 4709 11480 4743
rect 12173 4709 12207 4743
rect 12265 4709 12299 4743
rect 12817 4709 12851 4743
rect 13277 4709 13311 4743
rect 15945 4709 15979 4743
rect 17969 4709 18003 4743
rect 18337 4709 18371 4743
rect 1409 4641 1443 4675
rect 2237 4641 2271 4675
rect 2513 4641 2547 4675
rect 4629 4641 4663 4675
rect 6193 4641 6227 4675
rect 11713 4641 11747 4675
rect 14048 4641 14082 4675
rect 14381 4641 14415 4675
rect 15234 4641 15268 4675
rect 15577 4641 15611 4675
rect 15853 4641 15887 4675
rect 16129 4641 16163 4675
rect 16405 4641 16439 4675
rect 17601 4641 17635 4675
rect 18153 4641 18187 4675
rect 2053 4573 2087 4607
rect 2605 4573 2639 4607
rect 4813 4573 4847 4607
rect 5457 4573 5491 4607
rect 5641 4573 5675 4607
rect 6285 4573 6319 4607
rect 6469 4573 6503 4607
rect 13185 4573 13219 4607
rect 13553 4573 13587 4607
rect 14565 4573 14599 4607
rect 15025 4573 15059 4607
rect 17141 4573 17175 4607
rect 17233 4573 17267 4607
rect 5825 4505 5859 4539
rect 15669 4505 15703 4539
rect 16313 4505 16347 4539
rect 18521 4505 18555 4539
rect 10333 4437 10367 4471
rect 13001 4437 13035 4471
rect 14151 4437 14185 4471
rect 15163 4437 15197 4471
rect 15393 4437 15427 4471
rect 16589 4437 16623 4471
rect 17785 4437 17819 4471
rect 3341 4233 3375 4267
rect 5273 4233 5307 4267
rect 5733 4233 5767 4267
rect 6745 4233 6779 4267
rect 8769 4233 8803 4267
rect 8953 4233 8987 4267
rect 9689 4233 9723 4267
rect 3157 4165 3191 4199
rect 5365 4165 5399 4199
rect 15577 4165 15611 4199
rect 17417 4165 17451 4199
rect 5825 4097 5859 4131
rect 7389 4097 7423 4131
rect 9321 4097 9355 4131
rect 12357 4097 12391 4131
rect 14841 4097 14875 4131
rect 15025 4097 15059 4131
rect 1593 4029 1627 4063
rect 2697 4029 2731 4063
rect 2973 4029 3007 4063
rect 3893 4029 3927 4063
rect 6653 4029 6687 4063
rect 8861 4029 8895 4063
rect 9505 4029 9539 4063
rect 11529 4029 11563 4063
rect 13277 4029 13311 4063
rect 13553 4029 13587 4063
rect 13829 4029 13863 4063
rect 15761 4029 15795 4063
rect 15945 4029 15979 4063
rect 16589 4029 16623 4063
rect 16957 4029 16991 4063
rect 17233 4029 17267 4063
rect 17969 4029 18003 4063
rect 18337 4029 18371 4063
rect 1961 3961 1995 3995
rect 2329 3961 2363 3995
rect 4160 3961 4194 3995
rect 7656 3961 7690 3995
rect 11262 3961 11296 3995
rect 12449 3961 12483 3995
rect 13001 3961 13035 3995
rect 14197 3961 14231 3995
rect 14289 3961 14323 3995
rect 15117 3961 15151 3995
rect 17601 3961 17635 3995
rect 18153 3961 18187 3995
rect 18521 3961 18555 3995
rect 1501 3893 1535 3927
rect 1869 3893 1903 3927
rect 2237 3893 2271 3927
rect 2513 3893 2547 3927
rect 2789 3893 2823 3927
rect 3525 3893 3559 3927
rect 7113 3893 7147 3927
rect 10149 3893 10183 3927
rect 11713 3893 11747 3927
rect 11897 3893 11931 3927
rect 13093 3893 13127 3927
rect 13369 3893 13403 3927
rect 14013 3893 14047 3927
rect 16405 3893 16439 3927
rect 16773 3893 16807 3927
rect 17141 3893 17175 3927
rect 17693 3893 17727 3927
rect 2513 3689 2547 3723
rect 2789 3689 2823 3723
rect 8033 3689 8067 3723
rect 10241 3689 10275 3723
rect 10793 3689 10827 3723
rect 13461 3689 13495 3723
rect 14013 3689 14047 3723
rect 14933 3689 14967 3723
rect 15209 3689 15243 3723
rect 15761 3689 15795 3723
rect 2329 3621 2363 3655
rect 6898 3621 6932 3655
rect 12909 3621 12943 3655
rect 13001 3621 13035 3655
rect 16865 3621 16899 3655
rect 17233 3621 17267 3655
rect 17969 3621 18003 3655
rect 18337 3621 18371 3655
rect 1593 3553 1627 3587
rect 1961 3553 1995 3587
rect 2697 3553 2731 3587
rect 2973 3553 3007 3587
rect 3065 3553 3099 3587
rect 3525 3553 3559 3587
rect 3985 3553 4019 3587
rect 5448 3553 5482 3587
rect 8309 3553 8343 3587
rect 8528 3553 8562 3587
rect 10057 3553 10091 3587
rect 10241 3553 10275 3587
rect 10333 3553 10367 3587
rect 10885 3553 10919 3587
rect 11196 3553 11230 3587
rect 11621 3553 11655 3587
rect 11713 3553 11747 3587
rect 13220 3553 13254 3587
rect 13645 3553 13679 3587
rect 13921 3553 13955 3587
rect 14197 3553 14231 3587
rect 14508 3553 14542 3587
rect 14749 3553 14783 3587
rect 15025 3553 15059 3587
rect 15301 3553 15335 3587
rect 15577 3553 15611 3587
rect 15945 3553 15979 3587
rect 16221 3553 16255 3587
rect 16497 3553 16531 3587
rect 17601 3553 17635 3587
rect 5181 3485 5215 3519
rect 6653 3485 6687 3519
rect 11299 3485 11333 3519
rect 11989 3485 12023 3519
rect 14611 3485 14645 3519
rect 17049 3485 17083 3519
rect 3249 3417 3283 3451
rect 6561 3417 6595 3451
rect 11437 3417 11471 3451
rect 16129 3417 16163 3451
rect 17417 3417 17451 3451
rect 18153 3417 18187 3451
rect 1501 3349 1535 3383
rect 1869 3349 1903 3383
rect 2237 3349 2271 3383
rect 3341 3349 3375 3383
rect 3709 3349 3743 3383
rect 8125 3349 8159 3383
rect 8631 3349 8665 3383
rect 9873 3349 9907 3383
rect 10425 3349 10459 3383
rect 11069 3349 11103 3383
rect 11897 3349 11931 3383
rect 13323 3349 13357 3383
rect 13737 3349 13771 3383
rect 15485 3349 15519 3383
rect 16405 3349 16439 3383
rect 16681 3349 16715 3383
rect 17693 3349 17727 3383
rect 18429 3349 18463 3383
rect 2789 3145 2823 3179
rect 4629 3145 4663 3179
rect 7113 3145 7147 3179
rect 7757 3145 7791 3179
rect 10517 3145 10551 3179
rect 12679 3145 12713 3179
rect 12955 3145 12989 3179
rect 14933 3145 14967 3179
rect 16405 3145 16439 3179
rect 17049 3145 17083 3179
rect 18429 3145 18463 3179
rect 4261 3077 4295 3111
rect 6745 3077 6779 3111
rect 9137 3077 9171 3111
rect 15945 3077 15979 3111
rect 8585 3009 8619 3043
rect 10333 3009 10367 3043
rect 11805 3009 11839 3043
rect 13185 3009 13219 3043
rect 14289 3009 14323 3043
rect 15393 3009 15427 3043
rect 15577 3009 15611 3043
rect 15761 3009 15795 3043
rect 1593 2941 1627 2975
rect 1961 2941 1995 2975
rect 2697 2941 2731 2975
rect 2973 2941 3007 2975
rect 3249 2941 3283 2975
rect 3525 2941 3559 2975
rect 3801 2941 3835 2975
rect 4077 2941 4111 2975
rect 4353 2941 4387 2975
rect 4813 2941 4847 2975
rect 4905 2941 4939 2975
rect 6561 2941 6595 2975
rect 7389 2941 7423 2975
rect 7481 2941 7515 2975
rect 8309 2941 8343 2975
rect 9505 2941 9539 2975
rect 9873 2941 9907 2975
rect 10057 2941 10091 2975
rect 10793 2941 10827 2975
rect 10885 2941 10919 2975
rect 11069 2941 11103 2975
rect 12608 2941 12642 2975
rect 12852 2941 12886 2975
rect 14473 2941 14507 2975
rect 15117 2941 15151 2975
rect 16589 2941 16623 2975
rect 17141 2941 17175 2975
rect 17325 2941 17359 2975
rect 17601 2941 17635 2975
rect 17969 2941 18003 2975
rect 18337 2941 18371 2975
rect 1777 2873 1811 2907
rect 2329 2873 2363 2907
rect 8677 2873 8711 2907
rect 9689 2873 9723 2907
rect 11437 2873 11471 2907
rect 11897 2873 11931 2907
rect 12449 2873 12483 2907
rect 13277 2873 13311 2907
rect 14197 2873 14231 2907
rect 16773 2873 16807 2907
rect 17785 2873 17819 2907
rect 1501 2805 1535 2839
rect 2237 2805 2271 2839
rect 2513 2805 2547 2839
rect 3065 2805 3099 2839
rect 3341 2805 3375 2839
rect 3617 2805 3651 2839
rect 3893 2805 3927 2839
rect 4537 2805 4571 2839
rect 6929 2805 6963 2839
rect 7941 2805 7975 2839
rect 8125 2805 8159 2839
rect 9321 2805 9355 2839
rect 10241 2805 10275 2839
rect 11345 2805 11379 2839
rect 15301 2805 15335 2839
rect 18061 2805 18095 2839
rect 4721 2601 4755 2635
rect 5917 2601 5951 2635
rect 6377 2601 6411 2635
rect 14749 2601 14783 2635
rect 17417 2601 17451 2635
rect 1593 2533 1627 2567
rect 1961 2533 1995 2567
rect 2605 2533 2639 2567
rect 4077 2533 4111 2567
rect 4445 2533 4479 2567
rect 4813 2533 4847 2567
rect 5181 2533 5215 2567
rect 6745 2533 6779 2567
rect 7113 2533 7147 2567
rect 7481 2533 7515 2567
rect 7849 2533 7883 2567
rect 8309 2533 8343 2567
rect 9229 2533 9263 2567
rect 10149 2533 10183 2567
rect 10517 2533 10551 2567
rect 10609 2533 10643 2567
rect 11437 2533 11471 2567
rect 12081 2533 12115 2567
rect 13185 2533 13219 2567
rect 13277 2533 13311 2567
rect 14197 2533 14231 2567
rect 14933 2533 14967 2567
rect 15301 2533 15335 2567
rect 15393 2533 15427 2567
rect 16313 2533 16347 2567
rect 16589 2533 16623 2567
rect 16957 2533 16991 2567
rect 17601 2533 17635 2567
rect 18337 2533 18371 2567
rect 2329 2465 2363 2499
rect 2881 2465 2915 2499
rect 3341 2465 3375 2499
rect 3709 2465 3743 2499
rect 5549 2465 5583 2499
rect 5733 2465 5767 2499
rect 6009 2465 6043 2499
rect 6193 2465 6227 2499
rect 8861 2465 8895 2499
rect 14565 2465 14599 2499
rect 17233 2465 17267 2499
rect 17969 2465 18003 2499
rect 2145 2397 2179 2431
rect 4997 2397 5031 2431
rect 6929 2397 6963 2431
rect 10241 2397 10275 2431
rect 11989 2397 12023 2431
rect 12633 2397 12667 2431
rect 15117 2397 15151 2431
rect 1409 2329 1443 2363
rect 2697 2329 2731 2363
rect 3157 2329 3191 2363
rect 3893 2329 3927 2363
rect 4261 2329 4295 2363
rect 5365 2329 5399 2363
rect 6561 2329 6595 2363
rect 7297 2329 7331 2363
rect 7665 2329 7699 2363
rect 8125 2329 8159 2363
rect 8677 2329 8711 2363
rect 11069 2329 11103 2363
rect 16405 2329 16439 2363
rect 17785 2329 17819 2363
rect 18521 2329 18555 2363
rect 1869 2261 1903 2295
rect 3525 2261 3559 2295
rect 11345 2261 11379 2295
rect 14289 2261 14323 2295
rect 16865 2261 16899 2295
rect 18061 2261 18095 2295
<< metal1 >>
rect 290 15104 296 15156
rect 348 15144 354 15156
rect 3234 15144 3240 15156
rect 348 15116 3240 15144
rect 348 15104 354 15116
rect 3234 15104 3240 15116
rect 3292 15104 3298 15156
rect 8202 15104 8208 15156
rect 8260 15144 8266 15156
rect 15381 15147 15439 15153
rect 15381 15144 15393 15147
rect 8260 15116 15393 15144
rect 8260 15104 8266 15116
rect 15381 15113 15393 15116
rect 15427 15113 15439 15147
rect 15381 15107 15439 15113
rect 2682 15036 2688 15088
rect 2740 15076 2746 15088
rect 4246 15076 4252 15088
rect 2740 15048 4252 15076
rect 2740 15036 2746 15048
rect 4246 15036 4252 15048
rect 4304 15036 4310 15088
rect 4982 15036 4988 15088
rect 5040 15076 5046 15088
rect 15010 15076 15016 15088
rect 5040 15048 15016 15076
rect 5040 15036 5046 15048
rect 15010 15036 15016 15048
rect 15068 15036 15074 15088
rect 1578 14968 1584 15020
rect 1636 15008 1642 15020
rect 4522 15008 4528 15020
rect 1636 14980 4528 15008
rect 1636 14968 1642 14980
rect 4522 14968 4528 14980
rect 4580 14968 4586 15020
rect 10870 14968 10876 15020
rect 10928 15008 10934 15020
rect 18969 15011 19027 15017
rect 18969 15008 18981 15011
rect 10928 14980 18981 15008
rect 10928 14968 10934 14980
rect 18969 14977 18981 14980
rect 19015 14977 19027 15011
rect 18969 14971 19027 14977
rect 4706 14900 4712 14952
rect 4764 14940 4770 14952
rect 12710 14940 12716 14952
rect 4764 14912 12716 14940
rect 4764 14900 4770 14912
rect 12710 14900 12716 14912
rect 12768 14900 12774 14952
rect 13262 14900 13268 14952
rect 13320 14940 13326 14952
rect 15286 14940 15292 14952
rect 13320 14912 15292 14940
rect 13320 14900 13326 14912
rect 15286 14900 15292 14912
rect 15344 14900 15350 14952
rect 15381 14943 15439 14949
rect 15381 14909 15393 14943
rect 15427 14940 15439 14943
rect 17218 14940 17224 14952
rect 15427 14912 17224 14940
rect 15427 14909 15439 14912
rect 15381 14903 15439 14909
rect 17218 14900 17224 14912
rect 17276 14900 17282 14952
rect 1946 14832 1952 14884
rect 2004 14872 2010 14884
rect 7650 14872 7656 14884
rect 2004 14844 7656 14872
rect 2004 14832 2010 14844
rect 7650 14832 7656 14844
rect 7708 14832 7714 14884
rect 13538 14832 13544 14884
rect 13596 14872 13602 14884
rect 17678 14872 17684 14884
rect 13596 14844 17684 14872
rect 13596 14832 13602 14844
rect 17678 14832 17684 14844
rect 17736 14832 17742 14884
rect 13998 14764 14004 14816
rect 14056 14804 14062 14816
rect 17034 14804 17040 14816
rect 14056 14776 17040 14804
rect 14056 14764 14062 14776
rect 17034 14764 17040 14776
rect 17092 14764 17098 14816
rect 1104 14714 18860 14736
rect 1104 14662 6912 14714
rect 6964 14662 6976 14714
rect 7028 14662 7040 14714
rect 7092 14662 7104 14714
rect 7156 14662 12843 14714
rect 12895 14662 12907 14714
rect 12959 14662 12971 14714
rect 13023 14662 13035 14714
rect 13087 14662 18860 14714
rect 1104 14640 18860 14662
rect 1578 14600 1584 14612
rect 1539 14572 1584 14600
rect 1578 14560 1584 14572
rect 1636 14560 1642 14612
rect 1946 14600 1952 14612
rect 1907 14572 1952 14600
rect 1946 14560 1952 14572
rect 2004 14560 2010 14612
rect 2682 14600 2688 14612
rect 2643 14572 2688 14600
rect 2682 14560 2688 14572
rect 2740 14560 2746 14612
rect 4617 14603 4675 14609
rect 4617 14600 4629 14603
rect 3068 14572 4629 14600
rect 1854 14532 1860 14544
rect 1815 14504 1860 14532
rect 1854 14492 1860 14504
rect 1912 14492 1918 14544
rect 2225 14535 2283 14541
rect 2225 14501 2237 14535
rect 2271 14532 2283 14535
rect 2774 14532 2780 14544
rect 2271 14504 2780 14532
rect 2271 14501 2283 14504
rect 2225 14495 2283 14501
rect 2774 14492 2780 14504
rect 2832 14532 2838 14544
rect 3068 14532 3096 14572
rect 4617 14569 4629 14572
rect 4663 14569 4675 14603
rect 4617 14563 4675 14569
rect 8662 14560 8668 14612
rect 8720 14600 8726 14612
rect 8941 14603 8999 14609
rect 8941 14600 8953 14603
rect 8720 14572 8953 14600
rect 8720 14560 8726 14572
rect 3234 14532 3240 14544
rect 2832 14504 3096 14532
rect 3195 14504 3240 14532
rect 2832 14492 2838 14504
rect 3234 14492 3240 14504
rect 3292 14492 3298 14544
rect 3510 14492 3516 14544
rect 3568 14532 3574 14544
rect 3881 14535 3939 14541
rect 3881 14532 3893 14535
rect 3568 14504 3893 14532
rect 3568 14492 3574 14504
rect 3881 14501 3893 14504
rect 3927 14501 3939 14535
rect 3881 14495 3939 14501
rect 4154 14492 4160 14544
rect 4212 14532 4218 14544
rect 4249 14535 4307 14541
rect 4249 14532 4261 14535
rect 4212 14504 4261 14532
rect 4212 14492 4218 14504
rect 4249 14501 4261 14504
rect 4295 14501 4307 14535
rect 4798 14532 4804 14544
rect 4759 14504 4804 14532
rect 4249 14495 4307 14501
rect 4798 14492 4804 14504
rect 4856 14492 4862 14544
rect 4982 14532 4988 14544
rect 4943 14504 4988 14532
rect 4982 14492 4988 14504
rect 5040 14492 5046 14544
rect 5442 14532 5448 14544
rect 5403 14504 5448 14532
rect 5442 14492 5448 14504
rect 5500 14492 5506 14544
rect 6730 14532 6736 14544
rect 6691 14504 6736 14532
rect 6730 14492 6736 14504
rect 6788 14492 6794 14544
rect 7374 14492 7380 14544
rect 7432 14532 7438 14544
rect 7561 14535 7619 14541
rect 7561 14532 7573 14535
rect 7432 14504 7573 14532
rect 7432 14492 7438 14504
rect 7561 14501 7573 14504
rect 7607 14532 7619 14535
rect 7745 14535 7803 14541
rect 7745 14532 7757 14535
rect 7607 14504 7757 14532
rect 7607 14501 7619 14504
rect 7561 14495 7619 14501
rect 7745 14501 7757 14504
rect 7791 14501 7803 14535
rect 7745 14495 7803 14501
rect 1486 14464 1492 14476
rect 1447 14436 1492 14464
rect 1486 14424 1492 14436
rect 1544 14424 1550 14476
rect 2590 14464 2596 14476
rect 2551 14436 2596 14464
rect 2590 14424 2596 14436
rect 2648 14424 2654 14476
rect 3053 14467 3111 14473
rect 3053 14433 3065 14467
rect 3099 14464 3111 14467
rect 3142 14464 3148 14476
rect 3099 14436 3148 14464
rect 3099 14433 3111 14436
rect 3053 14427 3111 14433
rect 3142 14424 3148 14436
rect 3200 14424 3206 14476
rect 3418 14464 3424 14476
rect 3379 14436 3424 14464
rect 3418 14424 3424 14436
rect 3476 14424 3482 14476
rect 3602 14464 3608 14476
rect 3563 14436 3608 14464
rect 3602 14424 3608 14436
rect 3660 14424 3666 14476
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14433 4123 14467
rect 4065 14427 4123 14433
rect 4433 14467 4491 14473
rect 4433 14433 4445 14467
rect 4479 14464 4491 14467
rect 5534 14464 5540 14476
rect 4479 14436 5540 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 2409 14331 2467 14337
rect 2409 14297 2421 14331
rect 2455 14328 2467 14331
rect 2774 14328 2780 14340
rect 2455 14300 2780 14328
rect 2455 14297 2467 14300
rect 2409 14291 2467 14297
rect 2774 14288 2780 14300
rect 2832 14288 2838 14340
rect 3694 14328 3700 14340
rect 2884 14300 3700 14328
rect 2590 14220 2596 14272
rect 2648 14260 2654 14272
rect 2884 14260 2912 14300
rect 3694 14288 3700 14300
rect 3752 14288 3758 14340
rect 4080 14328 4108 14427
rect 5534 14424 5540 14436
rect 5592 14424 5598 14476
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14433 5687 14467
rect 5629 14427 5687 14433
rect 5644 14396 5672 14427
rect 5718 14424 5724 14476
rect 5776 14464 5782 14476
rect 5997 14467 6055 14473
rect 5997 14464 6009 14467
rect 5776 14436 6009 14464
rect 5776 14424 5782 14436
rect 5997 14433 6009 14436
rect 6043 14433 6055 14467
rect 5997 14427 6055 14433
rect 6086 14424 6092 14476
rect 6144 14464 6150 14476
rect 6365 14467 6423 14473
rect 6365 14464 6377 14467
rect 6144 14436 6377 14464
rect 6144 14424 6150 14436
rect 6365 14433 6377 14436
rect 6411 14464 6423 14467
rect 6549 14467 6607 14473
rect 6549 14464 6561 14467
rect 6411 14436 6561 14464
rect 6411 14433 6423 14436
rect 6365 14427 6423 14433
rect 6549 14433 6561 14436
rect 6595 14433 6607 14467
rect 6549 14427 6607 14433
rect 6638 14424 6644 14476
rect 6696 14464 6702 14476
rect 8864 14473 8892 14572
rect 8941 14569 8953 14572
rect 8987 14569 8999 14603
rect 8941 14563 8999 14569
rect 10137 14603 10195 14609
rect 10137 14569 10149 14603
rect 10183 14600 10195 14603
rect 11146 14600 11152 14612
rect 10183 14572 11152 14600
rect 10183 14569 10195 14572
rect 10137 14563 10195 14569
rect 11146 14560 11152 14572
rect 11204 14560 11210 14612
rect 11425 14603 11483 14609
rect 11425 14569 11437 14603
rect 11471 14569 11483 14603
rect 13262 14600 13268 14612
rect 13223 14572 13268 14600
rect 11425 14563 11483 14569
rect 11440 14532 11468 14563
rect 13262 14560 13268 14572
rect 13320 14560 13326 14612
rect 13538 14600 13544 14612
rect 13499 14572 13544 14600
rect 13538 14560 13544 14572
rect 13596 14560 13602 14612
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 14921 14603 14979 14609
rect 14921 14600 14933 14603
rect 13872 14572 14933 14600
rect 13872 14560 13878 14572
rect 14921 14569 14933 14572
rect 14967 14600 14979 14603
rect 17218 14600 17224 14612
rect 14967 14572 15516 14600
rect 17179 14572 17224 14600
rect 14967 14569 14979 14572
rect 14921 14563 14979 14569
rect 11606 14532 11612 14544
rect 11440 14504 11612 14532
rect 11606 14492 11612 14504
rect 11664 14492 11670 14544
rect 12434 14492 12440 14544
rect 12492 14532 12498 14544
rect 12710 14532 12716 14544
rect 12492 14504 12716 14532
rect 12492 14492 12498 14504
rect 12710 14492 12716 14504
rect 12768 14532 12774 14544
rect 13449 14535 13507 14541
rect 13449 14532 13461 14535
rect 12768 14504 13461 14532
rect 12768 14492 12774 14504
rect 13280 14476 13308 14504
rect 13449 14501 13461 14504
rect 13495 14501 13507 14535
rect 13998 14532 14004 14544
rect 13959 14504 14004 14532
rect 13449 14495 13507 14501
rect 13998 14492 14004 14504
rect 14056 14492 14062 14544
rect 14458 14492 14464 14544
rect 14516 14532 14522 14544
rect 14553 14535 14611 14541
rect 14553 14532 14565 14535
rect 14516 14504 14565 14532
rect 14516 14492 14522 14504
rect 14553 14501 14565 14504
rect 14599 14501 14611 14535
rect 15102 14532 15108 14544
rect 15063 14504 15108 14532
rect 14553 14495 14611 14501
rect 15102 14492 15108 14504
rect 15160 14492 15166 14544
rect 6917 14467 6975 14473
rect 6917 14464 6929 14467
rect 6696 14436 6929 14464
rect 6696 14424 6702 14436
rect 6917 14433 6929 14436
rect 6963 14433 6975 14467
rect 6917 14427 6975 14433
rect 8849 14467 8907 14473
rect 8849 14433 8861 14467
rect 8895 14433 8907 14467
rect 9306 14464 9312 14476
rect 9267 14436 9312 14464
rect 8849 14427 8907 14433
rect 9306 14424 9312 14436
rect 9364 14464 9370 14476
rect 9585 14467 9643 14473
rect 9585 14464 9597 14467
rect 9364 14436 9597 14464
rect 9364 14424 9370 14436
rect 9585 14433 9597 14436
rect 9631 14433 9643 14467
rect 9950 14464 9956 14476
rect 9911 14436 9956 14464
rect 9585 14427 9643 14433
rect 9950 14424 9956 14436
rect 10008 14464 10014 14476
rect 10229 14467 10287 14473
rect 10229 14464 10241 14467
rect 10008 14436 10241 14464
rect 10008 14424 10014 14436
rect 10229 14433 10241 14436
rect 10275 14433 10287 14467
rect 10594 14464 10600 14476
rect 10555 14436 10600 14464
rect 10229 14427 10287 14433
rect 10594 14424 10600 14436
rect 10652 14464 10658 14476
rect 10873 14467 10931 14473
rect 10873 14464 10885 14467
rect 10652 14436 10885 14464
rect 10652 14424 10658 14436
rect 10873 14433 10885 14436
rect 10919 14433 10931 14467
rect 11238 14464 11244 14476
rect 11199 14436 11244 14464
rect 10873 14427 10931 14433
rect 11238 14424 11244 14436
rect 11296 14464 11302 14476
rect 11517 14467 11575 14473
rect 11517 14464 11529 14467
rect 11296 14436 11529 14464
rect 11296 14424 11302 14436
rect 11517 14433 11529 14436
rect 11563 14433 11575 14467
rect 11882 14464 11888 14476
rect 11843 14436 11888 14464
rect 11517 14427 11575 14433
rect 11882 14424 11888 14436
rect 11940 14464 11946 14476
rect 12161 14467 12219 14473
rect 12161 14464 12173 14467
rect 11940 14436 12173 14464
rect 11940 14424 11946 14436
rect 12161 14433 12173 14436
rect 12207 14433 12219 14467
rect 12526 14464 12532 14476
rect 12487 14436 12532 14464
rect 12161 14427 12219 14433
rect 12526 14424 12532 14436
rect 12584 14464 12590 14476
rect 12805 14467 12863 14473
rect 12805 14464 12817 14467
rect 12584 14436 12817 14464
rect 12584 14424 12590 14436
rect 12805 14433 12817 14436
rect 12851 14433 12863 14467
rect 12805 14427 12863 14433
rect 13081 14467 13139 14473
rect 13081 14433 13093 14467
rect 13127 14464 13139 14467
rect 13170 14464 13176 14476
rect 13127 14436 13176 14464
rect 13127 14433 13139 14436
rect 13081 14427 13139 14433
rect 13170 14424 13176 14436
rect 13228 14424 13234 14476
rect 13262 14424 13268 14476
rect 13320 14424 13326 14476
rect 13814 14464 13820 14476
rect 13775 14436 13820 14464
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 14182 14464 14188 14476
rect 14143 14436 14188 14464
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 14274 14424 14280 14476
rect 14332 14464 14338 14476
rect 14737 14467 14795 14473
rect 14737 14464 14749 14467
rect 14332 14436 14749 14464
rect 14332 14424 14338 14436
rect 14737 14433 14749 14436
rect 14783 14433 14795 14467
rect 14737 14427 14795 14433
rect 14826 14424 14832 14476
rect 14884 14464 14890 14476
rect 15488 14473 15516 14572
rect 17218 14560 17224 14572
rect 17276 14560 17282 14612
rect 15746 14532 15752 14544
rect 15707 14504 15752 14532
rect 15746 14492 15752 14504
rect 15804 14492 15810 14544
rect 16114 14492 16120 14544
rect 16172 14532 16178 14544
rect 16761 14535 16819 14541
rect 16761 14532 16773 14535
rect 16172 14504 16773 14532
rect 16172 14492 16178 14504
rect 16761 14501 16773 14504
rect 16807 14501 16819 14535
rect 16942 14532 16948 14544
rect 16903 14504 16948 14532
rect 16761 14495 16819 14501
rect 16942 14492 16948 14504
rect 17000 14492 17006 14544
rect 17681 14535 17739 14541
rect 17681 14501 17693 14535
rect 17727 14532 17739 14535
rect 17770 14532 17776 14544
rect 17727 14504 17776 14532
rect 17727 14501 17739 14504
rect 17681 14495 17739 14501
rect 17770 14492 17776 14504
rect 17828 14492 17834 14544
rect 17862 14492 17868 14544
rect 17920 14532 17926 14544
rect 18049 14535 18107 14541
rect 18049 14532 18061 14535
rect 17920 14504 18061 14532
rect 17920 14492 17926 14504
rect 18049 14501 18061 14504
rect 18095 14501 18107 14535
rect 18049 14495 18107 14501
rect 15289 14467 15347 14473
rect 15289 14464 15301 14467
rect 14884 14436 15301 14464
rect 14884 14424 14890 14436
rect 15289 14433 15301 14436
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 15473 14467 15531 14473
rect 15473 14433 15485 14467
rect 15519 14433 15531 14467
rect 15473 14427 15531 14433
rect 15562 14424 15568 14476
rect 15620 14464 15626 14476
rect 15933 14467 15991 14473
rect 15933 14464 15945 14467
rect 15620 14436 15945 14464
rect 15620 14424 15626 14436
rect 15933 14433 15945 14436
rect 15979 14433 15991 14467
rect 15933 14427 15991 14433
rect 16574 14424 16580 14476
rect 16632 14464 16638 14476
rect 17402 14464 17408 14476
rect 16632 14436 16677 14464
rect 17363 14436 17408 14464
rect 16632 14424 16638 14436
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 18414 14464 18420 14476
rect 18375 14436 18420 14464
rect 18414 14424 18420 14436
rect 18472 14424 18478 14476
rect 15378 14396 15384 14408
rect 5644 14368 15384 14396
rect 15378 14356 15384 14368
rect 15436 14356 15442 14408
rect 16301 14399 16359 14405
rect 16301 14365 16313 14399
rect 16347 14396 16359 14399
rect 18432 14396 18460 14424
rect 16347 14368 18460 14396
rect 16347 14365 16359 14368
rect 16301 14359 16359 14365
rect 9493 14331 9551 14337
rect 4080 14300 9444 14328
rect 2648 14232 2912 14260
rect 2961 14263 3019 14269
rect 2648 14220 2654 14232
rect 2961 14229 2973 14263
rect 3007 14260 3019 14263
rect 3510 14260 3516 14272
rect 3007 14232 3516 14260
rect 3007 14229 3019 14232
rect 2961 14223 3019 14229
rect 3510 14220 3516 14232
rect 3568 14220 3574 14272
rect 5902 14260 5908 14272
rect 5863 14232 5908 14260
rect 5902 14220 5908 14232
rect 5960 14220 5966 14272
rect 5994 14220 6000 14272
rect 6052 14260 6058 14272
rect 6181 14263 6239 14269
rect 6181 14260 6193 14263
rect 6052 14232 6193 14260
rect 6052 14220 6058 14232
rect 6181 14229 6193 14232
rect 6227 14229 6239 14263
rect 6181 14223 6239 14229
rect 7469 14263 7527 14269
rect 7469 14229 7481 14263
rect 7515 14260 7527 14263
rect 8018 14260 8024 14272
rect 7515 14232 8024 14260
rect 7515 14229 7527 14232
rect 7469 14223 7527 14229
rect 8018 14220 8024 14232
rect 8076 14220 8082 14272
rect 8478 14220 8484 14272
rect 8536 14260 8542 14272
rect 8665 14263 8723 14269
rect 8665 14260 8677 14263
rect 8536 14232 8677 14260
rect 8536 14220 8542 14232
rect 8665 14229 8677 14232
rect 8711 14229 8723 14263
rect 9416 14260 9444 14300
rect 9493 14297 9505 14331
rect 9539 14328 9551 14331
rect 10502 14328 10508 14340
rect 9539 14300 10508 14328
rect 9539 14297 9551 14300
rect 9493 14291 9551 14297
rect 10502 14288 10508 14300
rect 10560 14288 10566 14340
rect 10612 14300 11284 14328
rect 10612 14260 10640 14300
rect 10778 14260 10784 14272
rect 9416 14232 10640 14260
rect 10739 14232 10784 14260
rect 8665 14223 8723 14229
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 11256 14260 11284 14300
rect 11330 14288 11336 14340
rect 11388 14328 11394 14340
rect 12069 14331 12127 14337
rect 12069 14328 12081 14331
rect 11388 14300 12081 14328
rect 11388 14288 11394 14300
rect 12069 14297 12081 14300
rect 12115 14297 12127 14331
rect 13446 14328 13452 14340
rect 12069 14291 12127 14297
rect 12406 14300 13452 14328
rect 12406 14260 12434 14300
rect 13446 14288 13452 14300
rect 13504 14288 13510 14340
rect 13630 14288 13636 14340
rect 13688 14328 13694 14340
rect 14274 14328 14280 14340
rect 13688 14300 14280 14328
rect 13688 14288 13694 14300
rect 14274 14288 14280 14300
rect 14332 14288 14338 14340
rect 14369 14331 14427 14337
rect 14369 14297 14381 14331
rect 14415 14328 14427 14331
rect 16390 14328 16396 14340
rect 14415 14300 16396 14328
rect 14415 14297 14427 14300
rect 14369 14291 14427 14297
rect 16390 14288 16396 14300
rect 16448 14288 16454 14340
rect 16758 14288 16764 14340
rect 16816 14328 16822 14340
rect 17865 14331 17923 14337
rect 17865 14328 17877 14331
rect 16816 14300 17877 14328
rect 16816 14288 16822 14300
rect 17865 14297 17877 14300
rect 17911 14297 17923 14331
rect 17865 14291 17923 14297
rect 18138 14288 18144 14340
rect 18196 14328 18202 14340
rect 18233 14331 18291 14337
rect 18233 14328 18245 14331
rect 18196 14300 18245 14328
rect 18196 14288 18202 14300
rect 18233 14297 18245 14300
rect 18279 14297 18291 14331
rect 18233 14291 18291 14297
rect 11256 14232 12434 14260
rect 12713 14263 12771 14269
rect 12713 14229 12725 14263
rect 12759 14260 12771 14263
rect 14458 14260 14464 14272
rect 12759 14232 14464 14260
rect 12759 14229 12771 14232
rect 12713 14223 12771 14229
rect 14458 14220 14464 14232
rect 14516 14220 14522 14272
rect 15470 14220 15476 14272
rect 15528 14260 15534 14272
rect 15657 14263 15715 14269
rect 15657 14260 15669 14263
rect 15528 14232 15669 14260
rect 15528 14220 15534 14232
rect 15657 14229 15669 14232
rect 15703 14229 15715 14263
rect 15657 14223 15715 14229
rect 16485 14263 16543 14269
rect 16485 14229 16497 14263
rect 16531 14260 16543 14263
rect 17310 14260 17316 14272
rect 16531 14232 17316 14260
rect 16531 14229 16543 14232
rect 16485 14223 16543 14229
rect 17310 14220 17316 14232
rect 17368 14220 17374 14272
rect 17589 14263 17647 14269
rect 17589 14229 17601 14263
rect 17635 14260 17647 14263
rect 17770 14260 17776 14272
rect 17635 14232 17776 14260
rect 17635 14229 17647 14232
rect 17589 14223 17647 14229
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 1104 14170 18860 14192
rect 1104 14118 3947 14170
rect 3999 14118 4011 14170
rect 4063 14118 4075 14170
rect 4127 14118 4139 14170
rect 4191 14118 9878 14170
rect 9930 14118 9942 14170
rect 9994 14118 10006 14170
rect 10058 14118 10070 14170
rect 10122 14118 15808 14170
rect 15860 14118 15872 14170
rect 15924 14118 15936 14170
rect 15988 14118 16000 14170
rect 16052 14118 18860 14170
rect 1104 14096 18860 14118
rect 1949 14059 2007 14065
rect 1949 14025 1961 14059
rect 1995 14056 2007 14059
rect 3418 14056 3424 14068
rect 1995 14028 3424 14056
rect 1995 14025 2007 14028
rect 1949 14019 2007 14025
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 3694 14016 3700 14068
rect 3752 14056 3758 14068
rect 4065 14059 4123 14065
rect 4065 14056 4077 14059
rect 3752 14028 4077 14056
rect 3752 14016 3758 14028
rect 4065 14025 4077 14028
rect 4111 14025 4123 14059
rect 4706 14056 4712 14068
rect 4667 14028 4712 14056
rect 4065 14019 4123 14025
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 6638 14056 6644 14068
rect 5592 14028 6132 14056
rect 6599 14028 6644 14056
rect 5592 14016 5598 14028
rect 2222 13988 2228 14000
rect 2183 13960 2228 13988
rect 2222 13948 2228 13960
rect 2280 13948 2286 14000
rect 2593 13991 2651 13997
rect 2593 13988 2605 13991
rect 2332 13960 2605 13988
rect 2332 13920 2360 13960
rect 2593 13957 2605 13960
rect 2639 13957 2651 13991
rect 2866 13988 2872 14000
rect 2827 13960 2872 13988
rect 2593 13951 2651 13957
rect 2866 13948 2872 13960
rect 2924 13948 2930 14000
rect 3237 13991 3295 13997
rect 3237 13988 3249 13991
rect 2976 13960 3249 13988
rect 2976 13920 3004 13960
rect 3237 13957 3249 13960
rect 3283 13957 3295 13991
rect 3237 13951 3295 13957
rect 3513 13991 3571 13997
rect 3513 13957 3525 13991
rect 3559 13957 3571 13991
rect 3513 13951 3571 13957
rect 3973 13991 4031 13997
rect 3973 13957 3985 13991
rect 4019 13988 4031 13991
rect 5810 13988 5816 14000
rect 4019 13960 5816 13988
rect 4019 13957 4031 13960
rect 3973 13951 4031 13957
rect 3528 13920 3556 13951
rect 5810 13948 5816 13960
rect 5868 13948 5874 14000
rect 4338 13920 4344 13932
rect 1596 13892 2360 13920
rect 2424 13892 3004 13920
rect 3037 13892 3556 13920
rect 3712 13892 4344 13920
rect 1596 13861 1624 13892
rect 2424 13861 2452 13892
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13821 1455 13855
rect 1397 13815 1455 13821
rect 1581 13855 1639 13861
rect 1581 13821 1593 13855
rect 1627 13821 1639 13855
rect 1581 13815 1639 13821
rect 1765 13855 1823 13861
rect 1765 13821 1777 13855
rect 1811 13852 1823 13855
rect 2409 13855 2467 13861
rect 1811 13824 2360 13852
rect 1811 13821 1823 13824
rect 1765 13815 1823 13821
rect 934 13744 940 13796
rect 992 13784 998 13796
rect 1412 13784 1440 13815
rect 992 13756 1440 13784
rect 992 13744 998 13756
rect 1486 13744 1492 13796
rect 1544 13784 1550 13796
rect 2041 13787 2099 13793
rect 2041 13784 2053 13787
rect 1544 13756 2053 13784
rect 1544 13744 1550 13756
rect 2041 13753 2053 13756
rect 2087 13753 2099 13787
rect 2332 13784 2360 13824
rect 2409 13821 2421 13855
rect 2455 13821 2467 13855
rect 2409 13815 2467 13821
rect 2777 13855 2835 13861
rect 2777 13821 2789 13855
rect 2823 13852 2835 13855
rect 2866 13852 2872 13864
rect 2823 13824 2872 13852
rect 2823 13821 2835 13824
rect 2777 13815 2835 13821
rect 2866 13812 2872 13824
rect 2924 13812 2930 13864
rect 3037 13861 3065 13892
rect 3037 13855 3111 13861
rect 3037 13824 3065 13855
rect 3053 13821 3065 13824
rect 3099 13821 3111 13855
rect 3053 13815 3111 13821
rect 3418 13812 3424 13864
rect 3476 13852 3482 13864
rect 3712 13861 3740 13892
rect 4338 13880 4344 13892
rect 4396 13880 4402 13932
rect 6104 13920 6132 14028
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 13170 14016 13176 14068
rect 13228 14056 13234 14068
rect 13725 14059 13783 14065
rect 13725 14056 13737 14059
rect 13228 14028 13737 14056
rect 13228 14016 13234 14028
rect 13725 14025 13737 14028
rect 13771 14025 13783 14059
rect 13725 14019 13783 14025
rect 14182 14016 14188 14068
rect 14240 14056 14246 14068
rect 14240 14028 14504 14056
rect 14240 14016 14246 14028
rect 6181 13991 6239 13997
rect 6181 13957 6193 13991
rect 6227 13988 6239 13991
rect 6730 13988 6736 14000
rect 6227 13960 6736 13988
rect 6227 13957 6239 13960
rect 6181 13951 6239 13957
rect 6730 13948 6736 13960
rect 6788 13948 6794 14000
rect 11146 13948 11152 14000
rect 11204 13988 11210 14000
rect 11790 13988 11796 14000
rect 11204 13960 11796 13988
rect 11204 13948 11210 13960
rect 11790 13948 11796 13960
rect 11848 13948 11854 14000
rect 13262 13988 13268 14000
rect 13223 13960 13268 13988
rect 13262 13948 13268 13960
rect 13320 13948 13326 14000
rect 13446 13988 13452 14000
rect 13407 13960 13452 13988
rect 13446 13948 13452 13960
rect 13504 13948 13510 14000
rect 14369 13991 14427 13997
rect 14369 13957 14381 13991
rect 14415 13957 14427 13991
rect 14476 13988 14504 14028
rect 15010 14016 15016 14068
rect 15068 14056 15074 14068
rect 15105 14059 15163 14065
rect 15105 14056 15117 14059
rect 15068 14028 15117 14056
rect 15068 14016 15074 14028
rect 15105 14025 15117 14028
rect 15151 14025 15163 14059
rect 15105 14019 15163 14025
rect 15378 14016 15384 14068
rect 15436 14056 15442 14068
rect 15565 14059 15623 14065
rect 15565 14056 15577 14059
rect 15436 14028 15577 14056
rect 15436 14016 15442 14028
rect 15565 14025 15577 14028
rect 15611 14025 15623 14059
rect 15565 14019 15623 14025
rect 16574 14016 16580 14068
rect 16632 14056 16638 14068
rect 16761 14059 16819 14065
rect 16632 14028 16677 14056
rect 16632 14016 16638 14028
rect 16761 14025 16773 14059
rect 16807 14056 16819 14059
rect 16942 14056 16948 14068
rect 16807 14028 16948 14056
rect 16807 14025 16819 14028
rect 16761 14019 16819 14025
rect 16942 14016 16948 14028
rect 17000 14016 17006 14068
rect 17681 14059 17739 14065
rect 17681 14025 17693 14059
rect 17727 14056 17739 14059
rect 18322 14056 18328 14068
rect 17727 14028 18328 14056
rect 17727 14025 17739 14028
rect 17681 14019 17739 14025
rect 18322 14016 18328 14028
rect 18380 14016 18386 14068
rect 15746 13988 15752 14000
rect 14476 13960 15752 13988
rect 14369 13951 14427 13957
rect 14384 13920 14412 13951
rect 15746 13948 15752 13960
rect 15804 13948 15810 14000
rect 17865 13991 17923 13997
rect 17865 13988 17877 13991
rect 16546 13960 17877 13988
rect 16546 13920 16574 13960
rect 17865 13957 17877 13960
rect 17911 13957 17923 13991
rect 17865 13951 17923 13957
rect 18233 13991 18291 13997
rect 18233 13957 18245 13991
rect 18279 13988 18291 13991
rect 18969 13991 19027 13997
rect 18969 13988 18981 13991
rect 18279 13960 18981 13988
rect 18279 13957 18291 13960
rect 18233 13951 18291 13957
rect 18969 13957 18981 13960
rect 19015 13957 19027 13991
rect 18969 13951 19027 13957
rect 6104 13892 14412 13920
rect 14476 13892 16574 13920
rect 17037 13923 17095 13929
rect 3697 13855 3755 13861
rect 3476 13824 3521 13852
rect 3476 13812 3482 13824
rect 3697 13821 3709 13855
rect 3743 13821 3755 13855
rect 3697 13815 3755 13821
rect 3786 13812 3792 13864
rect 3844 13852 3850 13864
rect 4249 13855 4307 13861
rect 4249 13852 4261 13855
rect 3844 13824 4261 13852
rect 3844 13812 3850 13824
rect 4249 13821 4261 13824
rect 4295 13821 4307 13855
rect 4249 13815 4307 13821
rect 4525 13855 4583 13861
rect 4525 13821 4537 13855
rect 4571 13852 4583 13855
rect 4614 13852 4620 13864
rect 4571 13824 4620 13852
rect 4571 13821 4583 13824
rect 4525 13815 4583 13821
rect 4614 13812 4620 13824
rect 4672 13852 4678 13864
rect 4672 13824 5948 13852
rect 4672 13812 4678 13824
rect 3234 13784 3240 13796
rect 2332 13756 3240 13784
rect 2041 13747 2099 13753
rect 3234 13744 3240 13756
rect 3292 13744 3298 13796
rect 5920 13784 5948 13824
rect 5994 13812 6000 13864
rect 6052 13852 6058 13864
rect 6052 13824 6097 13852
rect 6052 13812 6058 13824
rect 6178 13812 6184 13864
rect 6236 13852 6242 13864
rect 6457 13855 6515 13861
rect 6457 13852 6469 13855
rect 6236 13824 6469 13852
rect 6236 13812 6242 13824
rect 6457 13821 6469 13824
rect 6503 13821 6515 13855
rect 9490 13852 9496 13864
rect 6457 13815 6515 13821
rect 6564 13824 9496 13852
rect 6564 13784 6592 13824
rect 9490 13812 9496 13824
rect 9548 13852 9554 13864
rect 9548 13824 11652 13852
rect 9548 13812 9554 13824
rect 5920 13756 6592 13784
rect 11624 13784 11652 13824
rect 11698 13812 11704 13864
rect 11756 13852 11762 13864
rect 13630 13852 13636 13864
rect 11756 13824 13492 13852
rect 13591 13824 13636 13852
rect 11756 13812 11762 13824
rect 13464 13784 13492 13824
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 14476 13852 14504 13892
rect 17037 13889 17049 13923
rect 17083 13920 17095 13923
rect 17083 13892 18460 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 18432 13864 18460 13892
rect 13740 13824 14504 13852
rect 14553 13855 14611 13861
rect 13740 13784 13768 13824
rect 14553 13821 14565 13855
rect 14599 13852 14611 13855
rect 14826 13852 14832 13864
rect 14599 13824 14832 13852
rect 14599 13821 14611 13824
rect 14553 13815 14611 13821
rect 14826 13812 14832 13824
rect 14884 13812 14890 13864
rect 15289 13855 15347 13861
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 15562 13852 15568 13864
rect 15335 13824 15568 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 15562 13812 15568 13824
rect 15620 13812 15626 13864
rect 15746 13852 15752 13864
rect 15659 13824 15752 13852
rect 15746 13812 15752 13824
rect 15804 13852 15810 13864
rect 16206 13852 16212 13864
rect 15804 13824 16212 13852
rect 15804 13812 15810 13824
rect 16206 13812 16212 13824
rect 16264 13812 16270 13864
rect 16390 13852 16396 13864
rect 16351 13824 16396 13852
rect 16390 13812 16396 13824
rect 16448 13852 16454 13864
rect 17221 13855 17279 13861
rect 17221 13852 17233 13855
rect 16448 13824 17233 13852
rect 16448 13812 16454 13824
rect 17221 13821 17233 13824
rect 17267 13821 17279 13855
rect 17221 13815 17279 13821
rect 17405 13855 17463 13861
rect 17405 13821 17417 13855
rect 17451 13852 17463 13855
rect 18414 13852 18420 13864
rect 17451 13824 18276 13852
rect 18375 13824 18420 13852
rect 17451 13821 17463 13824
rect 17405 13815 17463 13821
rect 11624 13756 12434 13784
rect 13464 13756 13768 13784
rect 1670 13676 1676 13728
rect 1728 13716 1734 13728
rect 5902 13716 5908 13728
rect 1728 13688 5908 13716
rect 1728 13676 1734 13688
rect 5902 13676 5908 13688
rect 5960 13676 5966 13728
rect 12406 13716 12434 13756
rect 17034 13744 17040 13796
rect 17092 13784 17098 13796
rect 17589 13787 17647 13793
rect 17589 13784 17601 13787
rect 17092 13756 17601 13784
rect 17092 13744 17098 13756
rect 17589 13753 17601 13756
rect 17635 13753 17647 13787
rect 18049 13787 18107 13793
rect 18049 13784 18061 13787
rect 17589 13747 17647 13753
rect 17880 13756 18061 13784
rect 13814 13716 13820 13728
rect 12406 13688 13820 13716
rect 13814 13676 13820 13688
rect 13872 13716 13878 13728
rect 13909 13719 13967 13725
rect 13909 13716 13921 13719
rect 13872 13688 13921 13716
rect 13872 13676 13878 13688
rect 13909 13685 13921 13688
rect 13955 13685 13967 13719
rect 13909 13679 13967 13685
rect 17494 13676 17500 13728
rect 17552 13716 17558 13728
rect 17880 13716 17908 13756
rect 18049 13753 18061 13756
rect 18095 13753 18107 13787
rect 18248 13784 18276 13824
rect 18414 13812 18420 13824
rect 18472 13812 18478 13864
rect 18966 13852 18972 13864
rect 18524 13824 18972 13852
rect 18524 13784 18552 13824
rect 18966 13812 18972 13824
rect 19024 13812 19030 13864
rect 18248 13756 18552 13784
rect 18049 13747 18107 13753
rect 17552 13688 17908 13716
rect 17552 13676 17558 13688
rect 1104 13626 18860 13648
rect 1104 13574 6912 13626
rect 6964 13574 6976 13626
rect 7028 13574 7040 13626
rect 7092 13574 7104 13626
rect 7156 13574 12843 13626
rect 12895 13574 12907 13626
rect 12959 13574 12971 13626
rect 13023 13574 13035 13626
rect 13087 13574 18860 13626
rect 1104 13552 18860 13574
rect 2590 13472 2596 13524
rect 2648 13512 2654 13524
rect 2648 13484 3096 13512
rect 2648 13472 2654 13484
rect 1854 13444 1860 13456
rect 1815 13416 1860 13444
rect 1854 13404 1860 13416
rect 1912 13444 1918 13456
rect 2961 13447 3019 13453
rect 2961 13444 2973 13447
rect 1912 13416 2973 13444
rect 1912 13404 1918 13416
rect 2961 13413 2973 13416
rect 3007 13413 3019 13447
rect 2961 13407 3019 13413
rect 1486 13376 1492 13388
rect 1447 13348 1492 13376
rect 1486 13336 1492 13348
rect 1544 13336 1550 13388
rect 2130 13376 2136 13388
rect 2091 13348 2136 13376
rect 2130 13336 2136 13348
rect 2188 13336 2194 13388
rect 2590 13376 2596 13388
rect 2551 13348 2596 13376
rect 2590 13336 2596 13348
rect 2648 13336 2654 13388
rect 2682 13336 2688 13388
rect 2740 13385 2746 13388
rect 2740 13376 2752 13385
rect 3068 13376 3096 13484
rect 3142 13472 3148 13524
rect 3200 13472 3206 13524
rect 3326 13512 3332 13524
rect 3287 13484 3332 13512
rect 3326 13472 3332 13484
rect 3384 13472 3390 13524
rect 17034 13512 17040 13524
rect 12406 13484 17040 13512
rect 3160 13444 3188 13472
rect 3513 13447 3571 13453
rect 3513 13444 3525 13447
rect 3160 13416 3525 13444
rect 3513 13413 3525 13416
rect 3559 13413 3571 13447
rect 3513 13407 3571 13413
rect 3878 13404 3884 13456
rect 3936 13444 3942 13456
rect 11054 13444 11060 13456
rect 3936 13416 11060 13444
rect 3936 13404 3942 13416
rect 11054 13404 11060 13416
rect 11112 13444 11118 13456
rect 12406 13444 12434 13484
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 17221 13515 17279 13521
rect 17221 13481 17233 13515
rect 17267 13512 17279 13515
rect 17494 13512 17500 13524
rect 17267 13484 17500 13512
rect 17267 13481 17279 13484
rect 17221 13475 17279 13481
rect 17494 13472 17500 13484
rect 17552 13472 17558 13524
rect 17589 13515 17647 13521
rect 17589 13481 17601 13515
rect 17635 13512 17647 13515
rect 17862 13512 17868 13524
rect 17635 13484 17868 13512
rect 17635 13481 17647 13484
rect 17589 13475 17647 13481
rect 17862 13472 17868 13484
rect 17920 13472 17926 13524
rect 11112 13416 12434 13444
rect 17405 13447 17463 13453
rect 11112 13404 11118 13416
rect 17405 13413 17417 13447
rect 17451 13444 17463 13447
rect 17678 13444 17684 13456
rect 17451 13416 17684 13444
rect 17451 13413 17463 13416
rect 17405 13407 17463 13413
rect 17678 13404 17684 13416
rect 17736 13404 17742 13456
rect 18141 13447 18199 13453
rect 18141 13413 18153 13447
rect 18187 13444 18199 13447
rect 19610 13444 19616 13456
rect 18187 13416 19616 13444
rect 18187 13413 18199 13416
rect 18141 13407 18199 13413
rect 19610 13404 19616 13416
rect 19668 13404 19674 13456
rect 3145 13379 3203 13385
rect 3145 13376 3157 13379
rect 2740 13348 2785 13376
rect 3068 13348 3157 13376
rect 2740 13339 2752 13348
rect 3145 13345 3157 13348
rect 3191 13345 3203 13379
rect 3145 13339 3203 13345
rect 16853 13379 16911 13385
rect 16853 13345 16865 13379
rect 16899 13376 16911 13379
rect 17957 13379 18015 13385
rect 17957 13376 17969 13379
rect 16899 13348 17969 13376
rect 16899 13345 16911 13348
rect 16853 13339 16911 13345
rect 17957 13345 17969 13348
rect 18003 13345 18015 13379
rect 18414 13376 18420 13388
rect 18375 13348 18420 13376
rect 17957 13339 18015 13345
rect 2740 13336 2746 13339
rect 3878 13308 3884 13320
rect 3839 13280 3884 13308
rect 3878 13268 3884 13280
rect 3936 13268 3942 13320
rect 5718 13308 5724 13320
rect 4172 13280 5724 13308
rect 1670 13240 1676 13252
rect 1631 13212 1676 13240
rect 1670 13200 1676 13212
rect 1728 13200 1734 13252
rect 2317 13243 2375 13249
rect 2317 13209 2329 13243
rect 2363 13240 2375 13243
rect 2869 13243 2927 13249
rect 2363 13212 2774 13240
rect 2363 13209 2375 13212
rect 2317 13203 2375 13209
rect 1946 13172 1952 13184
rect 1907 13144 1952 13172
rect 1946 13132 1952 13144
rect 2004 13132 2010 13184
rect 2222 13132 2228 13184
rect 2280 13172 2286 13184
rect 2409 13175 2467 13181
rect 2409 13172 2421 13175
rect 2280 13144 2421 13172
rect 2280 13132 2286 13144
rect 2409 13141 2421 13144
rect 2455 13141 2467 13175
rect 2746 13172 2774 13212
rect 2869 13209 2881 13243
rect 2915 13240 2927 13243
rect 3234 13240 3240 13252
rect 2915 13212 3240 13240
rect 2915 13209 2927 13212
rect 2869 13203 2927 13209
rect 3234 13200 3240 13212
rect 3292 13200 3298 13252
rect 4172 13240 4200 13280
rect 5718 13268 5724 13280
rect 5776 13268 5782 13320
rect 4338 13240 4344 13252
rect 3344 13212 4200 13240
rect 4251 13212 4344 13240
rect 3344 13172 3372 13212
rect 4338 13200 4344 13212
rect 4396 13240 4402 13252
rect 14550 13240 14556 13252
rect 4396 13212 14556 13240
rect 4396 13200 4402 13212
rect 14550 13200 14556 13212
rect 14608 13240 14614 13252
rect 16868 13240 16896 13339
rect 18414 13336 18420 13348
rect 18472 13336 18478 13388
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13308 17831 13311
rect 18432 13308 18460 13336
rect 17819 13280 18460 13308
rect 17819 13277 17831 13280
rect 17773 13271 17831 13277
rect 14608 13212 16896 13240
rect 14608 13200 14614 13212
rect 16942 13200 16948 13252
rect 17000 13240 17006 13252
rect 18233 13243 18291 13249
rect 18233 13240 18245 13243
rect 17000 13212 18245 13240
rect 17000 13200 17006 13212
rect 18233 13209 18245 13212
rect 18279 13209 18291 13243
rect 18233 13203 18291 13209
rect 2746 13144 3372 13172
rect 2409 13135 2467 13141
rect 3418 13132 3424 13184
rect 3476 13172 3482 13184
rect 4157 13175 4215 13181
rect 4157 13172 4169 13175
rect 3476 13144 4169 13172
rect 3476 13132 3482 13144
rect 4157 13141 4169 13144
rect 4203 13172 4215 13175
rect 14182 13172 14188 13184
rect 4203 13144 14188 13172
rect 4203 13141 4215 13144
rect 4157 13135 4215 13141
rect 14182 13132 14188 13144
rect 14240 13172 14246 13184
rect 16390 13172 16396 13184
rect 14240 13144 16396 13172
rect 14240 13132 14246 13144
rect 16390 13132 16396 13144
rect 16448 13132 16454 13184
rect 1104 13082 18860 13104
rect 1104 13030 3947 13082
rect 3999 13030 4011 13082
rect 4063 13030 4075 13082
rect 4127 13030 4139 13082
rect 4191 13030 9878 13082
rect 9930 13030 9942 13082
rect 9994 13030 10006 13082
rect 10058 13030 10070 13082
rect 10122 13030 15808 13082
rect 15860 13030 15872 13082
rect 15924 13030 15936 13082
rect 15988 13030 16000 13082
rect 16052 13030 18860 13082
rect 1104 13008 18860 13030
rect 2682 12928 2688 12980
rect 2740 12968 2746 12980
rect 2958 12968 2964 12980
rect 2740 12940 2964 12968
rect 2740 12928 2746 12940
rect 2958 12928 2964 12940
rect 3016 12928 3022 12980
rect 3234 12928 3240 12980
rect 3292 12968 3298 12980
rect 12066 12968 12072 12980
rect 3292 12940 12072 12968
rect 3292 12928 3298 12940
rect 12066 12928 12072 12940
rect 12124 12928 12130 12980
rect 17402 12928 17408 12980
rect 17460 12968 17466 12980
rect 17497 12971 17555 12977
rect 17497 12968 17509 12971
rect 17460 12940 17509 12968
rect 17460 12928 17466 12940
rect 17497 12937 17509 12940
rect 17543 12937 17555 12971
rect 17497 12931 17555 12937
rect 1578 12860 1584 12912
rect 1636 12900 1642 12912
rect 3513 12903 3571 12909
rect 3513 12900 3525 12903
rect 1636 12872 3525 12900
rect 1636 12860 1642 12872
rect 3513 12869 3525 12872
rect 3559 12869 3571 12903
rect 3513 12863 3571 12869
rect 1504 12804 2268 12832
rect 1504 12776 1532 12804
rect 1486 12764 1492 12776
rect 1399 12736 1492 12764
rect 1486 12724 1492 12736
rect 1544 12724 1550 12776
rect 1673 12767 1731 12773
rect 1673 12733 1685 12767
rect 1719 12764 1731 12767
rect 2038 12764 2044 12776
rect 1719 12736 2044 12764
rect 1719 12733 1731 12736
rect 1673 12727 1731 12733
rect 2038 12724 2044 12736
rect 2096 12724 2102 12776
rect 2240 12764 2268 12804
rect 2590 12792 2596 12844
rect 2648 12832 2654 12844
rect 2685 12835 2743 12841
rect 2685 12832 2697 12835
rect 2648 12804 2697 12832
rect 2648 12792 2654 12804
rect 2685 12801 2697 12804
rect 2731 12801 2743 12835
rect 2685 12795 2743 12801
rect 2866 12792 2872 12844
rect 2924 12832 2930 12844
rect 3786 12832 3792 12844
rect 2924 12804 3792 12832
rect 2924 12792 2930 12804
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 16850 12792 16856 12844
rect 16908 12832 16914 12844
rect 18233 12835 18291 12841
rect 18233 12832 18245 12835
rect 16908 12804 18245 12832
rect 16908 12792 16914 12804
rect 18233 12801 18245 12804
rect 18279 12801 18291 12835
rect 18233 12795 18291 12801
rect 3329 12767 3387 12773
rect 3329 12764 3341 12767
rect 2240 12736 3341 12764
rect 3329 12733 3341 12736
rect 3375 12733 3387 12767
rect 3329 12727 3387 12733
rect 17773 12767 17831 12773
rect 17773 12733 17785 12767
rect 17819 12764 17831 12767
rect 18414 12764 18420 12776
rect 17819 12736 18420 12764
rect 17819 12733 17831 12736
rect 17773 12727 17831 12733
rect 18414 12724 18420 12736
rect 18472 12724 18478 12776
rect 1578 12656 1584 12708
rect 1636 12696 1642 12708
rect 1857 12699 1915 12705
rect 1857 12696 1869 12699
rect 1636 12668 1869 12696
rect 1636 12656 1642 12668
rect 1857 12665 1869 12668
rect 1903 12665 1915 12699
rect 1857 12659 1915 12665
rect 2501 12699 2559 12705
rect 2501 12665 2513 12699
rect 2547 12696 2559 12699
rect 3050 12696 3056 12708
rect 2547 12668 3056 12696
rect 2547 12665 2559 12668
rect 2501 12659 2559 12665
rect 3050 12656 3056 12668
rect 3108 12656 3114 12708
rect 17405 12699 17463 12705
rect 17405 12665 17417 12699
rect 17451 12696 17463 12699
rect 18046 12696 18052 12708
rect 17451 12668 18052 12696
rect 17451 12665 17463 12668
rect 17405 12659 17463 12665
rect 18046 12656 18052 12668
rect 18104 12656 18110 12708
rect 1762 12588 1768 12640
rect 1820 12628 1826 12640
rect 1949 12631 2007 12637
rect 1949 12628 1961 12631
rect 1820 12600 1961 12628
rect 1820 12588 1826 12600
rect 1949 12597 1961 12600
rect 1995 12597 2007 12631
rect 2130 12628 2136 12640
rect 2091 12600 2136 12628
rect 1949 12591 2007 12597
rect 2130 12588 2136 12600
rect 2188 12588 2194 12640
rect 2593 12631 2651 12637
rect 2593 12597 2605 12631
rect 2639 12628 2651 12631
rect 2866 12628 2872 12640
rect 2639 12600 2872 12628
rect 2639 12597 2651 12600
rect 2593 12591 2651 12597
rect 2866 12588 2872 12600
rect 2924 12588 2930 12640
rect 3234 12628 3240 12640
rect 3195 12600 3240 12628
rect 3234 12588 3240 12600
rect 3292 12588 3298 12640
rect 3786 12628 3792 12640
rect 3747 12600 3792 12628
rect 3786 12588 3792 12600
rect 3844 12588 3850 12640
rect 17494 12588 17500 12640
rect 17552 12628 17558 12640
rect 17957 12631 18015 12637
rect 17957 12628 17969 12631
rect 17552 12600 17969 12628
rect 17552 12588 17558 12600
rect 17957 12597 17969 12600
rect 18003 12597 18015 12631
rect 17957 12591 18015 12597
rect 1104 12538 18860 12560
rect 1104 12486 6912 12538
rect 6964 12486 6976 12538
rect 7028 12486 7040 12538
rect 7092 12486 7104 12538
rect 7156 12486 12843 12538
rect 12895 12486 12907 12538
rect 12959 12486 12971 12538
rect 13023 12486 13035 12538
rect 13087 12486 18860 12538
rect 1104 12464 18860 12486
rect 3050 12424 3056 12436
rect 3011 12396 3056 12424
rect 3050 12384 3056 12396
rect 3108 12384 3114 12436
rect 2682 12356 2688 12368
rect 2595 12328 2688 12356
rect 2682 12316 2688 12328
rect 2740 12356 2746 12368
rect 4157 12359 4215 12365
rect 4157 12356 4169 12359
rect 2740 12328 4169 12356
rect 2740 12316 2746 12328
rect 4157 12325 4169 12328
rect 4203 12356 4215 12359
rect 10870 12356 10876 12368
rect 4203 12328 10876 12356
rect 4203 12325 4215 12328
rect 4157 12319 4215 12325
rect 10870 12316 10876 12328
rect 10928 12316 10934 12368
rect 1394 12248 1400 12300
rect 1452 12288 1458 12300
rect 1489 12291 1547 12297
rect 1489 12288 1501 12291
rect 1452 12260 1501 12288
rect 1452 12248 1458 12260
rect 1489 12257 1501 12260
rect 1535 12257 1547 12291
rect 1854 12288 1860 12300
rect 1815 12260 1860 12288
rect 1489 12251 1547 12257
rect 1504 12220 1532 12251
rect 1854 12248 1860 12260
rect 1912 12248 1918 12300
rect 2593 12291 2651 12297
rect 2593 12257 2605 12291
rect 2639 12288 2651 12291
rect 3418 12288 3424 12300
rect 2639 12260 3424 12288
rect 2639 12257 2651 12260
rect 2593 12251 2651 12257
rect 3418 12248 3424 12260
rect 3476 12248 3482 12300
rect 4614 12248 4620 12300
rect 4672 12288 4678 12300
rect 4781 12291 4839 12297
rect 4781 12288 4793 12291
rect 4672 12260 4793 12288
rect 4672 12248 4678 12260
rect 4781 12257 4793 12260
rect 4827 12257 4839 12291
rect 4781 12251 4839 12257
rect 17589 12291 17647 12297
rect 17589 12257 17601 12291
rect 17635 12288 17647 12291
rect 18046 12288 18052 12300
rect 17635 12260 18052 12288
rect 17635 12257 17647 12260
rect 17589 12251 17647 12257
rect 18046 12248 18052 12260
rect 18104 12248 18110 12300
rect 18414 12288 18420 12300
rect 18375 12260 18420 12288
rect 18414 12248 18420 12260
rect 18472 12248 18478 12300
rect 2777 12223 2835 12229
rect 1504 12192 2544 12220
rect 1673 12155 1731 12161
rect 1673 12121 1685 12155
rect 1719 12152 1731 12155
rect 2406 12152 2412 12164
rect 1719 12124 2412 12152
rect 1719 12121 1731 12124
rect 1673 12115 1731 12121
rect 2406 12112 2412 12124
rect 2464 12112 2470 12164
rect 1946 12084 1952 12096
rect 1907 12056 1952 12084
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 2225 12087 2283 12093
rect 2225 12053 2237 12087
rect 2271 12084 2283 12087
rect 2314 12084 2320 12096
rect 2271 12056 2320 12084
rect 2271 12053 2283 12056
rect 2225 12047 2283 12053
rect 2314 12044 2320 12056
rect 2372 12044 2378 12096
rect 2516 12084 2544 12192
rect 2777 12189 2789 12223
rect 2823 12189 2835 12223
rect 3513 12223 3571 12229
rect 3513 12220 3525 12223
rect 2777 12183 2835 12189
rect 2976 12192 3525 12220
rect 2590 12112 2596 12164
rect 2648 12152 2654 12164
rect 2792 12152 2820 12183
rect 2866 12152 2872 12164
rect 2648 12124 2872 12152
rect 2648 12112 2654 12124
rect 2866 12112 2872 12124
rect 2924 12112 2930 12164
rect 2976 12084 3004 12192
rect 3513 12189 3525 12192
rect 3559 12189 3571 12223
rect 3513 12183 3571 12189
rect 4338 12180 4344 12232
rect 4396 12220 4402 12232
rect 4525 12223 4583 12229
rect 4525 12220 4537 12223
rect 4396 12192 4537 12220
rect 4396 12180 4402 12192
rect 4525 12189 4537 12192
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 17773 12223 17831 12229
rect 17773 12189 17785 12223
rect 17819 12220 17831 12223
rect 18432 12220 18460 12248
rect 17819 12192 18460 12220
rect 17819 12189 17831 12192
rect 17773 12183 17831 12189
rect 16574 12112 16580 12164
rect 16632 12152 16638 12164
rect 17865 12155 17923 12161
rect 17865 12152 17877 12155
rect 16632 12124 17877 12152
rect 16632 12112 16638 12124
rect 17865 12121 17877 12124
rect 17911 12121 17923 12155
rect 17865 12115 17923 12121
rect 3326 12084 3332 12096
rect 2516 12056 3004 12084
rect 3287 12056 3332 12084
rect 3326 12044 3332 12056
rect 3384 12044 3390 12096
rect 3510 12044 3516 12096
rect 3568 12084 3574 12096
rect 3786 12084 3792 12096
rect 3568 12056 3792 12084
rect 3568 12044 3574 12056
rect 3786 12044 3792 12056
rect 3844 12084 3850 12096
rect 3881 12087 3939 12093
rect 3881 12084 3893 12087
rect 3844 12056 3893 12084
rect 3844 12044 3850 12056
rect 3881 12053 3893 12056
rect 3927 12053 3939 12087
rect 3881 12047 3939 12053
rect 5905 12087 5963 12093
rect 5905 12053 5917 12087
rect 5951 12084 5963 12087
rect 6546 12084 6552 12096
rect 5951 12056 6552 12084
rect 5951 12053 5963 12056
rect 5905 12047 5963 12053
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 18325 12087 18383 12093
rect 18325 12053 18337 12087
rect 18371 12084 18383 12087
rect 18690 12084 18696 12096
rect 18371 12056 18696 12084
rect 18371 12053 18383 12056
rect 18325 12047 18383 12053
rect 18690 12044 18696 12056
rect 18748 12044 18754 12096
rect 1104 11994 18860 12016
rect 1104 11942 3947 11994
rect 3999 11942 4011 11994
rect 4063 11942 4075 11994
rect 4127 11942 4139 11994
rect 4191 11942 9878 11994
rect 9930 11942 9942 11994
rect 9994 11942 10006 11994
rect 10058 11942 10070 11994
rect 10122 11942 15808 11994
rect 15860 11942 15872 11994
rect 15924 11942 15936 11994
rect 15988 11942 16000 11994
rect 16052 11942 18860 11994
rect 1104 11920 18860 11942
rect 1946 11840 1952 11892
rect 2004 11880 2010 11892
rect 5721 11883 5779 11889
rect 5721 11880 5733 11883
rect 2004 11852 5733 11880
rect 2004 11840 2010 11852
rect 5721 11849 5733 11852
rect 5767 11880 5779 11883
rect 6270 11880 6276 11892
rect 5767 11852 6276 11880
rect 5767 11849 5779 11852
rect 5721 11843 5779 11849
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 2314 11744 2320 11756
rect 2275 11716 2320 11744
rect 2314 11704 2320 11716
rect 2372 11704 2378 11756
rect 2498 11744 2504 11756
rect 2459 11716 2504 11744
rect 2498 11704 2504 11716
rect 2556 11704 2562 11756
rect 15102 11744 15108 11756
rect 7484 11716 15108 11744
rect 1486 11676 1492 11688
rect 1447 11648 1492 11676
rect 1486 11636 1492 11648
rect 1544 11636 1550 11688
rect 2130 11636 2136 11688
rect 2188 11676 2194 11688
rect 2225 11679 2283 11685
rect 2225 11676 2237 11679
rect 2188 11648 2237 11676
rect 2188 11636 2194 11648
rect 2225 11645 2237 11648
rect 2271 11645 2283 11679
rect 2225 11639 2283 11645
rect 2777 11679 2835 11685
rect 2777 11645 2789 11679
rect 2823 11676 2835 11679
rect 4249 11679 4307 11685
rect 4249 11676 4261 11679
rect 2823 11648 4261 11676
rect 2823 11645 2835 11648
rect 2777 11639 2835 11645
rect 4249 11645 4261 11648
rect 4295 11676 4307 11679
rect 4338 11676 4344 11688
rect 4295 11648 4344 11676
rect 4295 11645 4307 11648
rect 4249 11639 4307 11645
rect 4338 11636 4344 11648
rect 4396 11676 4402 11688
rect 6273 11679 6331 11685
rect 6273 11676 6285 11679
rect 4396 11648 6285 11676
rect 4396 11636 4402 11648
rect 6273 11645 6285 11648
rect 6319 11676 6331 11679
rect 6457 11679 6515 11685
rect 6457 11676 6469 11679
rect 6319 11648 6469 11676
rect 6319 11645 6331 11648
rect 6273 11639 6331 11645
rect 6457 11645 6469 11648
rect 6503 11645 6515 11679
rect 6457 11639 6515 11645
rect 6546 11636 6552 11688
rect 6604 11676 6610 11688
rect 6713 11679 6771 11685
rect 6713 11676 6725 11679
rect 6604 11648 6725 11676
rect 6604 11636 6610 11648
rect 6713 11645 6725 11648
rect 6759 11645 6771 11679
rect 6713 11639 6771 11645
rect 2958 11568 2964 11620
rect 3016 11617 3022 11620
rect 3016 11611 3080 11617
rect 3016 11577 3034 11611
rect 3068 11577 3080 11611
rect 4494 11611 4552 11617
rect 4494 11608 4506 11611
rect 3016 11571 3080 11577
rect 4172 11580 4506 11608
rect 3016 11568 3022 11571
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 1857 11543 1915 11549
rect 1857 11509 1869 11543
rect 1903 11540 1915 11543
rect 1946 11540 1952 11552
rect 1903 11512 1952 11540
rect 1903 11509 1915 11512
rect 1857 11503 1915 11509
rect 1946 11500 1952 11512
rect 2004 11500 2010 11552
rect 2498 11500 2504 11552
rect 2556 11540 2562 11552
rect 4172 11549 4200 11580
rect 4494 11577 4506 11580
rect 4540 11577 4552 11611
rect 4494 11571 4552 11577
rect 4706 11568 4712 11620
rect 4764 11608 4770 11620
rect 7484 11608 7512 11716
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 7558 11636 7564 11688
rect 7616 11676 7622 11688
rect 7929 11679 7987 11685
rect 7929 11676 7941 11679
rect 7616 11648 7941 11676
rect 7616 11636 7622 11648
rect 7929 11645 7941 11648
rect 7975 11676 7987 11679
rect 8110 11676 8116 11688
rect 7975 11648 8116 11676
rect 7975 11645 7987 11648
rect 7929 11639 7987 11645
rect 8110 11636 8116 11648
rect 8168 11676 8174 11688
rect 9033 11679 9091 11685
rect 9033 11676 9045 11679
rect 8168 11648 9045 11676
rect 8168 11636 8174 11648
rect 9033 11645 9045 11648
rect 9079 11645 9091 11679
rect 17862 11676 17868 11688
rect 17823 11648 17868 11676
rect 9033 11639 9091 11645
rect 17862 11636 17868 11648
rect 17920 11636 17926 11688
rect 4764 11580 7512 11608
rect 8757 11611 8815 11617
rect 4764 11568 4770 11580
rect 8757 11577 8769 11611
rect 8803 11608 8815 11611
rect 8938 11608 8944 11620
rect 8803 11580 8944 11608
rect 8803 11577 8815 11580
rect 8757 11571 8815 11577
rect 8938 11568 8944 11580
rect 8996 11568 9002 11620
rect 17773 11611 17831 11617
rect 17773 11577 17785 11611
rect 17819 11608 17831 11611
rect 18414 11608 18420 11620
rect 17819 11580 18420 11608
rect 17819 11577 17831 11580
rect 17773 11571 17831 11577
rect 18414 11568 18420 11580
rect 18472 11568 18478 11620
rect 4157 11543 4215 11549
rect 4157 11540 4169 11543
rect 2556 11512 4169 11540
rect 2556 11500 2562 11512
rect 4157 11509 4169 11512
rect 4203 11509 4215 11543
rect 4157 11503 4215 11509
rect 4614 11500 4620 11552
rect 4672 11540 4678 11552
rect 5629 11543 5687 11549
rect 5629 11540 5641 11543
rect 4672 11512 5641 11540
rect 4672 11500 4678 11512
rect 5629 11509 5641 11512
rect 5675 11509 5687 11543
rect 5629 11503 5687 11509
rect 6273 11543 6331 11549
rect 6273 11509 6285 11543
rect 6319 11540 6331 11543
rect 7282 11540 7288 11552
rect 6319 11512 7288 11540
rect 6319 11509 6331 11512
rect 6273 11503 6331 11509
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 7834 11540 7840 11552
rect 7795 11512 7840 11540
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 17310 11500 17316 11552
rect 17368 11540 17374 11552
rect 17497 11543 17555 11549
rect 17497 11540 17509 11543
rect 17368 11512 17509 11540
rect 17368 11500 17374 11512
rect 17497 11509 17509 11512
rect 17543 11509 17555 11543
rect 17497 11503 17555 11509
rect 18049 11543 18107 11549
rect 18049 11509 18061 11543
rect 18095 11540 18107 11543
rect 18230 11540 18236 11552
rect 18095 11512 18236 11540
rect 18095 11509 18107 11512
rect 18049 11503 18107 11509
rect 18230 11500 18236 11512
rect 18288 11500 18294 11552
rect 18325 11543 18383 11549
rect 18325 11509 18337 11543
rect 18371 11540 18383 11543
rect 18782 11540 18788 11552
rect 18371 11512 18788 11540
rect 18371 11509 18383 11512
rect 18325 11503 18383 11509
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 1104 11450 18860 11472
rect 1104 11398 6912 11450
rect 6964 11398 6976 11450
rect 7028 11398 7040 11450
rect 7092 11398 7104 11450
rect 7156 11398 12843 11450
rect 12895 11398 12907 11450
rect 12959 11398 12971 11450
rect 13023 11398 13035 11450
rect 13087 11398 18860 11450
rect 1104 11376 18860 11398
rect 3145 11339 3203 11345
rect 3145 11305 3157 11339
rect 3191 11336 3203 11339
rect 3973 11339 4031 11345
rect 3973 11336 3985 11339
rect 3191 11308 3985 11336
rect 3191 11305 3203 11308
rect 3145 11299 3203 11305
rect 3973 11305 3985 11308
rect 4019 11336 4031 11339
rect 4706 11336 4712 11348
rect 4019 11308 4712 11336
rect 4019 11305 4031 11308
rect 3973 11299 4031 11305
rect 3160 11268 3188 11299
rect 4706 11296 4712 11308
rect 4764 11296 4770 11348
rect 5261 11339 5319 11345
rect 5261 11305 5273 11339
rect 5307 11336 5319 11339
rect 5813 11339 5871 11345
rect 5813 11336 5825 11339
rect 5307 11308 5825 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 5813 11305 5825 11308
rect 5859 11305 5871 11339
rect 5813 11299 5871 11305
rect 5902 11296 5908 11348
rect 5960 11336 5966 11348
rect 6454 11336 6460 11348
rect 5960 11308 6460 11336
rect 5960 11296 5966 11308
rect 6454 11296 6460 11308
rect 6512 11336 6518 11348
rect 17862 11336 17868 11348
rect 6512 11308 17868 11336
rect 6512 11296 6518 11308
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 18049 11339 18107 11345
rect 18049 11305 18061 11339
rect 18095 11336 18107 11339
rect 18598 11336 18604 11348
rect 18095 11308 18604 11336
rect 18095 11305 18107 11308
rect 18049 11299 18107 11305
rect 18598 11296 18604 11308
rect 18656 11296 18662 11348
rect 6638 11268 6644 11280
rect 2746 11240 3188 11268
rect 5920 11240 6644 11268
rect 1394 11160 1400 11212
rect 1452 11200 1458 11212
rect 1489 11203 1547 11209
rect 1489 11200 1501 11203
rect 1452 11172 1501 11200
rect 1452 11160 1458 11172
rect 1489 11169 1501 11172
rect 1535 11169 1547 11203
rect 2222 11200 2228 11212
rect 2183 11172 2228 11200
rect 1489 11163 1547 11169
rect 2222 11160 2228 11172
rect 2280 11160 2286 11212
rect 2406 11160 2412 11212
rect 2464 11200 2470 11212
rect 2746 11200 2774 11240
rect 2464 11172 2774 11200
rect 3053 11203 3111 11209
rect 2464 11160 2470 11172
rect 3053 11169 3065 11203
rect 3099 11200 3111 11203
rect 3099 11172 3188 11200
rect 3099 11169 3111 11172
rect 3053 11163 3111 11169
rect 2314 11132 2320 11144
rect 2275 11104 2320 11132
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 2498 11132 2504 11144
rect 2459 11104 2504 11132
rect 2498 11092 2504 11104
rect 2556 11092 2562 11144
rect 1673 11067 1731 11073
rect 1673 11033 1685 11067
rect 1719 11064 1731 11067
rect 3050 11064 3056 11076
rect 1719 11036 3056 11064
rect 1719 11033 1731 11036
rect 1673 11027 1731 11033
rect 3050 11024 3056 11036
rect 3108 11024 3114 11076
rect 1854 10996 1860 11008
rect 1815 10968 1860 10996
rect 1854 10956 1860 10968
rect 1912 10956 1918 11008
rect 2682 10996 2688 11008
rect 2643 10968 2688 10996
rect 2682 10956 2688 10968
rect 2740 10956 2746 11008
rect 3160 10996 3188 11172
rect 4522 11160 4528 11212
rect 4580 11200 4586 11212
rect 4893 11203 4951 11209
rect 4893 11200 4905 11203
rect 4580 11172 4905 11200
rect 4580 11160 4586 11172
rect 4893 11169 4905 11172
rect 4939 11200 4951 11203
rect 4982 11200 4988 11212
rect 4939 11172 4988 11200
rect 4939 11169 4951 11172
rect 4893 11163 4951 11169
rect 4982 11160 4988 11172
rect 5040 11200 5046 11212
rect 5353 11203 5411 11209
rect 5353 11200 5365 11203
rect 5040 11172 5365 11200
rect 5040 11160 5046 11172
rect 5353 11169 5365 11172
rect 5399 11169 5411 11203
rect 5353 11163 5411 11169
rect 3329 11135 3387 11141
rect 3329 11101 3341 11135
rect 3375 11132 3387 11135
rect 3418 11132 3424 11144
rect 3375 11104 3424 11132
rect 3375 11101 3387 11104
rect 3329 11095 3387 11101
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11132 5227 11135
rect 5920 11132 5948 11240
rect 6638 11228 6644 11240
rect 6696 11268 6702 11280
rect 7006 11268 7012 11280
rect 6696 11240 7012 11268
rect 6696 11228 6702 11240
rect 7006 11228 7012 11240
rect 7064 11268 7070 11280
rect 7834 11268 7840 11280
rect 7064 11240 7840 11268
rect 7064 11228 7070 11240
rect 7834 11228 7840 11240
rect 7892 11268 7898 11280
rect 7938 11271 7996 11277
rect 7938 11268 7950 11271
rect 7892 11240 7950 11268
rect 7892 11228 7898 11240
rect 7938 11237 7950 11240
rect 7984 11237 7996 11271
rect 7938 11231 7996 11237
rect 11548 11271 11606 11277
rect 11548 11237 11560 11271
rect 11594 11268 11606 11271
rect 11882 11268 11888 11280
rect 11594 11240 11888 11268
rect 11594 11237 11606 11240
rect 11548 11231 11606 11237
rect 11882 11228 11888 11240
rect 11940 11228 11946 11280
rect 11974 11228 11980 11280
rect 12032 11268 12038 11280
rect 17037 11271 17095 11277
rect 17037 11268 17049 11271
rect 12032 11240 17049 11268
rect 12032 11228 12038 11240
rect 17037 11237 17049 11240
rect 17083 11237 17095 11271
rect 17037 11231 17095 11237
rect 17313 11271 17371 11277
rect 17313 11237 17325 11271
rect 17359 11268 17371 11271
rect 17359 11240 18460 11268
rect 17359 11237 17371 11240
rect 17313 11231 17371 11237
rect 6181 11203 6239 11209
rect 6181 11200 6193 11203
rect 5215 11104 5948 11132
rect 6104 11172 6193 11200
rect 5215 11101 5227 11104
rect 5169 11095 5227 11101
rect 3510 11064 3516 11076
rect 3471 11036 3516 11064
rect 3510 11024 3516 11036
rect 3568 11024 3574 11076
rect 4157 11067 4215 11073
rect 4157 11064 4169 11067
rect 3620 11036 4169 11064
rect 3620 10996 3648 11036
rect 4157 11033 4169 11036
rect 4203 11064 4215 11067
rect 4706 11064 4712 11076
rect 4203 11036 4712 11064
rect 4203 11033 4215 11036
rect 4157 11027 4215 11033
rect 4706 11024 4712 11036
rect 4764 11024 4770 11076
rect 5552 11036 5856 11064
rect 3160 10968 3648 10996
rect 3694 10956 3700 11008
rect 3752 10996 3758 11008
rect 5552 10996 5580 11036
rect 5718 10996 5724 11008
rect 3752 10968 5580 10996
rect 5679 10968 5724 10996
rect 3752 10956 3758 10968
rect 5718 10956 5724 10968
rect 5776 10956 5782 11008
rect 5828 10996 5856 11036
rect 5902 11024 5908 11076
rect 5960 11064 5966 11076
rect 6104 11064 6132 11172
rect 6181 11169 6193 11172
rect 6227 11169 6239 11203
rect 6733 11203 6791 11209
rect 6733 11200 6745 11203
rect 6181 11163 6239 11169
rect 6380 11172 6745 11200
rect 6270 11132 6276 11144
rect 6231 11104 6276 11132
rect 6270 11092 6276 11104
rect 6328 11092 6334 11144
rect 6380 11064 6408 11172
rect 6733 11169 6745 11172
rect 6779 11169 6791 11203
rect 6733 11163 6791 11169
rect 7374 11160 7380 11212
rect 7432 11200 7438 11212
rect 8205 11203 8263 11209
rect 8205 11200 8217 11203
rect 7432 11172 8217 11200
rect 7432 11160 7438 11172
rect 8205 11169 8217 11172
rect 8251 11169 8263 11203
rect 8205 11163 8263 11169
rect 11698 11160 11704 11212
rect 11756 11200 11762 11212
rect 11793 11203 11851 11209
rect 11793 11200 11805 11203
rect 11756 11172 11805 11200
rect 11756 11160 11762 11172
rect 11793 11169 11805 11172
rect 11839 11200 11851 11203
rect 13538 11200 13544 11212
rect 13596 11209 13602 11212
rect 11839 11172 12434 11200
rect 13508 11172 13544 11200
rect 11839 11169 11851 11172
rect 11793 11163 11851 11169
rect 6457 11135 6515 11141
rect 6457 11101 6469 11135
rect 6503 11132 6515 11135
rect 6546 11132 6552 11144
rect 6503 11104 6552 11132
rect 6503 11101 6515 11104
rect 6457 11095 6515 11101
rect 6546 11092 6552 11104
rect 6604 11092 6610 11144
rect 11882 11092 11888 11144
rect 11940 11132 11946 11144
rect 12406 11132 12434 11172
rect 13538 11160 13544 11172
rect 13596 11163 13608 11209
rect 17052 11200 17080 11231
rect 18432 11209 18460 11240
rect 17865 11203 17923 11209
rect 17865 11200 17877 11203
rect 17052 11172 17877 11200
rect 17865 11169 17877 11172
rect 17911 11169 17923 11203
rect 17865 11163 17923 11169
rect 18417 11203 18475 11209
rect 18417 11169 18429 11203
rect 18463 11200 18475 11203
rect 18506 11200 18512 11212
rect 18463 11172 18512 11200
rect 18463 11169 18475 11172
rect 18417 11163 18475 11169
rect 13596 11160 13602 11163
rect 18506 11160 18512 11172
rect 18564 11160 18570 11212
rect 13817 11135 13875 11141
rect 11940 11104 12296 11132
rect 12406 11104 12664 11132
rect 11940 11092 11946 11104
rect 12268 11076 12296 11104
rect 5960 11036 6408 11064
rect 6656 11036 6960 11064
rect 5960 11024 5966 11036
rect 6656 10996 6684 11036
rect 6822 10996 6828 11008
rect 5828 10968 6684 10996
rect 6783 10968 6828 10996
rect 6822 10956 6828 10968
rect 6880 10956 6886 11008
rect 6932 10996 6960 11036
rect 9692 11036 10548 11064
rect 9692 10996 9720 11036
rect 6932 10968 9720 10996
rect 9766 10956 9772 11008
rect 9824 10996 9830 11008
rect 10318 10996 10324 11008
rect 9824 10968 10324 10996
rect 9824 10956 9830 10968
rect 10318 10956 10324 10968
rect 10376 10996 10382 11008
rect 10413 10999 10471 11005
rect 10413 10996 10425 10999
rect 10376 10968 10425 10996
rect 10376 10956 10382 10968
rect 10413 10965 10425 10968
rect 10459 10965 10471 10999
rect 10520 10996 10548 11036
rect 12250 11024 12256 11076
rect 12308 11064 12314 11076
rect 12437 11067 12495 11073
rect 12437 11064 12449 11067
rect 12308 11036 12449 11064
rect 12308 11024 12314 11036
rect 12437 11033 12449 11036
rect 12483 11033 12495 11067
rect 12437 11027 12495 11033
rect 11606 10996 11612 11008
rect 10520 10968 11612 10996
rect 10413 10959 10471 10965
rect 11606 10956 11612 10968
rect 11664 10956 11670 11008
rect 11882 10996 11888 11008
rect 11843 10968 11888 10996
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 12636 10996 12664 11104
rect 13817 11101 13829 11135
rect 13863 11101 13875 11135
rect 13817 11095 13875 11101
rect 13832 10996 13860 11095
rect 16022 11092 16028 11144
rect 16080 11132 16086 11144
rect 16298 11132 16304 11144
rect 16080 11104 16304 11132
rect 16080 11092 16086 11104
rect 16298 11092 16304 11104
rect 16356 11092 16362 11144
rect 17589 11135 17647 11141
rect 17589 11101 17601 11135
rect 17635 11132 17647 11135
rect 18046 11132 18052 11144
rect 17635 11104 18052 11132
rect 17635 11101 17647 11104
rect 17589 11095 17647 11101
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 14090 11024 14096 11076
rect 14148 11064 14154 11076
rect 17770 11064 17776 11076
rect 14148 11036 17632 11064
rect 17731 11036 17776 11064
rect 14148 11024 14154 11036
rect 14918 10996 14924 11008
rect 12636 10968 14924 10996
rect 14918 10956 14924 10968
rect 14976 10956 14982 11008
rect 16942 10996 16948 11008
rect 16855 10968 16948 10996
rect 16942 10956 16948 10968
rect 17000 10996 17006 11008
rect 17126 10996 17132 11008
rect 17000 10968 17132 10996
rect 17000 10956 17006 10968
rect 17126 10956 17132 10968
rect 17184 10956 17190 11008
rect 17604 10996 17632 11036
rect 17770 11024 17776 11036
rect 17828 11024 17834 11076
rect 18233 11067 18291 11073
rect 18233 11064 18245 11067
rect 17880 11036 18245 11064
rect 17880 10996 17908 11036
rect 18233 11033 18245 11036
rect 18279 11033 18291 11067
rect 18233 11027 18291 11033
rect 17604 10968 17908 10996
rect 1104 10906 18860 10928
rect 1104 10854 3947 10906
rect 3999 10854 4011 10906
rect 4063 10854 4075 10906
rect 4127 10854 4139 10906
rect 4191 10854 9878 10906
rect 9930 10854 9942 10906
rect 9994 10854 10006 10906
rect 10058 10854 10070 10906
rect 10122 10854 15808 10906
rect 15860 10854 15872 10906
rect 15924 10854 15936 10906
rect 15988 10854 16000 10906
rect 16052 10854 18860 10906
rect 1104 10832 18860 10854
rect 2222 10752 2228 10804
rect 2280 10792 2286 10804
rect 2501 10795 2559 10801
rect 2501 10792 2513 10795
rect 2280 10764 2513 10792
rect 2280 10752 2286 10764
rect 2501 10761 2513 10764
rect 2547 10761 2559 10795
rect 4157 10795 4215 10801
rect 4157 10792 4169 10795
rect 2501 10755 2559 10761
rect 2746 10764 4169 10792
rect 2130 10684 2136 10736
rect 2188 10724 2194 10736
rect 2746 10724 2774 10764
rect 4157 10761 4169 10764
rect 4203 10792 4215 10795
rect 11882 10792 11888 10804
rect 4203 10764 11888 10792
rect 4203 10761 4215 10764
rect 4157 10755 4215 10761
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 13538 10792 13544 10804
rect 13499 10764 13544 10792
rect 13538 10752 13544 10764
rect 13596 10752 13602 10804
rect 2188 10696 2774 10724
rect 2188 10684 2194 10696
rect 6086 10684 6092 10736
rect 6144 10724 6150 10736
rect 6181 10727 6239 10733
rect 6181 10724 6193 10727
rect 6144 10696 6193 10724
rect 6144 10684 6150 10696
rect 6181 10693 6193 10696
rect 6227 10693 6239 10727
rect 6181 10687 6239 10693
rect 6822 10684 6828 10736
rect 6880 10724 6886 10736
rect 6880 10696 7144 10724
rect 6880 10684 6886 10696
rect 1762 10616 1768 10668
rect 1820 10656 1826 10668
rect 1857 10659 1915 10665
rect 1857 10656 1869 10659
rect 1820 10628 1869 10656
rect 1820 10616 1826 10628
rect 1857 10625 1869 10628
rect 1903 10625 1915 10659
rect 1857 10619 1915 10625
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 2682 10656 2688 10668
rect 2087 10628 2688 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 4246 10616 4252 10668
rect 4304 10656 4310 10668
rect 5721 10659 5779 10665
rect 4304 10628 5672 10656
rect 4304 10616 4310 10628
rect 2130 10588 2136 10600
rect 2091 10560 2136 10588
rect 2130 10548 2136 10560
rect 2188 10548 2194 10600
rect 3326 10548 3332 10600
rect 3384 10588 3390 10600
rect 3706 10591 3764 10597
rect 3706 10588 3718 10591
rect 3384 10560 3718 10588
rect 3384 10548 3390 10560
rect 3706 10557 3718 10560
rect 3752 10557 3764 10591
rect 3706 10551 3764 10557
rect 3973 10591 4031 10597
rect 3973 10557 3985 10591
rect 4019 10588 4031 10591
rect 4338 10588 4344 10600
rect 4019 10560 4344 10588
rect 4019 10557 4031 10560
rect 3973 10551 4031 10557
rect 1486 10520 1492 10532
rect 1447 10492 1492 10520
rect 1486 10480 1492 10492
rect 1544 10520 1550 10532
rect 3418 10520 3424 10532
rect 1544 10492 3424 10520
rect 1544 10480 1550 10492
rect 3418 10480 3424 10492
rect 3476 10480 3482 10532
rect 3602 10480 3608 10532
rect 3660 10520 3666 10532
rect 3988 10520 4016 10551
rect 4338 10548 4344 10560
rect 4396 10548 4402 10600
rect 5442 10548 5448 10600
rect 5500 10588 5506 10600
rect 5537 10591 5595 10597
rect 5537 10588 5549 10591
rect 5500 10560 5549 10588
rect 5500 10548 5506 10560
rect 5537 10557 5549 10560
rect 5583 10557 5595 10591
rect 5644 10588 5672 10628
rect 5721 10625 5733 10659
rect 5767 10656 5779 10659
rect 5902 10656 5908 10668
rect 5767 10628 5908 10656
rect 5767 10625 5779 10628
rect 5721 10619 5779 10625
rect 5902 10616 5908 10628
rect 5960 10656 5966 10668
rect 6840 10656 6868 10684
rect 7006 10656 7012 10668
rect 5960 10628 6868 10656
rect 6967 10628 7012 10656
rect 5960 10616 5966 10628
rect 7006 10616 7012 10628
rect 7064 10616 7070 10668
rect 7116 10656 7144 10696
rect 7190 10684 7196 10736
rect 7248 10724 7254 10736
rect 7374 10724 7380 10736
rect 7248 10696 7380 10724
rect 7248 10684 7254 10696
rect 7374 10684 7380 10696
rect 7432 10684 7438 10736
rect 10244 10696 12204 10724
rect 10244 10656 10272 10696
rect 7116 10628 7512 10656
rect 6089 10591 6147 10597
rect 5644 10560 6040 10588
rect 5537 10551 5595 10557
rect 3660 10492 4016 10520
rect 4356 10520 4384 10548
rect 6012 10520 6040 10560
rect 6089 10557 6101 10591
rect 6135 10588 6147 10591
rect 6181 10591 6239 10597
rect 6181 10588 6193 10591
rect 6135 10560 6193 10588
rect 6135 10557 6147 10560
rect 6089 10551 6147 10557
rect 6181 10557 6193 10560
rect 6227 10557 6239 10591
rect 6181 10551 6239 10557
rect 6454 10548 6460 10600
rect 6512 10588 6518 10600
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 6512 10560 6837 10588
rect 6512 10548 6518 10560
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 6917 10591 6975 10597
rect 6917 10557 6929 10591
rect 6963 10588 6975 10591
rect 7190 10588 7196 10600
rect 6963 10560 7196 10588
rect 6963 10557 6975 10560
rect 6917 10551 6975 10557
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 7282 10548 7288 10600
rect 7340 10588 7346 10600
rect 7377 10591 7435 10597
rect 7377 10588 7389 10591
rect 7340 10560 7389 10588
rect 7340 10548 7346 10560
rect 7377 10557 7389 10560
rect 7423 10557 7435 10591
rect 7484 10588 7512 10628
rect 10152 10628 10272 10656
rect 7633 10591 7691 10597
rect 7633 10588 7645 10591
rect 7484 10560 7645 10588
rect 7377 10551 7435 10557
rect 7633 10557 7645 10560
rect 7679 10557 7691 10591
rect 10152 10588 10180 10628
rect 10318 10616 10324 10668
rect 10376 10656 10382 10668
rect 11333 10659 11391 10665
rect 11333 10656 11345 10659
rect 10376 10628 11345 10656
rect 10376 10616 10382 10628
rect 11333 10625 11345 10628
rect 11379 10625 11391 10659
rect 11333 10619 11391 10625
rect 7633 10551 7691 10557
rect 7760 10560 10180 10588
rect 10222 10591 10280 10597
rect 4356 10492 5948 10520
rect 6012 10492 6592 10520
rect 3660 10480 3666 10492
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 1762 10412 1768 10464
rect 1820 10452 1826 10464
rect 2590 10452 2596 10464
rect 1820 10424 2596 10452
rect 1820 10412 1826 10424
rect 2590 10412 2596 10424
rect 2648 10452 2654 10464
rect 2958 10452 2964 10464
rect 2648 10424 2964 10452
rect 2648 10412 2654 10424
rect 2958 10412 2964 10424
rect 3016 10412 3022 10464
rect 4890 10412 4896 10464
rect 4948 10452 4954 10464
rect 5077 10455 5135 10461
rect 5077 10452 5089 10455
rect 4948 10424 5089 10452
rect 4948 10412 4954 10424
rect 5077 10421 5089 10424
rect 5123 10421 5135 10455
rect 5077 10415 5135 10421
rect 5445 10455 5503 10461
rect 5445 10421 5457 10455
rect 5491 10452 5503 10455
rect 5718 10452 5724 10464
rect 5491 10424 5724 10452
rect 5491 10421 5503 10424
rect 5445 10415 5503 10421
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 5920 10461 5948 10492
rect 5905 10455 5963 10461
rect 5905 10421 5917 10455
rect 5951 10421 5963 10455
rect 5905 10415 5963 10421
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 6457 10455 6515 10461
rect 6457 10452 6469 10455
rect 6052 10424 6469 10452
rect 6052 10412 6058 10424
rect 6457 10421 6469 10424
rect 6503 10421 6515 10455
rect 6564 10452 6592 10492
rect 7760 10452 7788 10560
rect 10222 10557 10234 10591
rect 10268 10557 10280 10591
rect 10222 10551 10280 10557
rect 10413 10591 10471 10597
rect 10413 10557 10425 10591
rect 10459 10588 10471 10591
rect 10686 10588 10692 10600
rect 10459 10560 10692 10588
rect 10459 10557 10471 10560
rect 10413 10551 10471 10557
rect 9766 10480 9772 10532
rect 9824 10520 9830 10532
rect 9962 10523 10020 10529
rect 9962 10520 9974 10523
rect 9824 10492 9974 10520
rect 9824 10480 9830 10492
rect 9962 10489 9974 10492
rect 10008 10489 10020 10523
rect 10244 10520 10272 10551
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 11698 10588 11704 10600
rect 11072 10560 11704 10588
rect 11072 10520 11100 10560
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 12176 10588 12204 10696
rect 12250 10616 12256 10668
rect 12308 10656 12314 10668
rect 12345 10659 12403 10665
rect 12345 10656 12357 10659
rect 12308 10628 12357 10656
rect 12308 10616 12314 10628
rect 12345 10625 12357 10628
rect 12391 10625 12403 10659
rect 13262 10656 13268 10668
rect 13175 10628 13268 10656
rect 12345 10619 12403 10625
rect 13262 10616 13268 10628
rect 13320 10656 13326 10668
rect 13556 10656 13584 10752
rect 16758 10684 16764 10736
rect 16816 10724 16822 10736
rect 17218 10724 17224 10736
rect 16816 10696 17224 10724
rect 16816 10684 16822 10696
rect 17218 10684 17224 10696
rect 17276 10684 17282 10736
rect 14918 10656 14924 10668
rect 13320 10628 13584 10656
rect 14879 10628 14924 10656
rect 13320 10616 13326 10628
rect 14918 10616 14924 10628
rect 14976 10616 14982 10668
rect 16482 10616 16488 10668
rect 16540 10656 16546 10668
rect 17497 10659 17555 10665
rect 17497 10656 17509 10659
rect 16540 10628 17509 10656
rect 16540 10616 16546 10628
rect 17497 10625 17509 10628
rect 17543 10625 17555 10659
rect 17497 10619 17555 10625
rect 17770 10616 17776 10668
rect 17828 10656 17834 10668
rect 17828 10628 18460 10656
rect 17828 10616 17834 10628
rect 16577 10591 16635 10597
rect 16577 10588 16589 10591
rect 12176 10560 16589 10588
rect 16577 10557 16589 10560
rect 16623 10588 16635 10591
rect 16666 10588 16672 10600
rect 16623 10560 16672 10588
rect 16623 10557 16635 10560
rect 16577 10551 16635 10557
rect 16666 10548 16672 10560
rect 16724 10548 16730 10600
rect 16761 10591 16819 10597
rect 16761 10557 16773 10591
rect 16807 10588 16819 10591
rect 16807 10560 18092 10588
rect 16807 10557 16819 10560
rect 16761 10551 16819 10557
rect 10244 10492 11100 10520
rect 11149 10523 11207 10529
rect 9962 10483 10020 10489
rect 11149 10489 11161 10523
rect 11195 10520 11207 10523
rect 11195 10492 11836 10520
rect 11195 10489 11207 10492
rect 11149 10483 11207 10489
rect 8754 10452 8760 10464
rect 6564 10424 7788 10452
rect 8715 10424 8760 10452
rect 6457 10415 6515 10421
rect 8754 10412 8760 10424
rect 8812 10412 8818 10464
rect 8849 10455 8907 10461
rect 8849 10421 8861 10455
rect 8895 10452 8907 10455
rect 10134 10452 10140 10464
rect 8895 10424 10140 10452
rect 8895 10421 8907 10424
rect 8849 10415 8907 10421
rect 10134 10412 10140 10424
rect 10192 10412 10198 10464
rect 10410 10412 10416 10464
rect 10468 10452 10474 10464
rect 10781 10455 10839 10461
rect 10781 10452 10793 10455
rect 10468 10424 10793 10452
rect 10468 10412 10474 10424
rect 10781 10421 10793 10424
rect 10827 10421 10839 10455
rect 11238 10452 11244 10464
rect 11199 10424 11244 10452
rect 10781 10415 10839 10421
rect 11238 10412 11244 10424
rect 11296 10412 11302 10464
rect 11808 10461 11836 10492
rect 11882 10480 11888 10532
rect 11940 10520 11946 10532
rect 12161 10523 12219 10529
rect 12161 10520 12173 10523
rect 11940 10492 12173 10520
rect 11940 10480 11946 10492
rect 12161 10489 12173 10492
rect 12207 10489 12219 10523
rect 12161 10483 12219 10489
rect 12989 10523 13047 10529
rect 12989 10489 13001 10523
rect 13035 10520 13047 10523
rect 13354 10520 13360 10532
rect 13035 10492 13360 10520
rect 13035 10489 13047 10492
rect 12989 10483 13047 10489
rect 13354 10480 13360 10492
rect 13412 10520 13418 10532
rect 13412 10492 13768 10520
rect 13412 10480 13418 10492
rect 13740 10464 13768 10492
rect 13998 10480 14004 10532
rect 14056 10520 14062 10532
rect 14654 10523 14712 10529
rect 14654 10520 14666 10523
rect 14056 10492 14666 10520
rect 14056 10480 14062 10492
rect 14654 10489 14666 10492
rect 14700 10489 14712 10523
rect 14654 10483 14712 10489
rect 17313 10523 17371 10529
rect 17313 10489 17325 10523
rect 17359 10520 17371 10523
rect 17678 10520 17684 10532
rect 17359 10492 17684 10520
rect 17359 10489 17371 10492
rect 17313 10483 17371 10489
rect 17678 10480 17684 10492
rect 17736 10480 17742 10532
rect 17862 10520 17868 10532
rect 17823 10492 17868 10520
rect 17862 10480 17868 10492
rect 17920 10480 17926 10532
rect 18064 10529 18092 10560
rect 18432 10532 18460 10628
rect 18049 10523 18107 10529
rect 18049 10489 18061 10523
rect 18095 10520 18107 10523
rect 18138 10520 18144 10532
rect 18095 10492 18144 10520
rect 18095 10489 18107 10492
rect 18049 10483 18107 10489
rect 18138 10480 18144 10492
rect 18196 10480 18202 10532
rect 18414 10520 18420 10532
rect 18375 10492 18420 10520
rect 18414 10480 18420 10492
rect 18472 10480 18478 10532
rect 11793 10455 11851 10461
rect 11793 10421 11805 10455
rect 11839 10421 11851 10455
rect 11793 10415 11851 10421
rect 12253 10455 12311 10461
rect 12253 10421 12265 10455
rect 12299 10452 12311 10455
rect 12621 10455 12679 10461
rect 12621 10452 12633 10455
rect 12299 10424 12633 10452
rect 12299 10421 12311 10424
rect 12253 10415 12311 10421
rect 12621 10421 12633 10424
rect 12667 10421 12679 10455
rect 12621 10415 12679 10421
rect 13081 10455 13139 10461
rect 13081 10421 13093 10455
rect 13127 10452 13139 10455
rect 13170 10452 13176 10464
rect 13127 10424 13176 10452
rect 13127 10421 13139 10424
rect 13081 10415 13139 10421
rect 13170 10412 13176 10424
rect 13228 10412 13234 10464
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 16574 10452 16580 10464
rect 13780 10424 16580 10452
rect 13780 10412 13786 10424
rect 16574 10412 16580 10424
rect 16632 10412 16638 10464
rect 16942 10452 16948 10464
rect 16903 10424 16948 10452
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 17405 10455 17463 10461
rect 17405 10421 17417 10455
rect 17451 10452 17463 10455
rect 17586 10452 17592 10464
rect 17451 10424 17592 10452
rect 17451 10421 17463 10424
rect 17405 10415 17463 10421
rect 17586 10412 17592 10424
rect 17644 10412 17650 10464
rect 17770 10412 17776 10464
rect 17828 10452 17834 10464
rect 18325 10455 18383 10461
rect 18325 10452 18337 10455
rect 17828 10424 18337 10452
rect 17828 10412 17834 10424
rect 18325 10421 18337 10424
rect 18371 10421 18383 10455
rect 18325 10415 18383 10421
rect 1104 10362 18860 10384
rect 1104 10310 6912 10362
rect 6964 10310 6976 10362
rect 7028 10310 7040 10362
rect 7092 10310 7104 10362
rect 7156 10310 12843 10362
rect 12895 10310 12907 10362
rect 12959 10310 12971 10362
rect 13023 10310 13035 10362
rect 13087 10310 18860 10362
rect 1104 10288 18860 10310
rect 1854 10248 1860 10260
rect 1815 10220 1860 10248
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 1946 10208 1952 10260
rect 2004 10248 2010 10260
rect 2004 10220 2049 10248
rect 2004 10208 2010 10220
rect 2314 10208 2320 10260
rect 2372 10248 2378 10260
rect 2409 10251 2467 10257
rect 2409 10248 2421 10251
rect 2372 10220 2421 10248
rect 2372 10208 2378 10220
rect 2409 10217 2421 10220
rect 2455 10217 2467 10251
rect 2866 10248 2872 10260
rect 2827 10220 2872 10248
rect 2409 10211 2467 10217
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 3418 10248 3424 10260
rect 3379 10220 3424 10248
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 3510 10208 3516 10260
rect 3568 10248 3574 10260
rect 3694 10248 3700 10260
rect 3568 10220 3700 10248
rect 3568 10208 3574 10220
rect 3694 10208 3700 10220
rect 3752 10208 3758 10260
rect 4890 10248 4896 10260
rect 4851 10220 4896 10248
rect 4890 10208 4896 10220
rect 4948 10208 4954 10260
rect 5261 10251 5319 10257
rect 5261 10217 5273 10251
rect 5307 10217 5319 10251
rect 5261 10211 5319 10217
rect 5629 10251 5687 10257
rect 5629 10217 5641 10251
rect 5675 10248 5687 10251
rect 6089 10251 6147 10257
rect 6089 10248 6101 10251
rect 5675 10220 6101 10248
rect 5675 10217 5687 10220
rect 5629 10211 5687 10217
rect 6089 10217 6101 10220
rect 6135 10217 6147 10251
rect 6089 10211 6147 10217
rect 4614 10180 4620 10192
rect 1780 10152 4620 10180
rect 1780 10053 1808 10152
rect 4614 10140 4620 10152
rect 4672 10140 4678 10192
rect 4801 10183 4859 10189
rect 4801 10149 4813 10183
rect 4847 10180 4859 10183
rect 5276 10180 5304 10211
rect 6362 10208 6368 10260
rect 6420 10248 6426 10260
rect 6549 10251 6607 10257
rect 6549 10248 6561 10251
rect 6420 10220 6561 10248
rect 6420 10208 6426 10220
rect 6549 10217 6561 10220
rect 6595 10248 6607 10251
rect 8202 10248 8208 10260
rect 6595 10220 8208 10248
rect 6595 10217 6607 10220
rect 6549 10211 6607 10217
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 9861 10251 9919 10257
rect 9861 10217 9873 10251
rect 9907 10248 9919 10251
rect 10413 10251 10471 10257
rect 10413 10248 10425 10251
rect 9907 10220 10425 10248
rect 9907 10217 9919 10220
rect 9861 10211 9919 10217
rect 10413 10217 10425 10220
rect 10459 10217 10471 10251
rect 10870 10248 10876 10260
rect 10831 10220 10876 10248
rect 10413 10211 10471 10217
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 11241 10251 11299 10257
rect 11241 10217 11253 10251
rect 11287 10217 11299 10251
rect 11241 10211 11299 10217
rect 4847 10152 5304 10180
rect 5721 10183 5779 10189
rect 4847 10149 4859 10152
rect 4801 10143 4859 10149
rect 5721 10149 5733 10183
rect 5767 10180 5779 10183
rect 5994 10180 6000 10192
rect 5767 10152 6000 10180
rect 5767 10149 5779 10152
rect 5721 10143 5779 10149
rect 5994 10140 6000 10152
rect 6052 10140 6058 10192
rect 7806 10183 7864 10189
rect 7806 10180 7818 10183
rect 6380 10152 7818 10180
rect 2777 10115 2835 10121
rect 2777 10081 2789 10115
rect 2823 10112 2835 10115
rect 3694 10112 3700 10124
rect 2823 10084 3700 10112
rect 2823 10081 2835 10084
rect 2777 10075 2835 10081
rect 3694 10072 3700 10084
rect 3752 10072 3758 10124
rect 3878 10072 3884 10124
rect 3936 10112 3942 10124
rect 3973 10115 4031 10121
rect 3973 10112 3985 10115
rect 3936 10084 3985 10112
rect 3936 10072 3942 10084
rect 3973 10081 3985 10084
rect 4019 10112 4031 10115
rect 6380 10112 6408 10152
rect 7806 10149 7818 10152
rect 7852 10180 7864 10183
rect 8754 10180 8760 10192
rect 7852 10152 8760 10180
rect 7852 10149 7864 10152
rect 7806 10143 7864 10149
rect 8754 10140 8760 10152
rect 8812 10140 8818 10192
rect 9953 10183 10011 10189
rect 9953 10149 9965 10183
rect 9999 10180 10011 10183
rect 11256 10180 11284 10211
rect 11606 10208 11612 10260
rect 11664 10248 11670 10260
rect 11701 10251 11759 10257
rect 11701 10248 11713 10251
rect 11664 10220 11713 10248
rect 11664 10208 11670 10220
rect 11701 10217 11713 10220
rect 11747 10248 11759 10251
rect 12066 10248 12072 10260
rect 11747 10220 12072 10248
rect 11747 10217 11759 10220
rect 11701 10211 11759 10217
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 12342 10248 12348 10260
rect 12255 10220 12348 10248
rect 12342 10208 12348 10220
rect 12400 10248 12406 10260
rect 12897 10251 12955 10257
rect 12897 10248 12909 10251
rect 12400 10220 12909 10248
rect 12400 10208 12406 10220
rect 12897 10217 12909 10220
rect 12943 10248 12955 10251
rect 13538 10248 13544 10260
rect 12943 10220 13544 10248
rect 12943 10217 12955 10220
rect 12897 10211 12955 10217
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 13722 10248 13728 10260
rect 13683 10220 13728 10248
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 16482 10208 16488 10260
rect 16540 10248 16546 10260
rect 16577 10251 16635 10257
rect 16577 10248 16589 10251
rect 16540 10220 16589 10248
rect 16540 10208 16546 10220
rect 16577 10217 16589 10220
rect 16623 10217 16635 10251
rect 16577 10211 16635 10217
rect 16666 10208 16672 10260
rect 16724 10248 16730 10260
rect 17221 10251 17279 10257
rect 17221 10248 17233 10251
rect 16724 10220 17233 10248
rect 16724 10208 16730 10220
rect 17221 10217 17233 10220
rect 17267 10217 17279 10251
rect 17586 10248 17592 10260
rect 17547 10220 17592 10248
rect 17221 10211 17279 10217
rect 17586 10208 17592 10220
rect 17644 10208 17650 10260
rect 17678 10208 17684 10260
rect 17736 10248 17742 10260
rect 18046 10248 18052 10260
rect 17736 10220 17781 10248
rect 18007 10220 18052 10248
rect 17736 10208 17742 10220
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 17954 10180 17960 10192
rect 9999 10152 11284 10180
rect 11348 10152 17960 10180
rect 9999 10149 10011 10152
rect 9953 10143 10011 10149
rect 4019 10084 5028 10112
rect 4019 10081 4031 10084
rect 3973 10075 4031 10081
rect 1765 10047 1823 10053
rect 1765 10013 1777 10047
rect 1811 10013 1823 10047
rect 2958 10044 2964 10056
rect 2919 10016 2964 10044
rect 1765 10007 1823 10013
rect 2958 10004 2964 10016
rect 3016 10004 3022 10056
rect 3786 10004 3792 10056
rect 3844 10044 3850 10056
rect 3844 10016 4568 10044
rect 3844 10004 3850 10016
rect 2317 9979 2375 9985
rect 2317 9945 2329 9979
rect 2363 9976 2375 9979
rect 2363 9948 2544 9976
rect 2363 9945 2375 9948
rect 2317 9939 2375 9945
rect 1394 9908 1400 9920
rect 1355 9880 1400 9908
rect 1394 9868 1400 9880
rect 1452 9868 1458 9920
rect 2516 9908 2544 9948
rect 3050 9908 3056 9920
rect 2516 9880 3056 9908
rect 3050 9868 3056 9880
rect 3108 9868 3114 9920
rect 3234 9908 3240 9920
rect 3195 9880 3240 9908
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 4338 9868 4344 9920
rect 4396 9908 4402 9920
rect 4433 9911 4491 9917
rect 4433 9908 4445 9911
rect 4396 9880 4445 9908
rect 4396 9868 4402 9880
rect 4433 9877 4445 9880
rect 4479 9877 4491 9911
rect 4540 9908 4568 10016
rect 5000 9976 5028 10084
rect 5092 10084 6408 10112
rect 6457 10115 6515 10121
rect 5092 10053 5120 10084
rect 6457 10081 6469 10115
rect 6503 10112 6515 10115
rect 6917 10115 6975 10121
rect 6917 10112 6929 10115
rect 6503 10084 6929 10112
rect 6503 10081 6515 10084
rect 6457 10075 6515 10081
rect 6917 10081 6929 10084
rect 6963 10081 6975 10115
rect 6917 10075 6975 10081
rect 7282 10072 7288 10124
rect 7340 10112 7346 10124
rect 7561 10115 7619 10121
rect 7561 10112 7573 10115
rect 7340 10084 7573 10112
rect 7340 10072 7346 10084
rect 7561 10081 7573 10084
rect 7607 10081 7619 10115
rect 10686 10112 10692 10124
rect 7561 10075 7619 10081
rect 7668 10084 10692 10112
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10013 5135 10047
rect 5902 10044 5908 10056
rect 5863 10016 5908 10044
rect 5077 10007 5135 10013
rect 5902 10004 5908 10016
rect 5960 10004 5966 10056
rect 6638 10044 6644 10056
rect 6599 10016 6644 10044
rect 6638 10004 6644 10016
rect 6696 10004 6702 10056
rect 7668 10044 7696 10084
rect 10686 10072 10692 10084
rect 10744 10112 10750 10124
rect 10781 10115 10839 10121
rect 10781 10112 10793 10115
rect 10744 10084 10793 10112
rect 10744 10072 10750 10084
rect 10781 10081 10793 10084
rect 10827 10081 10839 10115
rect 11348 10112 11376 10152
rect 17954 10140 17960 10152
rect 18012 10140 18018 10192
rect 11606 10112 11612 10124
rect 10781 10075 10839 10081
rect 10980 10084 11376 10112
rect 11567 10084 11612 10112
rect 9766 10044 9772 10056
rect 6840 10016 7696 10044
rect 9727 10016 9772 10044
rect 6362 9976 6368 9988
rect 5000 9948 6368 9976
rect 6362 9936 6368 9948
rect 6420 9936 6426 9988
rect 6840 9908 6868 10016
rect 9766 10004 9772 10016
rect 9824 10004 9830 10056
rect 10980 9976 11008 10084
rect 11606 10072 11612 10084
rect 11664 10072 11670 10124
rect 11882 10072 11888 10124
rect 11940 10112 11946 10124
rect 12805 10115 12863 10121
rect 12805 10112 12817 10115
rect 11940 10084 12817 10112
rect 11940 10072 11946 10084
rect 12805 10081 12817 10084
rect 12851 10112 12863 10115
rect 12851 10084 13032 10112
rect 12851 10081 12863 10084
rect 12805 10075 12863 10081
rect 11057 10047 11115 10053
rect 11057 10013 11069 10047
rect 11103 10013 11115 10047
rect 11057 10007 11115 10013
rect 11793 10047 11851 10053
rect 11793 10013 11805 10047
rect 11839 10013 11851 10047
rect 11793 10007 11851 10013
rect 8496 9948 11008 9976
rect 11072 9976 11100 10007
rect 11698 9976 11704 9988
rect 11072 9948 11704 9976
rect 4540 9880 6868 9908
rect 4433 9871 4491 9877
rect 7190 9868 7196 9920
rect 7248 9908 7254 9920
rect 7285 9911 7343 9917
rect 7285 9908 7297 9911
rect 7248 9880 7297 9908
rect 7248 9868 7254 9880
rect 7285 9877 7297 9880
rect 7331 9908 7343 9911
rect 7374 9908 7380 9920
rect 7331 9880 7380 9908
rect 7331 9877 7343 9880
rect 7285 9871 7343 9877
rect 7374 9868 7380 9880
rect 7432 9908 7438 9920
rect 8496 9908 8524 9948
rect 11698 9936 11704 9948
rect 11756 9976 11762 9988
rect 11808 9976 11836 10007
rect 12250 9976 12256 9988
rect 11756 9948 12256 9976
rect 11756 9936 11762 9948
rect 12250 9936 12256 9948
rect 12308 9936 12314 9988
rect 7432 9880 8524 9908
rect 7432 9868 7438 9880
rect 8846 9868 8852 9920
rect 8904 9908 8910 9920
rect 8941 9911 8999 9917
rect 8941 9908 8953 9911
rect 8904 9880 8953 9908
rect 8904 9868 8910 9880
rect 8941 9877 8953 9880
rect 8987 9877 8999 9911
rect 10318 9908 10324 9920
rect 10279 9880 10324 9908
rect 8941 9871 8999 9877
rect 10318 9868 10324 9880
rect 10376 9868 10382 9920
rect 10870 9868 10876 9920
rect 10928 9908 10934 9920
rect 12069 9911 12127 9917
rect 12069 9908 12081 9911
rect 10928 9880 12081 9908
rect 10928 9868 10934 9880
rect 12069 9877 12081 9880
rect 12115 9877 12127 9911
rect 12069 9871 12127 9877
rect 12437 9911 12495 9917
rect 12437 9877 12449 9911
rect 12483 9908 12495 9911
rect 12526 9908 12532 9920
rect 12483 9880 12532 9908
rect 12483 9877 12495 9880
rect 12437 9871 12495 9877
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 13004 9908 13032 10084
rect 14918 10072 14924 10124
rect 14976 10112 14982 10124
rect 15197 10115 15255 10121
rect 15197 10112 15209 10115
rect 14976 10084 15209 10112
rect 14976 10072 14982 10084
rect 15197 10081 15209 10084
rect 15243 10081 15255 10115
rect 15197 10075 15255 10081
rect 15464 10115 15522 10121
rect 15464 10081 15476 10115
rect 15510 10112 15522 10115
rect 17586 10112 17592 10124
rect 15510 10084 17592 10112
rect 15510 10081 15522 10084
rect 15464 10075 15522 10081
rect 13081 10047 13139 10053
rect 13081 10013 13093 10047
rect 13127 10044 13139 10047
rect 13262 10044 13268 10056
rect 13127 10016 13268 10044
rect 13127 10013 13139 10016
rect 13081 10007 13139 10013
rect 13262 10004 13268 10016
rect 13320 10004 13326 10056
rect 13170 9936 13176 9988
rect 13228 9976 13234 9988
rect 13357 9979 13415 9985
rect 13357 9976 13369 9979
rect 13228 9948 13369 9976
rect 13228 9936 13234 9948
rect 13357 9945 13369 9948
rect 13403 9976 13415 9979
rect 13814 9976 13820 9988
rect 13403 9948 13820 9976
rect 13403 9945 13415 9948
rect 13357 9939 13415 9945
rect 13814 9936 13820 9948
rect 13872 9936 13878 9988
rect 13541 9911 13599 9917
rect 13541 9908 13553 9911
rect 13004 9880 13553 9908
rect 13541 9877 13553 9880
rect 13587 9908 13599 9911
rect 13906 9908 13912 9920
rect 13587 9880 13912 9908
rect 13587 9877 13599 9880
rect 13541 9871 13599 9877
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 15212 9908 15240 10075
rect 16960 10053 16988 10084
rect 17586 10072 17592 10084
rect 17644 10112 17650 10124
rect 18141 10115 18199 10121
rect 17644 10084 18092 10112
rect 17644 10072 17650 10084
rect 16945 10047 17003 10053
rect 16945 10013 16957 10047
rect 16991 10013 17003 10047
rect 17126 10044 17132 10056
rect 17087 10016 17132 10044
rect 16945 10007 17003 10013
rect 17126 10004 17132 10016
rect 17184 10004 17190 10056
rect 18064 10044 18092 10084
rect 18141 10081 18153 10115
rect 18187 10112 18199 10115
rect 18187 10084 18368 10112
rect 18187 10081 18199 10084
rect 18141 10075 18199 10081
rect 18233 10047 18291 10053
rect 18233 10044 18245 10047
rect 18064 10016 18245 10044
rect 18233 10013 18245 10016
rect 18279 10013 18291 10047
rect 18233 10007 18291 10013
rect 17310 9976 17316 9988
rect 16132 9948 17316 9976
rect 16132 9920 16160 9948
rect 17310 9936 17316 9948
rect 17368 9976 17374 9988
rect 18340 9976 18368 10084
rect 17368 9948 18368 9976
rect 17368 9936 17374 9948
rect 15378 9908 15384 9920
rect 15212 9880 15384 9908
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 16114 9868 16120 9920
rect 16172 9868 16178 9920
rect 16758 9908 16764 9920
rect 16719 9880 16764 9908
rect 16758 9868 16764 9880
rect 16816 9868 16822 9920
rect 1104 9818 18860 9840
rect 1104 9766 3947 9818
rect 3999 9766 4011 9818
rect 4063 9766 4075 9818
rect 4127 9766 4139 9818
rect 4191 9766 9878 9818
rect 9930 9766 9942 9818
rect 9994 9766 10006 9818
rect 10058 9766 10070 9818
rect 10122 9766 15808 9818
rect 15860 9766 15872 9818
rect 15924 9766 15936 9818
rect 15988 9766 16000 9818
rect 16052 9766 18860 9818
rect 1104 9744 18860 9766
rect 1578 9664 1584 9716
rect 1636 9704 1642 9716
rect 5442 9704 5448 9716
rect 1636 9676 5304 9704
rect 5403 9676 5448 9704
rect 1636 9664 1642 9676
rect 3510 9636 3516 9648
rect 2332 9608 3516 9636
rect 1765 9503 1823 9509
rect 1765 9469 1777 9503
rect 1811 9500 1823 9503
rect 2130 9500 2136 9512
rect 1811 9472 2136 9500
rect 1811 9469 1823 9472
rect 1765 9463 1823 9469
rect 2130 9460 2136 9472
rect 2188 9460 2194 9512
rect 2332 9509 2360 9608
rect 3510 9596 3516 9608
rect 3568 9596 3574 9648
rect 5276 9636 5304 9676
rect 5442 9664 5448 9676
rect 5500 9664 5506 9716
rect 5718 9664 5724 9716
rect 5776 9704 5782 9716
rect 7190 9704 7196 9716
rect 5776 9676 7196 9704
rect 5776 9664 5782 9676
rect 7190 9664 7196 9676
rect 7248 9664 7254 9716
rect 8662 9664 8668 9716
rect 8720 9704 8726 9716
rect 8849 9707 8907 9713
rect 8849 9704 8861 9707
rect 8720 9676 8861 9704
rect 8720 9664 8726 9676
rect 8849 9673 8861 9676
rect 8895 9704 8907 9707
rect 8941 9707 8999 9713
rect 8941 9704 8953 9707
rect 8895 9676 8953 9704
rect 8895 9673 8907 9676
rect 8849 9667 8907 9673
rect 8941 9673 8953 9676
rect 8987 9673 8999 9707
rect 9122 9704 9128 9716
rect 9083 9676 9128 9704
rect 8941 9667 8999 9673
rect 9122 9664 9128 9676
rect 9180 9664 9186 9716
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 9824 9676 10640 9704
rect 9824 9664 9830 9676
rect 5994 9636 6000 9648
rect 3620 9608 4108 9636
rect 5276 9608 6000 9636
rect 3326 9528 3332 9580
rect 3384 9568 3390 9580
rect 3421 9571 3479 9577
rect 3421 9568 3433 9571
rect 3384 9540 3433 9568
rect 3384 9528 3390 9540
rect 3421 9537 3433 9540
rect 3467 9568 3479 9571
rect 3620 9568 3648 9608
rect 3467 9540 3648 9568
rect 4080 9568 4108 9608
rect 5994 9596 6000 9608
rect 6052 9596 6058 9648
rect 6638 9636 6644 9648
rect 6104 9608 6644 9636
rect 6104 9577 6132 9608
rect 6638 9596 6644 9608
rect 6696 9596 6702 9648
rect 7377 9639 7435 9645
rect 7377 9605 7389 9639
rect 7423 9636 7435 9639
rect 8202 9636 8208 9648
rect 7423 9608 8208 9636
rect 7423 9605 7435 9608
rect 7377 9599 7435 9605
rect 8202 9596 8208 9608
rect 8260 9596 8266 9648
rect 8294 9596 8300 9648
rect 8352 9636 8358 9648
rect 10134 9636 10140 9648
rect 8352 9608 10140 9636
rect 8352 9596 8358 9608
rect 10134 9596 10140 9608
rect 10192 9596 10198 9648
rect 10226 9596 10232 9648
rect 10284 9636 10290 9648
rect 10612 9636 10640 9676
rect 10686 9664 10692 9716
rect 10744 9704 10750 9716
rect 16390 9704 16396 9716
rect 10744 9676 16396 9704
rect 10744 9664 10750 9676
rect 16390 9664 16396 9676
rect 16448 9664 16454 9716
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 17770 9704 17776 9716
rect 16632 9676 17776 9704
rect 16632 9664 16638 9676
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 15654 9636 15660 9648
rect 10284 9608 10548 9636
rect 10612 9608 12388 9636
rect 15615 9608 15660 9636
rect 10284 9596 10290 9608
rect 4249 9571 4307 9577
rect 4249 9568 4261 9571
rect 4080 9540 4261 9568
rect 3467 9537 3479 9540
rect 3421 9531 3479 9537
rect 4249 9537 4261 9540
rect 4295 9537 4307 9571
rect 4249 9531 4307 9537
rect 6089 9571 6147 9577
rect 6089 9537 6101 9571
rect 6135 9537 6147 9571
rect 6089 9531 6147 9537
rect 6546 9528 6552 9580
rect 6604 9568 6610 9580
rect 7009 9571 7067 9577
rect 7009 9568 7021 9571
rect 6604 9540 7021 9568
rect 6604 9528 6610 9540
rect 7009 9537 7021 9540
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 8846 9528 8852 9580
rect 8904 9568 8910 9580
rect 9677 9571 9735 9577
rect 9677 9568 9689 9571
rect 8904 9540 9689 9568
rect 8904 9528 8910 9540
rect 9677 9537 9689 9540
rect 9723 9537 9735 9571
rect 10410 9568 10416 9580
rect 10371 9540 10416 9568
rect 9677 9531 9735 9537
rect 10410 9528 10416 9540
rect 10468 9528 10474 9580
rect 10520 9577 10548 9608
rect 10505 9571 10563 9577
rect 10505 9537 10517 9571
rect 10551 9537 10563 9571
rect 10505 9531 10563 9537
rect 11057 9571 11115 9577
rect 11057 9537 11069 9571
rect 11103 9568 11115 9571
rect 11606 9568 11612 9580
rect 11103 9540 11612 9568
rect 11103 9537 11115 9540
rect 11057 9531 11115 9537
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 12066 9568 12072 9580
rect 12027 9540 12072 9568
rect 12066 9528 12072 9540
rect 12124 9528 12130 9580
rect 12360 9577 12388 9608
rect 15654 9596 15660 9608
rect 15712 9596 15718 9648
rect 15841 9639 15899 9645
rect 15841 9605 15853 9639
rect 15887 9636 15899 9639
rect 18046 9636 18052 9648
rect 15887 9608 18052 9636
rect 15887 9605 15899 9608
rect 15841 9599 15899 9605
rect 18046 9596 18052 9608
rect 18104 9596 18110 9648
rect 12345 9571 12403 9577
rect 12345 9537 12357 9571
rect 12391 9568 12403 9571
rect 13081 9571 13139 9577
rect 12391 9540 12940 9568
rect 12391 9537 12403 9540
rect 12345 9531 12403 9537
rect 2309 9503 2367 9509
rect 2309 9469 2321 9503
rect 2355 9469 2367 9503
rect 2309 9463 2367 9469
rect 2409 9503 2467 9509
rect 2409 9469 2421 9503
rect 2455 9500 2467 9503
rect 3786 9500 3792 9512
rect 2455 9472 3792 9500
rect 2455 9469 2467 9472
rect 2409 9463 2467 9469
rect 3786 9460 3792 9472
rect 3844 9460 3850 9512
rect 4062 9500 4068 9512
rect 4023 9472 4068 9500
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 4709 9503 4767 9509
rect 4709 9469 4721 9503
rect 4755 9500 4767 9503
rect 8202 9500 8208 9512
rect 4755 9472 8208 9500
rect 4755 9469 4767 9472
rect 4709 9463 4767 9469
rect 8202 9460 8208 9472
rect 8260 9460 8266 9512
rect 9398 9460 9404 9512
rect 9456 9500 9462 9512
rect 9493 9503 9551 9509
rect 9493 9500 9505 9503
rect 9456 9472 9505 9500
rect 9456 9460 9462 9472
rect 9493 9469 9505 9472
rect 9539 9500 9551 9503
rect 9858 9500 9864 9512
rect 9539 9472 9864 9500
rect 9539 9469 9551 9472
rect 9493 9463 9551 9469
rect 9858 9460 9864 9472
rect 9916 9460 9922 9512
rect 10318 9500 10324 9512
rect 10279 9472 10324 9500
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 10962 9460 10968 9512
rect 11020 9500 11026 9512
rect 12618 9500 12624 9512
rect 11020 9472 12624 9500
rect 11020 9460 11026 9472
rect 12618 9460 12624 9472
rect 12676 9460 12682 9512
rect 12912 9509 12940 9540
rect 13081 9537 13093 9571
rect 13127 9568 13139 9571
rect 13262 9568 13268 9580
rect 13127 9540 13268 9568
rect 13127 9537 13139 9540
rect 13081 9531 13139 9537
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 16482 9568 16488 9580
rect 15304 9540 16488 9568
rect 12897 9503 12955 9509
rect 12897 9469 12909 9503
rect 12943 9500 12955 9503
rect 14366 9500 14372 9512
rect 12943 9472 14372 9500
rect 12943 9469 12955 9472
rect 12897 9463 12955 9469
rect 14366 9460 14372 9472
rect 14424 9460 14430 9512
rect 15125 9503 15183 9509
rect 15125 9469 15137 9503
rect 15171 9500 15183 9503
rect 15304 9500 15332 9540
rect 16482 9528 16488 9540
rect 16540 9528 16546 9580
rect 17402 9568 17408 9580
rect 16592 9540 17408 9568
rect 15171 9472 15332 9500
rect 15171 9469 15183 9472
rect 15125 9463 15183 9469
rect 15378 9460 15384 9512
rect 15436 9500 15442 9512
rect 16592 9500 16620 9540
rect 17402 9528 17408 9540
rect 17460 9528 17466 9580
rect 17586 9568 17592 9580
rect 17547 9540 17592 9568
rect 17586 9528 17592 9540
rect 17644 9528 17650 9580
rect 15436 9472 15481 9500
rect 15580 9472 16620 9500
rect 15436 9460 15442 9472
rect 1486 9432 1492 9444
rect 1447 9404 1492 9432
rect 1486 9392 1492 9404
rect 1544 9432 1550 9444
rect 2685 9435 2743 9441
rect 2685 9432 2697 9435
rect 1544 9404 2697 9432
rect 1544 9392 1550 9404
rect 2685 9401 2697 9404
rect 2731 9401 2743 9435
rect 2685 9395 2743 9401
rect 3237 9435 3295 9441
rect 3237 9401 3249 9435
rect 3283 9432 3295 9435
rect 3970 9432 3976 9444
rect 3283 9404 3976 9432
rect 3283 9401 3295 9404
rect 3237 9395 3295 9401
rect 3970 9392 3976 9404
rect 4028 9392 4034 9444
rect 4614 9432 4620 9444
rect 4356 9404 4620 9432
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 1946 9364 1952 9376
rect 1907 9336 1952 9364
rect 1946 9324 1952 9336
rect 2004 9324 2010 9376
rect 2130 9364 2136 9376
rect 2091 9336 2136 9364
rect 2130 9324 2136 9336
rect 2188 9324 2194 9376
rect 2590 9364 2596 9376
rect 2551 9336 2596 9364
rect 2590 9324 2596 9336
rect 2648 9324 2654 9376
rect 2866 9364 2872 9376
rect 2827 9336 2872 9364
rect 2866 9324 2872 9336
rect 2924 9324 2930 9376
rect 3329 9367 3387 9373
rect 3329 9333 3341 9367
rect 3375 9364 3387 9367
rect 3418 9364 3424 9376
rect 3375 9336 3424 9364
rect 3375 9333 3387 9336
rect 3329 9327 3387 9333
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 3694 9364 3700 9376
rect 3655 9336 3700 9364
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 4157 9367 4215 9373
rect 4157 9333 4169 9367
rect 4203 9364 4215 9367
rect 4356 9364 4384 9404
rect 4614 9392 4620 9404
rect 4672 9392 4678 9444
rect 5813 9435 5871 9441
rect 5813 9401 5825 9435
rect 5859 9432 5871 9435
rect 5859 9404 6316 9432
rect 5859 9401 5871 9404
rect 5813 9395 5871 9401
rect 4203 9336 4384 9364
rect 4203 9333 4215 9336
rect 4157 9327 4215 9333
rect 4430 9324 4436 9376
rect 4488 9364 4494 9376
rect 4525 9367 4583 9373
rect 4525 9364 4537 9367
rect 4488 9336 4537 9364
rect 4488 9324 4494 9336
rect 4525 9333 4537 9336
rect 4571 9333 4583 9367
rect 4890 9364 4896 9376
rect 4851 9336 4896 9364
rect 4525 9327 4583 9333
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 5902 9364 5908 9376
rect 5863 9336 5908 9364
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 6288 9364 6316 9404
rect 6362 9392 6368 9444
rect 6420 9432 6426 9444
rect 6730 9432 6736 9444
rect 6420 9404 6736 9432
rect 6420 9392 6426 9404
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 6825 9435 6883 9441
rect 6825 9401 6837 9435
rect 6871 9432 6883 9435
rect 7374 9432 7380 9444
rect 6871 9404 7380 9432
rect 6871 9401 6883 9404
rect 6825 9395 6883 9401
rect 7374 9392 7380 9404
rect 7432 9432 7438 9444
rect 7469 9435 7527 9441
rect 7469 9432 7481 9435
rect 7432 9404 7481 9432
rect 7432 9392 7438 9404
rect 7469 9401 7481 9404
rect 7515 9432 7527 9435
rect 10686 9432 10692 9444
rect 7515 9404 10692 9432
rect 7515 9401 7527 9404
rect 7469 9395 7527 9401
rect 10686 9392 10692 9404
rect 10744 9392 10750 9444
rect 13262 9432 13268 9444
rect 10980 9404 13268 9432
rect 6457 9367 6515 9373
rect 6457 9364 6469 9367
rect 6288 9336 6469 9364
rect 6457 9333 6469 9336
rect 6503 9333 6515 9367
rect 6457 9327 6515 9333
rect 6638 9324 6644 9376
rect 6696 9364 6702 9376
rect 6917 9367 6975 9373
rect 6917 9364 6929 9367
rect 6696 9336 6929 9364
rect 6696 9324 6702 9336
rect 6917 9333 6929 9336
rect 6963 9364 6975 9367
rect 8294 9364 8300 9376
rect 6963 9336 8300 9364
rect 6963 9333 6975 9336
rect 6917 9327 6975 9333
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 8849 9367 8907 9373
rect 8849 9333 8861 9367
rect 8895 9364 8907 9367
rect 9585 9367 9643 9373
rect 9585 9364 9597 9367
rect 8895 9336 9597 9364
rect 8895 9333 8907 9336
rect 8849 9327 8907 9333
rect 9585 9333 9597 9336
rect 9631 9333 9643 9367
rect 9585 9327 9643 9333
rect 9674 9324 9680 9376
rect 9732 9364 9738 9376
rect 9953 9367 10011 9373
rect 9953 9364 9965 9367
rect 9732 9336 9965 9364
rect 9732 9324 9738 9336
rect 9953 9333 9965 9336
rect 9999 9333 10011 9367
rect 9953 9327 10011 9333
rect 10134 9324 10140 9376
rect 10192 9364 10198 9376
rect 10980 9364 11008 9404
rect 13262 9392 13268 9404
rect 13320 9392 13326 9444
rect 13541 9435 13599 9441
rect 13541 9401 13553 9435
rect 13587 9432 13599 9435
rect 14734 9432 14740 9444
rect 13587 9404 14740 9432
rect 13587 9401 13599 9404
rect 13541 9395 13599 9401
rect 10192 9336 11008 9364
rect 10192 9324 10198 9336
rect 11054 9324 11060 9376
rect 11112 9364 11118 9376
rect 11149 9367 11207 9373
rect 11149 9364 11161 9367
rect 11112 9336 11161 9364
rect 11112 9324 11118 9336
rect 11149 9333 11161 9336
rect 11195 9333 11207 9367
rect 11149 9327 11207 9333
rect 11330 9324 11336 9376
rect 11388 9364 11394 9376
rect 11882 9364 11888 9376
rect 11388 9336 11888 9364
rect 11388 9324 11394 9336
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 12434 9364 12440 9376
rect 12395 9336 12440 9364
rect 12434 9324 12440 9336
rect 12492 9324 12498 9376
rect 12618 9324 12624 9376
rect 12676 9364 12682 9376
rect 12805 9367 12863 9373
rect 12805 9364 12817 9367
rect 12676 9336 12817 9364
rect 12676 9324 12682 9336
rect 12805 9333 12817 9336
rect 12851 9364 12863 9367
rect 13556 9364 13584 9395
rect 14734 9392 14740 9404
rect 14792 9392 14798 9444
rect 15010 9392 15016 9444
rect 15068 9432 15074 9444
rect 15580 9432 15608 9472
rect 16758 9460 16764 9512
rect 16816 9500 16822 9512
rect 16816 9472 18460 9500
rect 16816 9460 16822 9472
rect 18432 9444 18460 9472
rect 15068 9404 15608 9432
rect 16301 9435 16359 9441
rect 15068 9392 15074 9404
rect 16301 9401 16313 9435
rect 16347 9432 16359 9435
rect 17310 9432 17316 9444
rect 16347 9404 16988 9432
rect 17271 9404 17316 9432
rect 16347 9401 16359 9404
rect 16301 9395 16359 9401
rect 13998 9364 14004 9376
rect 12851 9336 13584 9364
rect 13959 9336 14004 9364
rect 12851 9333 12863 9336
rect 12805 9327 12863 9333
rect 13998 9324 14004 9336
rect 14056 9324 14062 9376
rect 15930 9364 15936 9376
rect 15891 9336 15936 9364
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 16206 9324 16212 9376
rect 16264 9364 16270 9376
rect 16960 9373 16988 9404
rect 17310 9392 17316 9404
rect 17368 9392 17374 9444
rect 17862 9432 17868 9444
rect 17823 9404 17868 9432
rect 17862 9392 17868 9404
rect 17920 9392 17926 9444
rect 18046 9432 18052 9444
rect 18007 9404 18052 9432
rect 18046 9392 18052 9404
rect 18104 9392 18110 9444
rect 18138 9392 18144 9444
rect 18196 9432 18202 9444
rect 18233 9435 18291 9441
rect 18233 9432 18245 9435
rect 18196 9404 18245 9432
rect 18196 9392 18202 9404
rect 18233 9401 18245 9404
rect 18279 9401 18291 9435
rect 18414 9432 18420 9444
rect 18375 9404 18420 9432
rect 18233 9395 18291 9401
rect 18414 9392 18420 9404
rect 18472 9392 18478 9444
rect 16393 9367 16451 9373
rect 16393 9364 16405 9367
rect 16264 9336 16405 9364
rect 16264 9324 16270 9336
rect 16393 9333 16405 9336
rect 16439 9333 16451 9367
rect 16393 9327 16451 9333
rect 16945 9367 17003 9373
rect 16945 9333 16957 9367
rect 16991 9333 17003 9367
rect 16945 9327 17003 9333
rect 17402 9324 17408 9376
rect 17460 9364 17466 9376
rect 17460 9336 17505 9364
rect 17460 9324 17466 9336
rect 1104 9274 18860 9296
rect 1104 9222 6912 9274
rect 6964 9222 6976 9274
rect 7028 9222 7040 9274
rect 7092 9222 7104 9274
rect 7156 9222 12843 9274
rect 12895 9222 12907 9274
rect 12959 9222 12971 9274
rect 13023 9222 13035 9274
rect 13087 9222 18860 9274
rect 1104 9200 18860 9222
rect 3237 9163 3295 9169
rect 3237 9129 3249 9163
rect 3283 9160 3295 9163
rect 3326 9160 3332 9172
rect 3283 9132 3332 9160
rect 3283 9129 3295 9132
rect 3237 9123 3295 9129
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 3510 9120 3516 9172
rect 3568 9160 3574 9172
rect 3605 9163 3663 9169
rect 3605 9160 3617 9163
rect 3568 9132 3617 9160
rect 3568 9120 3574 9132
rect 3605 9129 3617 9132
rect 3651 9160 3663 9163
rect 4614 9160 4620 9172
rect 3651 9132 4620 9160
rect 3651 9129 3663 9132
rect 3605 9123 3663 9129
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 4706 9120 4712 9172
rect 4764 9160 4770 9172
rect 4890 9160 4896 9172
rect 4764 9132 4896 9160
rect 4764 9120 4770 9132
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 5813 9163 5871 9169
rect 5813 9129 5825 9163
rect 5859 9160 5871 9163
rect 5902 9160 5908 9172
rect 5859 9132 5908 9160
rect 5859 9129 5871 9132
rect 5813 9123 5871 9129
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 5994 9120 6000 9172
rect 6052 9160 6058 9172
rect 7742 9160 7748 9172
rect 6052 9132 7748 9160
rect 6052 9120 6058 9132
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 9950 9120 9956 9172
rect 10008 9160 10014 9172
rect 10045 9163 10103 9169
rect 10045 9160 10057 9163
rect 10008 9132 10057 9160
rect 10008 9120 10014 9132
rect 10045 9129 10057 9132
rect 10091 9129 10103 9163
rect 10962 9160 10968 9172
rect 10923 9132 10968 9160
rect 10045 9123 10103 9129
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 11238 9120 11244 9172
rect 11296 9160 11302 9172
rect 11977 9163 12035 9169
rect 11977 9160 11989 9163
rect 11296 9132 11989 9160
rect 11296 9120 11302 9132
rect 11977 9129 11989 9132
rect 12023 9129 12035 9163
rect 12434 9160 12440 9172
rect 12395 9132 12440 9160
rect 11977 9123 12035 9129
rect 12434 9120 12440 9132
rect 12492 9120 12498 9172
rect 12989 9163 13047 9169
rect 12989 9129 13001 9163
rect 13035 9160 13047 9163
rect 13081 9163 13139 9169
rect 13081 9160 13093 9163
rect 13035 9132 13093 9160
rect 13035 9129 13047 9132
rect 12989 9123 13047 9129
rect 13081 9129 13093 9132
rect 13127 9160 13139 9163
rect 14642 9160 14648 9172
rect 13127 9132 14648 9160
rect 13127 9129 13139 9132
rect 13081 9123 13139 9129
rect 14642 9120 14648 9132
rect 14700 9160 14706 9172
rect 15378 9160 15384 9172
rect 14700 9132 15384 9160
rect 14700 9120 14706 9132
rect 15378 9120 15384 9132
rect 15436 9120 15442 9172
rect 15565 9163 15623 9169
rect 15565 9129 15577 9163
rect 15611 9160 15623 9163
rect 15930 9160 15936 9172
rect 15611 9132 15936 9160
rect 15611 9129 15623 9132
rect 15565 9123 15623 9129
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 16206 9160 16212 9172
rect 16167 9132 16212 9160
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 16577 9163 16635 9169
rect 16577 9129 16589 9163
rect 16623 9160 16635 9163
rect 17037 9163 17095 9169
rect 17037 9160 17049 9163
rect 16623 9132 17049 9160
rect 16623 9129 16635 9132
rect 16577 9123 16635 9129
rect 17037 9129 17049 9132
rect 17083 9129 17095 9163
rect 17037 9123 17095 9129
rect 17405 9163 17463 9169
rect 17405 9129 17417 9163
rect 17451 9160 17463 9163
rect 17770 9160 17776 9172
rect 17451 9132 17776 9160
rect 17451 9129 17463 9132
rect 17405 9123 17463 9129
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 1578 9052 1584 9104
rect 1636 9092 1642 9104
rect 5350 9092 5356 9104
rect 1636 9064 5356 9092
rect 1636 9052 1642 9064
rect 5350 9052 5356 9064
rect 5408 9092 5414 9104
rect 5629 9095 5687 9101
rect 5629 9092 5641 9095
rect 5408 9064 5641 9092
rect 5408 9052 5414 9064
rect 5629 9061 5641 9064
rect 5675 9092 5687 9095
rect 6273 9095 6331 9101
rect 6273 9092 6285 9095
rect 5675 9064 6285 9092
rect 5675 9061 5687 9064
rect 5629 9055 5687 9061
rect 6273 9061 6285 9064
rect 6319 9061 6331 9095
rect 6638 9092 6644 9104
rect 6599 9064 6644 9092
rect 6273 9055 6331 9061
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 7552 9095 7610 9101
rect 7552 9061 7564 9095
rect 7598 9092 7610 9095
rect 8757 9095 8815 9101
rect 8757 9092 8769 9095
rect 7598 9064 8769 9092
rect 7598 9061 7610 9064
rect 7552 9055 7610 9061
rect 8757 9061 8769 9064
rect 8803 9092 8815 9095
rect 8846 9092 8852 9104
rect 8803 9064 8852 9092
rect 8803 9061 8815 9064
rect 8757 9055 8815 9061
rect 8846 9052 8852 9064
rect 8904 9052 8910 9104
rect 10980 9092 11008 9120
rect 12250 9092 12256 9104
rect 9977 9064 11008 9092
rect 11072 9064 12256 9092
rect 1394 9024 1400 9036
rect 1355 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 8984 1458 9036
rect 1670 8984 1676 9036
rect 1728 9024 1734 9036
rect 2113 9027 2171 9033
rect 2113 9024 2125 9027
rect 1728 8996 2125 9024
rect 1728 8984 1734 8996
rect 2113 8993 2125 8996
rect 2159 8993 2171 9027
rect 2113 8987 2171 8993
rect 2406 8984 2412 9036
rect 2464 9024 2470 9036
rect 6181 9027 6239 9033
rect 2464 8996 6132 9024
rect 2464 8984 2470 8996
rect 1854 8956 1860 8968
rect 1815 8928 1860 8956
rect 1854 8916 1860 8928
rect 1912 8916 1918 8968
rect 3418 8956 3424 8968
rect 3379 8928 3424 8956
rect 3418 8916 3424 8928
rect 3476 8916 3482 8968
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 3436 8820 3464 8916
rect 3970 8888 3976 8900
rect 3931 8860 3976 8888
rect 3970 8848 3976 8860
rect 4028 8848 4034 8900
rect 6104 8888 6132 8996
rect 6181 8993 6193 9027
rect 6227 9024 6239 9027
rect 6362 9024 6368 9036
rect 6227 8996 6368 9024
rect 6227 8993 6239 8996
rect 6181 8987 6239 8993
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 7282 9024 7288 9036
rect 7243 8996 7288 9024
rect 7282 8984 7288 8996
rect 7340 9024 7346 9036
rect 7834 9024 7840 9036
rect 7340 8996 7840 9024
rect 7340 8984 7346 8996
rect 7834 8984 7840 8996
rect 7892 8984 7898 9036
rect 9582 9024 9588 9036
rect 9495 8996 9588 9024
rect 9582 8984 9588 8996
rect 9640 9024 9646 9036
rect 9977 9024 10005 9064
rect 9640 8996 10005 9024
rect 9640 8984 9646 8996
rect 10318 8984 10324 9036
rect 10376 9024 10382 9036
rect 10413 9027 10471 9033
rect 10413 9024 10425 9027
rect 10376 8996 10425 9024
rect 10376 8984 10382 8996
rect 10413 8993 10425 8996
rect 10459 8993 10471 9027
rect 10413 8987 10471 8993
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 9024 10563 9027
rect 10962 9024 10968 9036
rect 10551 8996 10968 9024
rect 10551 8993 10563 8996
rect 10505 8987 10563 8993
rect 10962 8984 10968 8996
rect 11020 9024 11026 9036
rect 11072 9024 11100 9064
rect 12250 9052 12256 9064
rect 12308 9052 12314 9104
rect 12345 9095 12403 9101
rect 12345 9061 12357 9095
rect 12391 9092 12403 9095
rect 12526 9092 12532 9104
rect 12391 9064 12532 9092
rect 12391 9061 12403 9064
rect 12345 9055 12403 9061
rect 12526 9052 12532 9064
rect 12584 9052 12590 9104
rect 13262 9052 13268 9104
rect 13320 9092 13326 9104
rect 13633 9095 13691 9101
rect 13633 9092 13645 9095
rect 13320 9064 13645 9092
rect 13320 9052 13326 9064
rect 13633 9061 13645 9064
rect 13679 9092 13691 9095
rect 15654 9092 15660 9104
rect 13679 9064 15660 9092
rect 13679 9061 13691 9064
rect 13633 9055 13691 9061
rect 15654 9052 15660 9064
rect 15712 9052 15718 9104
rect 16117 9095 16175 9101
rect 16117 9061 16129 9095
rect 16163 9092 16175 9095
rect 16163 9064 18460 9092
rect 16163 9061 16175 9064
rect 16117 9055 16175 9061
rect 18432 9036 18460 9064
rect 11020 8996 11100 9024
rect 11020 8984 11026 8996
rect 11882 8984 11888 9036
rect 11940 9024 11946 9036
rect 12805 9027 12863 9033
rect 12805 9024 12817 9027
rect 11940 8996 12817 9024
rect 11940 8984 11946 8996
rect 12805 8993 12817 8996
rect 12851 8993 12863 9027
rect 12805 8987 12863 8993
rect 13541 9027 13599 9033
rect 13541 8993 13553 9027
rect 13587 8993 13599 9027
rect 13541 8987 13599 8993
rect 15473 9027 15531 9033
rect 15473 8993 15485 9027
rect 15519 9024 15531 9027
rect 16942 9024 16948 9036
rect 15519 8996 16948 9024
rect 15519 8993 15531 8996
rect 15473 8987 15531 8993
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8956 6515 8959
rect 6546 8956 6552 8968
rect 6503 8928 6552 8956
rect 6503 8925 6515 8928
rect 6457 8919 6515 8925
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8720 8928 8953 8956
rect 8720 8916 8726 8928
rect 8941 8925 8953 8928
rect 8987 8956 8999 8959
rect 9677 8959 9735 8965
rect 9677 8956 9689 8959
rect 8987 8928 9689 8956
rect 8987 8925 8999 8928
rect 8941 8919 8999 8925
rect 9677 8925 9689 8928
rect 9723 8956 9735 8959
rect 9766 8956 9772 8968
rect 9723 8928 9772 8956
rect 9723 8925 9735 8928
rect 9677 8919 9735 8925
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 10597 8959 10655 8965
rect 10597 8925 10609 8959
rect 10643 8925 10655 8959
rect 10597 8919 10655 8925
rect 8757 8891 8815 8897
rect 6104 8860 7328 8888
rect 3786 8820 3792 8832
rect 1627 8792 3792 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 3786 8780 3792 8792
rect 3844 8780 3850 8832
rect 7300 8820 7328 8860
rect 8757 8857 8769 8891
rect 8803 8888 8815 8891
rect 9876 8888 9904 8919
rect 10612 8888 10640 8919
rect 11606 8916 11612 8968
rect 11664 8956 11670 8968
rect 12529 8959 12587 8965
rect 12529 8956 12541 8959
rect 11664 8928 12541 8956
rect 11664 8916 11670 8928
rect 12529 8925 12541 8928
rect 12575 8925 12587 8959
rect 13556 8956 13584 8987
rect 16942 8984 16948 8996
rect 17000 8984 17006 9036
rect 17678 9024 17684 9036
rect 17052 8996 17684 9024
rect 12529 8919 12587 8925
rect 12636 8928 13584 8956
rect 8803 8860 10640 8888
rect 8803 8857 8815 8860
rect 8757 8851 8815 8857
rect 10686 8848 10692 8900
rect 10744 8888 10750 8900
rect 12636 8888 12664 8928
rect 10744 8860 12664 8888
rect 10744 8848 10750 8860
rect 12802 8848 12808 8900
rect 12860 8888 12866 8900
rect 13173 8891 13231 8897
rect 13173 8888 13185 8891
rect 12860 8860 13185 8888
rect 12860 8848 12866 8860
rect 13173 8857 13185 8860
rect 13219 8857 13231 8891
rect 13556 8888 13584 8928
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 13780 8928 13825 8956
rect 13780 8916 13786 8928
rect 13998 8916 14004 8968
rect 14056 8956 14062 8968
rect 15657 8959 15715 8965
rect 15657 8956 15669 8959
rect 14056 8928 15669 8956
rect 14056 8916 14062 8928
rect 15657 8925 15669 8928
rect 15703 8925 15715 8959
rect 16482 8956 16488 8968
rect 15657 8919 15715 8925
rect 15764 8928 16488 8956
rect 14093 8891 14151 8897
rect 14093 8888 14105 8891
rect 13556 8860 14105 8888
rect 13173 8851 13231 8857
rect 14093 8857 14105 8860
rect 14139 8888 14151 8891
rect 15013 8891 15071 8897
rect 15013 8888 15025 8891
rect 14139 8860 15025 8888
rect 14139 8857 14151 8860
rect 14093 8851 14151 8857
rect 15013 8857 15025 8860
rect 15059 8888 15071 8891
rect 15764 8888 15792 8928
rect 16482 8916 16488 8928
rect 16540 8916 16546 8968
rect 16666 8956 16672 8968
rect 16627 8928 16672 8956
rect 16666 8916 16672 8928
rect 16724 8916 16730 8968
rect 16853 8959 16911 8965
rect 16853 8925 16865 8959
rect 16899 8956 16911 8959
rect 17052 8956 17080 8996
rect 17678 8984 17684 8996
rect 17736 8984 17742 9036
rect 17865 9027 17923 9033
rect 17865 8993 17877 9027
rect 17911 8993 17923 9027
rect 18414 9024 18420 9036
rect 18375 8996 18420 9024
rect 17865 8987 17923 8993
rect 16899 8928 17080 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 15059 8860 15792 8888
rect 15059 8857 15071 8860
rect 15013 8851 15071 8857
rect 16206 8848 16212 8900
rect 16264 8888 16270 8900
rect 16868 8888 16896 8919
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 17497 8959 17555 8965
rect 17497 8956 17509 8959
rect 17368 8928 17509 8956
rect 17368 8916 17374 8928
rect 17497 8925 17509 8928
rect 17543 8925 17555 8959
rect 17497 8919 17555 8925
rect 17586 8916 17592 8968
rect 17644 8956 17650 8968
rect 17644 8928 17689 8956
rect 17644 8916 17650 8928
rect 16264 8860 16896 8888
rect 16264 8848 16270 8860
rect 8018 8820 8024 8832
rect 7300 8792 8024 8820
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 8662 8820 8668 8832
rect 8623 8792 8668 8820
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 9030 8780 9036 8832
rect 9088 8820 9094 8832
rect 9217 8823 9275 8829
rect 9217 8820 9229 8823
rect 9088 8792 9229 8820
rect 9088 8780 9094 8792
rect 9217 8789 9229 8792
rect 9263 8789 9275 8823
rect 9217 8783 9275 8789
rect 9306 8780 9312 8832
rect 9364 8820 9370 8832
rect 9674 8820 9680 8832
rect 9364 8792 9680 8820
rect 9364 8780 9370 8792
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 10410 8780 10416 8832
rect 10468 8820 10474 8832
rect 11057 8823 11115 8829
rect 11057 8820 11069 8823
rect 10468 8792 11069 8820
rect 10468 8780 10474 8792
rect 11057 8789 11069 8792
rect 11103 8820 11115 8823
rect 11330 8820 11336 8832
rect 11103 8792 11336 8820
rect 11103 8789 11115 8792
rect 11057 8783 11115 8789
rect 11330 8780 11336 8792
rect 11388 8780 11394 8832
rect 11698 8780 11704 8832
rect 11756 8820 11762 8832
rect 12342 8820 12348 8832
rect 11756 8792 12348 8820
rect 11756 8780 11762 8792
rect 12342 8780 12348 8792
rect 12400 8820 12406 8832
rect 13081 8823 13139 8829
rect 13081 8820 13093 8823
rect 12400 8792 13093 8820
rect 12400 8780 12406 8792
rect 13081 8789 13093 8792
rect 13127 8789 13139 8823
rect 13081 8783 13139 8789
rect 13262 8780 13268 8832
rect 13320 8820 13326 8832
rect 13538 8820 13544 8832
rect 13320 8792 13544 8820
rect 13320 8780 13326 8792
rect 13538 8780 13544 8792
rect 13596 8780 13602 8832
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 13998 8820 14004 8832
rect 13872 8792 14004 8820
rect 13872 8780 13878 8792
rect 13998 8780 14004 8792
rect 14056 8780 14062 8832
rect 14918 8780 14924 8832
rect 14976 8820 14982 8832
rect 15105 8823 15163 8829
rect 15105 8820 15117 8823
rect 14976 8792 15117 8820
rect 14976 8780 14982 8792
rect 15105 8789 15117 8792
rect 15151 8789 15163 8823
rect 15105 8783 15163 8789
rect 16390 8780 16396 8832
rect 16448 8820 16454 8832
rect 17880 8820 17908 8987
rect 18414 8984 18420 8996
rect 18472 8984 18478 9036
rect 18230 8956 18236 8968
rect 18191 8928 18236 8956
rect 18230 8916 18236 8928
rect 18288 8916 18294 8968
rect 16448 8792 17908 8820
rect 18049 8823 18107 8829
rect 16448 8780 16454 8792
rect 18049 8789 18061 8823
rect 18095 8820 18107 8823
rect 18230 8820 18236 8832
rect 18095 8792 18236 8820
rect 18095 8789 18107 8792
rect 18049 8783 18107 8789
rect 18230 8780 18236 8792
rect 18288 8780 18294 8832
rect 1104 8730 18860 8752
rect 1104 8678 3947 8730
rect 3999 8678 4011 8730
rect 4063 8678 4075 8730
rect 4127 8678 4139 8730
rect 4191 8678 9878 8730
rect 9930 8678 9942 8730
rect 9994 8678 10006 8730
rect 10058 8678 10070 8730
rect 10122 8678 15808 8730
rect 15860 8678 15872 8730
rect 15924 8678 15936 8730
rect 15988 8678 16000 8730
rect 16052 8678 18860 8730
rect 1104 8656 18860 8678
rect 2590 8576 2596 8628
rect 2648 8616 2654 8628
rect 3329 8619 3387 8625
rect 3329 8616 3341 8619
rect 2648 8588 3341 8616
rect 2648 8576 2654 8588
rect 3329 8585 3341 8588
rect 3375 8585 3387 8619
rect 3329 8579 3387 8585
rect 3418 8576 3424 8628
rect 3476 8616 3482 8628
rect 3513 8619 3571 8625
rect 3513 8616 3525 8619
rect 3476 8588 3525 8616
rect 3476 8576 3482 8588
rect 3513 8585 3525 8588
rect 3559 8616 3571 8619
rect 5994 8616 6000 8628
rect 3559 8588 6000 8616
rect 3559 8585 3571 8588
rect 3513 8579 3571 8585
rect 5994 8576 6000 8588
rect 6052 8576 6058 8628
rect 6362 8576 6368 8628
rect 6420 8616 6426 8628
rect 13814 8616 13820 8628
rect 6420 8588 13820 8616
rect 6420 8576 6426 8588
rect 13814 8576 13820 8588
rect 13872 8576 13878 8628
rect 16025 8619 16083 8625
rect 16025 8585 16037 8619
rect 16071 8616 16083 8619
rect 16206 8616 16212 8628
rect 16071 8588 16212 8616
rect 16071 8585 16083 8588
rect 16025 8579 16083 8585
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 16390 8576 16396 8628
rect 16448 8616 16454 8628
rect 16577 8619 16635 8625
rect 16577 8616 16589 8619
rect 16448 8588 16589 8616
rect 16448 8576 16454 8588
rect 16577 8585 16589 8588
rect 16623 8585 16635 8619
rect 16577 8579 16635 8585
rect 16666 8576 16672 8628
rect 16724 8616 16730 8628
rect 17037 8619 17095 8625
rect 17037 8616 17049 8619
rect 16724 8588 17049 8616
rect 16724 8576 16730 8588
rect 17037 8585 17049 8588
rect 17083 8585 17095 8619
rect 17037 8579 17095 8585
rect 2958 8548 2964 8560
rect 2919 8520 2964 8548
rect 2958 8508 2964 8520
rect 3016 8508 3022 8560
rect 6086 8548 6092 8560
rect 6047 8520 6092 8548
rect 6086 8508 6092 8520
rect 6144 8508 6150 8560
rect 6457 8551 6515 8557
rect 6457 8517 6469 8551
rect 6503 8517 6515 8551
rect 8018 8548 8024 8560
rect 7979 8520 8024 8548
rect 6457 8511 6515 8517
rect 5442 8480 5448 8492
rect 4908 8452 5448 8480
rect 1854 8372 1860 8424
rect 1912 8412 1918 8424
rect 2869 8415 2927 8421
rect 2869 8412 2881 8415
rect 1912 8384 2881 8412
rect 1912 8372 1918 8384
rect 2869 8381 2881 8384
rect 2915 8412 2927 8415
rect 3602 8412 3608 8424
rect 2915 8384 3608 8412
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 3602 8372 3608 8384
rect 3660 8412 3666 8424
rect 4729 8415 4787 8421
rect 3660 8384 4660 8412
rect 3660 8372 3666 8384
rect 2624 8347 2682 8353
rect 2624 8313 2636 8347
rect 2670 8344 2682 8347
rect 2958 8344 2964 8356
rect 2670 8316 2964 8344
rect 2670 8313 2682 8316
rect 2624 8307 2682 8313
rect 2958 8304 2964 8316
rect 3016 8304 3022 8356
rect 3145 8347 3203 8353
rect 3145 8313 3157 8347
rect 3191 8313 3203 8347
rect 4632 8344 4660 8384
rect 4729 8381 4741 8415
rect 4775 8412 4787 8415
rect 4908 8412 4936 8452
rect 5442 8440 5448 8452
rect 5500 8480 5506 8492
rect 5813 8483 5871 8489
rect 5813 8480 5825 8483
rect 5500 8452 5825 8480
rect 5500 8440 5506 8452
rect 5813 8449 5825 8452
rect 5859 8480 5871 8483
rect 6472 8480 6500 8511
rect 8018 8508 8024 8520
rect 8076 8508 8082 8560
rect 8662 8508 8668 8560
rect 8720 8548 8726 8560
rect 9950 8548 9956 8560
rect 8720 8520 9168 8548
rect 9911 8520 9956 8548
rect 8720 8508 8726 8520
rect 7834 8480 7840 8492
rect 5859 8452 6500 8480
rect 7795 8452 7840 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 9030 8480 9036 8492
rect 8991 8452 9036 8480
rect 9030 8440 9036 8452
rect 9088 8440 9094 8492
rect 9140 8489 9168 8520
rect 9950 8508 9956 8520
rect 10008 8508 10014 8560
rect 11517 8551 11575 8557
rect 11517 8517 11529 8551
rect 11563 8517 11575 8551
rect 11517 8511 11575 8517
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8449 9183 8483
rect 11532 8480 11560 8511
rect 13446 8508 13452 8560
rect 13504 8548 13510 8560
rect 13630 8548 13636 8560
rect 13504 8520 13636 8548
rect 13504 8508 13510 8520
rect 13630 8508 13636 8520
rect 13688 8508 13694 8560
rect 16301 8551 16359 8557
rect 16301 8548 16313 8551
rect 15672 8520 16313 8548
rect 13722 8480 13728 8492
rect 11532 8452 11836 8480
rect 13683 8452 13728 8480
rect 9125 8443 9183 8449
rect 4775 8384 4936 8412
rect 4985 8415 5043 8421
rect 4775 8381 4787 8384
rect 4729 8375 4787 8381
rect 4985 8381 4997 8415
rect 5031 8381 5043 8415
rect 4985 8375 5043 8381
rect 6273 8415 6331 8421
rect 6273 8381 6285 8415
rect 6319 8412 6331 8415
rect 7282 8412 7288 8424
rect 6319 8384 7288 8412
rect 6319 8381 6331 8384
rect 6273 8375 6331 8381
rect 5000 8344 5028 8375
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8412 8999 8415
rect 9306 8412 9312 8424
rect 8987 8384 9312 8412
rect 8987 8381 8999 8384
rect 8941 8375 8999 8381
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 10137 8415 10195 8421
rect 10137 8381 10149 8415
rect 10183 8412 10195 8415
rect 11698 8412 11704 8424
rect 10183 8384 11704 8412
rect 10183 8381 10195 8384
rect 10137 8375 10195 8381
rect 11698 8372 11704 8384
rect 11756 8372 11762 8424
rect 11808 8412 11836 8452
rect 13722 8440 13728 8452
rect 13780 8440 13786 8492
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 14700 8452 14745 8480
rect 14700 8440 14706 8452
rect 11957 8415 12015 8421
rect 11957 8412 11969 8415
rect 11808 8384 11969 8412
rect 11957 8381 11969 8384
rect 12003 8412 12015 8415
rect 13740 8412 13768 8440
rect 15672 8412 15700 8520
rect 16301 8517 16313 8520
rect 16347 8548 16359 8551
rect 16942 8548 16948 8560
rect 16347 8520 16948 8548
rect 16347 8517 16359 8520
rect 16301 8511 16359 8517
rect 16942 8508 16948 8520
rect 17000 8508 17006 8560
rect 15838 8440 15844 8492
rect 15896 8480 15902 8492
rect 16117 8483 16175 8489
rect 16117 8480 16129 8483
rect 15896 8452 16129 8480
rect 15896 8440 15902 8452
rect 16117 8449 16129 8452
rect 16163 8449 16175 8483
rect 16117 8443 16175 8449
rect 16206 8440 16212 8492
rect 16264 8480 16270 8492
rect 17586 8480 17592 8492
rect 16264 8452 17592 8480
rect 16264 8440 16270 8452
rect 17586 8440 17592 8452
rect 17644 8440 17650 8492
rect 18138 8480 18144 8492
rect 17788 8452 18144 8480
rect 12003 8384 13768 8412
rect 14844 8384 15700 8412
rect 12003 8381 12015 8384
rect 11957 8375 12015 8381
rect 4632 8316 5028 8344
rect 5537 8347 5595 8353
rect 3145 8307 3203 8313
rect 5537 8313 5549 8347
rect 5583 8344 5595 8347
rect 6546 8344 6552 8356
rect 5583 8316 6552 8344
rect 5583 8313 5595 8316
rect 5537 8307 5595 8313
rect 1489 8279 1547 8285
rect 1489 8245 1501 8279
rect 1535 8276 1547 8279
rect 1578 8276 1584 8288
rect 1535 8248 1584 8276
rect 1535 8245 1547 8248
rect 1489 8239 1547 8245
rect 1578 8236 1584 8248
rect 1636 8236 1642 8288
rect 3160 8276 3188 8307
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 7558 8304 7564 8356
rect 7616 8353 7622 8356
rect 7616 8344 7628 8353
rect 7616 8316 7661 8344
rect 7616 8307 7628 8316
rect 7616 8304 7622 8307
rect 7742 8304 7748 8356
rect 7800 8344 7806 8356
rect 7800 8316 10180 8344
rect 7800 8304 7806 8316
rect 3329 8279 3387 8285
rect 3329 8276 3341 8279
rect 3160 8248 3341 8276
rect 3329 8245 3341 8248
rect 3375 8245 3387 8279
rect 3602 8276 3608 8288
rect 3563 8248 3608 8276
rect 3329 8239 3387 8245
rect 3602 8236 3608 8248
rect 3660 8236 3666 8288
rect 5166 8276 5172 8288
rect 5127 8248 5172 8276
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 5626 8236 5632 8288
rect 5684 8276 5690 8288
rect 5684 8248 5729 8276
rect 5684 8236 5690 8248
rect 6270 8236 6276 8288
rect 6328 8276 6334 8288
rect 8202 8276 8208 8288
rect 6328 8248 8208 8276
rect 6328 8236 6334 8248
rect 8202 8236 8208 8248
rect 8260 8236 8266 8288
rect 8294 8236 8300 8288
rect 8352 8276 8358 8288
rect 8573 8279 8631 8285
rect 8573 8276 8585 8279
rect 8352 8248 8585 8276
rect 8352 8236 8358 8248
rect 8573 8245 8585 8248
rect 8619 8245 8631 8279
rect 10152 8276 10180 8316
rect 10226 8304 10232 8356
rect 10284 8344 10290 8356
rect 10382 8347 10440 8353
rect 10382 8344 10394 8347
rect 10284 8316 10394 8344
rect 10284 8304 10290 8316
rect 10382 8313 10394 8316
rect 10428 8313 10440 8347
rect 13633 8347 13691 8353
rect 13633 8344 13645 8347
rect 10382 8307 10440 8313
rect 10520 8316 13645 8344
rect 10520 8276 10548 8316
rect 13633 8313 13645 8316
rect 13679 8344 13691 8347
rect 14001 8347 14059 8353
rect 14001 8344 14013 8347
rect 13679 8316 14013 8344
rect 13679 8313 13691 8316
rect 13633 8307 13691 8313
rect 14001 8313 14013 8316
rect 14047 8344 14059 8347
rect 14844 8344 14872 8384
rect 15746 8372 15752 8424
rect 15804 8412 15810 8424
rect 17405 8415 17463 8421
rect 17405 8412 17417 8415
rect 15804 8384 17417 8412
rect 15804 8372 15810 8384
rect 17405 8381 17417 8384
rect 17451 8412 17463 8415
rect 17788 8412 17816 8452
rect 18138 8440 18144 8452
rect 18196 8440 18202 8492
rect 17451 8384 17816 8412
rect 17865 8415 17923 8421
rect 17451 8381 17463 8384
rect 17405 8375 17463 8381
rect 17865 8381 17877 8415
rect 17911 8381 17923 8415
rect 18322 8412 18328 8424
rect 18283 8384 18328 8412
rect 17865 8375 17923 8381
rect 14047 8316 14872 8344
rect 14912 8347 14970 8353
rect 14047 8313 14059 8316
rect 14001 8307 14059 8313
rect 14912 8313 14924 8347
rect 14958 8344 14970 8347
rect 15654 8344 15660 8356
rect 14958 8316 15660 8344
rect 14958 8313 14970 8316
rect 14912 8307 14970 8313
rect 15654 8304 15660 8316
rect 15712 8304 15718 8356
rect 16758 8344 16764 8356
rect 16719 8316 16764 8344
rect 16758 8304 16764 8316
rect 16816 8344 16822 8356
rect 16816 8316 16896 8344
rect 16816 8304 16822 8316
rect 10152 8248 10548 8276
rect 8573 8239 8631 8245
rect 11790 8236 11796 8288
rect 11848 8276 11854 8288
rect 11974 8276 11980 8288
rect 11848 8248 11980 8276
rect 11848 8236 11854 8248
rect 11974 8236 11980 8248
rect 12032 8236 12038 8288
rect 12710 8236 12716 8288
rect 12768 8276 12774 8288
rect 13081 8279 13139 8285
rect 13081 8276 13093 8279
rect 12768 8248 13093 8276
rect 12768 8236 12774 8248
rect 13081 8245 13093 8248
rect 13127 8245 13139 8279
rect 13081 8239 13139 8245
rect 13170 8236 13176 8288
rect 13228 8276 13234 8288
rect 13541 8279 13599 8285
rect 13228 8248 13273 8276
rect 13228 8236 13234 8248
rect 13541 8245 13553 8279
rect 13587 8276 13599 8279
rect 13814 8276 13820 8288
rect 13587 8248 13820 8276
rect 13587 8245 13599 8248
rect 13541 8239 13599 8245
rect 13814 8236 13820 8248
rect 13872 8276 13878 8288
rect 15746 8276 15752 8288
rect 13872 8248 15752 8276
rect 13872 8236 13878 8248
rect 15746 8236 15752 8248
rect 15804 8236 15810 8288
rect 15838 8236 15844 8288
rect 15896 8276 15902 8288
rect 16666 8276 16672 8288
rect 15896 8248 16672 8276
rect 15896 8236 15902 8248
rect 16666 8236 16672 8248
rect 16724 8236 16730 8288
rect 16868 8276 16896 8316
rect 16942 8304 16948 8356
rect 17000 8344 17006 8356
rect 17497 8347 17555 8353
rect 17497 8344 17509 8347
rect 17000 8316 17509 8344
rect 17000 8304 17006 8316
rect 17497 8313 17509 8316
rect 17543 8344 17555 8347
rect 17770 8344 17776 8356
rect 17543 8316 17776 8344
rect 17543 8313 17555 8316
rect 17497 8307 17555 8313
rect 17770 8304 17776 8316
rect 17828 8304 17834 8356
rect 17880 8276 17908 8375
rect 18322 8372 18328 8384
rect 18380 8372 18386 8424
rect 18506 8344 18512 8356
rect 18467 8316 18512 8344
rect 18506 8304 18512 8316
rect 18564 8304 18570 8356
rect 18046 8276 18052 8288
rect 16868 8248 17908 8276
rect 18007 8248 18052 8276
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 1104 8186 18860 8208
rect 1104 8134 6912 8186
rect 6964 8134 6976 8186
rect 7028 8134 7040 8186
rect 7092 8134 7104 8186
rect 7156 8134 12843 8186
rect 12895 8134 12907 8186
rect 12959 8134 12971 8186
rect 13023 8134 13035 8186
rect 13087 8134 18860 8186
rect 1104 8112 18860 8134
rect 1854 8072 1860 8084
rect 1815 8044 1860 8072
rect 1854 8032 1860 8044
rect 1912 8032 1918 8084
rect 2501 8075 2559 8081
rect 2501 8041 2513 8075
rect 2547 8072 2559 8075
rect 2961 8075 3019 8081
rect 2961 8072 2973 8075
rect 2547 8044 2973 8072
rect 2547 8041 2559 8044
rect 2501 8035 2559 8041
rect 2961 8041 2973 8044
rect 3007 8041 3019 8075
rect 3418 8072 3424 8084
rect 3379 8044 3424 8072
rect 2961 8035 3019 8041
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 4246 8072 4252 8084
rect 4207 8044 4252 8072
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 5074 8032 5080 8084
rect 5132 8072 5138 8084
rect 5169 8075 5227 8081
rect 5169 8072 5181 8075
rect 5132 8044 5181 8072
rect 5132 8032 5138 8044
rect 5169 8041 5181 8044
rect 5215 8072 5227 8075
rect 5258 8072 5264 8084
rect 5215 8044 5264 8072
rect 5215 8041 5227 8044
rect 5169 8035 5227 8041
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 5350 8032 5356 8084
rect 5408 8032 5414 8084
rect 5626 8032 5632 8084
rect 5684 8072 5690 8084
rect 5721 8075 5779 8081
rect 5721 8072 5733 8075
rect 5684 8044 5733 8072
rect 5684 8032 5690 8044
rect 5721 8041 5733 8044
rect 5767 8041 5779 8075
rect 6546 8072 6552 8084
rect 6507 8044 6552 8072
rect 5721 8035 5779 8041
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 6638 8032 6644 8084
rect 6696 8072 6702 8084
rect 6917 8075 6975 8081
rect 6696 8044 6868 8072
rect 6696 8032 6702 8044
rect 1581 8007 1639 8013
rect 1581 7973 1593 8007
rect 1627 8004 1639 8007
rect 2866 8004 2872 8016
rect 1627 7976 2872 8004
rect 1627 7973 1639 7976
rect 1581 7967 1639 7973
rect 2866 7964 2872 7976
rect 2924 7964 2930 8016
rect 5368 8004 5396 8032
rect 5810 8004 5816 8016
rect 5368 7976 5816 8004
rect 5810 7964 5816 7976
rect 5868 8004 5874 8016
rect 6181 8007 6239 8013
rect 6181 8004 6193 8007
rect 5868 7976 6193 8004
rect 5868 7964 5874 7976
rect 6181 7973 6193 7976
rect 6227 8004 6239 8007
rect 6840 8004 6868 8044
rect 6917 8041 6929 8075
rect 6963 8072 6975 8075
rect 7374 8072 7380 8084
rect 6963 8044 7380 8072
rect 6963 8041 6975 8044
rect 6917 8035 6975 8041
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 7745 8075 7803 8081
rect 7745 8041 7757 8075
rect 7791 8072 7803 8075
rect 8205 8075 8263 8081
rect 8205 8072 8217 8075
rect 7791 8044 8217 8072
rect 7791 8041 7803 8044
rect 7745 8035 7803 8041
rect 8205 8041 8217 8044
rect 8251 8041 8263 8075
rect 8205 8035 8263 8041
rect 8665 8075 8723 8081
rect 8665 8041 8677 8075
rect 8711 8072 8723 8075
rect 9122 8072 9128 8084
rect 8711 8044 9128 8072
rect 8711 8041 8723 8044
rect 8665 8035 8723 8041
rect 9122 8032 9128 8044
rect 9180 8032 9186 8084
rect 9306 8032 9312 8084
rect 9364 8072 9370 8084
rect 16298 8072 16304 8084
rect 9364 8044 16160 8072
rect 16259 8044 16304 8072
rect 9364 8032 9370 8044
rect 7009 8007 7067 8013
rect 7009 8004 7021 8007
rect 6227 7976 6684 8004
rect 6840 7976 7021 8004
rect 6227 7973 6239 7976
rect 6181 7967 6239 7973
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7936 2007 7939
rect 2130 7936 2136 7948
rect 1995 7908 2136 7936
rect 1995 7905 2007 7908
rect 1949 7899 2007 7905
rect 2130 7896 2136 7908
rect 2188 7896 2194 7948
rect 3329 7939 3387 7945
rect 3329 7905 3341 7939
rect 3375 7936 3387 7939
rect 3418 7936 3424 7948
rect 3375 7908 3424 7936
rect 3375 7905 3387 7908
rect 3329 7899 3387 7905
rect 3418 7896 3424 7908
rect 3476 7896 3482 7948
rect 3694 7896 3700 7948
rect 3752 7936 3758 7948
rect 4341 7939 4399 7945
rect 4341 7936 4353 7939
rect 3752 7908 4353 7936
rect 3752 7896 3758 7908
rect 4341 7905 4353 7908
rect 4387 7936 4399 7939
rect 5350 7936 5356 7948
rect 4387 7908 5356 7936
rect 4387 7905 4399 7908
rect 4341 7899 4399 7905
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 5626 7896 5632 7948
rect 5684 7936 5690 7948
rect 6089 7939 6147 7945
rect 6089 7936 6101 7939
rect 5684 7908 6101 7936
rect 5684 7896 5690 7908
rect 6089 7905 6101 7908
rect 6135 7936 6147 7939
rect 6362 7936 6368 7948
rect 6135 7908 6368 7936
rect 6135 7905 6147 7908
rect 6089 7899 6147 7905
rect 6362 7896 6368 7908
rect 6420 7896 6426 7948
rect 6656 7936 6684 7976
rect 7009 7973 7021 7976
rect 7055 7973 7067 8007
rect 7009 7967 7067 7973
rect 7837 8007 7895 8013
rect 7837 7973 7849 8007
rect 7883 8004 7895 8007
rect 8294 8004 8300 8016
rect 7883 7976 8300 8004
rect 7883 7973 7895 7976
rect 7837 7967 7895 7973
rect 8294 7964 8300 7976
rect 8352 7964 8358 8016
rect 11974 8004 11980 8016
rect 8588 7976 11980 8004
rect 7742 7936 7748 7948
rect 6656 7908 7748 7936
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 8110 7896 8116 7948
rect 8168 7936 8174 7948
rect 8588 7945 8616 7976
rect 11974 7964 11980 7976
rect 12032 7964 12038 8016
rect 12100 8007 12158 8013
rect 12100 7973 12112 8007
rect 12146 8004 12158 8007
rect 12710 8004 12716 8016
rect 12146 7976 12716 8004
rect 12146 7973 12158 7976
rect 12100 7967 12158 7973
rect 12710 7964 12716 7976
rect 12768 7964 12774 8016
rect 12986 8004 12992 8016
rect 12899 7976 12992 8004
rect 12986 7964 12992 7976
rect 13044 8004 13050 8016
rect 13722 8004 13728 8016
rect 13044 7976 13216 8004
rect 13044 7964 13050 7976
rect 8573 7939 8631 7945
rect 8573 7936 8585 7939
rect 8168 7908 8585 7936
rect 8168 7896 8174 7908
rect 8573 7905 8585 7908
rect 8619 7905 8631 7939
rect 8573 7899 8631 7905
rect 8938 7896 8944 7948
rect 8996 7936 9002 7948
rect 9125 7939 9183 7945
rect 9125 7936 9137 7939
rect 8996 7908 9137 7936
rect 8996 7896 9002 7908
rect 9125 7905 9137 7908
rect 9171 7905 9183 7939
rect 9125 7899 9183 7905
rect 9398 7896 9404 7948
rect 9456 7936 9462 7948
rect 13078 7936 13084 7948
rect 9456 7908 13084 7936
rect 9456 7896 9462 7908
rect 13078 7896 13084 7908
rect 13136 7896 13142 7948
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7837 2651 7871
rect 2593 7831 2651 7837
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7868 2743 7871
rect 2958 7868 2964 7880
rect 2731 7840 2964 7868
rect 2731 7837 2743 7840
rect 2685 7831 2743 7837
rect 2608 7800 2636 7831
rect 2958 7828 2964 7840
rect 3016 7868 3022 7880
rect 3510 7868 3516 7880
rect 3016 7840 3516 7868
rect 3016 7828 3022 7840
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7868 3663 7871
rect 4525 7871 4583 7877
rect 3651 7840 4292 7868
rect 3651 7837 3663 7840
rect 3605 7831 3663 7837
rect 3881 7803 3939 7809
rect 3881 7800 3893 7803
rect 2608 7772 3893 7800
rect 3881 7769 3893 7772
rect 3927 7769 3939 7803
rect 4264 7800 4292 7840
rect 4525 7837 4537 7871
rect 4571 7837 4583 7871
rect 5258 7868 5264 7880
rect 5219 7840 5264 7868
rect 4525 7831 4583 7837
rect 4540 7800 4568 7831
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 5442 7868 5448 7880
rect 5403 7840 5448 7868
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 6270 7868 6276 7880
rect 6231 7840 6276 7868
rect 6270 7828 6276 7840
rect 6328 7868 6334 7880
rect 7098 7868 7104 7880
rect 6328 7840 7104 7868
rect 6328 7828 6334 7840
rect 7098 7828 7104 7840
rect 7156 7868 7162 7880
rect 7558 7868 7564 7880
rect 7156 7840 7564 7868
rect 7156 7828 7162 7840
rect 7558 7828 7564 7840
rect 7616 7828 7622 7880
rect 8021 7871 8079 7877
rect 8021 7837 8033 7871
rect 8067 7868 8079 7871
rect 8386 7868 8392 7880
rect 8067 7840 8392 7868
rect 8067 7837 8079 7840
rect 8021 7831 8079 7837
rect 8386 7828 8392 7840
rect 8444 7828 8450 7880
rect 8662 7828 8668 7880
rect 8720 7868 8726 7880
rect 8757 7871 8815 7877
rect 8757 7868 8769 7871
rect 8720 7840 8769 7868
rect 8720 7828 8726 7840
rect 8757 7837 8769 7840
rect 8803 7837 8815 7871
rect 12342 7868 12348 7880
rect 12303 7840 12348 7868
rect 8757 7831 8815 7837
rect 12342 7828 12348 7840
rect 12400 7828 12406 7880
rect 5460 7800 5488 7828
rect 4264 7772 5488 7800
rect 3881 7763 3939 7769
rect 7282 7760 7288 7812
rect 7340 7800 7346 7812
rect 10413 7803 10471 7809
rect 10413 7800 10425 7803
rect 7340 7772 10425 7800
rect 7340 7760 7346 7772
rect 10413 7769 10425 7772
rect 10459 7800 10471 7803
rect 12802 7800 12808 7812
rect 10459 7772 11468 7800
rect 12763 7772 12808 7800
rect 10459 7769 10471 7772
rect 10413 7763 10471 7769
rect 1486 7732 1492 7744
rect 1447 7704 1492 7732
rect 1486 7692 1492 7704
rect 1544 7692 1550 7744
rect 2133 7735 2191 7741
rect 2133 7701 2145 7735
rect 2179 7732 2191 7735
rect 2406 7732 2412 7744
rect 2179 7704 2412 7732
rect 2179 7701 2191 7704
rect 2133 7695 2191 7701
rect 2406 7692 2412 7704
rect 2464 7692 2470 7744
rect 4614 7692 4620 7744
rect 4672 7732 4678 7744
rect 4801 7735 4859 7741
rect 4801 7732 4813 7735
rect 4672 7704 4813 7732
rect 4672 7692 4678 7704
rect 4801 7701 4813 7704
rect 4847 7701 4859 7735
rect 4801 7695 4859 7701
rect 7377 7735 7435 7741
rect 7377 7701 7389 7735
rect 7423 7732 7435 7735
rect 7742 7732 7748 7744
rect 7423 7704 7748 7732
rect 7423 7701 7435 7704
rect 7377 7695 7435 7701
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 10965 7735 11023 7741
rect 10965 7701 10977 7735
rect 11011 7732 11023 7735
rect 11054 7732 11060 7744
rect 11011 7704 11060 7732
rect 11011 7701 11023 7704
rect 10965 7695 11023 7701
rect 11054 7692 11060 7704
rect 11112 7692 11118 7744
rect 11440 7732 11468 7772
rect 12802 7760 12808 7772
rect 12860 7760 12866 7812
rect 13188 7800 13216 7976
rect 13280 7976 13728 8004
rect 13280 7877 13308 7976
rect 13722 7964 13728 7976
rect 13780 7964 13786 8016
rect 14001 8007 14059 8013
rect 14001 7973 14013 8007
rect 14047 8004 14059 8007
rect 14090 8004 14096 8016
rect 14047 7976 14096 8004
rect 14047 7973 14059 7976
rect 14001 7967 14059 7973
rect 13449 7939 13507 7945
rect 13449 7905 13461 7939
rect 13495 7936 13507 7939
rect 13814 7936 13820 7948
rect 13495 7908 13820 7936
rect 13495 7905 13507 7908
rect 13449 7899 13507 7905
rect 13814 7896 13820 7908
rect 13872 7936 13878 7948
rect 14016 7936 14044 7967
rect 14090 7964 14096 7976
rect 14148 7964 14154 8016
rect 14829 8007 14887 8013
rect 14829 7973 14841 8007
rect 14875 8004 14887 8007
rect 15378 8004 15384 8016
rect 14875 7976 15384 8004
rect 14875 7973 14887 7976
rect 14829 7967 14887 7973
rect 15378 7964 15384 7976
rect 15436 7964 15442 8016
rect 13872 7908 14044 7936
rect 13872 7896 13878 7908
rect 14642 7896 14648 7948
rect 14700 7936 14706 7948
rect 14921 7939 14979 7945
rect 14921 7936 14933 7939
rect 14700 7908 14933 7936
rect 14700 7896 14706 7908
rect 14921 7905 14933 7908
rect 14967 7905 14979 7939
rect 14921 7899 14979 7905
rect 15188 7939 15246 7945
rect 15188 7905 15200 7939
rect 15234 7936 15246 7939
rect 15654 7936 15660 7948
rect 15234 7908 15660 7936
rect 15234 7905 15246 7908
rect 15188 7899 15246 7905
rect 15654 7896 15660 7908
rect 15712 7896 15718 7948
rect 13265 7871 13323 7877
rect 13265 7837 13277 7871
rect 13311 7837 13323 7871
rect 13265 7831 13323 7837
rect 13357 7871 13415 7877
rect 13357 7837 13369 7871
rect 13403 7868 13415 7871
rect 16132 7868 16160 8044
rect 16298 8032 16304 8044
rect 16356 8032 16362 8084
rect 16666 8032 16672 8084
rect 16724 8072 16730 8084
rect 16761 8075 16819 8081
rect 16761 8072 16773 8075
rect 16724 8044 16773 8072
rect 16724 8032 16730 8044
rect 16761 8041 16773 8044
rect 16807 8041 16819 8075
rect 16942 8072 16948 8084
rect 16903 8044 16948 8072
rect 16761 8035 16819 8041
rect 16776 8004 16804 8035
rect 16942 8032 16948 8044
rect 17000 8032 17006 8084
rect 17129 8075 17187 8081
rect 17129 8041 17141 8075
rect 17175 8072 17187 8075
rect 17402 8072 17408 8084
rect 17175 8044 17408 8072
rect 17175 8041 17187 8044
rect 17129 8035 17187 8041
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 17497 8075 17555 8081
rect 17497 8041 17509 8075
rect 17543 8072 17555 8075
rect 17954 8072 17960 8084
rect 17543 8044 17960 8072
rect 17543 8041 17555 8044
rect 17497 8035 17555 8041
rect 17954 8032 17960 8044
rect 18012 8072 18018 8084
rect 18690 8072 18696 8084
rect 18012 8044 18696 8072
rect 18012 8032 18018 8044
rect 18690 8032 18696 8044
rect 18748 8032 18754 8084
rect 17310 8004 17316 8016
rect 16776 7976 17316 8004
rect 17310 7964 17316 7976
rect 17368 7964 17374 8016
rect 18230 7964 18236 8016
rect 18288 8004 18294 8016
rect 18325 8007 18383 8013
rect 18325 8004 18337 8007
rect 18288 7976 18337 8004
rect 18288 7964 18294 7976
rect 18325 7973 18337 7976
rect 18371 7973 18383 8007
rect 18325 7967 18383 7973
rect 17589 7939 17647 7945
rect 17589 7936 17601 7939
rect 17420 7908 17601 7936
rect 17126 7868 17132 7880
rect 13403 7840 14688 7868
rect 16132 7840 17132 7868
rect 13403 7837 13415 7840
rect 13357 7831 13415 7837
rect 13372 7800 13400 7831
rect 14660 7812 14688 7840
rect 17126 7828 17132 7840
rect 17184 7828 17190 7880
rect 17420 7868 17448 7908
rect 17589 7905 17601 7908
rect 17635 7905 17647 7939
rect 17589 7899 17647 7905
rect 17770 7896 17776 7948
rect 17828 7936 17834 7948
rect 18141 7939 18199 7945
rect 18141 7936 18153 7939
rect 17828 7908 18153 7936
rect 17828 7896 17834 7908
rect 18141 7905 18153 7908
rect 18187 7905 18199 7939
rect 18141 7899 18199 7905
rect 17678 7868 17684 7880
rect 17236 7840 17448 7868
rect 17639 7840 17684 7868
rect 13188 7772 13400 7800
rect 14642 7760 14648 7812
rect 14700 7760 14706 7812
rect 17236 7800 17264 7840
rect 17678 7828 17684 7840
rect 17736 7828 17742 7880
rect 18506 7800 18512 7812
rect 16776 7772 17264 7800
rect 18467 7772 18512 7800
rect 16776 7744 16804 7772
rect 18506 7760 18512 7772
rect 18564 7760 18570 7812
rect 11698 7732 11704 7744
rect 11440 7704 11704 7732
rect 11698 7692 11704 7704
rect 11756 7692 11762 7744
rect 13538 7692 13544 7744
rect 13596 7732 13602 7744
rect 13817 7735 13875 7741
rect 13817 7732 13829 7735
rect 13596 7704 13829 7732
rect 13596 7692 13602 7704
rect 13817 7701 13829 7704
rect 13863 7701 13875 7735
rect 13817 7695 13875 7701
rect 14366 7692 14372 7744
rect 14424 7732 14430 7744
rect 16298 7732 16304 7744
rect 14424 7704 16304 7732
rect 14424 7692 14430 7704
rect 16298 7692 16304 7704
rect 16356 7692 16362 7744
rect 16482 7732 16488 7744
rect 16443 7704 16488 7732
rect 16482 7692 16488 7704
rect 16540 7692 16546 7744
rect 16669 7735 16727 7741
rect 16669 7701 16681 7735
rect 16715 7732 16727 7735
rect 16758 7732 16764 7744
rect 16715 7704 16764 7732
rect 16715 7701 16727 7704
rect 16669 7695 16727 7701
rect 16758 7692 16764 7704
rect 16816 7692 16822 7744
rect 17957 7735 18015 7741
rect 17957 7701 17969 7735
rect 18003 7732 18015 7735
rect 18414 7732 18420 7744
rect 18003 7704 18420 7732
rect 18003 7701 18015 7704
rect 17957 7695 18015 7701
rect 18414 7692 18420 7704
rect 18472 7692 18478 7744
rect 1104 7642 18860 7664
rect 1104 7590 3947 7642
rect 3999 7590 4011 7642
rect 4063 7590 4075 7642
rect 4127 7590 4139 7642
rect 4191 7590 9878 7642
rect 9930 7590 9942 7642
rect 9994 7590 10006 7642
rect 10058 7590 10070 7642
rect 10122 7590 15808 7642
rect 15860 7590 15872 7642
rect 15924 7590 15936 7642
rect 15988 7590 16000 7642
rect 16052 7590 18860 7642
rect 1104 7568 18860 7590
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 2096 7500 3157 7528
rect 2096 7488 2102 7500
rect 3145 7497 3157 7500
rect 3191 7497 3203 7531
rect 3145 7491 3203 7497
rect 3326 7488 3332 7540
rect 3384 7528 3390 7540
rect 3973 7531 4031 7537
rect 3973 7528 3985 7531
rect 3384 7500 3985 7528
rect 3384 7488 3390 7500
rect 3973 7497 3985 7500
rect 4019 7497 4031 7531
rect 5074 7528 5080 7540
rect 5035 7500 5080 7528
rect 3973 7491 4031 7497
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 5258 7488 5264 7540
rect 5316 7528 5322 7540
rect 6457 7531 6515 7537
rect 6457 7528 6469 7531
rect 5316 7500 6469 7528
rect 5316 7488 5322 7500
rect 6457 7497 6469 7500
rect 6503 7497 6515 7531
rect 6457 7491 6515 7497
rect 6638 7488 6644 7540
rect 6696 7488 6702 7540
rect 11882 7528 11888 7540
rect 7576 7500 11560 7528
rect 11843 7500 11888 7528
rect 2866 7460 2872 7472
rect 2827 7432 2872 7460
rect 2866 7420 2872 7432
rect 2924 7420 2930 7472
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 2133 7395 2191 7401
rect 2133 7392 2145 7395
rect 1636 7364 2145 7392
rect 1636 7352 1642 7364
rect 2133 7361 2145 7364
rect 2179 7361 2191 7395
rect 2958 7392 2964 7404
rect 2133 7355 2191 7361
rect 2240 7364 2964 7392
rect 1394 7324 1400 7336
rect 1355 7296 1400 7324
rect 1394 7284 1400 7296
rect 1452 7284 1458 7336
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7324 2007 7327
rect 2240 7324 2268 7364
rect 2958 7352 2964 7364
rect 3016 7352 3022 7404
rect 3344 7392 3372 7488
rect 3418 7420 3424 7472
rect 3476 7460 3482 7472
rect 3881 7463 3939 7469
rect 3476 7432 3556 7460
rect 3476 7420 3482 7432
rect 3528 7401 3556 7432
rect 3881 7429 3893 7463
rect 3927 7460 3939 7463
rect 4246 7460 4252 7472
rect 3927 7432 4252 7460
rect 3927 7429 3939 7432
rect 3881 7423 3939 7429
rect 4246 7420 4252 7432
rect 4304 7420 4310 7472
rect 5629 7463 5687 7469
rect 5629 7429 5641 7463
rect 5675 7460 5687 7463
rect 5810 7460 5816 7472
rect 5675 7432 5816 7460
rect 5675 7429 5687 7432
rect 5629 7423 5687 7429
rect 5810 7420 5816 7432
rect 5868 7420 5874 7472
rect 6273 7463 6331 7469
rect 6273 7429 6285 7463
rect 6319 7460 6331 7463
rect 6656 7460 6684 7488
rect 6319 7432 6684 7460
rect 6319 7429 6331 7432
rect 6273 7423 6331 7429
rect 3068 7364 3372 7392
rect 3513 7395 3571 7401
rect 2406 7324 2412 7336
rect 1995 7296 2268 7324
rect 2367 7296 2412 7324
rect 1995 7293 2007 7296
rect 1949 7287 2007 7293
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 3068 7333 3096 7364
rect 3513 7361 3525 7395
rect 3559 7361 3571 7395
rect 3513 7355 3571 7361
rect 3602 7352 3608 7404
rect 3660 7392 3666 7404
rect 4801 7395 4859 7401
rect 4801 7392 4813 7395
rect 3660 7364 4813 7392
rect 3660 7352 3666 7364
rect 4801 7361 4813 7364
rect 4847 7361 4859 7395
rect 5350 7392 5356 7404
rect 5311 7364 5356 7392
rect 4801 7355 4859 7361
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 6638 7392 6644 7404
rect 6012 7364 6644 7392
rect 3053 7327 3111 7333
rect 3053 7293 3065 7327
rect 3099 7293 3111 7327
rect 3053 7287 3111 7293
rect 3329 7327 3387 7333
rect 3329 7293 3341 7327
rect 3375 7324 3387 7327
rect 4614 7324 4620 7336
rect 3375 7296 4476 7324
rect 4575 7296 4620 7324
rect 3375 7293 3387 7296
rect 3329 7287 3387 7293
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 2317 7259 2375 7265
rect 1627 7228 1808 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 1780 7197 1808 7228
rect 2317 7225 2329 7259
rect 2363 7256 2375 7259
rect 4448 7256 4476 7296
rect 4614 7284 4620 7296
rect 4672 7284 4678 7336
rect 4709 7327 4767 7333
rect 4709 7293 4721 7327
rect 4755 7324 4767 7327
rect 5166 7324 5172 7336
rect 4755 7296 5172 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 5166 7284 5172 7296
rect 5224 7284 5230 7336
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 6012 7333 6040 7364
rect 6638 7352 6644 7364
rect 6696 7352 6702 7404
rect 7098 7392 7104 7404
rect 7059 7364 7104 7392
rect 7098 7352 7104 7364
rect 7156 7352 7162 7404
rect 7576 7333 7604 7500
rect 10045 7463 10103 7469
rect 10045 7429 10057 7463
rect 10091 7429 10103 7463
rect 10045 7423 10103 7429
rect 8386 7392 8392 7404
rect 8347 7364 8392 7392
rect 8386 7352 8392 7364
rect 8444 7352 8450 7404
rect 5997 7327 6055 7333
rect 5997 7324 6009 7327
rect 5592 7296 6009 7324
rect 5592 7284 5598 7296
rect 5997 7293 6009 7296
rect 6043 7293 6055 7327
rect 7561 7327 7619 7333
rect 7561 7324 7573 7327
rect 5997 7287 6055 7293
rect 6840 7296 7573 7324
rect 5626 7256 5632 7268
rect 2363 7228 4292 7256
rect 4448 7228 5632 7256
rect 2363 7225 2375 7228
rect 2317 7219 2375 7225
rect 1765 7191 1823 7197
rect 1765 7157 1777 7191
rect 1811 7157 1823 7191
rect 1765 7151 1823 7157
rect 2777 7191 2835 7197
rect 2777 7157 2789 7191
rect 2823 7188 2835 7191
rect 3234 7188 3240 7200
rect 2823 7160 3240 7188
rect 2823 7157 2835 7160
rect 2777 7151 2835 7157
rect 3234 7148 3240 7160
rect 3292 7148 3298 7200
rect 4264 7197 4292 7228
rect 5626 7216 5632 7228
rect 5684 7216 5690 7268
rect 6362 7216 6368 7268
rect 6420 7256 6426 7268
rect 6840 7265 6868 7296
rect 7561 7293 7573 7296
rect 7607 7293 7619 7327
rect 7561 7287 7619 7293
rect 8570 7284 8576 7336
rect 8628 7324 8634 7336
rect 8665 7327 8723 7333
rect 8665 7324 8677 7327
rect 8628 7296 8677 7324
rect 8628 7284 8634 7296
rect 8665 7293 8677 7296
rect 8711 7293 8723 7327
rect 8665 7287 8723 7293
rect 9306 7284 9312 7336
rect 9364 7324 9370 7336
rect 10060 7324 10088 7423
rect 10134 7420 10140 7472
rect 10192 7460 10198 7472
rect 11532 7460 11560 7500
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 12342 7528 12348 7540
rect 12084 7500 12348 7528
rect 12084 7460 12112 7500
rect 12342 7488 12348 7500
rect 12400 7488 12406 7540
rect 12986 7528 12992 7540
rect 12452 7500 12992 7528
rect 10192 7432 10237 7460
rect 11532 7432 12112 7460
rect 10192 7420 10198 7432
rect 12158 7420 12164 7472
rect 12216 7460 12222 7472
rect 12216 7432 12261 7460
rect 12216 7420 12222 7432
rect 9364 7296 10088 7324
rect 9364 7284 9370 7296
rect 6825 7259 6883 7265
rect 6825 7256 6837 7259
rect 6420 7228 6837 7256
rect 6420 7216 6426 7228
rect 6825 7225 6837 7228
rect 6871 7225 6883 7259
rect 6825 7219 6883 7225
rect 6932 7228 8432 7256
rect 4249 7191 4307 7197
rect 4249 7157 4261 7191
rect 4295 7157 4307 7191
rect 4249 7151 4307 7157
rect 6638 7148 6644 7200
rect 6696 7188 6702 7200
rect 6932 7197 6960 7228
rect 6917 7191 6975 7197
rect 6917 7188 6929 7191
rect 6696 7160 6929 7188
rect 6696 7148 6702 7160
rect 6917 7157 6929 7160
rect 6963 7157 6975 7191
rect 7374 7188 7380 7200
rect 7335 7160 7380 7188
rect 6917 7151 6975 7157
rect 7374 7148 7380 7160
rect 7432 7148 7438 7200
rect 7650 7148 7656 7200
rect 7708 7188 7714 7200
rect 7745 7191 7803 7197
rect 7745 7188 7757 7191
rect 7708 7160 7757 7188
rect 7708 7148 7714 7160
rect 7745 7157 7757 7160
rect 7791 7157 7803 7191
rect 8110 7188 8116 7200
rect 8071 7160 8116 7188
rect 7745 7151 7803 7157
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 8202 7148 8208 7200
rect 8260 7188 8266 7200
rect 8404 7188 8432 7228
rect 8754 7216 8760 7268
rect 8812 7256 8818 7268
rect 8910 7259 8968 7265
rect 8910 7256 8922 7259
rect 8812 7228 8922 7256
rect 8812 7216 8818 7228
rect 8910 7225 8922 7228
rect 8956 7225 8968 7259
rect 10060 7256 10088 7296
rect 10962 7284 10968 7336
rect 11020 7324 11026 7336
rect 11517 7327 11575 7333
rect 11517 7324 11529 7327
rect 11020 7296 11529 7324
rect 11020 7284 11026 7296
rect 11517 7293 11529 7296
rect 11563 7293 11575 7327
rect 11698 7324 11704 7336
rect 11659 7296 11704 7324
rect 11517 7287 11575 7293
rect 11698 7284 11704 7296
rect 11756 7284 11762 7336
rect 12452 7324 12480 7500
rect 12986 7488 12992 7500
rect 13044 7488 13050 7540
rect 13262 7488 13268 7540
rect 13320 7528 13326 7540
rect 13320 7500 13860 7528
rect 13320 7488 13326 7500
rect 13832 7472 13860 7500
rect 15194 7488 15200 7540
rect 15252 7488 15258 7540
rect 15378 7488 15384 7540
rect 15436 7528 15442 7540
rect 17954 7528 17960 7540
rect 15436 7500 17960 7528
rect 15436 7488 15442 7500
rect 17954 7488 17960 7500
rect 18012 7488 18018 7540
rect 12710 7420 12716 7472
rect 12768 7460 12774 7472
rect 12768 7432 13676 7460
rect 12768 7420 12774 7432
rect 12820 7401 12848 7432
rect 12805 7395 12863 7401
rect 12805 7361 12817 7395
rect 12851 7361 12863 7395
rect 12805 7355 12863 7361
rect 13078 7352 13084 7404
rect 13136 7392 13142 7404
rect 13538 7392 13544 7404
rect 13136 7364 13308 7392
rect 13499 7364 13544 7392
rect 13136 7352 13142 7364
rect 12618 7324 12624 7336
rect 11900 7296 12480 7324
rect 12579 7296 12624 7324
rect 11250 7259 11308 7265
rect 11250 7256 11262 7259
rect 10060 7228 11262 7256
rect 8910 7219 8968 7225
rect 11250 7225 11262 7228
rect 11296 7225 11308 7259
rect 11250 7219 11308 7225
rect 11900 7188 11928 7296
rect 12618 7284 12624 7296
rect 12676 7284 12682 7336
rect 12713 7327 12771 7333
rect 12713 7293 12725 7327
rect 12759 7324 12771 7327
rect 13170 7324 13176 7336
rect 12759 7296 13176 7324
rect 12759 7293 12771 7296
rect 12713 7287 12771 7293
rect 13170 7284 13176 7296
rect 13228 7284 13234 7336
rect 13280 7324 13308 7364
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 13648 7401 13676 7432
rect 13814 7420 13820 7472
rect 13872 7420 13878 7472
rect 15212 7460 15240 7488
rect 15841 7463 15899 7469
rect 15841 7460 15853 7463
rect 15212 7432 15853 7460
rect 15841 7429 15853 7432
rect 15887 7429 15899 7463
rect 15841 7423 15899 7429
rect 17497 7463 17555 7469
rect 17497 7429 17509 7463
rect 17543 7460 17555 7463
rect 18322 7460 18328 7472
rect 17543 7432 18328 7460
rect 17543 7429 17555 7432
rect 17497 7423 17555 7429
rect 18322 7420 18328 7432
rect 18380 7420 18386 7472
rect 13633 7395 13691 7401
rect 13633 7361 13645 7395
rect 13679 7361 13691 7395
rect 16393 7395 16451 7401
rect 16393 7392 16405 7395
rect 13633 7355 13691 7361
rect 15580 7364 16405 7392
rect 14277 7327 14335 7333
rect 13280 7296 14136 7324
rect 11974 7216 11980 7268
rect 12032 7256 12038 7268
rect 12032 7228 12388 7256
rect 12032 7216 12038 7228
rect 8260 7160 8305 7188
rect 8404 7160 11928 7188
rect 8260 7148 8266 7160
rect 12066 7148 12072 7200
rect 12124 7188 12130 7200
rect 12253 7191 12311 7197
rect 12253 7188 12265 7191
rect 12124 7160 12265 7188
rect 12124 7148 12130 7160
rect 12253 7157 12265 7160
rect 12299 7157 12311 7191
rect 12360 7188 12388 7228
rect 12802 7216 12808 7268
rect 12860 7256 12866 7268
rect 13449 7259 13507 7265
rect 13449 7256 13461 7259
rect 12860 7228 13461 7256
rect 12860 7216 12866 7228
rect 13449 7225 13461 7228
rect 13495 7256 13507 7259
rect 13998 7256 14004 7268
rect 13495 7228 14004 7256
rect 13495 7225 13507 7228
rect 13449 7219 13507 7225
rect 13998 7216 14004 7228
rect 14056 7216 14062 7268
rect 14108 7256 14136 7296
rect 14277 7293 14289 7327
rect 14323 7324 14335 7327
rect 14366 7324 14372 7336
rect 14323 7296 14372 7324
rect 14323 7293 14335 7296
rect 14277 7287 14335 7293
rect 14366 7284 14372 7296
rect 14424 7284 14430 7336
rect 15378 7324 15384 7336
rect 14476 7296 15384 7324
rect 14476 7256 14504 7296
rect 15378 7284 15384 7296
rect 15436 7284 15442 7336
rect 14108 7228 14504 7256
rect 14544 7259 14602 7265
rect 14544 7225 14556 7259
rect 14590 7225 14602 7259
rect 15580 7256 15608 7364
rect 16393 7361 16405 7364
rect 16439 7361 16451 7395
rect 18138 7392 18144 7404
rect 18099 7364 18144 7392
rect 16393 7355 16451 7361
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 15654 7284 15660 7336
rect 15712 7284 15718 7336
rect 15838 7284 15844 7336
rect 15896 7324 15902 7336
rect 16482 7324 16488 7336
rect 15896 7296 16488 7324
rect 15896 7284 15902 7296
rect 16482 7284 16488 7296
rect 16540 7284 16546 7336
rect 16666 7324 16672 7336
rect 16627 7296 16672 7324
rect 16666 7284 16672 7296
rect 16724 7324 16730 7336
rect 17313 7327 17371 7333
rect 17313 7324 17325 7327
rect 16724 7296 17325 7324
rect 16724 7284 16730 7296
rect 17313 7293 17325 7296
rect 17359 7293 17371 7327
rect 17313 7287 17371 7293
rect 17402 7284 17408 7336
rect 17460 7324 17466 7336
rect 17589 7327 17647 7333
rect 17589 7324 17601 7327
rect 17460 7296 17601 7324
rect 17460 7284 17466 7296
rect 17589 7293 17601 7296
rect 17635 7293 17647 7327
rect 17589 7287 17647 7293
rect 17957 7327 18015 7333
rect 17957 7293 17969 7327
rect 18003 7324 18015 7327
rect 18046 7324 18052 7336
rect 18003 7296 18052 7324
rect 18003 7293 18015 7296
rect 17957 7287 18015 7293
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 14544 7219 14602 7225
rect 15396 7228 15608 7256
rect 13081 7191 13139 7197
rect 13081 7188 13093 7191
rect 12360 7160 13093 7188
rect 12253 7151 12311 7157
rect 13081 7157 13093 7160
rect 13127 7157 13139 7191
rect 13081 7151 13139 7157
rect 13630 7148 13636 7200
rect 13688 7188 13694 7200
rect 13909 7191 13967 7197
rect 13909 7188 13921 7191
rect 13688 7160 13921 7188
rect 13688 7148 13694 7160
rect 13909 7157 13921 7160
rect 13955 7157 13967 7191
rect 14559 7188 14587 7219
rect 15396 7200 15424 7228
rect 15378 7188 15384 7200
rect 14559 7160 15384 7188
rect 13909 7151 13967 7157
rect 15378 7148 15384 7160
rect 15436 7148 15442 7200
rect 15672 7197 15700 7284
rect 16209 7259 16267 7265
rect 16209 7225 16221 7259
rect 16255 7256 16267 7259
rect 17218 7256 17224 7268
rect 16255 7228 17224 7256
rect 16255 7225 16267 7228
rect 16209 7219 16267 7225
rect 17218 7216 17224 7228
rect 17276 7216 17282 7268
rect 17494 7216 17500 7268
rect 17552 7256 17558 7268
rect 18325 7259 18383 7265
rect 18325 7256 18337 7259
rect 17552 7228 18337 7256
rect 17552 7216 17558 7228
rect 18325 7225 18337 7228
rect 18371 7225 18383 7259
rect 18506 7256 18512 7268
rect 18467 7228 18512 7256
rect 18325 7219 18383 7225
rect 18506 7216 18512 7228
rect 18564 7216 18570 7268
rect 15657 7191 15715 7197
rect 15657 7157 15669 7191
rect 15703 7157 15715 7191
rect 15657 7151 15715 7157
rect 16298 7148 16304 7200
rect 16356 7188 16362 7200
rect 17126 7188 17132 7200
rect 16356 7160 16401 7188
rect 17087 7160 17132 7188
rect 16356 7148 16362 7160
rect 17126 7148 17132 7160
rect 17184 7148 17190 7200
rect 17770 7188 17776 7200
rect 17731 7160 17776 7188
rect 17770 7148 17776 7160
rect 17828 7148 17834 7200
rect 1104 7098 18860 7120
rect 1104 7046 6912 7098
rect 6964 7046 6976 7098
rect 7028 7046 7040 7098
rect 7092 7046 7104 7098
rect 7156 7046 12843 7098
rect 12895 7046 12907 7098
rect 12959 7046 12971 7098
rect 13023 7046 13035 7098
rect 13087 7046 18860 7098
rect 1104 7024 18860 7046
rect 3513 6987 3571 6993
rect 3513 6984 3525 6987
rect 2884 6956 3525 6984
rect 2498 6876 2504 6928
rect 2556 6916 2562 6928
rect 2774 6916 2780 6928
rect 2556 6888 2780 6916
rect 2556 6876 2562 6888
rect 2774 6876 2780 6888
rect 2832 6876 2838 6928
rect 1581 6851 1639 6857
rect 1581 6817 1593 6851
rect 1627 6817 1639 6851
rect 1762 6848 1768 6860
rect 1723 6820 1768 6848
rect 1581 6811 1639 6817
rect 1596 6780 1624 6811
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 2884 6857 2912 6956
rect 3513 6953 3525 6956
rect 3559 6984 3571 6987
rect 5721 6987 5779 6993
rect 3559 6956 5672 6984
rect 3559 6953 3571 6956
rect 3513 6947 3571 6953
rect 2958 6876 2964 6928
rect 3016 6916 3022 6928
rect 3329 6919 3387 6925
rect 3329 6916 3341 6919
rect 3016 6888 3341 6916
rect 3016 6876 3022 6888
rect 3329 6885 3341 6888
rect 3375 6916 3387 6919
rect 5644 6916 5672 6956
rect 5721 6953 5733 6987
rect 5767 6984 5779 6987
rect 6270 6984 6276 6996
rect 5767 6956 6276 6984
rect 5767 6953 5779 6956
rect 5721 6947 5779 6953
rect 6270 6944 6276 6956
rect 6328 6944 6334 6996
rect 7742 6984 7748 6996
rect 7703 6956 7748 6984
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 8113 6987 8171 6993
rect 8113 6953 8125 6987
rect 8159 6984 8171 6987
rect 8202 6984 8208 6996
rect 8159 6956 8208 6984
rect 8159 6953 8171 6956
rect 8113 6947 8171 6953
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 8294 6944 8300 6996
rect 8352 6984 8358 6996
rect 11238 6984 11244 6996
rect 8352 6956 11244 6984
rect 8352 6944 8358 6956
rect 11238 6944 11244 6956
rect 11296 6944 11302 6996
rect 11974 6984 11980 6996
rect 11935 6956 11980 6984
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 12805 6987 12863 6993
rect 12805 6984 12817 6987
rect 12400 6956 12817 6984
rect 12400 6944 12406 6956
rect 12805 6953 12817 6956
rect 12851 6953 12863 6987
rect 13630 6984 13636 6996
rect 13591 6956 13636 6984
rect 12805 6947 12863 6953
rect 13630 6944 13636 6956
rect 13688 6944 13694 6996
rect 15010 6984 15016 6996
rect 13740 6956 15016 6984
rect 7374 6916 7380 6928
rect 3375 6888 5212 6916
rect 5644 6888 7380 6916
rect 3375 6885 3387 6888
rect 3329 6879 3387 6885
rect 1949 6851 2007 6857
rect 1949 6817 1961 6851
rect 1995 6848 2007 6851
rect 2317 6851 2375 6857
rect 1995 6820 2268 6848
rect 1995 6817 2007 6820
rect 1949 6811 2007 6817
rect 1596 6752 2176 6780
rect 2148 6721 2176 6752
rect 2133 6715 2191 6721
rect 2133 6681 2145 6715
rect 2179 6681 2191 6715
rect 2133 6675 2191 6681
rect 1486 6644 1492 6656
rect 1447 6616 1492 6644
rect 1486 6604 1492 6616
rect 1544 6604 1550 6656
rect 2240 6644 2268 6820
rect 2317 6817 2329 6851
rect 2363 6817 2375 6851
rect 2317 6811 2375 6817
rect 2593 6851 2651 6857
rect 2593 6817 2605 6851
rect 2639 6817 2651 6851
rect 2593 6811 2651 6817
rect 2869 6851 2927 6857
rect 2869 6817 2881 6851
rect 2915 6817 2927 6851
rect 2869 6811 2927 6817
rect 2332 6712 2360 6811
rect 2608 6780 2636 6811
rect 3510 6808 3516 6860
rect 3568 6848 3574 6860
rect 4597 6851 4655 6857
rect 4597 6848 4609 6851
rect 3568 6820 4609 6848
rect 3568 6808 3574 6820
rect 4597 6817 4609 6820
rect 4643 6817 4655 6851
rect 5184 6848 5212 6888
rect 7374 6876 7380 6888
rect 7432 6876 7438 6928
rect 7650 6916 7656 6928
rect 7611 6888 7656 6916
rect 7650 6876 7656 6888
rect 7708 6876 7714 6928
rect 8481 6919 8539 6925
rect 8481 6916 8493 6919
rect 8220 6888 8493 6916
rect 8220 6860 8248 6888
rect 8481 6885 8493 6888
rect 8527 6885 8539 6919
rect 8481 6879 8539 6885
rect 11054 6876 11060 6928
rect 11112 6876 11118 6928
rect 11149 6919 11207 6925
rect 11149 6885 11161 6919
rect 11195 6916 11207 6919
rect 12897 6919 12955 6925
rect 11195 6888 12296 6916
rect 11195 6885 11207 6888
rect 11149 6879 11207 6885
rect 6914 6848 6920 6860
rect 5184 6820 6920 6848
rect 4597 6811 4655 6817
rect 6914 6808 6920 6820
rect 6972 6808 6978 6860
rect 7193 6851 7251 6857
rect 7193 6817 7205 6851
rect 7239 6848 7251 6851
rect 7558 6848 7564 6860
rect 7239 6820 7564 6848
rect 7239 6817 7251 6820
rect 7193 6811 7251 6817
rect 7558 6808 7564 6820
rect 7616 6848 7622 6860
rect 8202 6848 8208 6860
rect 7616 6820 8208 6848
rect 7616 6808 7622 6820
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 8573 6851 8631 6857
rect 8573 6817 8585 6851
rect 8619 6848 8631 6851
rect 8941 6851 8999 6857
rect 8941 6848 8953 6851
rect 8619 6820 8953 6848
rect 8619 6817 8631 6820
rect 8573 6811 8631 6817
rect 8941 6817 8953 6820
rect 8987 6817 8999 6851
rect 11072 6848 11100 6876
rect 11882 6848 11888 6860
rect 8941 6811 8999 6817
rect 10980 6820 11888 6848
rect 2608 6752 3740 6780
rect 2961 6715 3019 6721
rect 2961 6712 2973 6715
rect 2332 6684 2973 6712
rect 2961 6681 2973 6684
rect 3007 6712 3019 6715
rect 3602 6712 3608 6724
rect 3007 6684 3608 6712
rect 3007 6681 3019 6684
rect 2961 6675 3019 6681
rect 3602 6672 3608 6684
rect 3660 6672 3666 6724
rect 2409 6647 2467 6653
rect 2409 6644 2421 6647
rect 2240 6616 2421 6644
rect 2409 6613 2421 6616
rect 2455 6613 2467 6647
rect 2409 6607 2467 6613
rect 2498 6604 2504 6656
rect 2556 6644 2562 6656
rect 2685 6647 2743 6653
rect 2685 6644 2697 6647
rect 2556 6616 2697 6644
rect 2556 6604 2562 6616
rect 2685 6613 2697 6616
rect 2731 6613 2743 6647
rect 2685 6607 2743 6613
rect 3237 6647 3295 6653
rect 3237 6613 3249 6647
rect 3283 6644 3295 6647
rect 3712 6644 3740 6752
rect 4246 6740 4252 6792
rect 4304 6780 4310 6792
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 4304 6752 4353 6780
rect 4304 6740 4310 6752
rect 4341 6749 4353 6752
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6780 6423 6783
rect 6822 6780 6828 6792
rect 6411 6752 6828 6780
rect 6411 6749 6423 6752
rect 6365 6743 6423 6749
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 7944 6712 7972 6743
rect 8294 6740 8300 6792
rect 8352 6780 8358 6792
rect 8588 6780 8616 6811
rect 8754 6780 8760 6792
rect 8352 6752 8616 6780
rect 8715 6752 8760 6780
rect 8352 6740 8358 6752
rect 8754 6740 8760 6752
rect 8812 6740 8818 6792
rect 9122 6780 9128 6792
rect 9083 6752 9128 6780
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 10980 6789 11008 6820
rect 11882 6808 11888 6820
rect 11940 6848 11946 6860
rect 11940 6820 12204 6848
rect 11940 6808 11946 6820
rect 10965 6783 11023 6789
rect 10965 6749 10977 6783
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6749 11115 6783
rect 12066 6780 12072 6792
rect 12027 6752 12072 6780
rect 11057 6743 11115 6749
rect 10134 6712 10140 6724
rect 7944 6684 10140 6712
rect 10134 6672 10140 6684
rect 10192 6672 10198 6724
rect 11072 6712 11100 6743
rect 12066 6740 12072 6752
rect 12124 6740 12130 6792
rect 12176 6789 12204 6820
rect 12161 6783 12219 6789
rect 12161 6749 12173 6783
rect 12207 6749 12219 6783
rect 12268 6780 12296 6888
rect 12897 6885 12909 6919
rect 12943 6916 12955 6919
rect 13262 6916 13268 6928
rect 12943 6888 13268 6916
rect 12943 6885 12955 6888
rect 12897 6879 12955 6885
rect 13262 6876 13268 6888
rect 13320 6916 13326 6928
rect 13740 6916 13768 6956
rect 15010 6944 15016 6956
rect 15068 6944 15074 6996
rect 15378 6944 15384 6996
rect 15436 6984 15442 6996
rect 15749 6987 15807 6993
rect 15749 6984 15761 6987
rect 15436 6956 15761 6984
rect 15436 6944 15442 6956
rect 15749 6953 15761 6956
rect 15795 6984 15807 6987
rect 16114 6984 16120 6996
rect 15795 6956 16120 6984
rect 15795 6953 15807 6956
rect 15749 6947 15807 6953
rect 16114 6944 16120 6956
rect 16172 6944 16178 6996
rect 16298 6944 16304 6996
rect 16356 6984 16362 6996
rect 16393 6987 16451 6993
rect 16393 6984 16405 6987
rect 16356 6956 16405 6984
rect 16356 6944 16362 6956
rect 16393 6953 16405 6956
rect 16439 6953 16451 6987
rect 16393 6947 16451 6953
rect 16574 6944 16580 6996
rect 16632 6984 16638 6996
rect 16853 6987 16911 6993
rect 16853 6984 16865 6987
rect 16632 6956 16865 6984
rect 16632 6944 16638 6956
rect 16853 6953 16865 6956
rect 16899 6984 16911 6987
rect 16942 6984 16948 6996
rect 16899 6956 16948 6984
rect 16899 6953 16911 6956
rect 16853 6947 16911 6953
rect 16942 6944 16948 6956
rect 17000 6944 17006 6996
rect 17126 6944 17132 6996
rect 17184 6984 17190 6996
rect 17589 6987 17647 6993
rect 17589 6984 17601 6987
rect 17184 6956 17601 6984
rect 17184 6944 17190 6956
rect 17589 6953 17601 6956
rect 17635 6953 17647 6987
rect 17589 6947 17647 6953
rect 13320 6888 13768 6916
rect 13320 6876 13326 6888
rect 13814 6876 13820 6928
rect 13872 6916 13878 6928
rect 16025 6919 16083 6925
rect 16025 6916 16037 6919
rect 13872 6888 16037 6916
rect 13872 6876 13878 6888
rect 16025 6885 16037 6888
rect 16071 6916 16083 6919
rect 17310 6916 17316 6928
rect 16071 6888 17316 6916
rect 16071 6885 16083 6888
rect 16025 6879 16083 6885
rect 17310 6876 17316 6888
rect 17368 6876 17374 6928
rect 13725 6851 13783 6857
rect 13004 6820 13676 6848
rect 12268 6752 12572 6780
rect 12161 6743 12219 6749
rect 12437 6715 12495 6721
rect 12437 6712 12449 6715
rect 11072 6684 12449 6712
rect 12437 6681 12449 6684
rect 12483 6681 12495 6715
rect 12544 6712 12572 6752
rect 12802 6740 12808 6792
rect 12860 6780 12866 6792
rect 13004 6789 13032 6820
rect 12989 6783 13047 6789
rect 12989 6780 13001 6783
rect 12860 6752 13001 6780
rect 12860 6740 12866 6752
rect 12989 6749 13001 6752
rect 13035 6749 13047 6783
rect 12989 6743 13047 6749
rect 13078 6740 13084 6792
rect 13136 6780 13142 6792
rect 13648 6780 13676 6820
rect 13725 6817 13737 6851
rect 13771 6848 13783 6851
rect 14185 6851 14243 6857
rect 14185 6848 14197 6851
rect 13771 6820 14197 6848
rect 13771 6817 13783 6820
rect 13725 6811 13783 6817
rect 14185 6817 14197 6820
rect 14231 6848 14243 6851
rect 14274 6848 14280 6860
rect 14231 6820 14280 6848
rect 14231 6817 14243 6820
rect 14185 6811 14243 6817
rect 14274 6808 14280 6820
rect 14332 6808 14338 6860
rect 14636 6851 14694 6857
rect 14636 6817 14648 6851
rect 14682 6848 14694 6851
rect 15378 6848 15384 6860
rect 14682 6820 15384 6848
rect 14682 6817 14694 6820
rect 14636 6811 14694 6817
rect 15378 6808 15384 6820
rect 15436 6808 15442 6860
rect 15746 6808 15752 6860
rect 15804 6848 15810 6860
rect 15841 6851 15899 6857
rect 15841 6848 15853 6851
rect 15804 6820 15853 6848
rect 15804 6808 15810 6820
rect 15841 6817 15853 6820
rect 15887 6848 15899 6851
rect 16574 6848 16580 6860
rect 15887 6820 16580 6848
rect 15887 6817 15899 6820
rect 15841 6811 15899 6817
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 16666 6808 16672 6860
rect 16724 6848 16730 6860
rect 16761 6851 16819 6857
rect 16761 6848 16773 6851
rect 16724 6820 16773 6848
rect 16724 6808 16730 6820
rect 16761 6817 16773 6820
rect 16807 6817 16819 6851
rect 18322 6848 18328 6860
rect 16761 6811 16819 6817
rect 17052 6820 17816 6848
rect 18283 6820 18328 6848
rect 13817 6783 13875 6789
rect 13817 6780 13829 6783
rect 13136 6752 13400 6780
rect 13648 6752 13829 6780
rect 13136 6740 13142 6752
rect 13265 6715 13323 6721
rect 13265 6712 13277 6715
rect 12544 6684 13277 6712
rect 12437 6675 12495 6681
rect 13265 6681 13277 6684
rect 13311 6681 13323 6715
rect 13372 6712 13400 6752
rect 13817 6749 13829 6752
rect 13863 6749 13875 6783
rect 14366 6780 14372 6792
rect 14327 6752 14372 6780
rect 13817 6743 13875 6749
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 16942 6780 16948 6792
rect 15396 6752 16948 6780
rect 13372 6684 13952 6712
rect 13265 6675 13323 6681
rect 5258 6644 5264 6656
rect 3283 6616 5264 6644
rect 3283 6613 3295 6616
rect 3237 6607 3295 6613
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 7285 6647 7343 6653
rect 7285 6613 7297 6647
rect 7331 6644 7343 6647
rect 7466 6644 7472 6656
rect 7331 6616 7472 6644
rect 7331 6613 7343 6616
rect 7285 6607 7343 6613
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 8941 6647 8999 6653
rect 8941 6613 8953 6647
rect 8987 6644 8999 6647
rect 9493 6647 9551 6653
rect 9493 6644 9505 6647
rect 8987 6616 9505 6644
rect 8987 6613 8999 6616
rect 8941 6607 8999 6613
rect 9493 6613 9505 6616
rect 9539 6644 9551 6647
rect 11330 6644 11336 6656
rect 9539 6616 11336 6644
rect 9539 6613 9551 6616
rect 9493 6607 9551 6613
rect 11330 6604 11336 6616
rect 11388 6604 11394 6656
rect 11514 6644 11520 6656
rect 11475 6616 11520 6644
rect 11514 6604 11520 6616
rect 11572 6604 11578 6656
rect 11609 6647 11667 6653
rect 11609 6613 11621 6647
rect 11655 6644 11667 6647
rect 11974 6644 11980 6656
rect 11655 6616 11980 6644
rect 11655 6613 11667 6616
rect 11609 6607 11667 6613
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 13924 6644 13952 6684
rect 15396 6644 15424 6752
rect 16942 6740 16948 6752
rect 17000 6740 17006 6792
rect 17052 6789 17080 6820
rect 17037 6783 17095 6789
rect 17037 6749 17049 6783
rect 17083 6749 17095 6783
rect 17037 6743 17095 6749
rect 16482 6672 16488 6724
rect 16540 6712 16546 6724
rect 17052 6712 17080 6743
rect 17126 6740 17132 6792
rect 17184 6780 17190 6792
rect 17788 6789 17816 6820
rect 18322 6808 18328 6820
rect 18380 6808 18386 6860
rect 17681 6783 17739 6789
rect 17681 6780 17693 6783
rect 17184 6752 17693 6780
rect 17184 6740 17190 6752
rect 17681 6749 17693 6752
rect 17727 6749 17739 6783
rect 17681 6743 17739 6749
rect 17773 6783 17831 6789
rect 17773 6749 17785 6783
rect 17819 6749 17831 6783
rect 17773 6743 17831 6749
rect 17218 6712 17224 6724
rect 16540 6684 17080 6712
rect 17179 6684 17224 6712
rect 16540 6672 16546 6684
rect 17218 6672 17224 6684
rect 17276 6672 17282 6724
rect 18506 6712 18512 6724
rect 18467 6684 18512 6712
rect 18506 6672 18512 6684
rect 18564 6672 18570 6724
rect 13924 6616 15424 6644
rect 16301 6647 16359 6653
rect 16301 6613 16313 6647
rect 16347 6644 16359 6647
rect 16390 6644 16396 6656
rect 16347 6616 16396 6644
rect 16347 6613 16359 6616
rect 16301 6607 16359 6613
rect 16390 6604 16396 6616
rect 16448 6644 16454 6656
rect 16666 6644 16672 6656
rect 16448 6616 16672 6644
rect 16448 6604 16454 6616
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 18046 6644 18052 6656
rect 18007 6616 18052 6644
rect 18046 6604 18052 6616
rect 18104 6604 18110 6656
rect 1104 6554 18860 6576
rect 1104 6502 3947 6554
rect 3999 6502 4011 6554
rect 4063 6502 4075 6554
rect 4127 6502 4139 6554
rect 4191 6502 9878 6554
rect 9930 6502 9942 6554
rect 9994 6502 10006 6554
rect 10058 6502 10070 6554
rect 10122 6502 15808 6554
rect 15860 6502 15872 6554
rect 15924 6502 15936 6554
rect 15988 6502 16000 6554
rect 16052 6502 18860 6554
rect 1104 6480 18860 6502
rect 3510 6440 3516 6452
rect 3471 6412 3516 6440
rect 3510 6400 3516 6412
rect 3568 6400 3574 6452
rect 3602 6400 3608 6452
rect 3660 6440 3666 6452
rect 7834 6440 7840 6452
rect 3660 6412 7840 6440
rect 3660 6400 3666 6412
rect 7834 6400 7840 6412
rect 7892 6400 7898 6452
rect 8021 6443 8079 6449
rect 8021 6409 8033 6443
rect 8067 6440 8079 6443
rect 8110 6440 8116 6452
rect 8067 6412 8116 6440
rect 8067 6409 8079 6412
rect 8021 6403 8079 6409
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 10778 6440 10784 6452
rect 8220 6412 10784 6440
rect 4890 6332 4896 6384
rect 4948 6372 4954 6384
rect 5261 6375 5319 6381
rect 5261 6372 5273 6375
rect 4948 6344 5273 6372
rect 4948 6332 4954 6344
rect 5261 6341 5273 6344
rect 5307 6372 5319 6375
rect 5810 6372 5816 6384
rect 5307 6344 5816 6372
rect 5307 6341 5319 6344
rect 5261 6335 5319 6341
rect 5810 6332 5816 6344
rect 5868 6372 5874 6384
rect 7650 6372 7656 6384
rect 5868 6344 7656 6372
rect 5868 6332 5874 6344
rect 7650 6332 7656 6344
rect 7708 6332 7714 6384
rect 3418 6304 3424 6316
rect 3379 6276 3424 6304
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 4982 6304 4988 6316
rect 4816 6276 4988 6304
rect 1946 6236 1952 6248
rect 1907 6208 1952 6236
rect 1946 6196 1952 6208
rect 2004 6196 2010 6248
rect 3165 6239 3223 6245
rect 3165 6205 3177 6239
rect 3211 6236 3223 6239
rect 4816 6236 4844 6276
rect 4982 6264 4988 6276
rect 5040 6304 5046 6316
rect 6089 6307 6147 6313
rect 6089 6304 6101 6307
rect 5040 6276 6101 6304
rect 5040 6264 5046 6276
rect 6089 6273 6101 6276
rect 6135 6304 6147 6307
rect 7009 6307 7067 6313
rect 7009 6304 7021 6307
rect 6135 6276 7021 6304
rect 6135 6273 6147 6276
rect 6089 6267 6147 6273
rect 7009 6273 7021 6276
rect 7055 6273 7067 6307
rect 8220 6304 8248 6412
rect 10778 6400 10784 6412
rect 10836 6400 10842 6452
rect 14737 6443 14795 6449
rect 14737 6440 14749 6443
rect 10888 6412 14749 6440
rect 8386 6332 8392 6384
rect 8444 6372 8450 6384
rect 9217 6375 9275 6381
rect 9217 6372 9229 6375
rect 8444 6344 9229 6372
rect 8444 6332 8450 6344
rect 9217 6341 9229 6344
rect 9263 6341 9275 6375
rect 10686 6372 10692 6384
rect 10647 6344 10692 6372
rect 9217 6335 9275 6341
rect 10686 6332 10692 6344
rect 10744 6332 10750 6384
rect 7009 6267 7067 6273
rect 7300 6276 8248 6304
rect 8665 6307 8723 6313
rect 3211 6208 4844 6236
rect 4886 6239 4944 6245
rect 3211 6205 3223 6208
rect 3165 6199 3223 6205
rect 4886 6205 4898 6239
rect 4932 6236 4944 6239
rect 5534 6236 5540 6248
rect 4932 6208 5540 6236
rect 4932 6205 4944 6208
rect 4886 6199 4944 6205
rect 1581 6171 1639 6177
rect 1581 6137 1593 6171
rect 1627 6168 1639 6171
rect 4626 6171 4684 6177
rect 4626 6168 4638 6171
rect 1627 6140 1808 6168
rect 1627 6137 1639 6140
rect 1581 6131 1639 6137
rect 1486 6100 1492 6112
rect 1447 6072 1492 6100
rect 1486 6060 1492 6072
rect 1544 6060 1550 6112
rect 1780 6109 1808 6140
rect 3344 6140 4638 6168
rect 3344 6112 3372 6140
rect 4626 6137 4638 6140
rect 4672 6137 4684 6171
rect 4626 6131 4684 6137
rect 1765 6103 1823 6109
rect 1765 6069 1777 6103
rect 1811 6069 1823 6103
rect 1765 6063 1823 6069
rect 2041 6103 2099 6109
rect 2041 6069 2053 6103
rect 2087 6100 2099 6103
rect 3326 6100 3332 6112
rect 2087 6072 3332 6100
rect 2087 6069 2099 6072
rect 2041 6063 2099 6069
rect 3326 6060 3332 6072
rect 3384 6060 3390 6112
rect 3418 6060 3424 6112
rect 3476 6100 3482 6112
rect 4246 6100 4252 6112
rect 3476 6072 4252 6100
rect 3476 6060 3482 6072
rect 4246 6060 4252 6072
rect 4304 6100 4310 6112
rect 4901 6100 4929 6199
rect 5534 6196 5540 6208
rect 5592 6196 5598 6248
rect 5810 6236 5816 6248
rect 5771 6208 5816 6236
rect 5810 6196 5816 6208
rect 5868 6196 5874 6248
rect 6822 6236 6828 6248
rect 6783 6208 6828 6236
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7300 6245 7328 6276
rect 8665 6273 8677 6307
rect 8711 6304 8723 6307
rect 8754 6304 8760 6316
rect 8711 6276 8760 6304
rect 8711 6273 8723 6276
rect 8665 6267 8723 6273
rect 8754 6264 8760 6276
rect 8812 6264 8818 6316
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 6972 6208 7297 6236
rect 6972 6196 6978 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 8389 6239 8447 6245
rect 8389 6205 8401 6239
rect 8435 6236 8447 6239
rect 9122 6236 9128 6248
rect 8435 6208 9128 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 9122 6196 9128 6208
rect 9180 6196 9186 6248
rect 10318 6196 10324 6248
rect 10376 6245 10382 6248
rect 10376 6236 10388 6245
rect 10597 6239 10655 6245
rect 10376 6208 10421 6236
rect 10376 6199 10388 6208
rect 10597 6205 10609 6239
rect 10643 6236 10655 6239
rect 10778 6236 10784 6248
rect 10643 6208 10784 6236
rect 10643 6205 10655 6208
rect 10597 6199 10655 6205
rect 10376 6196 10382 6199
rect 10778 6196 10784 6208
rect 10836 6196 10842 6248
rect 10888 6245 10916 6412
rect 14737 6409 14749 6412
rect 14783 6409 14795 6443
rect 14737 6403 14795 6409
rect 16393 6443 16451 6449
rect 16393 6409 16405 6443
rect 16439 6440 16451 6443
rect 17129 6443 17187 6449
rect 17129 6440 17141 6443
rect 16439 6412 17141 6440
rect 16439 6409 16451 6412
rect 16393 6403 16451 6409
rect 17129 6409 17141 6412
rect 17175 6409 17187 6443
rect 17494 6440 17500 6452
rect 17455 6412 17500 6440
rect 17129 6403 17187 6409
rect 17494 6400 17500 6412
rect 17552 6400 17558 6452
rect 13170 6372 13176 6384
rect 12728 6344 13176 6372
rect 10873 6239 10931 6245
rect 10873 6205 10885 6239
rect 10919 6205 10931 6239
rect 10873 6199 10931 6205
rect 11330 6196 11336 6248
rect 11388 6236 11394 6248
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 11388 6208 11713 6236
rect 11388 6196 11394 6208
rect 11701 6205 11713 6208
rect 11747 6205 11759 6239
rect 12728 6236 12756 6344
rect 13170 6332 13176 6344
rect 13228 6332 13234 6384
rect 16850 6332 16856 6384
rect 16908 6372 16914 6384
rect 16945 6375 17003 6381
rect 16945 6372 16957 6375
rect 16908 6344 16957 6372
rect 16908 6332 16914 6344
rect 16945 6341 16957 6344
rect 16991 6372 17003 6375
rect 17402 6372 17408 6384
rect 16991 6344 17408 6372
rect 16991 6341 17003 6344
rect 16945 6335 17003 6341
rect 17402 6332 17408 6344
rect 17460 6332 17466 6384
rect 15381 6307 15439 6313
rect 15381 6273 15393 6307
rect 15427 6304 15439 6307
rect 15654 6304 15660 6316
rect 15427 6276 15660 6304
rect 15427 6273 15439 6276
rect 15381 6267 15439 6273
rect 15654 6264 15660 6276
rect 15712 6264 15718 6316
rect 16114 6304 16120 6316
rect 16075 6276 16120 6304
rect 16114 6264 16120 6276
rect 16172 6264 16178 6316
rect 16666 6304 16672 6316
rect 16627 6276 16672 6304
rect 16666 6264 16672 6276
rect 16724 6304 16730 6316
rect 16724 6276 17632 6304
rect 16724 6264 16730 6276
rect 13170 6236 13176 6248
rect 11701 6199 11759 6205
rect 11808 6208 12756 6236
rect 13131 6208 13176 6236
rect 5258 6128 5264 6180
rect 5316 6168 5322 6180
rect 11808 6168 11836 6208
rect 13170 6196 13176 6208
rect 13228 6196 13234 6248
rect 15105 6239 15163 6245
rect 15105 6205 15117 6239
rect 15151 6236 15163 6239
rect 15194 6236 15200 6248
rect 15151 6208 15200 6236
rect 15151 6205 15163 6208
rect 15105 6199 15163 6205
rect 15194 6196 15200 6208
rect 15252 6196 15258 6248
rect 16022 6196 16028 6248
rect 16080 6236 16086 6248
rect 16393 6239 16451 6245
rect 16393 6236 16405 6239
rect 16080 6208 16405 6236
rect 16080 6196 16086 6208
rect 16393 6205 16405 6208
rect 16439 6205 16451 6239
rect 16393 6199 16451 6205
rect 16574 6196 16580 6248
rect 16632 6236 16638 6248
rect 17604 6245 17632 6276
rect 17313 6239 17371 6245
rect 17313 6236 17325 6239
rect 16632 6208 17325 6236
rect 16632 6196 16638 6208
rect 17313 6205 17325 6208
rect 17359 6205 17371 6239
rect 17313 6199 17371 6205
rect 17589 6239 17647 6245
rect 17589 6205 17601 6239
rect 17635 6205 17647 6239
rect 17589 6199 17647 6205
rect 17678 6196 17684 6248
rect 17736 6236 17742 6248
rect 17865 6239 17923 6245
rect 17865 6236 17877 6239
rect 17736 6208 17877 6236
rect 17736 6196 17742 6208
rect 17865 6205 17877 6208
rect 17911 6236 17923 6239
rect 18046 6236 18052 6248
rect 17911 6208 18052 6236
rect 17911 6205 17923 6208
rect 17865 6199 17923 6205
rect 18046 6196 18052 6208
rect 18104 6196 18110 6248
rect 5316 6140 11836 6168
rect 5316 6128 5322 6140
rect 11882 6128 11888 6180
rect 11940 6177 11946 6180
rect 11940 6171 12004 6177
rect 11940 6137 11958 6171
rect 11992 6137 12004 6171
rect 12986 6168 12992 6180
rect 11940 6131 12004 6137
rect 12084 6140 12992 6168
rect 11940 6128 11946 6131
rect 5442 6100 5448 6112
rect 4304 6072 4929 6100
rect 5403 6072 5448 6100
rect 4304 6060 4310 6072
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 5905 6103 5963 6109
rect 5905 6069 5917 6103
rect 5951 6100 5963 6103
rect 5994 6100 6000 6112
rect 5951 6072 6000 6100
rect 5951 6069 5963 6072
rect 5905 6063 5963 6069
rect 5994 6060 6000 6072
rect 6052 6060 6058 6112
rect 6454 6100 6460 6112
rect 6415 6072 6460 6100
rect 6454 6060 6460 6072
rect 6512 6060 6518 6112
rect 7834 6060 7840 6112
rect 7892 6100 7898 6112
rect 8481 6103 8539 6109
rect 8481 6100 8493 6103
rect 7892 6072 8493 6100
rect 7892 6060 7898 6072
rect 8481 6069 8493 6072
rect 8527 6100 8539 6103
rect 8849 6103 8907 6109
rect 8849 6100 8861 6103
rect 8527 6072 8861 6100
rect 8527 6069 8539 6072
rect 8481 6063 8539 6069
rect 8849 6069 8861 6072
rect 8895 6100 8907 6103
rect 12084 6100 12112 6140
rect 12986 6128 12992 6140
rect 13044 6128 13050 6180
rect 13418 6171 13476 6177
rect 13418 6137 13430 6171
rect 13464 6137 13476 6171
rect 17218 6168 17224 6180
rect 13418 6131 13476 6137
rect 14660 6140 17224 6168
rect 8895 6072 12112 6100
rect 8895 6069 8907 6072
rect 8849 6063 8907 6069
rect 12342 6060 12348 6112
rect 12400 6100 12406 6112
rect 13081 6103 13139 6109
rect 13081 6100 13093 6103
rect 12400 6072 13093 6100
rect 12400 6060 12406 6072
rect 13081 6069 13093 6072
rect 13127 6100 13139 6103
rect 13433 6100 13461 6131
rect 14660 6112 14688 6140
rect 17218 6128 17224 6140
rect 17276 6128 17282 6180
rect 18325 6171 18383 6177
rect 18325 6168 18337 6171
rect 17788 6140 18337 6168
rect 13127 6072 13461 6100
rect 14553 6103 14611 6109
rect 13127 6069 13139 6072
rect 13081 6063 13139 6069
rect 14553 6069 14565 6103
rect 14599 6100 14611 6103
rect 14642 6100 14648 6112
rect 14599 6072 14648 6100
rect 14599 6069 14611 6072
rect 14553 6063 14611 6069
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 15197 6103 15255 6109
rect 15197 6069 15209 6103
rect 15243 6100 15255 6103
rect 15565 6103 15623 6109
rect 15565 6100 15577 6103
rect 15243 6072 15577 6100
rect 15243 6069 15255 6072
rect 15197 6063 15255 6069
rect 15565 6069 15577 6072
rect 15611 6069 15623 6103
rect 15565 6063 15623 6069
rect 15838 6060 15844 6112
rect 15896 6100 15902 6112
rect 15933 6103 15991 6109
rect 15933 6100 15945 6103
rect 15896 6072 15945 6100
rect 15896 6060 15902 6072
rect 15933 6069 15945 6072
rect 15979 6069 15991 6103
rect 15933 6063 15991 6069
rect 16025 6103 16083 6109
rect 16025 6069 16037 6103
rect 16071 6100 16083 6103
rect 16114 6100 16120 6112
rect 16071 6072 16120 6100
rect 16071 6069 16083 6072
rect 16025 6063 16083 6069
rect 16114 6060 16120 6072
rect 16172 6060 16178 6112
rect 16390 6060 16396 6112
rect 16448 6100 16454 6112
rect 16485 6103 16543 6109
rect 16485 6100 16497 6103
rect 16448 6072 16497 6100
rect 16448 6060 16454 6072
rect 16485 6069 16497 6072
rect 16531 6100 16543 6103
rect 16574 6100 16580 6112
rect 16531 6072 16580 6100
rect 16531 6069 16543 6072
rect 16485 6063 16543 6069
rect 16574 6060 16580 6072
rect 16632 6060 16638 6112
rect 17788 6109 17816 6140
rect 18325 6137 18337 6140
rect 18371 6137 18383 6171
rect 18506 6168 18512 6180
rect 18467 6140 18512 6168
rect 18325 6131 18383 6137
rect 18506 6128 18512 6140
rect 18564 6128 18570 6180
rect 17773 6103 17831 6109
rect 17773 6069 17785 6103
rect 17819 6069 17831 6103
rect 17773 6063 17831 6069
rect 18049 6103 18107 6109
rect 18049 6069 18061 6103
rect 18095 6100 18107 6103
rect 18230 6100 18236 6112
rect 18095 6072 18236 6100
rect 18095 6069 18107 6072
rect 18049 6063 18107 6069
rect 18230 6060 18236 6072
rect 18288 6060 18294 6112
rect 1104 6010 18860 6032
rect 1104 5958 6912 6010
rect 6964 5958 6976 6010
rect 7028 5958 7040 6010
rect 7092 5958 7104 6010
rect 7156 5958 12843 6010
rect 12895 5958 12907 6010
rect 12959 5958 12971 6010
rect 13023 5958 13035 6010
rect 13087 5958 18860 6010
rect 1104 5936 18860 5958
rect 1765 5899 1823 5905
rect 1765 5896 1777 5899
rect 1596 5868 1777 5896
rect 1596 5837 1624 5868
rect 1765 5865 1777 5868
rect 1811 5865 1823 5899
rect 1765 5859 1823 5865
rect 1946 5856 1952 5908
rect 2004 5896 2010 5908
rect 2501 5899 2559 5905
rect 2501 5896 2513 5899
rect 2004 5868 2513 5896
rect 2004 5856 2010 5868
rect 2501 5865 2513 5868
rect 2547 5896 2559 5899
rect 2685 5899 2743 5905
rect 2685 5896 2697 5899
rect 2547 5868 2697 5896
rect 2547 5865 2559 5868
rect 2501 5859 2559 5865
rect 2685 5865 2697 5868
rect 2731 5865 2743 5899
rect 2685 5859 2743 5865
rect 3329 5899 3387 5905
rect 3329 5865 3341 5899
rect 3375 5896 3387 5899
rect 3881 5899 3939 5905
rect 3881 5896 3893 5899
rect 3375 5868 3893 5896
rect 3375 5865 3387 5868
rect 3329 5859 3387 5865
rect 3881 5865 3893 5868
rect 3927 5865 3939 5899
rect 4246 5896 4252 5908
rect 4207 5868 4252 5896
rect 3881 5859 3939 5865
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 5169 5899 5227 5905
rect 5169 5865 5181 5899
rect 5215 5896 5227 5899
rect 5442 5896 5448 5908
rect 5215 5868 5448 5896
rect 5215 5865 5227 5868
rect 5169 5859 5227 5865
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 5994 5856 6000 5908
rect 6052 5896 6058 5908
rect 6365 5899 6423 5905
rect 6365 5896 6377 5899
rect 6052 5868 6377 5896
rect 6052 5856 6058 5868
rect 6365 5865 6377 5868
rect 6411 5896 6423 5899
rect 7282 5896 7288 5908
rect 6411 5868 7288 5896
rect 6411 5865 6423 5868
rect 6365 5859 6423 5865
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 10778 5856 10784 5908
rect 10836 5896 10842 5908
rect 10962 5896 10968 5908
rect 10836 5868 10968 5896
rect 10836 5856 10842 5868
rect 10962 5856 10968 5868
rect 11020 5896 11026 5908
rect 11330 5896 11336 5908
rect 11020 5868 11336 5896
rect 11020 5856 11026 5868
rect 11330 5856 11336 5868
rect 11388 5856 11394 5908
rect 11514 5856 11520 5908
rect 11572 5896 11578 5908
rect 11885 5899 11943 5905
rect 11885 5896 11897 5899
rect 11572 5868 11897 5896
rect 11572 5856 11578 5868
rect 11885 5865 11897 5868
rect 11931 5865 11943 5899
rect 11885 5859 11943 5865
rect 13173 5899 13231 5905
rect 13173 5865 13185 5899
rect 13219 5896 13231 5899
rect 15654 5896 15660 5908
rect 13219 5868 15660 5896
rect 13219 5865 13231 5868
rect 13173 5859 13231 5865
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 15838 5896 15844 5908
rect 15799 5868 15844 5896
rect 15838 5856 15844 5868
rect 15896 5856 15902 5908
rect 16022 5856 16028 5908
rect 16080 5896 16086 5908
rect 18046 5896 18052 5908
rect 16080 5868 17908 5896
rect 18007 5868 18052 5896
rect 16080 5856 16086 5868
rect 1581 5831 1639 5837
rect 1581 5797 1593 5831
rect 1627 5797 1639 5831
rect 2409 5831 2467 5837
rect 2409 5828 2421 5831
rect 1581 5791 1639 5797
rect 1964 5800 2421 5828
rect 1964 5769 1992 5800
rect 2409 5797 2421 5800
rect 2455 5828 2467 5831
rect 2590 5828 2596 5840
rect 2455 5800 2596 5828
rect 2455 5797 2467 5800
rect 2409 5791 2467 5797
rect 2590 5788 2596 5800
rect 2648 5788 2654 5840
rect 2774 5788 2780 5840
rect 2832 5828 2838 5840
rect 4264 5828 4292 5856
rect 2832 5800 4292 5828
rect 5077 5831 5135 5837
rect 2832 5788 2838 5800
rect 5077 5797 5089 5831
rect 5123 5828 5135 5831
rect 6454 5828 6460 5840
rect 5123 5800 6460 5828
rect 5123 5797 5135 5800
rect 5077 5791 5135 5797
rect 6454 5788 6460 5800
rect 6512 5788 6518 5840
rect 17129 5831 17187 5837
rect 17129 5797 17141 5831
rect 17175 5828 17187 5831
rect 17310 5828 17316 5840
rect 17175 5800 17316 5828
rect 17175 5797 17187 5800
rect 17129 5791 17187 5797
rect 17310 5788 17316 5800
rect 17368 5788 17374 5840
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5729 2007 5763
rect 1949 5723 2007 5729
rect 2225 5763 2283 5769
rect 2225 5729 2237 5763
rect 2271 5760 2283 5763
rect 2866 5760 2872 5772
rect 2271 5732 2872 5760
rect 2271 5729 2283 5732
rect 2225 5723 2283 5729
rect 2866 5720 2872 5732
rect 2924 5720 2930 5772
rect 3326 5720 3332 5772
rect 3384 5760 3390 5772
rect 4341 5763 4399 5769
rect 3384 5732 3556 5760
rect 3384 5720 3390 5732
rect 3418 5692 3424 5704
rect 3379 5664 3424 5692
rect 3418 5652 3424 5664
rect 3476 5652 3482 5704
rect 3528 5701 3556 5732
rect 4341 5729 4353 5763
rect 4387 5760 4399 5763
rect 5810 5760 5816 5772
rect 4387 5732 5816 5760
rect 4387 5729 4399 5732
rect 4341 5723 4399 5729
rect 5810 5720 5816 5732
rect 5868 5720 5874 5772
rect 5997 5763 6055 5769
rect 5997 5729 6009 5763
rect 6043 5760 6055 5763
rect 6086 5760 6092 5772
rect 6043 5732 6092 5760
rect 6043 5729 6055 5732
rect 5997 5723 6055 5729
rect 6086 5720 6092 5732
rect 6144 5720 6150 5772
rect 6730 5720 6736 5772
rect 6788 5760 6794 5772
rect 7377 5763 7435 5769
rect 7377 5760 7389 5763
rect 6788 5732 7389 5760
rect 6788 5720 6794 5732
rect 7377 5729 7389 5732
rect 7423 5760 7435 5763
rect 7926 5760 7932 5772
rect 7423 5732 7932 5760
rect 7423 5729 7435 5732
rect 7377 5723 7435 5729
rect 7926 5720 7932 5732
rect 7984 5760 7990 5772
rect 8846 5760 8852 5772
rect 7984 5732 8852 5760
rect 7984 5720 7990 5732
rect 8846 5720 8852 5732
rect 8904 5720 8910 5772
rect 9122 5720 9128 5772
rect 9180 5760 9186 5772
rect 9180 5732 9225 5760
rect 9180 5720 9186 5732
rect 12250 5720 12256 5772
rect 12308 5760 12314 5772
rect 12345 5763 12403 5769
rect 12345 5760 12357 5763
rect 12308 5732 12357 5760
rect 12308 5720 12314 5732
rect 12345 5729 12357 5732
rect 12391 5729 12403 5763
rect 13262 5760 13268 5772
rect 13223 5732 13268 5760
rect 12345 5723 12403 5729
rect 13262 5720 13268 5732
rect 13320 5720 13326 5772
rect 13906 5720 13912 5772
rect 13964 5760 13970 5772
rect 14642 5769 14648 5772
rect 14093 5763 14151 5769
rect 14093 5760 14105 5763
rect 13964 5732 14105 5760
rect 13964 5720 13970 5732
rect 14093 5729 14105 5732
rect 14139 5729 14151 5763
rect 14636 5760 14648 5769
rect 14603 5732 14648 5760
rect 14093 5723 14151 5729
rect 14636 5723 14648 5732
rect 14642 5720 14648 5723
rect 14700 5720 14706 5772
rect 15654 5720 15660 5772
rect 15712 5760 15718 5772
rect 16022 5760 16028 5772
rect 15712 5732 16028 5760
rect 15712 5720 15718 5732
rect 16022 5720 16028 5732
rect 16080 5760 16086 5772
rect 16209 5763 16267 5769
rect 16209 5760 16221 5763
rect 16080 5732 16221 5760
rect 16080 5720 16086 5732
rect 16209 5729 16221 5732
rect 16255 5729 16267 5763
rect 16209 5723 16267 5729
rect 16301 5763 16359 5769
rect 16301 5729 16313 5763
rect 16347 5760 16359 5763
rect 16574 5760 16580 5772
rect 16347 5732 16580 5760
rect 16347 5729 16359 5732
rect 16301 5723 16359 5729
rect 16574 5720 16580 5732
rect 16632 5720 16638 5772
rect 17037 5763 17095 5769
rect 17037 5729 17049 5763
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 3513 5695 3571 5701
rect 3513 5661 3525 5695
rect 3559 5661 3571 5695
rect 3513 5655 3571 5661
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5692 4583 5695
rect 4982 5692 4988 5704
rect 4571 5664 4988 5692
rect 4571 5661 4583 5664
rect 4525 5655 4583 5661
rect 2685 5627 2743 5633
rect 2685 5593 2697 5627
rect 2731 5624 2743 5627
rect 3528 5624 3556 5655
rect 4982 5652 4988 5664
rect 5040 5652 5046 5704
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5661 5319 5695
rect 5261 5655 5319 5661
rect 5276 5624 5304 5655
rect 5350 5652 5356 5704
rect 5408 5692 5414 5704
rect 11514 5692 11520 5704
rect 5408 5664 11520 5692
rect 5408 5652 5414 5664
rect 11514 5652 11520 5664
rect 11572 5652 11578 5704
rect 11974 5692 11980 5704
rect 11935 5664 11980 5692
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 12161 5695 12219 5701
rect 12161 5661 12173 5695
rect 12207 5661 12219 5695
rect 13170 5692 13176 5704
rect 12161 5655 12219 5661
rect 12544 5664 13176 5692
rect 5994 5624 6000 5636
rect 2731 5596 3464 5624
rect 3528 5596 5304 5624
rect 5368 5596 6000 5624
rect 2731 5593 2743 5596
rect 2685 5587 2743 5593
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 1578 5516 1584 5568
rect 1636 5556 1642 5568
rect 2041 5559 2099 5565
rect 2041 5556 2053 5559
rect 1636 5528 2053 5556
rect 1636 5516 1642 5528
rect 2041 5525 2053 5528
rect 2087 5525 2099 5559
rect 2958 5556 2964 5568
rect 2919 5528 2964 5556
rect 2041 5519 2099 5525
rect 2958 5516 2964 5528
rect 3016 5516 3022 5568
rect 3436 5556 3464 5596
rect 4246 5556 4252 5568
rect 3436 5528 4252 5556
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 4706 5556 4712 5568
rect 4667 5528 4712 5556
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 4798 5516 4804 5568
rect 4856 5556 4862 5568
rect 5368 5556 5396 5596
rect 5994 5584 6000 5596
rect 6052 5584 6058 5636
rect 6917 5627 6975 5633
rect 6917 5593 6929 5627
rect 6963 5624 6975 5627
rect 7926 5624 7932 5636
rect 6963 5596 7932 5624
rect 6963 5593 6975 5596
rect 6917 5587 6975 5593
rect 7926 5584 7932 5596
rect 7984 5584 7990 5636
rect 12066 5624 12072 5636
rect 8036 5596 12072 5624
rect 4856 5528 5396 5556
rect 4856 5516 4862 5528
rect 5534 5516 5540 5568
rect 5592 5556 5598 5568
rect 6181 5559 6239 5565
rect 6181 5556 6193 5559
rect 5592 5528 6193 5556
rect 5592 5516 5598 5528
rect 6181 5525 6193 5528
rect 6227 5556 6239 5559
rect 6270 5556 6276 5568
rect 6227 5528 6276 5556
rect 6227 5525 6239 5528
rect 6181 5519 6239 5525
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 7285 5559 7343 5565
rect 7285 5525 7297 5559
rect 7331 5556 7343 5559
rect 7374 5556 7380 5568
rect 7331 5528 7380 5556
rect 7331 5525 7343 5528
rect 7285 5519 7343 5525
rect 7374 5516 7380 5528
rect 7432 5516 7438 5568
rect 7650 5516 7656 5568
rect 7708 5556 7714 5568
rect 8036 5556 8064 5596
rect 12066 5584 12072 5596
rect 12124 5584 12130 5636
rect 12176 5624 12204 5655
rect 12342 5624 12348 5636
rect 12176 5596 12348 5624
rect 12342 5584 12348 5596
rect 12400 5584 12406 5636
rect 12434 5584 12440 5636
rect 12492 5624 12498 5636
rect 12544 5633 12572 5664
rect 13170 5652 13176 5664
rect 13228 5692 13234 5704
rect 14366 5692 14372 5704
rect 13228 5664 14372 5692
rect 13228 5652 13234 5664
rect 14366 5652 14372 5664
rect 14424 5652 14430 5704
rect 16393 5695 16451 5701
rect 16393 5661 16405 5695
rect 16439 5692 16451 5695
rect 16482 5692 16488 5704
rect 16439 5664 16488 5692
rect 16439 5661 16451 5664
rect 16393 5655 16451 5661
rect 12529 5627 12587 5633
rect 12529 5624 12541 5627
rect 12492 5596 12541 5624
rect 12492 5584 12498 5596
rect 12529 5593 12541 5596
rect 12575 5593 12587 5627
rect 12529 5587 12587 5593
rect 15378 5584 15384 5636
rect 15436 5624 15442 5636
rect 15749 5627 15807 5633
rect 15749 5624 15761 5627
rect 15436 5596 15761 5624
rect 15436 5584 15442 5596
rect 15749 5593 15761 5596
rect 15795 5624 15807 5627
rect 16408 5624 16436 5655
rect 16482 5652 16488 5664
rect 16540 5652 16546 5704
rect 17052 5692 17080 5723
rect 17402 5720 17408 5772
rect 17460 5760 17466 5772
rect 17880 5769 17908 5868
rect 18046 5856 18052 5868
rect 18104 5856 18110 5908
rect 18230 5788 18236 5840
rect 18288 5828 18294 5840
rect 18325 5831 18383 5837
rect 18325 5828 18337 5831
rect 18288 5800 18337 5828
rect 18288 5788 18294 5800
rect 18325 5797 18337 5800
rect 18371 5797 18383 5831
rect 18325 5791 18383 5797
rect 17589 5763 17647 5769
rect 17589 5760 17601 5763
rect 17460 5732 17601 5760
rect 17460 5720 17466 5732
rect 17589 5729 17601 5732
rect 17635 5729 17647 5763
rect 17589 5723 17647 5729
rect 17865 5763 17923 5769
rect 17865 5729 17877 5763
rect 17911 5729 17923 5763
rect 17865 5723 17923 5729
rect 16592 5664 17080 5692
rect 15795 5596 16436 5624
rect 15795 5593 15807 5596
rect 15749 5587 15807 5593
rect 7708 5528 8064 5556
rect 7708 5516 7714 5528
rect 9306 5516 9312 5568
rect 9364 5556 9370 5568
rect 9582 5556 9588 5568
rect 9364 5528 9409 5556
rect 9543 5528 9588 5556
rect 9364 5516 9370 5528
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 10318 5516 10324 5568
rect 10376 5556 10382 5568
rect 11517 5559 11575 5565
rect 11517 5556 11529 5559
rect 10376 5528 11529 5556
rect 10376 5516 10382 5528
rect 11517 5525 11529 5528
rect 11563 5525 11575 5559
rect 11517 5519 11575 5525
rect 11606 5516 11612 5568
rect 11664 5556 11670 5568
rect 13173 5559 13231 5565
rect 13173 5556 13185 5559
rect 11664 5528 13185 5556
rect 11664 5516 11670 5528
rect 13173 5525 13185 5528
rect 13219 5525 13231 5559
rect 13173 5519 13231 5525
rect 13906 5516 13912 5568
rect 13964 5556 13970 5568
rect 16592 5556 16620 5664
rect 17218 5652 17224 5704
rect 17276 5692 17282 5704
rect 17276 5664 17321 5692
rect 17276 5652 17282 5664
rect 18506 5624 18512 5636
rect 18467 5596 18512 5624
rect 18506 5584 18512 5596
rect 18564 5584 18570 5636
rect 13964 5528 16620 5556
rect 16669 5559 16727 5565
rect 13964 5516 13970 5528
rect 16669 5525 16681 5559
rect 16715 5556 16727 5559
rect 16758 5556 16764 5568
rect 16715 5528 16764 5556
rect 16715 5525 16727 5528
rect 16669 5519 16727 5525
rect 16758 5516 16764 5528
rect 16816 5516 16822 5568
rect 17773 5559 17831 5565
rect 17773 5525 17785 5559
rect 17819 5556 17831 5559
rect 17954 5556 17960 5568
rect 17819 5528 17960 5556
rect 17819 5525 17831 5528
rect 17773 5519 17831 5525
rect 17954 5516 17960 5528
rect 18012 5516 18018 5568
rect 1104 5466 18860 5488
rect 1104 5414 3947 5466
rect 3999 5414 4011 5466
rect 4063 5414 4075 5466
rect 4127 5414 4139 5466
rect 4191 5414 9878 5466
rect 9930 5414 9942 5466
rect 9994 5414 10006 5466
rect 10058 5414 10070 5466
rect 10122 5414 15808 5466
rect 15860 5414 15872 5466
rect 15924 5414 15936 5466
rect 15988 5414 16000 5466
rect 16052 5414 18860 5466
rect 1104 5392 18860 5414
rect 2866 5352 2872 5364
rect 2827 5324 2872 5352
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 3418 5312 3424 5364
rect 3476 5352 3482 5364
rect 3697 5355 3755 5361
rect 3697 5352 3709 5355
rect 3476 5324 3709 5352
rect 3476 5312 3482 5324
rect 3697 5321 3709 5324
rect 3743 5321 3755 5355
rect 3697 5315 3755 5321
rect 4893 5355 4951 5361
rect 4893 5321 4905 5355
rect 4939 5352 4951 5355
rect 4982 5352 4988 5364
rect 4939 5324 4988 5352
rect 4939 5321 4951 5324
rect 4893 5315 4951 5321
rect 2409 5287 2467 5293
rect 2409 5253 2421 5287
rect 2455 5253 2467 5287
rect 2409 5247 2467 5253
rect 2777 5287 2835 5293
rect 2777 5253 2789 5287
rect 2823 5284 2835 5287
rect 4798 5284 4804 5296
rect 2823 5256 4804 5284
rect 2823 5253 2835 5256
rect 2777 5247 2835 5253
rect 2424 5216 2452 5247
rect 2792 5216 2820 5247
rect 4798 5244 4804 5256
rect 4856 5244 4862 5296
rect 1596 5188 2452 5216
rect 2516 5188 2820 5216
rect 1394 5148 1400 5160
rect 1355 5120 1400 5148
rect 1394 5108 1400 5120
rect 1452 5108 1458 5160
rect 1596 5157 1624 5188
rect 1581 5151 1639 5157
rect 1581 5117 1593 5151
rect 1627 5117 1639 5151
rect 1581 5111 1639 5117
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5148 2375 5151
rect 2516 5148 2544 5188
rect 2958 5176 2964 5228
rect 3016 5216 3022 5228
rect 3329 5219 3387 5225
rect 3329 5216 3341 5219
rect 3016 5188 3341 5216
rect 3016 5176 3022 5188
rect 3329 5185 3341 5188
rect 3375 5185 3387 5219
rect 3510 5216 3516 5228
rect 3471 5188 3516 5216
rect 3329 5179 3387 5185
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5216 4399 5219
rect 4908 5216 4936 5315
rect 4982 5312 4988 5324
rect 5040 5312 5046 5364
rect 5258 5312 5264 5364
rect 5316 5352 5322 5364
rect 5316 5324 8984 5352
rect 5316 5312 5322 5324
rect 8956 5284 8984 5324
rect 9306 5312 9312 5364
rect 9364 5352 9370 5364
rect 9401 5355 9459 5361
rect 9401 5352 9413 5355
rect 9364 5324 9413 5352
rect 9364 5312 9370 5324
rect 9401 5321 9413 5324
rect 9447 5321 9459 5355
rect 10873 5355 10931 5361
rect 9401 5315 9459 5321
rect 9508 5324 10824 5352
rect 9508 5284 9536 5324
rect 8956 5256 9536 5284
rect 10796 5284 10824 5324
rect 10873 5321 10885 5355
rect 10919 5352 10931 5355
rect 11238 5352 11244 5364
rect 10919 5324 11244 5352
rect 10919 5321 10931 5324
rect 10873 5315 10931 5321
rect 11238 5312 11244 5324
rect 11296 5312 11302 5364
rect 11330 5312 11336 5364
rect 11388 5352 11394 5364
rect 14553 5355 14611 5361
rect 14553 5352 14565 5355
rect 11388 5324 14565 5352
rect 11388 5312 11394 5324
rect 14553 5321 14565 5324
rect 14599 5352 14611 5355
rect 14642 5352 14648 5364
rect 14599 5324 14648 5352
rect 14599 5321 14611 5324
rect 14553 5315 14611 5321
rect 14642 5312 14648 5324
rect 14700 5312 14706 5364
rect 14829 5355 14887 5361
rect 14829 5321 14841 5355
rect 14875 5352 14887 5355
rect 15013 5355 15071 5361
rect 15013 5352 15025 5355
rect 14875 5324 15025 5352
rect 14875 5321 14887 5324
rect 14829 5315 14887 5321
rect 15013 5321 15025 5324
rect 15059 5352 15071 5355
rect 15102 5352 15108 5364
rect 15059 5324 15108 5352
rect 15059 5321 15071 5324
rect 15013 5315 15071 5321
rect 15102 5312 15108 5324
rect 15160 5352 15166 5364
rect 15378 5352 15384 5364
rect 15160 5324 15384 5352
rect 15160 5312 15166 5324
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 15654 5352 15660 5364
rect 15615 5324 15660 5352
rect 15654 5312 15660 5324
rect 15712 5312 15718 5364
rect 16025 5355 16083 5361
rect 16025 5321 16037 5355
rect 16071 5352 16083 5355
rect 16114 5352 16120 5364
rect 16071 5324 16120 5352
rect 16071 5321 16083 5324
rect 16025 5315 16083 5321
rect 16114 5312 16120 5324
rect 16172 5312 16178 5364
rect 16298 5312 16304 5364
rect 16356 5352 16362 5364
rect 16356 5324 17172 5352
rect 16356 5312 16362 5324
rect 11882 5284 11888 5296
rect 10796 5256 11888 5284
rect 11882 5244 11888 5256
rect 11940 5244 11946 5296
rect 12437 5287 12495 5293
rect 12437 5253 12449 5287
rect 12483 5284 12495 5287
rect 15289 5287 15347 5293
rect 15289 5284 15301 5287
rect 12483 5256 15301 5284
rect 12483 5253 12495 5256
rect 12437 5247 12495 5253
rect 15289 5253 15301 5256
rect 15335 5284 15347 5287
rect 16390 5284 16396 5296
rect 15335 5256 16396 5284
rect 15335 5253 15347 5256
rect 15289 5247 15347 5253
rect 16390 5244 16396 5256
rect 16448 5244 16454 5296
rect 4387 5188 4936 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 9306 5176 9312 5228
rect 9364 5216 9370 5228
rect 9364 5188 9628 5216
rect 9364 5176 9370 5188
rect 2363 5120 2544 5148
rect 2593 5151 2651 5157
rect 2363 5117 2375 5120
rect 2317 5111 2375 5117
rect 2593 5117 2605 5151
rect 2639 5117 2651 5151
rect 2593 5111 2651 5117
rect 3237 5151 3295 5157
rect 3237 5117 3249 5151
rect 3283 5148 3295 5151
rect 4706 5148 4712 5160
rect 3283 5120 4712 5148
rect 3283 5117 3295 5120
rect 3237 5111 3295 5117
rect 1946 5080 1952 5092
rect 1907 5052 1952 5080
rect 1946 5040 1952 5052
rect 2004 5040 2010 5092
rect 2608 5080 2636 5111
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 6270 5148 6276 5160
rect 6183 5120 6276 5148
rect 6270 5108 6276 5120
rect 6328 5108 6334 5160
rect 7581 5151 7639 5157
rect 7581 5117 7593 5151
rect 7627 5148 7639 5151
rect 7742 5148 7748 5160
rect 7627 5120 7748 5148
rect 7627 5117 7639 5120
rect 7581 5111 7639 5117
rect 7742 5108 7748 5120
rect 7800 5108 7806 5160
rect 7837 5151 7895 5157
rect 7837 5117 7849 5151
rect 7883 5148 7895 5151
rect 8021 5151 8079 5157
rect 8021 5148 8033 5151
rect 7883 5120 8033 5148
rect 7883 5117 7895 5120
rect 7837 5111 7895 5117
rect 8021 5117 8033 5120
rect 8067 5148 8079 5151
rect 8570 5148 8576 5160
rect 8067 5120 8576 5148
rect 8067 5117 8079 5120
rect 8021 5111 8079 5117
rect 2866 5080 2872 5092
rect 2608 5052 2872 5080
rect 2866 5040 2872 5052
rect 2924 5080 2930 5092
rect 3694 5080 3700 5092
rect 2924 5052 3700 5080
rect 2924 5040 2930 5052
rect 3694 5040 3700 5052
rect 3752 5040 3758 5092
rect 4065 5083 4123 5089
rect 4065 5049 4077 5083
rect 4111 5080 4123 5083
rect 4982 5080 4988 5092
rect 4111 5052 4988 5080
rect 4111 5049 4123 5052
rect 4065 5043 4123 5049
rect 4982 5040 4988 5052
rect 5040 5040 5046 5092
rect 5442 5040 5448 5092
rect 5500 5080 5506 5092
rect 6006 5083 6064 5089
rect 6006 5080 6018 5083
rect 5500 5052 6018 5080
rect 5500 5040 5506 5052
rect 6006 5049 6018 5052
rect 6052 5080 6064 5083
rect 6288 5080 6316 5108
rect 7374 5080 7380 5092
rect 6052 5052 6132 5080
rect 6288 5052 7380 5080
rect 6052 5049 6064 5052
rect 6006 5043 6064 5049
rect 6104 5024 6132 5052
rect 7374 5040 7380 5052
rect 7432 5080 7438 5092
rect 7852 5080 7880 5111
rect 8570 5108 8576 5120
rect 8628 5108 8634 5160
rect 9493 5151 9551 5157
rect 9493 5117 9505 5151
rect 9539 5117 9551 5151
rect 9600 5148 9628 5188
rect 10594 5176 10600 5228
rect 10652 5216 10658 5228
rect 13262 5216 13268 5228
rect 10652 5188 13268 5216
rect 10652 5176 10658 5188
rect 13262 5176 13268 5188
rect 13320 5176 13326 5228
rect 13998 5216 14004 5228
rect 13911 5188 14004 5216
rect 13998 5176 14004 5188
rect 14056 5216 14062 5228
rect 15933 5219 15991 5225
rect 14056 5188 15884 5216
rect 14056 5176 14062 5188
rect 9749 5151 9807 5157
rect 9749 5148 9761 5151
rect 9600 5120 9761 5148
rect 9493 5111 9551 5117
rect 9749 5117 9761 5120
rect 9795 5117 9807 5151
rect 10962 5148 10968 5160
rect 10923 5120 10968 5148
rect 9749 5111 9807 5117
rect 7432 5052 7880 5080
rect 8288 5083 8346 5089
rect 7432 5040 7438 5052
rect 8288 5049 8300 5083
rect 8334 5080 8346 5083
rect 8754 5080 8760 5092
rect 8334 5052 8760 5080
rect 8334 5049 8346 5052
rect 8288 5043 8346 5049
rect 8754 5040 8760 5052
rect 8812 5040 8818 5092
rect 9508 5080 9536 5111
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 12526 5108 12532 5160
rect 12584 5148 12590 5160
rect 12656 5151 12714 5157
rect 12656 5148 12668 5151
rect 12584 5120 12668 5148
rect 12584 5108 12590 5120
rect 12656 5117 12668 5120
rect 12702 5117 12714 5151
rect 13814 5148 13820 5160
rect 13775 5120 13820 5148
rect 12656 5111 12714 5117
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 14090 5108 14096 5160
rect 14148 5148 14154 5160
rect 14461 5151 14519 5157
rect 14461 5148 14473 5151
rect 14148 5120 14473 5148
rect 14148 5108 14154 5120
rect 14461 5117 14473 5120
rect 14507 5148 14519 5151
rect 14642 5148 14648 5160
rect 14507 5120 14648 5148
rect 14507 5117 14519 5120
rect 14461 5111 14519 5117
rect 14642 5108 14648 5120
rect 14700 5108 14706 5160
rect 15286 5108 15292 5160
rect 15344 5148 15350 5160
rect 15654 5148 15660 5160
rect 15344 5120 15660 5148
rect 15344 5108 15350 5120
rect 15654 5108 15660 5120
rect 15712 5108 15718 5160
rect 10778 5080 10784 5092
rect 9508 5052 10784 5080
rect 10778 5040 10784 5052
rect 10836 5040 10842 5092
rect 12437 5083 12495 5089
rect 12437 5080 12449 5083
rect 10980 5052 12449 5080
rect 1854 5012 1860 5024
rect 1815 4984 1860 5012
rect 1854 4972 1860 4984
rect 1912 4972 1918 5024
rect 2130 5012 2136 5024
rect 2091 4984 2136 5012
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 4154 4972 4160 5024
rect 4212 5012 4218 5024
rect 4212 4984 4257 5012
rect 4212 4972 4218 4984
rect 6086 4972 6092 5024
rect 6144 4972 6150 5024
rect 6178 4972 6184 5024
rect 6236 5012 6242 5024
rect 6457 5015 6515 5021
rect 6457 5012 6469 5015
rect 6236 4984 6469 5012
rect 6236 4972 6242 4984
rect 6457 4981 6469 4984
rect 6503 4981 6515 5015
rect 6457 4975 6515 4981
rect 6546 4972 6552 5024
rect 6604 5012 6610 5024
rect 8662 5012 8668 5024
rect 6604 4984 8668 5012
rect 6604 4972 6610 4984
rect 8662 4972 8668 4984
rect 8720 5012 8726 5024
rect 10980 5012 11008 5052
rect 12437 5049 12449 5052
rect 12483 5049 12495 5083
rect 12437 5043 12495 5049
rect 12611 5052 13860 5080
rect 8720 4984 11008 5012
rect 8720 4972 8726 4984
rect 11054 4972 11060 5024
rect 11112 5012 11118 5024
rect 11425 5015 11483 5021
rect 11425 5012 11437 5015
rect 11112 4984 11437 5012
rect 11112 4972 11118 4984
rect 11425 4981 11437 4984
rect 11471 5012 11483 5015
rect 12611 5012 12639 5052
rect 13832 5024 13860 5052
rect 15194 5040 15200 5092
rect 15252 5080 15258 5092
rect 15473 5083 15531 5089
rect 15473 5080 15485 5083
rect 15252 5052 15485 5080
rect 15252 5040 15258 5052
rect 15473 5049 15485 5052
rect 15519 5080 15531 5083
rect 15746 5080 15752 5092
rect 15519 5052 15752 5080
rect 15519 5049 15531 5052
rect 15473 5043 15531 5049
rect 15746 5040 15752 5052
rect 15804 5040 15810 5092
rect 15856 5080 15884 5188
rect 15933 5185 15945 5219
rect 15979 5216 15991 5219
rect 16298 5216 16304 5228
rect 15979 5188 16304 5216
rect 15979 5185 15991 5188
rect 15933 5179 15991 5185
rect 16298 5176 16304 5188
rect 16356 5176 16362 5228
rect 16482 5176 16488 5228
rect 16540 5216 16546 5228
rect 16577 5219 16635 5225
rect 16577 5216 16589 5219
rect 16540 5188 16589 5216
rect 16540 5176 16546 5188
rect 16577 5185 16589 5188
rect 16623 5185 16635 5219
rect 16577 5179 16635 5185
rect 17144 5160 17172 5324
rect 17218 5176 17224 5228
rect 17276 5216 17282 5228
rect 17497 5219 17555 5225
rect 17497 5216 17509 5219
rect 17276 5188 17509 5216
rect 17276 5176 17282 5188
rect 17497 5185 17509 5188
rect 17543 5185 17555 5219
rect 18506 5216 18512 5228
rect 18467 5188 18512 5216
rect 17497 5179 17555 5185
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 16393 5151 16451 5157
rect 16393 5117 16405 5151
rect 16439 5148 16451 5151
rect 16666 5148 16672 5160
rect 16439 5120 16672 5148
rect 16439 5117 16451 5120
rect 16393 5111 16451 5117
rect 16666 5108 16672 5120
rect 16724 5108 16730 5160
rect 17126 5148 17132 5160
rect 17039 5120 17132 5148
rect 17126 5108 17132 5120
rect 17184 5148 17190 5160
rect 17405 5151 17463 5157
rect 17405 5148 17417 5151
rect 17184 5120 17417 5148
rect 17184 5108 17190 5120
rect 17405 5117 17417 5120
rect 17451 5117 17463 5151
rect 17862 5148 17868 5160
rect 17823 5120 17868 5148
rect 17405 5111 17463 5117
rect 17862 5108 17868 5120
rect 17920 5108 17926 5160
rect 18325 5151 18383 5157
rect 18325 5117 18337 5151
rect 18371 5148 18383 5151
rect 18598 5148 18604 5160
rect 18371 5120 18604 5148
rect 18371 5117 18383 5120
rect 18325 5111 18383 5117
rect 18598 5108 18604 5120
rect 18656 5108 18662 5160
rect 16758 5080 16764 5092
rect 15856 5052 16764 5080
rect 16758 5040 16764 5052
rect 16816 5040 16822 5092
rect 16850 5040 16856 5092
rect 16908 5080 16914 5092
rect 17313 5083 17371 5089
rect 17313 5080 17325 5083
rect 16908 5052 17325 5080
rect 16908 5040 16914 5052
rect 17313 5049 17325 5052
rect 17359 5049 17371 5083
rect 17313 5043 17371 5049
rect 11471 4984 12639 5012
rect 11471 4981 11483 4984
rect 11425 4975 11483 4981
rect 12710 4972 12716 5024
rect 12768 5021 12774 5024
rect 12768 5015 12817 5021
rect 12768 4981 12771 5015
rect 12805 4981 12817 5015
rect 12768 4975 12817 4981
rect 12768 4972 12774 4975
rect 13814 4972 13820 5024
rect 13872 4972 13878 5024
rect 13998 4972 14004 5024
rect 14056 5012 14062 5024
rect 14093 5015 14151 5021
rect 14093 5012 14105 5015
rect 14056 4984 14105 5012
rect 14056 4972 14062 4984
rect 14093 4981 14105 4984
rect 14139 4981 14151 5015
rect 15102 5012 15108 5024
rect 15015 4984 15108 5012
rect 14093 4975 14151 4981
rect 15102 4972 15108 4984
rect 15160 5012 15166 5024
rect 16114 5012 16120 5024
rect 15160 4984 16120 5012
rect 15160 4972 15166 4984
rect 16114 4972 16120 4984
rect 16172 4972 16178 5024
rect 16485 5015 16543 5021
rect 16485 4981 16497 5015
rect 16531 5012 16543 5015
rect 16945 5015 17003 5021
rect 16945 5012 16957 5015
rect 16531 4984 16957 5012
rect 16531 4981 16543 4984
rect 16485 4975 16543 4981
rect 16945 4981 16957 4984
rect 16991 4981 17003 5015
rect 16945 4975 17003 4981
rect 18049 5015 18107 5021
rect 18049 4981 18061 5015
rect 18095 5012 18107 5015
rect 18230 5012 18236 5024
rect 18095 4984 18236 5012
rect 18095 4981 18107 4984
rect 18049 4975 18107 4981
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 1104 4922 18860 4944
rect 1104 4870 6912 4922
rect 6964 4870 6976 4922
rect 7028 4870 7040 4922
rect 7092 4870 7104 4922
rect 7156 4870 12843 4922
rect 12895 4870 12907 4922
rect 12959 4870 12971 4922
rect 13023 4870 13035 4922
rect 13087 4870 18860 4922
rect 1104 4848 18860 4870
rect 1946 4768 1952 4820
rect 2004 4808 2010 4820
rect 2317 4811 2375 4817
rect 2317 4808 2329 4811
rect 2004 4780 2329 4808
rect 2004 4768 2010 4780
rect 2317 4777 2329 4780
rect 2363 4777 2375 4811
rect 2866 4808 2872 4820
rect 2827 4780 2872 4808
rect 2317 4771 2375 4777
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 3786 4768 3792 4820
rect 3844 4808 3850 4820
rect 3973 4811 4031 4817
rect 3973 4808 3985 4811
rect 3844 4780 3985 4808
rect 3844 4768 3850 4780
rect 3973 4777 3985 4780
rect 4019 4777 4031 4811
rect 4154 4808 4160 4820
rect 4115 4780 4160 4808
rect 3973 4771 4031 4777
rect 4154 4768 4160 4780
rect 4212 4768 4218 4820
rect 4522 4808 4528 4820
rect 4483 4780 4528 4808
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 4982 4808 4988 4820
rect 4943 4780 4988 4808
rect 4982 4768 4988 4780
rect 5040 4768 5046 4820
rect 5074 4768 5080 4820
rect 5132 4808 5138 4820
rect 5353 4811 5411 4817
rect 5353 4808 5365 4811
rect 5132 4780 5365 4808
rect 5132 4768 5138 4780
rect 5353 4777 5365 4780
rect 5399 4808 5411 4811
rect 6641 4811 6699 4817
rect 6641 4808 6653 4811
rect 5399 4780 6653 4808
rect 5399 4777 5411 4780
rect 5353 4771 5411 4777
rect 6641 4777 6653 4780
rect 6687 4777 6699 4811
rect 6641 4771 6699 4777
rect 6917 4811 6975 4817
rect 6917 4777 6929 4811
rect 6963 4808 6975 4811
rect 9490 4808 9496 4820
rect 6963 4780 9496 4808
rect 6963 4777 6975 4780
rect 6917 4771 6975 4777
rect 1581 4743 1639 4749
rect 1581 4709 1593 4743
rect 1627 4740 1639 4743
rect 2130 4740 2136 4752
rect 1627 4712 2136 4740
rect 1627 4709 1639 4712
rect 1581 4703 1639 4709
rect 2130 4700 2136 4712
rect 2188 4700 2194 4752
rect 3053 4743 3111 4749
rect 3053 4740 3065 4743
rect 2516 4712 3065 4740
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 2516 4681 2544 4712
rect 3053 4709 3065 4712
rect 3099 4740 3111 4743
rect 6546 4740 6552 4752
rect 3099 4712 6552 4740
rect 3099 4709 3111 4712
rect 3053 4703 3111 4709
rect 6546 4700 6552 4712
rect 6604 4700 6610 4752
rect 2225 4675 2283 4681
rect 2225 4641 2237 4675
rect 2271 4641 2283 4675
rect 2225 4635 2283 4641
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4641 2559 4675
rect 2501 4635 2559 4641
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4573 2099 4607
rect 2240 4604 2268 4635
rect 3786 4632 3792 4684
rect 3844 4672 3850 4684
rect 4617 4675 4675 4681
rect 4617 4672 4629 4675
rect 3844 4644 4629 4672
rect 3844 4632 3850 4644
rect 4617 4641 4629 4644
rect 4663 4641 4675 4675
rect 4617 4635 4675 4641
rect 4706 4632 4712 4684
rect 4764 4672 4770 4684
rect 4764 4644 5028 4672
rect 4764 4632 4770 4644
rect 2593 4607 2651 4613
rect 2593 4604 2605 4607
rect 2240 4576 2605 4604
rect 2041 4567 2099 4573
rect 2593 4573 2605 4576
rect 2639 4604 2651 4607
rect 4801 4607 4859 4613
rect 2639 4576 4568 4604
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 2056 4468 2084 4567
rect 3142 4468 3148 4480
rect 2056 4440 3148 4468
rect 3142 4428 3148 4440
rect 3200 4428 3206 4480
rect 4540 4468 4568 4576
rect 4801 4573 4813 4607
rect 4847 4573 4859 4607
rect 5000 4604 5028 4644
rect 5994 4632 6000 4684
rect 6052 4672 6058 4684
rect 6181 4675 6239 4681
rect 6181 4672 6193 4675
rect 6052 4644 6193 4672
rect 6052 4632 6058 4644
rect 6181 4641 6193 4644
rect 6227 4672 6239 4675
rect 6932 4672 6960 4771
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 12526 4808 12532 4820
rect 9640 4780 12532 4808
rect 9640 4768 9646 4780
rect 10778 4700 10784 4752
rect 10836 4700 10842 4752
rect 11238 4700 11244 4752
rect 11296 4740 11302 4752
rect 11434 4743 11492 4749
rect 11434 4740 11446 4743
rect 11296 4712 11446 4740
rect 11296 4700 11302 4712
rect 11434 4709 11446 4712
rect 11480 4709 11492 4743
rect 11434 4703 11492 4709
rect 11606 4700 11612 4752
rect 11664 4740 11670 4752
rect 12268 4749 12296 4780
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 12710 4768 12716 4820
rect 12768 4808 12774 4820
rect 12768 4780 13308 4808
rect 12768 4768 12774 4780
rect 12161 4743 12219 4749
rect 12161 4740 12173 4743
rect 11664 4712 12173 4740
rect 11664 4700 11670 4712
rect 12161 4709 12173 4712
rect 12207 4709 12219 4743
rect 12161 4703 12219 4709
rect 12253 4743 12311 4749
rect 12253 4709 12265 4743
rect 12299 4709 12311 4743
rect 12253 4703 12311 4709
rect 12805 4743 12863 4749
rect 12805 4709 12817 4743
rect 12851 4740 12863 4743
rect 13170 4740 13176 4752
rect 12851 4712 13176 4740
rect 12851 4709 12863 4712
rect 12805 4703 12863 4709
rect 13170 4700 13176 4712
rect 13228 4700 13234 4752
rect 13280 4749 13308 4780
rect 13354 4768 13360 4820
rect 13412 4808 13418 4820
rect 13412 4780 16436 4808
rect 13412 4768 13418 4780
rect 13265 4743 13323 4749
rect 13265 4709 13277 4743
rect 13311 4709 13323 4743
rect 13265 4703 13323 4709
rect 14642 4700 14648 4752
rect 14700 4740 14706 4752
rect 15933 4743 15991 4749
rect 15933 4740 15945 4743
rect 14700 4712 15945 4740
rect 14700 4700 14706 4712
rect 6227 4644 6960 4672
rect 10796 4672 10824 4700
rect 11701 4675 11759 4681
rect 11701 4672 11713 4675
rect 10796 4644 11713 4672
rect 6227 4641 6239 4644
rect 6181 4635 6239 4641
rect 11701 4641 11713 4644
rect 11747 4641 11759 4675
rect 11701 4635 11759 4641
rect 5166 4604 5172 4616
rect 5000 4576 5172 4604
rect 4801 4567 4859 4573
rect 4816 4536 4844 4567
rect 5166 4564 5172 4576
rect 5224 4604 5230 4616
rect 5445 4607 5503 4613
rect 5445 4604 5457 4607
rect 5224 4576 5457 4604
rect 5224 4564 5230 4576
rect 5445 4573 5457 4576
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4573 5687 4607
rect 6270 4604 6276 4616
rect 6231 4576 6276 4604
rect 5629 4567 5687 4573
rect 5534 4536 5540 4548
rect 4816 4508 5540 4536
rect 5534 4496 5540 4508
rect 5592 4536 5598 4548
rect 5644 4536 5672 4567
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 6457 4607 6515 4613
rect 6457 4573 6469 4607
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 5810 4536 5816 4548
rect 5592 4508 5672 4536
rect 5771 4508 5816 4536
rect 5592 4496 5598 4508
rect 5810 4496 5816 4508
rect 5868 4496 5874 4548
rect 6086 4496 6092 4548
rect 6144 4536 6150 4548
rect 6472 4536 6500 4567
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 10594 4604 10600 4616
rect 6604 4576 10600 4604
rect 6604 4564 6610 4576
rect 10594 4564 10600 4576
rect 10652 4564 10658 4616
rect 11716 4604 11744 4635
rect 13814 4632 13820 4684
rect 13872 4672 13878 4684
rect 14036 4675 14094 4681
rect 14036 4672 14048 4675
rect 13872 4644 14048 4672
rect 13872 4632 13878 4644
rect 14036 4641 14048 4644
rect 14082 4641 14094 4675
rect 14036 4635 14094 4641
rect 14369 4675 14427 4681
rect 14369 4641 14381 4675
rect 14415 4672 14427 4675
rect 14458 4672 14464 4684
rect 14415 4644 14464 4672
rect 14415 4641 14427 4644
rect 14369 4635 14427 4641
rect 12434 4604 12440 4616
rect 11716 4576 12440 4604
rect 7558 4536 7564 4548
rect 6144 4508 6500 4536
rect 6564 4508 7564 4536
rect 6144 4496 6150 4508
rect 6564 4468 6592 4508
rect 7558 4496 7564 4508
rect 7616 4496 7622 4548
rect 4540 4440 6592 4468
rect 10321 4471 10379 4477
rect 10321 4437 10333 4471
rect 10367 4468 10379 4471
rect 10410 4468 10416 4480
rect 10367 4440 10416 4468
rect 10367 4437 10379 4440
rect 10321 4431 10379 4437
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 10778 4428 10784 4480
rect 10836 4468 10842 4480
rect 10962 4468 10968 4480
rect 10836 4440 10968 4468
rect 10836 4428 10842 4440
rect 10962 4428 10968 4440
rect 11020 4428 11026 4480
rect 11514 4428 11520 4480
rect 11572 4468 11578 4480
rect 11716 4468 11744 4576
rect 12434 4564 12440 4576
rect 12492 4564 12498 4616
rect 13173 4607 13231 4613
rect 13173 4573 13185 4607
rect 13219 4573 13231 4607
rect 13538 4604 13544 4616
rect 13499 4576 13544 4604
rect 13173 4567 13231 4573
rect 13188 4536 13216 4567
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 14051 4604 14079 4635
rect 14458 4632 14464 4644
rect 14516 4632 14522 4684
rect 15102 4632 15108 4684
rect 15160 4672 15166 4684
rect 15580 4681 15608 4712
rect 15933 4709 15945 4712
rect 15979 4709 15991 4743
rect 15933 4703 15991 4709
rect 15222 4675 15280 4681
rect 15222 4672 15234 4675
rect 15160 4644 15234 4672
rect 15160 4632 15166 4644
rect 15222 4641 15234 4644
rect 15268 4641 15280 4675
rect 15222 4635 15280 4641
rect 15565 4675 15623 4681
rect 15565 4641 15577 4675
rect 15611 4641 15623 4675
rect 15565 4635 15623 4641
rect 15746 4632 15752 4684
rect 15804 4672 15810 4684
rect 15841 4675 15899 4681
rect 15841 4672 15853 4675
rect 15804 4644 15853 4672
rect 15804 4632 15810 4644
rect 15841 4641 15853 4644
rect 15887 4641 15899 4675
rect 15841 4635 15899 4641
rect 16117 4675 16175 4681
rect 16117 4641 16129 4675
rect 16163 4641 16175 4675
rect 16117 4635 16175 4641
rect 14553 4607 14611 4613
rect 14553 4604 14565 4607
rect 14051 4576 14565 4604
rect 14553 4573 14565 4576
rect 14599 4573 14611 4607
rect 14553 4567 14611 4573
rect 15013 4607 15071 4613
rect 15013 4573 15025 4607
rect 15059 4604 15071 4607
rect 16132 4604 16160 4635
rect 16298 4632 16304 4684
rect 16356 4632 16362 4684
rect 16408 4681 16436 4780
rect 16574 4768 16580 4820
rect 16632 4808 16638 4820
rect 16669 4811 16727 4817
rect 16669 4808 16681 4811
rect 16632 4780 16681 4808
rect 16632 4768 16638 4780
rect 16669 4777 16681 4780
rect 16715 4777 16727 4811
rect 17034 4808 17040 4820
rect 16947 4780 17040 4808
rect 16669 4771 16727 4777
rect 17034 4768 17040 4780
rect 17092 4808 17098 4820
rect 18782 4808 18788 4820
rect 17092 4780 18788 4808
rect 17092 4768 17098 4780
rect 18782 4768 18788 4780
rect 18840 4768 18846 4820
rect 16482 4700 16488 4752
rect 16540 4740 16546 4752
rect 17310 4740 17316 4752
rect 16540 4712 17316 4740
rect 16540 4700 16546 4712
rect 17310 4700 17316 4712
rect 17368 4700 17374 4752
rect 17954 4740 17960 4752
rect 17915 4712 17960 4740
rect 17954 4700 17960 4712
rect 18012 4700 18018 4752
rect 18046 4700 18052 4752
rect 18104 4740 18110 4752
rect 18325 4743 18383 4749
rect 18325 4740 18337 4743
rect 18104 4712 18337 4740
rect 18104 4700 18110 4712
rect 18325 4709 18337 4712
rect 18371 4709 18383 4743
rect 18325 4703 18383 4709
rect 16393 4675 16451 4681
rect 16393 4641 16405 4675
rect 16439 4641 16451 4675
rect 16393 4635 16451 4641
rect 16942 4632 16948 4684
rect 17000 4672 17006 4684
rect 17589 4675 17647 4681
rect 17589 4672 17601 4675
rect 17000 4644 17601 4672
rect 17000 4632 17006 4644
rect 17589 4641 17601 4644
rect 17635 4641 17647 4675
rect 18138 4672 18144 4684
rect 18099 4644 18144 4672
rect 17589 4635 17647 4641
rect 18138 4632 18144 4644
rect 18196 4632 18202 4684
rect 16316 4604 16344 4632
rect 17129 4607 17187 4613
rect 17129 4604 17141 4607
rect 15059 4576 16160 4604
rect 16224 4576 17141 4604
rect 15059 4573 15071 4576
rect 15013 4567 15071 4573
rect 13906 4536 13912 4548
rect 13188 4508 13912 4536
rect 13906 4496 13912 4508
rect 13964 4496 13970 4548
rect 15286 4496 15292 4548
rect 15344 4536 15350 4548
rect 15657 4539 15715 4545
rect 15657 4536 15669 4539
rect 15344 4508 15669 4536
rect 15344 4496 15350 4508
rect 15657 4505 15669 4508
rect 15703 4505 15715 4539
rect 15657 4499 15715 4505
rect 15746 4496 15752 4548
rect 15804 4536 15810 4548
rect 16224 4536 16252 4576
rect 17129 4573 17141 4576
rect 17175 4573 17187 4607
rect 17129 4567 17187 4573
rect 17218 4564 17224 4616
rect 17276 4604 17282 4616
rect 17276 4576 17321 4604
rect 17276 4564 17282 4576
rect 15804 4508 16252 4536
rect 16301 4539 16359 4545
rect 15804 4496 15810 4508
rect 16301 4505 16313 4539
rect 16347 4536 16359 4539
rect 17034 4536 17040 4548
rect 16347 4508 17040 4536
rect 16347 4505 16359 4508
rect 16301 4499 16359 4505
rect 17034 4496 17040 4508
rect 17092 4496 17098 4548
rect 18506 4536 18512 4548
rect 18467 4508 18512 4536
rect 18506 4496 18512 4508
rect 18564 4496 18570 4548
rect 11572 4440 11744 4468
rect 11572 4428 11578 4440
rect 11882 4428 11888 4480
rect 11940 4468 11946 4480
rect 12989 4471 13047 4477
rect 12989 4468 13001 4471
rect 11940 4440 13001 4468
rect 11940 4428 11946 4440
rect 12989 4437 13001 4440
rect 13035 4468 13047 4471
rect 13446 4468 13452 4480
rect 13035 4440 13452 4468
rect 13035 4437 13047 4440
rect 12989 4431 13047 4437
rect 13446 4428 13452 4440
rect 13504 4428 13510 4480
rect 14139 4471 14197 4477
rect 14139 4437 14151 4471
rect 14185 4468 14197 4471
rect 14274 4468 14280 4480
rect 14185 4440 14280 4468
rect 14185 4437 14197 4440
rect 14139 4431 14197 4437
rect 14274 4428 14280 4440
rect 14332 4428 14338 4480
rect 15194 4477 15200 4480
rect 15151 4471 15200 4477
rect 15151 4437 15163 4471
rect 15197 4437 15200 4471
rect 15151 4431 15200 4437
rect 15194 4428 15200 4431
rect 15252 4428 15258 4480
rect 15378 4468 15384 4480
rect 15339 4440 15384 4468
rect 15378 4428 15384 4440
rect 15436 4428 15442 4480
rect 16574 4468 16580 4480
rect 16535 4440 16580 4468
rect 16574 4428 16580 4440
rect 16632 4428 16638 4480
rect 17773 4471 17831 4477
rect 17773 4437 17785 4471
rect 17819 4468 17831 4471
rect 17954 4468 17960 4480
rect 17819 4440 17960 4468
rect 17819 4437 17831 4440
rect 17773 4431 17831 4437
rect 17954 4428 17960 4440
rect 18012 4428 18018 4480
rect 1104 4378 18860 4400
rect 1104 4326 3947 4378
rect 3999 4326 4011 4378
rect 4063 4326 4075 4378
rect 4127 4326 4139 4378
rect 4191 4326 9878 4378
rect 9930 4326 9942 4378
rect 9994 4326 10006 4378
rect 10058 4326 10070 4378
rect 10122 4326 15808 4378
rect 15860 4326 15872 4378
rect 15924 4326 15936 4378
rect 15988 4326 16000 4378
rect 16052 4326 18860 4378
rect 1104 4304 18860 4326
rect 2682 4224 2688 4276
rect 2740 4264 2746 4276
rect 3329 4267 3387 4273
rect 3329 4264 3341 4267
rect 2740 4236 3341 4264
rect 2740 4224 2746 4236
rect 3329 4233 3341 4236
rect 3375 4264 3387 4267
rect 3602 4264 3608 4276
rect 3375 4236 3608 4264
rect 3375 4233 3387 4236
rect 3329 4227 3387 4233
rect 3602 4224 3608 4236
rect 3660 4224 3666 4276
rect 4522 4264 4528 4276
rect 3896 4236 4528 4264
rect 3145 4199 3203 4205
rect 3145 4165 3157 4199
rect 3191 4196 3203 4199
rect 3896 4196 3924 4236
rect 4522 4224 4528 4236
rect 4580 4264 4586 4276
rect 5261 4267 5319 4273
rect 4580 4236 5120 4264
rect 4580 4224 4586 4236
rect 3191 4168 3924 4196
rect 3191 4165 3203 4168
rect 3145 4159 3203 4165
rect 1581 4063 1639 4069
rect 1581 4029 1593 4063
rect 1627 4060 1639 4063
rect 2498 4060 2504 4072
rect 1627 4032 2504 4060
rect 1627 4029 1639 4032
rect 1581 4023 1639 4029
rect 2498 4020 2504 4032
rect 2556 4020 2562 4072
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4029 2743 4063
rect 2685 4023 2743 4029
rect 2961 4063 3019 4069
rect 2961 4029 2973 4063
rect 3007 4060 3019 4063
rect 3160 4060 3188 4159
rect 5092 4128 5120 4236
rect 5261 4233 5273 4267
rect 5307 4264 5319 4267
rect 5442 4264 5448 4276
rect 5307 4236 5448 4264
rect 5307 4233 5319 4236
rect 5261 4227 5319 4233
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 5721 4267 5779 4273
rect 5721 4233 5733 4267
rect 5767 4264 5779 4267
rect 6270 4264 6276 4276
rect 5767 4236 6276 4264
rect 5767 4233 5779 4236
rect 5721 4227 5779 4233
rect 6270 4224 6276 4236
rect 6328 4224 6334 4276
rect 6546 4224 6552 4276
rect 6604 4264 6610 4276
rect 6733 4267 6791 4273
rect 6733 4264 6745 4267
rect 6604 4236 6745 4264
rect 6604 4224 6610 4236
rect 6733 4233 6745 4236
rect 6779 4233 6791 4267
rect 8754 4264 8760 4276
rect 8715 4236 8760 4264
rect 6733 4227 6791 4233
rect 8754 4224 8760 4236
rect 8812 4264 8818 4276
rect 8941 4267 8999 4273
rect 8941 4264 8953 4267
rect 8812 4236 8953 4264
rect 8812 4224 8818 4236
rect 8941 4233 8953 4236
rect 8987 4233 8999 4267
rect 8941 4227 8999 4233
rect 9677 4267 9735 4273
rect 9677 4233 9689 4267
rect 9723 4264 9735 4267
rect 10594 4264 10600 4276
rect 9723 4236 10600 4264
rect 9723 4233 9735 4236
rect 9677 4227 9735 4233
rect 10594 4224 10600 4236
rect 10652 4224 10658 4276
rect 11146 4224 11152 4276
rect 11204 4264 11210 4276
rect 11204 4236 11560 4264
rect 11204 4224 11210 4236
rect 5166 4156 5172 4208
rect 5224 4196 5230 4208
rect 5353 4199 5411 4205
rect 5353 4196 5365 4199
rect 5224 4168 5365 4196
rect 5224 4156 5230 4168
rect 5353 4165 5365 4168
rect 5399 4165 5411 4199
rect 5353 4159 5411 4165
rect 5813 4131 5871 4137
rect 5813 4128 5825 4131
rect 5092 4100 5825 4128
rect 5813 4097 5825 4100
rect 5859 4097 5871 4131
rect 7374 4128 7380 4140
rect 7335 4100 7380 4128
rect 5813 4091 5871 4097
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4128 9367 4131
rect 9398 4128 9404 4140
rect 9355 4100 9404 4128
rect 9355 4097 9367 4100
rect 9309 4091 9367 4097
rect 9398 4088 9404 4100
rect 9456 4128 9462 4140
rect 11532 4128 11560 4236
rect 12342 4224 12348 4276
rect 12400 4264 12406 4276
rect 15102 4264 15108 4276
rect 12400 4236 15108 4264
rect 12400 4224 12406 4236
rect 15102 4224 15108 4236
rect 15160 4264 15166 4276
rect 15160 4236 15884 4264
rect 15160 4224 15166 4236
rect 15562 4196 15568 4208
rect 15523 4168 15568 4196
rect 15562 4156 15568 4168
rect 15620 4156 15626 4208
rect 15856 4196 15884 4236
rect 16114 4224 16120 4276
rect 16172 4264 16178 4276
rect 16942 4264 16948 4276
rect 16172 4236 16948 4264
rect 16172 4224 16178 4236
rect 16942 4224 16948 4236
rect 17000 4224 17006 4276
rect 15930 4196 15936 4208
rect 15856 4168 15936 4196
rect 15930 4156 15936 4168
rect 15988 4156 15994 4208
rect 17405 4199 17463 4205
rect 17405 4165 17417 4199
rect 17451 4165 17463 4199
rect 17405 4159 17463 4165
rect 9456 4100 10548 4128
rect 11532 4100 11652 4128
rect 9456 4088 9462 4100
rect 3007 4032 3188 4060
rect 3881 4063 3939 4069
rect 3007 4029 3019 4032
rect 2961 4023 3019 4029
rect 3881 4029 3893 4063
rect 3927 4060 3939 4063
rect 5166 4060 5172 4072
rect 3927 4032 5172 4060
rect 3927 4029 3939 4032
rect 3881 4023 3939 4029
rect 1946 3992 1952 4004
rect 1907 3964 1952 3992
rect 1946 3952 1952 3964
rect 2004 3952 2010 4004
rect 2317 3995 2375 4001
rect 2317 3961 2329 3995
rect 2363 3961 2375 3995
rect 2700 3992 2728 4023
rect 5166 4020 5172 4032
rect 5224 4020 5230 4072
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4060 6699 4063
rect 6730 4060 6736 4072
rect 6687 4032 6736 4060
rect 6687 4029 6699 4032
rect 6641 4023 6699 4029
rect 6730 4020 6736 4032
rect 6788 4020 6794 4072
rect 8846 4060 8852 4072
rect 7484 4032 8156 4060
rect 8807 4032 8852 4060
rect 4148 3995 4206 4001
rect 2700 3964 3556 3992
rect 2317 3955 2375 3961
rect 1486 3924 1492 3936
rect 1447 3896 1492 3924
rect 1486 3884 1492 3896
rect 1544 3884 1550 3936
rect 1854 3924 1860 3936
rect 1815 3896 1860 3924
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 2222 3924 2228 3936
rect 2183 3896 2228 3924
rect 2222 3884 2228 3896
rect 2280 3884 2286 3936
rect 2332 3924 2360 3955
rect 2501 3927 2559 3933
rect 2501 3924 2513 3927
rect 2332 3896 2513 3924
rect 2501 3893 2513 3896
rect 2547 3893 2559 3927
rect 2501 3887 2559 3893
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 3528 3933 3556 3964
rect 4148 3961 4160 3995
rect 4194 3992 4206 3995
rect 4614 3992 4620 4004
rect 4194 3964 4620 3992
rect 4194 3961 4206 3964
rect 4148 3955 4206 3961
rect 4614 3952 4620 3964
rect 4672 3952 4678 4004
rect 7484 3992 7512 4032
rect 4724 3964 7512 3992
rect 7644 3995 7702 4001
rect 3513 3927 3571 3933
rect 2832 3896 2877 3924
rect 2832 3884 2838 3896
rect 3513 3893 3525 3927
rect 3559 3924 3571 3927
rect 3602 3924 3608 3936
rect 3559 3896 3608 3924
rect 3559 3893 3571 3896
rect 3513 3887 3571 3893
rect 3602 3884 3608 3896
rect 3660 3884 3666 3936
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 4724 3924 4752 3964
rect 7644 3961 7656 3995
rect 7690 3992 7702 3995
rect 8018 3992 8024 4004
rect 7690 3964 8024 3992
rect 7690 3961 7702 3964
rect 7644 3955 7702 3961
rect 8018 3952 8024 3964
rect 8076 3952 8082 4004
rect 8128 3992 8156 4032
rect 8846 4020 8852 4032
rect 8904 4020 8910 4072
rect 9490 4060 9496 4072
rect 9451 4032 9496 4060
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 10318 4060 10324 4072
rect 9600 4032 10324 4060
rect 9600 3992 9628 4032
rect 10318 4020 10324 4032
rect 10376 4020 10382 4072
rect 10520 4060 10548 4100
rect 11514 4060 11520 4072
rect 10520 4032 11376 4060
rect 11475 4032 11520 4060
rect 8128 3964 9628 3992
rect 10410 3952 10416 4004
rect 10468 3992 10474 4004
rect 11250 3995 11308 4001
rect 11250 3992 11262 3995
rect 10468 3964 11262 3992
rect 10468 3952 10474 3964
rect 11250 3961 11262 3964
rect 11296 3961 11308 3995
rect 11348 3992 11376 4032
rect 11514 4020 11520 4032
rect 11572 4020 11578 4072
rect 11624 4060 11652 4100
rect 11698 4088 11704 4140
rect 11756 4128 11762 4140
rect 12345 4131 12403 4137
rect 12345 4128 12357 4131
rect 11756 4100 12357 4128
rect 11756 4088 11762 4100
rect 12345 4097 12357 4100
rect 12391 4097 12403 4131
rect 12345 4091 12403 4097
rect 12710 4088 12716 4140
rect 12768 4128 12774 4140
rect 14826 4128 14832 4140
rect 12768 4100 13308 4128
rect 14787 4100 14832 4128
rect 12768 4088 12774 4100
rect 11974 4060 11980 4072
rect 11624 4032 11980 4060
rect 11974 4020 11980 4032
rect 12032 4020 12038 4072
rect 13280 4069 13308 4100
rect 14826 4088 14832 4100
rect 14884 4088 14890 4140
rect 15013 4131 15071 4137
rect 15013 4097 15025 4131
rect 15059 4128 15071 4131
rect 15378 4128 15384 4140
rect 15059 4100 15384 4128
rect 15059 4097 15071 4100
rect 15013 4091 15071 4097
rect 15378 4088 15384 4100
rect 15436 4088 15442 4140
rect 15654 4088 15660 4140
rect 15712 4128 15718 4140
rect 17310 4128 17316 4140
rect 15712 4100 17316 4128
rect 15712 4088 15718 4100
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 17420 4128 17448 4159
rect 18046 4128 18052 4140
rect 17420 4100 18052 4128
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4060 13323 4063
rect 13541 4063 13599 4069
rect 13541 4060 13553 4063
rect 13311 4032 13553 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 13541 4029 13553 4032
rect 13587 4029 13599 4063
rect 13541 4023 13599 4029
rect 13817 4063 13875 4069
rect 13817 4029 13829 4063
rect 13863 4060 13875 4063
rect 13998 4060 14004 4072
rect 13863 4032 14004 4060
rect 13863 4029 13875 4032
rect 13817 4023 13875 4029
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 15746 4060 15752 4072
rect 15707 4032 15752 4060
rect 15746 4020 15752 4032
rect 15804 4020 15810 4072
rect 15930 4060 15936 4072
rect 15891 4032 15936 4060
rect 15930 4020 15936 4032
rect 15988 4020 15994 4072
rect 16577 4063 16635 4069
rect 16577 4029 16589 4063
rect 16623 4060 16635 4063
rect 16758 4060 16764 4072
rect 16623 4032 16764 4060
rect 16623 4029 16635 4032
rect 16577 4023 16635 4029
rect 16758 4020 16764 4032
rect 16816 4020 16822 4072
rect 16942 4060 16948 4072
rect 16903 4032 16948 4060
rect 16942 4020 16948 4032
rect 17000 4020 17006 4072
rect 17126 4020 17132 4072
rect 17184 4060 17190 4072
rect 17221 4063 17279 4069
rect 17221 4060 17233 4063
rect 17184 4032 17233 4060
rect 17184 4020 17190 4032
rect 17221 4029 17233 4032
rect 17267 4029 17279 4063
rect 17957 4063 18015 4069
rect 17957 4060 17969 4063
rect 17221 4023 17279 4029
rect 17420 4032 17969 4060
rect 12434 3992 12440 4004
rect 11348 3964 12440 3992
rect 11250 3955 11308 3961
rect 12434 3952 12440 3964
rect 12492 3952 12498 4004
rect 12989 3995 13047 4001
rect 12989 3961 13001 3995
rect 13035 3992 13047 3995
rect 13630 3992 13636 4004
rect 13035 3964 13636 3992
rect 13035 3961 13047 3964
rect 12989 3955 13047 3961
rect 13630 3952 13636 3964
rect 13688 3952 13694 4004
rect 14185 3995 14243 4001
rect 14185 3961 14197 3995
rect 14231 3961 14243 3995
rect 14185 3955 14243 3961
rect 3844 3896 4752 3924
rect 3844 3884 3850 3896
rect 4798 3884 4804 3936
rect 4856 3924 4862 3936
rect 5994 3924 6000 3936
rect 4856 3896 6000 3924
rect 4856 3884 4862 3896
rect 5994 3884 6000 3896
rect 6052 3884 6058 3936
rect 7101 3927 7159 3933
rect 7101 3893 7113 3927
rect 7147 3924 7159 3927
rect 7742 3924 7748 3936
rect 7147 3896 7748 3924
rect 7147 3893 7159 3896
rect 7101 3887 7159 3893
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 8110 3884 8116 3936
rect 8168 3924 8174 3936
rect 10137 3927 10195 3933
rect 10137 3924 10149 3927
rect 8168 3896 10149 3924
rect 8168 3884 8174 3896
rect 10137 3893 10149 3896
rect 10183 3924 10195 3927
rect 10226 3924 10232 3936
rect 10183 3896 10232 3924
rect 10183 3893 10195 3896
rect 10137 3887 10195 3893
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 10594 3884 10600 3936
rect 10652 3924 10658 3936
rect 11330 3924 11336 3936
rect 10652 3896 11336 3924
rect 10652 3884 10658 3896
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 11606 3884 11612 3936
rect 11664 3924 11670 3936
rect 11701 3927 11759 3933
rect 11701 3924 11713 3927
rect 11664 3896 11713 3924
rect 11664 3884 11670 3896
rect 11701 3893 11713 3896
rect 11747 3893 11759 3927
rect 11882 3924 11888 3936
rect 11843 3896 11888 3924
rect 11701 3887 11759 3893
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 13081 3927 13139 3933
rect 13081 3893 13093 3927
rect 13127 3924 13139 3927
rect 13170 3924 13176 3936
rect 13127 3896 13176 3924
rect 13127 3893 13139 3896
rect 13081 3887 13139 3893
rect 13170 3884 13176 3896
rect 13228 3884 13234 3936
rect 13354 3924 13360 3936
rect 13315 3896 13360 3924
rect 13354 3884 13360 3896
rect 13412 3884 13418 3936
rect 14001 3927 14059 3933
rect 14001 3893 14013 3927
rect 14047 3924 14059 3927
rect 14200 3924 14228 3955
rect 14274 3952 14280 4004
rect 14332 3992 14338 4004
rect 15105 3995 15163 4001
rect 14332 3964 14377 3992
rect 14332 3952 14338 3964
rect 15105 3961 15117 3995
rect 15151 3992 15163 3995
rect 15194 3992 15200 4004
rect 15151 3964 15200 3992
rect 15151 3961 15163 3964
rect 15105 3955 15163 3961
rect 15194 3952 15200 3964
rect 15252 3952 15258 4004
rect 17420 3992 17448 4032
rect 17957 4029 17969 4032
rect 18003 4029 18015 4063
rect 17957 4023 18015 4029
rect 18230 4020 18236 4072
rect 18288 4060 18294 4072
rect 18325 4063 18383 4069
rect 18325 4060 18337 4063
rect 18288 4032 18337 4060
rect 18288 4020 18294 4032
rect 18325 4029 18337 4032
rect 18371 4029 18383 4063
rect 18325 4023 18383 4029
rect 16776 3964 17448 3992
rect 17589 3995 17647 4001
rect 14047 3896 14228 3924
rect 14047 3893 14059 3896
rect 14001 3887 14059 3893
rect 15010 3884 15016 3936
rect 15068 3924 15074 3936
rect 16776 3933 16804 3964
rect 17589 3961 17601 3995
rect 17635 3961 17647 3995
rect 18138 3992 18144 4004
rect 18099 3964 18144 3992
rect 17589 3955 17647 3961
rect 16393 3927 16451 3933
rect 16393 3924 16405 3927
rect 15068 3896 16405 3924
rect 15068 3884 15074 3896
rect 16393 3893 16405 3896
rect 16439 3893 16451 3927
rect 16393 3887 16451 3893
rect 16761 3927 16819 3933
rect 16761 3893 16773 3927
rect 16807 3893 16819 3927
rect 17126 3924 17132 3936
rect 17087 3896 17132 3924
rect 16761 3887 16819 3893
rect 17126 3884 17132 3896
rect 17184 3884 17190 3936
rect 17310 3884 17316 3936
rect 17368 3924 17374 3936
rect 17604 3924 17632 3955
rect 18138 3952 18144 3964
rect 18196 3952 18202 4004
rect 18506 3992 18512 4004
rect 18467 3964 18512 3992
rect 18506 3952 18512 3964
rect 18564 3952 18570 4004
rect 17368 3896 17632 3924
rect 17681 3927 17739 3933
rect 17368 3884 17374 3896
rect 17681 3893 17693 3927
rect 17727 3924 17739 3927
rect 19150 3924 19156 3936
rect 17727 3896 19156 3924
rect 17727 3893 17739 3896
rect 17681 3887 17739 3893
rect 19150 3884 19156 3896
rect 19208 3884 19214 3936
rect 1104 3834 18860 3856
rect 1104 3782 6912 3834
rect 6964 3782 6976 3834
rect 7028 3782 7040 3834
rect 7092 3782 7104 3834
rect 7156 3782 12843 3834
rect 12895 3782 12907 3834
rect 12959 3782 12971 3834
rect 13023 3782 13035 3834
rect 13087 3782 18860 3834
rect 1104 3760 18860 3782
rect 1946 3680 1952 3732
rect 2004 3720 2010 3732
rect 2501 3723 2559 3729
rect 2501 3720 2513 3723
rect 2004 3692 2513 3720
rect 2004 3680 2010 3692
rect 2501 3689 2513 3692
rect 2547 3689 2559 3723
rect 2501 3683 2559 3689
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3689 2835 3723
rect 2777 3683 2835 3689
rect 2317 3655 2375 3661
rect 2317 3621 2329 3655
rect 2363 3652 2375 3655
rect 2792 3652 2820 3683
rect 3602 3680 3608 3732
rect 3660 3720 3666 3732
rect 8018 3720 8024 3732
rect 3660 3692 7604 3720
rect 7979 3692 8024 3720
rect 3660 3680 3666 3692
rect 2363 3624 2820 3652
rect 3068 3624 6316 3652
rect 2363 3621 2375 3624
rect 2317 3615 2375 3621
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3553 1639 3587
rect 1946 3584 1952 3596
rect 1907 3556 1952 3584
rect 1581 3547 1639 3553
rect 1596 3516 1624 3547
rect 1946 3544 1952 3556
rect 2004 3544 2010 3596
rect 2682 3584 2688 3596
rect 2643 3556 2688 3584
rect 2682 3544 2688 3556
rect 2740 3544 2746 3596
rect 3068 3593 3096 3624
rect 2961 3587 3019 3593
rect 2961 3553 2973 3587
rect 3007 3553 3019 3587
rect 2961 3547 3019 3553
rect 3053 3587 3111 3593
rect 3053 3553 3065 3587
rect 3099 3553 3111 3587
rect 3053 3547 3111 3553
rect 2866 3516 2872 3528
rect 1596 3488 2872 3516
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 2976 3516 3004 3547
rect 3142 3544 3148 3596
rect 3200 3584 3206 3596
rect 3513 3587 3571 3593
rect 3513 3584 3525 3587
rect 3200 3556 3525 3584
rect 3200 3544 3206 3556
rect 3513 3553 3525 3556
rect 3559 3553 3571 3587
rect 3513 3547 3571 3553
rect 3973 3587 4031 3593
rect 3973 3553 3985 3587
rect 4019 3584 4031 3587
rect 5258 3584 5264 3596
rect 4019 3556 5264 3584
rect 4019 3553 4031 3556
rect 3973 3547 4031 3553
rect 3988 3516 4016 3547
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 5436 3587 5494 3593
rect 5436 3553 5448 3587
rect 5482 3584 5494 3587
rect 6178 3584 6184 3596
rect 5482 3556 6184 3584
rect 5482 3553 5494 3556
rect 5436 3547 5494 3553
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 6288 3584 6316 3624
rect 6546 3612 6552 3664
rect 6604 3652 6610 3664
rect 6886 3655 6944 3661
rect 6886 3652 6898 3655
rect 6604 3624 6898 3652
rect 6604 3612 6610 3624
rect 6886 3621 6898 3624
rect 6932 3621 6944 3655
rect 6886 3615 6944 3621
rect 7466 3584 7472 3596
rect 6288 3556 7472 3584
rect 7466 3544 7472 3556
rect 7524 3544 7530 3596
rect 7576 3584 7604 3692
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 10229 3723 10287 3729
rect 10229 3720 10241 3723
rect 8904 3692 10241 3720
rect 8904 3680 8910 3692
rect 10229 3689 10241 3692
rect 10275 3689 10287 3723
rect 10229 3683 10287 3689
rect 10781 3723 10839 3729
rect 10781 3689 10793 3723
rect 10827 3689 10839 3723
rect 13449 3723 13507 3729
rect 13449 3720 13461 3723
rect 10781 3683 10839 3689
rect 13004 3692 13461 3720
rect 7926 3612 7932 3664
rect 7984 3652 7990 3664
rect 10594 3652 10600 3664
rect 7984 3624 8432 3652
rect 7984 3612 7990 3624
rect 8202 3584 8208 3596
rect 7576 3556 8208 3584
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 8297 3587 8355 3593
rect 8297 3553 8309 3587
rect 8343 3553 8355 3587
rect 8404 3584 8432 3624
rect 9048 3624 10600 3652
rect 8516 3587 8574 3593
rect 8516 3584 8528 3587
rect 8404 3556 8528 3584
rect 8297 3547 8355 3553
rect 8516 3553 8528 3556
rect 8562 3553 8574 3587
rect 8516 3547 8574 3553
rect 5166 3516 5172 3528
rect 2976 3488 4016 3516
rect 5079 3488 5172 3516
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 6641 3519 6699 3525
rect 6641 3485 6653 3519
rect 6687 3485 6699 3519
rect 6641 3479 6699 3485
rect 3237 3451 3295 3457
rect 3237 3417 3249 3451
rect 3283 3448 3295 3451
rect 4982 3448 4988 3460
rect 3283 3420 4988 3448
rect 3283 3417 3295 3420
rect 3237 3411 3295 3417
rect 4982 3408 4988 3420
rect 5040 3408 5046 3460
rect 1394 3340 1400 3392
rect 1452 3380 1458 3392
rect 1489 3383 1547 3389
rect 1489 3380 1501 3383
rect 1452 3352 1501 3380
rect 1452 3340 1458 3352
rect 1489 3349 1501 3352
rect 1535 3349 1547 3383
rect 1854 3380 1860 3392
rect 1815 3352 1860 3380
rect 1489 3343 1547 3349
rect 1854 3340 1860 3352
rect 1912 3340 1918 3392
rect 2222 3380 2228 3392
rect 2183 3352 2228 3380
rect 2222 3340 2228 3352
rect 2280 3340 2286 3392
rect 3326 3340 3332 3392
rect 3384 3380 3390 3392
rect 3694 3380 3700 3392
rect 3384 3352 3429 3380
rect 3607 3352 3700 3380
rect 3384 3340 3390 3352
rect 3694 3340 3700 3352
rect 3752 3380 3758 3392
rect 4798 3380 4804 3392
rect 3752 3352 4804 3380
rect 3752 3340 3758 3352
rect 4798 3340 4804 3352
rect 4856 3340 4862 3392
rect 5184 3380 5212 3476
rect 6546 3448 6552 3460
rect 6507 3420 6552 3448
rect 6546 3408 6552 3420
rect 6604 3408 6610 3460
rect 6656 3380 6684 3479
rect 7834 3476 7840 3528
rect 7892 3516 7898 3528
rect 8312 3516 8340 3547
rect 9048 3516 9076 3624
rect 10594 3612 10600 3624
rect 10652 3612 10658 3664
rect 10796 3652 10824 3683
rect 12342 3652 12348 3664
rect 10796 3624 12348 3652
rect 10045 3587 10103 3593
rect 10045 3553 10057 3587
rect 10091 3553 10103 3587
rect 10045 3547 10103 3553
rect 10229 3587 10287 3593
rect 10229 3553 10241 3587
rect 10275 3584 10287 3587
rect 10321 3587 10379 3593
rect 10321 3584 10333 3587
rect 10275 3556 10333 3584
rect 10275 3553 10287 3556
rect 10229 3547 10287 3553
rect 10321 3553 10333 3556
rect 10367 3584 10379 3587
rect 10778 3584 10784 3596
rect 10367 3556 10784 3584
rect 10367 3553 10379 3556
rect 10321 3547 10379 3553
rect 7892 3488 9076 3516
rect 10060 3516 10088 3547
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 10888 3593 10916 3624
rect 12342 3612 12348 3624
rect 12400 3612 12406 3664
rect 12526 3612 12532 3664
rect 12584 3652 12590 3664
rect 13004 3661 13032 3692
rect 13449 3689 13461 3692
rect 13495 3689 13507 3723
rect 13449 3683 13507 3689
rect 13906 3680 13912 3732
rect 13964 3720 13970 3732
rect 14001 3723 14059 3729
rect 14001 3720 14013 3723
rect 13964 3692 14013 3720
rect 13964 3680 13970 3692
rect 14001 3689 14013 3692
rect 14047 3689 14059 3723
rect 14001 3683 14059 3689
rect 14921 3723 14979 3729
rect 14921 3689 14933 3723
rect 14967 3689 14979 3723
rect 14921 3683 14979 3689
rect 15197 3723 15255 3729
rect 15197 3689 15209 3723
rect 15243 3720 15255 3723
rect 15654 3720 15660 3732
rect 15243 3692 15660 3720
rect 15243 3689 15255 3692
rect 15197 3683 15255 3689
rect 12897 3655 12955 3661
rect 12897 3652 12909 3655
rect 12584 3624 12909 3652
rect 12584 3612 12590 3624
rect 12897 3621 12909 3624
rect 12943 3621 12955 3655
rect 12897 3615 12955 3621
rect 12989 3655 13047 3661
rect 12989 3621 13001 3655
rect 13035 3621 13047 3655
rect 14936 3652 14964 3683
rect 15654 3680 15660 3692
rect 15712 3680 15718 3732
rect 15749 3723 15807 3729
rect 15749 3689 15761 3723
rect 15795 3720 15807 3723
rect 16942 3720 16948 3732
rect 15795 3692 16948 3720
rect 15795 3689 15807 3692
rect 15749 3683 15807 3689
rect 16942 3680 16948 3692
rect 17000 3680 17006 3732
rect 17126 3680 17132 3732
rect 17184 3720 17190 3732
rect 17184 3692 18368 3720
rect 17184 3680 17190 3692
rect 16853 3655 16911 3661
rect 16853 3652 16865 3655
rect 14936 3624 16865 3652
rect 12989 3615 13047 3621
rect 16853 3621 16865 3624
rect 16899 3621 16911 3655
rect 16853 3615 16911 3621
rect 17034 3612 17040 3664
rect 17092 3652 17098 3664
rect 17221 3655 17279 3661
rect 17221 3652 17233 3655
rect 17092 3624 17233 3652
rect 17092 3612 17098 3624
rect 17221 3621 17233 3624
rect 17267 3621 17279 3655
rect 17954 3652 17960 3664
rect 17915 3624 17960 3652
rect 17221 3615 17279 3621
rect 17954 3612 17960 3624
rect 18012 3612 18018 3664
rect 18340 3661 18368 3692
rect 18325 3655 18383 3661
rect 18325 3621 18337 3655
rect 18371 3621 18383 3655
rect 18325 3615 18383 3621
rect 10873 3587 10931 3593
rect 10873 3553 10885 3587
rect 10919 3553 10931 3587
rect 10873 3547 10931 3553
rect 10962 3544 10968 3596
rect 11020 3584 11026 3596
rect 11184 3587 11242 3593
rect 11184 3584 11196 3587
rect 11020 3556 11196 3584
rect 11020 3544 11026 3556
rect 11184 3553 11196 3556
rect 11230 3553 11242 3587
rect 11606 3584 11612 3596
rect 11567 3556 11612 3584
rect 11184 3547 11242 3553
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 11698 3544 11704 3596
rect 11756 3584 11762 3596
rect 11882 3584 11888 3596
rect 11756 3556 11888 3584
rect 11756 3544 11762 3556
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 13208 3587 13266 3593
rect 13208 3553 13220 3587
rect 13254 3553 13266 3587
rect 13208 3547 13266 3553
rect 11054 3516 11060 3528
rect 10060 3488 11060 3516
rect 7892 3476 7898 3488
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 11287 3519 11345 3525
rect 11287 3485 11299 3519
rect 11333 3516 11345 3519
rect 11974 3516 11980 3528
rect 11333 3488 11836 3516
rect 11935 3488 11980 3516
rect 11333 3485 11345 3488
rect 11287 3479 11345 3485
rect 7742 3408 7748 3460
rect 7800 3448 7806 3460
rect 11422 3448 11428 3460
rect 7800 3420 11192 3448
rect 11383 3420 11428 3448
rect 7800 3408 7806 3420
rect 7374 3380 7380 3392
rect 5184 3352 7380 3380
rect 7374 3340 7380 3352
rect 7432 3340 7438 3392
rect 8113 3383 8171 3389
rect 8113 3349 8125 3383
rect 8159 3380 8171 3383
rect 8294 3380 8300 3392
rect 8159 3352 8300 3380
rect 8159 3349 8171 3352
rect 8113 3343 8171 3349
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 8619 3383 8677 3389
rect 8619 3349 8631 3383
rect 8665 3380 8677 3383
rect 9674 3380 9680 3392
rect 8665 3352 9680 3380
rect 8665 3349 8677 3352
rect 8619 3343 8677 3349
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 9766 3340 9772 3392
rect 9824 3380 9830 3392
rect 9861 3383 9919 3389
rect 9861 3380 9873 3383
rect 9824 3352 9873 3380
rect 9824 3340 9830 3352
rect 9861 3349 9873 3352
rect 9907 3349 9919 3383
rect 10410 3380 10416 3392
rect 10371 3352 10416 3380
rect 9861 3343 9919 3349
rect 10410 3340 10416 3352
rect 10468 3340 10474 3392
rect 11054 3380 11060 3392
rect 11015 3352 11060 3380
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 11164 3380 11192 3420
rect 11422 3408 11428 3420
rect 11480 3408 11486 3460
rect 11808 3448 11836 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 12434 3476 12440 3528
rect 12492 3516 12498 3528
rect 13223 3516 13251 3547
rect 13354 3544 13360 3596
rect 13412 3584 13418 3596
rect 13633 3587 13691 3593
rect 13633 3584 13645 3587
rect 13412 3556 13645 3584
rect 13412 3544 13418 3556
rect 13633 3553 13645 3556
rect 13679 3553 13691 3587
rect 13906 3584 13912 3596
rect 13867 3556 13912 3584
rect 13633 3547 13691 3553
rect 13906 3544 13912 3556
rect 13964 3544 13970 3596
rect 14185 3587 14243 3593
rect 14185 3553 14197 3587
rect 14231 3553 14243 3587
rect 14185 3547 14243 3553
rect 12492 3488 13251 3516
rect 12492 3476 12498 3488
rect 12066 3448 12072 3460
rect 11808 3420 12072 3448
rect 12066 3408 12072 3420
rect 12124 3408 12130 3460
rect 12158 3408 12164 3460
rect 12216 3448 12222 3460
rect 13372 3448 13400 3544
rect 13814 3476 13820 3528
rect 13872 3516 13878 3528
rect 14200 3516 14228 3547
rect 14458 3544 14464 3596
rect 14516 3593 14522 3596
rect 14516 3587 14554 3593
rect 14542 3553 14554 3587
rect 14734 3584 14740 3596
rect 14695 3556 14740 3584
rect 14516 3547 14554 3553
rect 14516 3544 14522 3547
rect 14734 3544 14740 3556
rect 14792 3544 14798 3596
rect 15010 3584 15016 3596
rect 14971 3556 15016 3584
rect 15010 3544 15016 3556
rect 15068 3544 15074 3596
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3553 15347 3587
rect 15289 3547 15347 3553
rect 15565 3587 15623 3593
rect 15565 3553 15577 3587
rect 15611 3553 15623 3587
rect 15565 3547 15623 3553
rect 13872 3488 14228 3516
rect 14599 3519 14657 3525
rect 13872 3476 13878 3488
rect 14599 3485 14611 3519
rect 14645 3516 14657 3519
rect 15194 3516 15200 3528
rect 14645 3488 15200 3516
rect 14645 3485 14657 3488
rect 14599 3479 14657 3485
rect 15194 3476 15200 3488
rect 15252 3476 15258 3528
rect 12216 3420 13400 3448
rect 12216 3408 12222 3420
rect 13630 3408 13636 3460
rect 13688 3448 13694 3460
rect 15304 3448 15332 3547
rect 15580 3460 15608 3547
rect 15654 3544 15660 3596
rect 15712 3584 15718 3596
rect 15933 3587 15991 3593
rect 15933 3584 15945 3587
rect 15712 3556 15945 3584
rect 15712 3544 15718 3556
rect 15933 3553 15945 3556
rect 15979 3553 15991 3587
rect 15933 3547 15991 3553
rect 16209 3587 16267 3593
rect 16209 3553 16221 3587
rect 16255 3584 16267 3587
rect 16298 3584 16304 3596
rect 16255 3556 16304 3584
rect 16255 3553 16267 3556
rect 16209 3547 16267 3553
rect 16298 3544 16304 3556
rect 16356 3544 16362 3596
rect 16390 3544 16396 3596
rect 16448 3584 16454 3596
rect 16485 3587 16543 3593
rect 16485 3584 16497 3587
rect 16448 3556 16497 3584
rect 16448 3544 16454 3556
rect 16485 3553 16497 3556
rect 16531 3553 16543 3587
rect 17589 3587 17647 3593
rect 17589 3584 17601 3587
rect 16485 3547 16543 3553
rect 16592 3556 17601 3584
rect 16592 3516 16620 3556
rect 17589 3553 17601 3556
rect 17635 3553 17647 3587
rect 19610 3584 19616 3596
rect 17589 3547 17647 3553
rect 17880 3556 19616 3584
rect 16040 3488 16620 3516
rect 17037 3519 17095 3525
rect 13688 3420 15332 3448
rect 13688 3408 13694 3420
rect 15562 3408 15568 3460
rect 15620 3408 15626 3460
rect 11606 3380 11612 3392
rect 11164 3352 11612 3380
rect 11606 3340 11612 3352
rect 11664 3340 11670 3392
rect 11885 3383 11943 3389
rect 11885 3349 11897 3383
rect 11931 3380 11943 3383
rect 11974 3380 11980 3392
rect 11931 3352 11980 3380
rect 11931 3349 11943 3352
rect 11885 3343 11943 3349
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 13262 3340 13268 3392
rect 13320 3389 13326 3392
rect 13320 3383 13369 3389
rect 13320 3349 13323 3383
rect 13357 3349 13369 3383
rect 13722 3380 13728 3392
rect 13683 3352 13728 3380
rect 13320 3343 13369 3349
rect 13320 3340 13326 3343
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 15473 3383 15531 3389
rect 15473 3349 15485 3383
rect 15519 3380 15531 3383
rect 16040 3380 16068 3488
rect 17037 3485 17049 3519
rect 17083 3516 17095 3519
rect 17880 3516 17908 3556
rect 19610 3544 19616 3556
rect 19668 3544 19674 3596
rect 18598 3516 18604 3528
rect 17083 3488 17908 3516
rect 17972 3488 18604 3516
rect 17083 3485 17095 3488
rect 17037 3479 17095 3485
rect 16117 3451 16175 3457
rect 16117 3417 16129 3451
rect 16163 3448 16175 3451
rect 17218 3448 17224 3460
rect 16163 3420 17224 3448
rect 16163 3417 16175 3420
rect 16117 3411 16175 3417
rect 17218 3408 17224 3420
rect 17276 3408 17282 3460
rect 17405 3451 17463 3457
rect 17405 3417 17417 3451
rect 17451 3448 17463 3451
rect 17972 3448 18000 3488
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 18138 3448 18144 3460
rect 17451 3420 18000 3448
rect 18099 3420 18144 3448
rect 17451 3417 17463 3420
rect 17405 3411 17463 3417
rect 18138 3408 18144 3420
rect 18196 3408 18202 3460
rect 16390 3380 16396 3392
rect 15519 3352 16068 3380
rect 16351 3352 16396 3380
rect 15519 3349 15531 3352
rect 15473 3343 15531 3349
rect 16390 3340 16396 3352
rect 16448 3340 16454 3392
rect 16666 3380 16672 3392
rect 16627 3352 16672 3380
rect 16666 3340 16672 3352
rect 16724 3340 16730 3392
rect 17586 3340 17592 3392
rect 17644 3380 17650 3392
rect 17681 3383 17739 3389
rect 17681 3380 17693 3383
rect 17644 3352 17693 3380
rect 17644 3340 17650 3352
rect 17681 3349 17693 3352
rect 17727 3349 17739 3383
rect 17681 3343 17739 3349
rect 17862 3340 17868 3392
rect 17920 3380 17926 3392
rect 18417 3383 18475 3389
rect 18417 3380 18429 3383
rect 17920 3352 18429 3380
rect 17920 3340 17926 3352
rect 18417 3349 18429 3352
rect 18463 3349 18475 3383
rect 18417 3343 18475 3349
rect 1104 3290 18860 3312
rect 1104 3238 3947 3290
rect 3999 3238 4011 3290
rect 4063 3238 4075 3290
rect 4127 3238 4139 3290
rect 4191 3238 9878 3290
rect 9930 3238 9942 3290
rect 9994 3238 10006 3290
rect 10058 3238 10070 3290
rect 10122 3238 15808 3290
rect 15860 3238 15872 3290
rect 15924 3238 15936 3290
rect 15988 3238 16000 3290
rect 16052 3238 18860 3290
rect 1104 3216 18860 3238
rect 1946 3136 1952 3188
rect 2004 3176 2010 3188
rect 2777 3179 2835 3185
rect 2777 3176 2789 3179
rect 2004 3148 2789 3176
rect 2004 3136 2010 3148
rect 2777 3145 2789 3148
rect 2823 3145 2835 3179
rect 2777 3139 2835 3145
rect 2958 3136 2964 3188
rect 3016 3176 3022 3188
rect 3694 3176 3700 3188
rect 3016 3148 3700 3176
rect 3016 3136 3022 3148
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 4614 3176 4620 3188
rect 4575 3148 4620 3176
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 6178 3136 6184 3188
rect 6236 3176 6242 3188
rect 7101 3179 7159 3185
rect 7101 3176 7113 3179
rect 6236 3148 7113 3176
rect 6236 3136 6242 3148
rect 7101 3145 7113 3148
rect 7147 3145 7159 3179
rect 7101 3139 7159 3145
rect 7745 3179 7803 3185
rect 7745 3145 7757 3179
rect 7791 3176 7803 3179
rect 8018 3176 8024 3188
rect 7791 3148 8024 3176
rect 7791 3145 7803 3148
rect 7745 3139 7803 3145
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 10410 3176 10416 3188
rect 9140 3148 10416 3176
rect 1670 3068 1676 3120
rect 1728 3108 1734 3120
rect 4154 3108 4160 3120
rect 1728 3080 4160 3108
rect 1728 3068 1734 3080
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 4249 3111 4307 3117
rect 4249 3077 4261 3111
rect 4295 3108 4307 3111
rect 5074 3108 5080 3120
rect 4295 3080 5080 3108
rect 4295 3077 4307 3080
rect 4249 3071 4307 3077
rect 2774 3040 2780 3052
rect 1596 3012 2780 3040
rect 1596 2981 1624 3012
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 3050 3000 3056 3052
rect 3108 3040 3114 3052
rect 3108 3012 3556 3040
rect 3108 3000 3114 3012
rect 1581 2975 1639 2981
rect 1581 2941 1593 2975
rect 1627 2941 1639 2975
rect 1581 2935 1639 2941
rect 1949 2975 2007 2981
rect 1949 2941 1961 2975
rect 1995 2972 2007 2975
rect 2038 2972 2044 2984
rect 1995 2944 2044 2972
rect 1995 2941 2007 2944
rect 1949 2935 2007 2941
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 2130 2932 2136 2984
rect 2188 2972 2194 2984
rect 2188 2944 2452 2972
rect 2188 2932 2194 2944
rect 1762 2904 1768 2916
rect 1723 2876 1768 2904
rect 1762 2864 1768 2876
rect 1820 2864 1826 2916
rect 2314 2904 2320 2916
rect 2275 2876 2320 2904
rect 2314 2864 2320 2876
rect 2372 2864 2378 2916
rect 2424 2904 2452 2944
rect 2590 2932 2596 2984
rect 2648 2972 2654 2984
rect 2685 2975 2743 2981
rect 2685 2972 2697 2975
rect 2648 2944 2697 2972
rect 2648 2932 2654 2944
rect 2685 2941 2697 2944
rect 2731 2941 2743 2975
rect 2958 2972 2964 2984
rect 2919 2944 2964 2972
rect 2685 2935 2743 2941
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 3234 2972 3240 2984
rect 3195 2944 3240 2972
rect 3234 2932 3240 2944
rect 3292 2932 3298 2984
rect 3528 2981 3556 3012
rect 3694 3000 3700 3052
rect 3752 3040 3758 3052
rect 4264 3040 4292 3071
rect 5074 3068 5080 3080
rect 5132 3068 5138 3120
rect 6733 3111 6791 3117
rect 6733 3077 6745 3111
rect 6779 3108 6791 3111
rect 7466 3108 7472 3120
rect 6779 3080 7472 3108
rect 6779 3077 6791 3080
rect 6733 3071 6791 3077
rect 7466 3068 7472 3080
rect 7524 3068 7530 3120
rect 8478 3068 8484 3120
rect 8536 3068 8542 3120
rect 9140 3117 9168 3148
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 10505 3179 10563 3185
rect 10505 3145 10517 3179
rect 10551 3145 10563 3179
rect 10505 3139 10563 3145
rect 9125 3111 9183 3117
rect 9125 3077 9137 3111
rect 9171 3077 9183 3111
rect 9125 3071 9183 3077
rect 9674 3068 9680 3120
rect 9732 3108 9738 3120
rect 10134 3108 10140 3120
rect 9732 3080 10140 3108
rect 9732 3068 9738 3080
rect 10134 3068 10140 3080
rect 10192 3068 10198 3120
rect 10226 3068 10232 3120
rect 10284 3108 10290 3120
rect 10520 3108 10548 3139
rect 12526 3136 12532 3188
rect 12584 3176 12590 3188
rect 12986 3185 12992 3188
rect 12667 3179 12725 3185
rect 12667 3176 12679 3179
rect 12584 3148 12679 3176
rect 12584 3136 12590 3148
rect 12667 3145 12679 3148
rect 12713 3145 12725 3179
rect 12667 3139 12725 3145
rect 12943 3179 12992 3185
rect 12943 3145 12955 3179
rect 12989 3145 12992 3179
rect 12943 3139 12992 3145
rect 12986 3136 12992 3139
rect 13044 3136 13050 3188
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 14921 3179 14979 3185
rect 13872 3148 14679 3176
rect 13872 3136 13878 3148
rect 10284 3080 10548 3108
rect 10612 3080 14587 3108
rect 10284 3068 10290 3080
rect 3752 3012 4292 3040
rect 3752 3000 3758 3012
rect 6822 3000 6828 3052
rect 6880 3040 6886 3052
rect 6880 3012 7236 3040
rect 6880 3000 6886 3012
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2941 3571 2975
rect 3786 2972 3792 2984
rect 3747 2944 3792 2972
rect 3513 2935 3571 2941
rect 3786 2932 3792 2944
rect 3844 2932 3850 2984
rect 4062 2972 4068 2984
rect 4023 2944 4068 2972
rect 4062 2932 4068 2944
rect 4120 2932 4126 2984
rect 4338 2972 4344 2984
rect 4299 2944 4344 2972
rect 4338 2932 4344 2944
rect 4396 2932 4402 2984
rect 4614 2932 4620 2984
rect 4672 2972 4678 2984
rect 4801 2975 4859 2981
rect 4801 2972 4813 2975
rect 4672 2944 4813 2972
rect 4672 2932 4678 2944
rect 4801 2941 4813 2944
rect 4847 2972 4859 2975
rect 4893 2975 4951 2981
rect 4893 2972 4905 2975
rect 4847 2944 4905 2972
rect 4847 2941 4859 2944
rect 4801 2935 4859 2941
rect 4893 2941 4905 2944
rect 4939 2941 4951 2975
rect 4893 2935 4951 2941
rect 6549 2975 6607 2981
rect 6549 2941 6561 2975
rect 6595 2972 6607 2975
rect 7208 2972 7236 3012
rect 7282 3000 7288 3052
rect 7340 3040 7346 3052
rect 7926 3040 7932 3052
rect 7340 3012 7932 3040
rect 7340 3000 7346 3012
rect 7926 3000 7932 3012
rect 7984 3040 7990 3052
rect 8496 3040 8524 3068
rect 8573 3043 8631 3049
rect 8573 3040 8585 3043
rect 7984 3012 8432 3040
rect 8496 3012 8585 3040
rect 7984 3000 7990 3012
rect 7377 2975 7435 2981
rect 7377 2972 7389 2975
rect 6595 2944 6960 2972
rect 7208 2944 7389 2972
rect 6595 2941 6607 2944
rect 6549 2935 6607 2941
rect 4246 2904 4252 2916
rect 2424 2876 4252 2904
rect 4246 2864 4252 2876
rect 4304 2864 4310 2916
rect 6932 2904 6960 2944
rect 7377 2941 7389 2944
rect 7423 2972 7435 2975
rect 7469 2975 7527 2981
rect 7469 2972 7481 2975
rect 7423 2944 7481 2972
rect 7423 2941 7435 2944
rect 7377 2935 7435 2941
rect 7469 2941 7481 2944
rect 7515 2941 7527 2975
rect 7469 2935 7527 2941
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 8297 2975 8355 2981
rect 8297 2972 8309 2975
rect 7800 2944 8309 2972
rect 7800 2932 7806 2944
rect 8297 2941 8309 2944
rect 8343 2941 8355 2975
rect 8297 2935 8355 2941
rect 8404 2904 8432 3012
rect 8573 3009 8585 3012
rect 8619 3009 8631 3043
rect 8573 3003 8631 3009
rect 10321 3043 10379 3049
rect 10321 3009 10333 3043
rect 10367 3009 10379 3043
rect 10321 3003 10379 3009
rect 9398 2932 9404 2984
rect 9456 2972 9462 2984
rect 9493 2975 9551 2981
rect 9493 2972 9505 2975
rect 9456 2944 9505 2972
rect 9456 2932 9462 2944
rect 9493 2941 9505 2944
rect 9539 2941 9551 2975
rect 9493 2935 9551 2941
rect 9766 2932 9772 2984
rect 9824 2972 9830 2984
rect 9861 2975 9919 2981
rect 9861 2972 9873 2975
rect 9824 2944 9873 2972
rect 9824 2932 9830 2944
rect 9861 2941 9873 2944
rect 9907 2941 9919 2975
rect 9861 2935 9919 2941
rect 10045 2975 10103 2981
rect 10045 2941 10057 2975
rect 10091 2972 10103 2975
rect 10336 2972 10364 3003
rect 10410 3000 10416 3052
rect 10468 3040 10474 3052
rect 10612 3040 10640 3080
rect 11790 3040 11796 3052
rect 10468 3012 10640 3040
rect 11751 3012 11796 3040
rect 10468 3000 10474 3012
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13722 3040 13728 3052
rect 13219 3012 13728 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 10594 2972 10600 2984
rect 10091 2944 10600 2972
rect 10091 2941 10103 2944
rect 10045 2935 10103 2941
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 10778 2972 10784 2984
rect 10739 2944 10784 2972
rect 10778 2932 10784 2944
rect 10836 2932 10842 2984
rect 10870 2932 10876 2984
rect 10928 2972 10934 2984
rect 11054 2972 11060 2984
rect 10928 2944 10973 2972
rect 11015 2944 11060 2972
rect 10928 2932 10934 2944
rect 11054 2932 11060 2944
rect 11112 2932 11118 2984
rect 12596 2975 12654 2981
rect 12596 2941 12608 2975
rect 12642 2972 12654 2975
rect 12642 2941 12664 2972
rect 12596 2935 12664 2941
rect 8665 2907 8723 2913
rect 8665 2904 8677 2907
rect 6932 2876 8248 2904
rect 8404 2876 8677 2904
rect 1302 2796 1308 2848
rect 1360 2836 1366 2848
rect 1489 2839 1547 2845
rect 1489 2836 1501 2839
rect 1360 2808 1501 2836
rect 1360 2796 1366 2808
rect 1489 2805 1501 2808
rect 1535 2805 1547 2839
rect 2222 2836 2228 2848
rect 2183 2808 2228 2836
rect 1489 2799 1547 2805
rect 2222 2796 2228 2808
rect 2280 2796 2286 2848
rect 2498 2836 2504 2848
rect 2459 2808 2504 2836
rect 2498 2796 2504 2808
rect 2556 2796 2562 2848
rect 3050 2836 3056 2848
rect 3011 2808 3056 2836
rect 3050 2796 3056 2808
rect 3108 2796 3114 2848
rect 3142 2796 3148 2848
rect 3200 2836 3206 2848
rect 3329 2839 3387 2845
rect 3329 2836 3341 2839
rect 3200 2808 3341 2836
rect 3200 2796 3206 2808
rect 3329 2805 3341 2808
rect 3375 2805 3387 2839
rect 3602 2836 3608 2848
rect 3563 2808 3608 2836
rect 3329 2799 3387 2805
rect 3602 2796 3608 2808
rect 3660 2796 3666 2848
rect 3878 2836 3884 2848
rect 3839 2808 3884 2836
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 4522 2836 4528 2848
rect 4483 2808 4528 2836
rect 4522 2796 4528 2808
rect 4580 2796 4586 2848
rect 6932 2845 6960 2876
rect 6917 2839 6975 2845
rect 6917 2805 6929 2839
rect 6963 2805 6975 2839
rect 6917 2799 6975 2805
rect 7834 2796 7840 2848
rect 7892 2836 7898 2848
rect 7929 2839 7987 2845
rect 7929 2836 7941 2839
rect 7892 2808 7941 2836
rect 7892 2796 7898 2808
rect 7929 2805 7941 2808
rect 7975 2805 7987 2839
rect 8110 2836 8116 2848
rect 8071 2808 8116 2836
rect 7929 2799 7987 2805
rect 8110 2796 8116 2808
rect 8168 2796 8174 2848
rect 8220 2836 8248 2876
rect 8665 2873 8677 2876
rect 8711 2873 8723 2907
rect 9674 2904 9680 2916
rect 8665 2867 8723 2873
rect 8772 2876 9444 2904
rect 9635 2876 9680 2904
rect 8772 2836 8800 2876
rect 9306 2836 9312 2848
rect 8220 2808 8800 2836
rect 9267 2808 9312 2836
rect 9306 2796 9312 2808
rect 9364 2796 9370 2848
rect 9416 2836 9444 2876
rect 9674 2864 9680 2876
rect 9732 2864 9738 2916
rect 11425 2907 11483 2913
rect 11425 2904 11437 2907
rect 10428 2876 11437 2904
rect 9766 2836 9772 2848
rect 9416 2808 9772 2836
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 10229 2839 10287 2845
rect 10229 2805 10241 2839
rect 10275 2836 10287 2839
rect 10428 2836 10456 2876
rect 11425 2873 11437 2876
rect 11471 2873 11483 2907
rect 11425 2867 11483 2873
rect 11606 2864 11612 2916
rect 11664 2904 11670 2916
rect 11885 2907 11943 2913
rect 11885 2904 11897 2907
rect 11664 2876 11897 2904
rect 11664 2864 11670 2876
rect 11885 2873 11897 2876
rect 11931 2873 11943 2907
rect 11885 2867 11943 2873
rect 10275 2808 10456 2836
rect 10275 2805 10287 2808
rect 10229 2799 10287 2805
rect 10594 2796 10600 2848
rect 10652 2836 10658 2848
rect 11333 2839 11391 2845
rect 11333 2836 11345 2839
rect 10652 2808 11345 2836
rect 10652 2796 10658 2808
rect 11333 2805 11345 2808
rect 11379 2805 11391 2839
rect 11900 2836 11928 2867
rect 12434 2864 12440 2916
rect 12492 2904 12498 2916
rect 12492 2876 12537 2904
rect 12492 2864 12498 2876
rect 12636 2836 12664 2935
rect 12802 2932 12808 2984
rect 12860 2981 12866 2984
rect 12860 2975 12898 2981
rect 12886 2972 12898 2975
rect 14461 2975 14519 2981
rect 14461 2972 14473 2975
rect 12886 2944 13032 2972
rect 12886 2941 12898 2944
rect 12860 2935 12898 2941
rect 12860 2932 12866 2935
rect 11900 2808 12664 2836
rect 13004 2836 13032 2944
rect 14016 2944 14473 2972
rect 13262 2864 13268 2916
rect 13320 2904 13326 2916
rect 13320 2876 13365 2904
rect 13320 2864 13326 2876
rect 14016 2836 14044 2944
rect 14461 2941 14473 2944
rect 14507 2941 14519 2975
rect 14559 2972 14587 3080
rect 14651 3040 14679 3148
rect 14921 3145 14933 3179
rect 14967 3176 14979 3179
rect 15654 3176 15660 3188
rect 14967 3148 15660 3176
rect 14967 3145 14979 3148
rect 14921 3139 14979 3145
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 16393 3179 16451 3185
rect 16393 3145 16405 3179
rect 16439 3176 16451 3179
rect 16482 3176 16488 3188
rect 16439 3148 16488 3176
rect 16439 3145 16451 3148
rect 16393 3139 16451 3145
rect 16482 3136 16488 3148
rect 16540 3176 16546 3188
rect 16850 3176 16856 3188
rect 16540 3148 16856 3176
rect 16540 3136 16546 3148
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 17037 3179 17095 3185
rect 17037 3145 17049 3179
rect 17083 3176 17095 3179
rect 17126 3176 17132 3188
rect 17083 3148 17132 3176
rect 17083 3145 17095 3148
rect 17037 3139 17095 3145
rect 17126 3136 17132 3148
rect 17184 3136 17190 3188
rect 17678 3136 17684 3188
rect 17736 3176 17742 3188
rect 18417 3179 18475 3185
rect 18417 3176 18429 3179
rect 17736 3148 18429 3176
rect 17736 3136 17742 3148
rect 18417 3145 18429 3148
rect 18463 3145 18475 3179
rect 18417 3139 18475 3145
rect 14734 3068 14740 3120
rect 14792 3108 14798 3120
rect 15933 3111 15991 3117
rect 15933 3108 15945 3111
rect 14792 3080 15945 3108
rect 14792 3068 14798 3080
rect 15933 3077 15945 3080
rect 15979 3077 15991 3111
rect 15933 3071 15991 3077
rect 16666 3068 16672 3120
rect 16724 3108 16730 3120
rect 16724 3080 17724 3108
rect 16724 3068 16730 3080
rect 15381 3043 15439 3049
rect 15381 3040 15393 3043
rect 14651 3012 15393 3040
rect 15381 3009 15393 3012
rect 15427 3009 15439 3043
rect 15381 3003 15439 3009
rect 15470 3000 15476 3052
rect 15528 3040 15534 3052
rect 15565 3043 15623 3049
rect 15565 3040 15577 3043
rect 15528 3012 15577 3040
rect 15528 3000 15534 3012
rect 15565 3009 15577 3012
rect 15611 3009 15623 3043
rect 15746 3040 15752 3052
rect 15707 3012 15752 3040
rect 15565 3003 15623 3009
rect 15746 3000 15752 3012
rect 15804 3000 15810 3052
rect 16390 3000 16396 3052
rect 16448 3040 16454 3052
rect 16448 3012 17632 3040
rect 16448 3000 16454 3012
rect 15105 2975 15163 2981
rect 15105 2972 15117 2975
rect 14559 2944 15117 2972
rect 14461 2935 14519 2941
rect 15105 2941 15117 2944
rect 15151 2941 15163 2975
rect 16574 2972 16580 2984
rect 16535 2944 16580 2972
rect 15105 2935 15163 2941
rect 16574 2932 16580 2944
rect 16632 2932 16638 2984
rect 17126 2972 17132 2984
rect 17087 2944 17132 2972
rect 17126 2932 17132 2944
rect 17184 2932 17190 2984
rect 17218 2932 17224 2984
rect 17276 2972 17282 2984
rect 17604 2981 17632 3012
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 17276 2944 17325 2972
rect 17276 2932 17282 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 17589 2975 17647 2981
rect 17589 2941 17601 2975
rect 17635 2941 17647 2975
rect 17696 2972 17724 3080
rect 17770 3000 17776 3052
rect 17828 3040 17834 3052
rect 17828 3012 18368 3040
rect 17828 3000 17834 3012
rect 18340 2981 18368 3012
rect 17957 2975 18015 2981
rect 17957 2972 17969 2975
rect 17696 2944 17969 2972
rect 17589 2935 17647 2941
rect 17957 2941 17969 2944
rect 18003 2941 18015 2975
rect 17957 2935 18015 2941
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2941 18383 2975
rect 18325 2935 18383 2941
rect 14185 2907 14243 2913
rect 14185 2873 14197 2907
rect 14231 2904 14243 2907
rect 14550 2904 14556 2916
rect 14231 2876 14556 2904
rect 14231 2873 14243 2876
rect 14185 2867 14243 2873
rect 14550 2864 14556 2876
rect 14608 2864 14614 2916
rect 16482 2904 16488 2916
rect 15304 2876 16488 2904
rect 15304 2845 15332 2876
rect 16482 2864 16488 2876
rect 16540 2864 16546 2916
rect 16758 2904 16764 2916
rect 16719 2876 16764 2904
rect 16758 2864 16764 2876
rect 16816 2864 16822 2916
rect 17770 2864 17776 2916
rect 17828 2904 17834 2916
rect 17828 2876 17873 2904
rect 17828 2864 17834 2876
rect 13004 2808 14044 2836
rect 15289 2839 15347 2845
rect 11333 2799 11391 2805
rect 15289 2805 15301 2839
rect 15335 2805 15347 2839
rect 15289 2799 15347 2805
rect 17402 2796 17408 2848
rect 17460 2836 17466 2848
rect 18049 2839 18107 2845
rect 18049 2836 18061 2839
rect 17460 2808 18061 2836
rect 17460 2796 17466 2808
rect 18049 2805 18061 2808
rect 18095 2805 18107 2839
rect 18049 2799 18107 2805
rect 1104 2746 18860 2768
rect 1104 2694 6912 2746
rect 6964 2694 6976 2746
rect 7028 2694 7040 2746
rect 7092 2694 7104 2746
rect 7156 2694 12843 2746
rect 12895 2694 12907 2746
rect 12959 2694 12971 2746
rect 13023 2694 13035 2746
rect 13087 2694 18860 2746
rect 1104 2672 18860 2694
rect 3050 2632 3056 2644
rect 1964 2604 3056 2632
rect 1578 2564 1584 2576
rect 1539 2536 1584 2564
rect 1578 2524 1584 2536
rect 1636 2524 1642 2576
rect 1964 2573 1992 2604
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 4154 2592 4160 2644
rect 4212 2632 4218 2644
rect 4709 2635 4767 2641
rect 4709 2632 4721 2635
rect 4212 2604 4721 2632
rect 4212 2592 4218 2604
rect 4709 2601 4721 2604
rect 4755 2601 4767 2635
rect 4709 2595 4767 2601
rect 5718 2592 5724 2644
rect 5776 2632 5782 2644
rect 5905 2635 5963 2641
rect 5905 2632 5917 2635
rect 5776 2604 5917 2632
rect 5776 2592 5782 2604
rect 5905 2601 5917 2604
rect 5951 2601 5963 2635
rect 5905 2595 5963 2601
rect 6365 2635 6423 2641
rect 6365 2601 6377 2635
rect 6411 2632 6423 2635
rect 6411 2604 7144 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 1949 2567 2007 2573
rect 1949 2533 1961 2567
rect 1995 2533 2007 2567
rect 2590 2564 2596 2576
rect 2551 2536 2596 2564
rect 1949 2527 2007 2533
rect 2590 2524 2596 2536
rect 2648 2524 2654 2576
rect 3142 2564 3148 2576
rect 2792 2536 3148 2564
rect 2317 2499 2375 2505
rect 2317 2465 2329 2499
rect 2363 2496 2375 2499
rect 2792 2496 2820 2536
rect 3142 2524 3148 2536
rect 3200 2524 3206 2576
rect 3602 2564 3608 2576
rect 3252 2536 3608 2564
rect 2363 2468 2820 2496
rect 2869 2499 2927 2505
rect 2363 2465 2375 2468
rect 2317 2459 2375 2465
rect 2869 2465 2881 2499
rect 2915 2496 2927 2499
rect 3252 2496 3280 2536
rect 3602 2524 3608 2536
rect 3660 2524 3666 2576
rect 3878 2524 3884 2576
rect 3936 2564 3942 2576
rect 4065 2567 4123 2573
rect 4065 2564 4077 2567
rect 3936 2536 4077 2564
rect 3936 2524 3942 2536
rect 4065 2533 4077 2536
rect 4111 2533 4123 2567
rect 4430 2564 4436 2576
rect 4391 2536 4436 2564
rect 4065 2527 4123 2533
rect 4430 2524 4436 2536
rect 4488 2524 4494 2576
rect 4522 2524 4528 2576
rect 4580 2564 4586 2576
rect 4801 2567 4859 2573
rect 4801 2564 4813 2567
rect 4580 2536 4813 2564
rect 4580 2524 4586 2536
rect 4801 2533 4813 2536
rect 4847 2533 4859 2567
rect 4801 2527 4859 2533
rect 4982 2524 4988 2576
rect 5040 2564 5046 2576
rect 5169 2567 5227 2573
rect 5169 2564 5181 2567
rect 5040 2536 5181 2564
rect 5040 2524 5046 2536
rect 5169 2533 5181 2536
rect 5215 2533 5227 2567
rect 5169 2527 5227 2533
rect 6638 2524 6644 2576
rect 6696 2564 6702 2576
rect 7116 2573 7144 2604
rect 9766 2592 9772 2644
rect 9824 2632 9830 2644
rect 10962 2632 10968 2644
rect 9824 2604 10968 2632
rect 9824 2592 9830 2604
rect 6733 2567 6791 2573
rect 6733 2564 6745 2567
rect 6696 2536 6745 2564
rect 6696 2524 6702 2536
rect 6733 2533 6745 2536
rect 6779 2533 6791 2567
rect 6733 2527 6791 2533
rect 7101 2567 7159 2573
rect 7101 2533 7113 2567
rect 7147 2533 7159 2567
rect 7466 2564 7472 2576
rect 7427 2536 7472 2564
rect 7101 2527 7159 2533
rect 7466 2524 7472 2536
rect 7524 2524 7530 2576
rect 7837 2567 7895 2573
rect 7837 2533 7849 2567
rect 7883 2564 7895 2567
rect 8110 2564 8116 2576
rect 7883 2536 8116 2564
rect 7883 2533 7895 2536
rect 7837 2527 7895 2533
rect 8110 2524 8116 2536
rect 8168 2524 8174 2576
rect 8294 2564 8300 2576
rect 8255 2536 8300 2564
rect 8294 2524 8300 2536
rect 8352 2524 8358 2576
rect 9214 2564 9220 2576
rect 9175 2536 9220 2564
rect 9214 2524 9220 2536
rect 9272 2524 9278 2576
rect 10134 2564 10140 2576
rect 10095 2536 10140 2564
rect 10134 2524 10140 2536
rect 10192 2524 10198 2576
rect 10502 2564 10508 2576
rect 10463 2536 10508 2564
rect 10502 2524 10508 2536
rect 10560 2524 10566 2576
rect 10612 2573 10640 2604
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 14737 2635 14795 2641
rect 12492 2604 14596 2632
rect 12492 2592 12498 2604
rect 10597 2567 10655 2573
rect 10597 2533 10609 2567
rect 10643 2564 10655 2567
rect 10643 2536 10677 2564
rect 10643 2533 10655 2536
rect 10597 2527 10655 2533
rect 11330 2524 11336 2576
rect 11388 2564 11394 2576
rect 11425 2567 11483 2573
rect 11425 2564 11437 2567
rect 11388 2536 11437 2564
rect 11388 2524 11394 2536
rect 11425 2533 11437 2536
rect 11471 2533 11483 2567
rect 12066 2564 12072 2576
rect 12027 2536 12072 2564
rect 11425 2527 11483 2533
rect 12066 2524 12072 2536
rect 12124 2524 12130 2576
rect 13170 2564 13176 2576
rect 13131 2536 13176 2564
rect 13170 2524 13176 2536
rect 13228 2524 13234 2576
rect 13265 2567 13323 2573
rect 13265 2533 13277 2567
rect 13311 2564 13323 2567
rect 13446 2564 13452 2576
rect 13311 2536 13452 2564
rect 13311 2533 13323 2536
rect 13265 2527 13323 2533
rect 13446 2524 13452 2536
rect 13504 2524 13510 2576
rect 14182 2564 14188 2576
rect 14143 2536 14188 2564
rect 14182 2524 14188 2536
rect 14240 2524 14246 2576
rect 2915 2468 3280 2496
rect 3329 2499 3387 2505
rect 2915 2465 2927 2468
rect 2869 2459 2927 2465
rect 3329 2465 3341 2499
rect 3375 2496 3387 2499
rect 3418 2496 3424 2508
rect 3375 2468 3424 2496
rect 3375 2465 3387 2468
rect 3329 2459 3387 2465
rect 3418 2456 3424 2468
rect 3476 2456 3482 2508
rect 3694 2496 3700 2508
rect 3655 2468 3700 2496
rect 3694 2456 3700 2468
rect 3752 2456 3758 2508
rect 4246 2456 4252 2508
rect 4304 2496 4310 2508
rect 5537 2499 5595 2505
rect 4304 2468 5028 2496
rect 4304 2456 4310 2468
rect 1118 2388 1124 2440
rect 1176 2428 1182 2440
rect 5000 2437 5028 2468
rect 5537 2465 5549 2499
rect 5583 2465 5595 2499
rect 5537 2459 5595 2465
rect 2133 2431 2191 2437
rect 2133 2428 2145 2431
rect 1176 2400 2145 2428
rect 1176 2388 1182 2400
rect 2133 2397 2145 2400
rect 2179 2397 2191 2431
rect 2133 2391 2191 2397
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2397 5043 2431
rect 4985 2391 5043 2397
rect 198 2320 204 2372
rect 256 2360 262 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 256 2332 1409 2360
rect 256 2320 262 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 2682 2360 2688 2372
rect 2643 2332 2688 2360
rect 1397 2323 1455 2329
rect 2682 2320 2688 2332
rect 2740 2320 2746 2372
rect 3142 2360 3148 2372
rect 3103 2332 3148 2360
rect 3142 2320 3148 2332
rect 3200 2320 3206 2372
rect 3602 2320 3608 2372
rect 3660 2360 3666 2372
rect 3881 2363 3939 2369
rect 3881 2360 3893 2363
rect 3660 2332 3893 2360
rect 3660 2320 3666 2332
rect 3881 2329 3893 2332
rect 3927 2329 3939 2363
rect 4246 2360 4252 2372
rect 4207 2332 4252 2360
rect 3881 2323 3939 2329
rect 4246 2320 4252 2332
rect 4304 2320 4310 2372
rect 5166 2320 5172 2372
rect 5224 2360 5230 2372
rect 5353 2363 5411 2369
rect 5353 2360 5365 2363
rect 5224 2332 5365 2360
rect 5224 2320 5230 2332
rect 5353 2329 5365 2332
rect 5399 2329 5411 2363
rect 5353 2323 5411 2329
rect 658 2252 664 2304
rect 716 2292 722 2304
rect 1857 2295 1915 2301
rect 1857 2292 1869 2295
rect 716 2264 1869 2292
rect 716 2252 722 2264
rect 1857 2261 1869 2264
rect 1903 2261 1915 2295
rect 1857 2255 1915 2261
rect 2866 2252 2872 2304
rect 2924 2292 2930 2304
rect 3513 2295 3571 2301
rect 3513 2292 3525 2295
rect 2924 2264 3525 2292
rect 2924 2252 2930 2264
rect 3513 2261 3525 2264
rect 3559 2261 3571 2295
rect 5552 2292 5580 2459
rect 5626 2456 5632 2508
rect 5684 2496 5690 2508
rect 5721 2499 5779 2505
rect 5721 2496 5733 2499
rect 5684 2468 5733 2496
rect 5684 2456 5690 2468
rect 5721 2465 5733 2468
rect 5767 2496 5779 2499
rect 5997 2499 6055 2505
rect 5997 2496 6009 2499
rect 5767 2468 6009 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 5997 2465 6009 2468
rect 6043 2465 6055 2499
rect 5997 2459 6055 2465
rect 6181 2499 6239 2505
rect 6181 2465 6193 2499
rect 6227 2496 6239 2499
rect 7282 2496 7288 2508
rect 6227 2468 7288 2496
rect 6227 2465 6239 2468
rect 6181 2459 6239 2465
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 8849 2499 8907 2505
rect 8849 2465 8861 2499
rect 8895 2496 8907 2499
rect 9306 2496 9312 2508
rect 8895 2468 9312 2496
rect 8895 2465 8907 2468
rect 8849 2459 8907 2465
rect 9306 2456 9312 2468
rect 9364 2456 9370 2508
rect 14568 2505 14596 2604
rect 14737 2601 14749 2635
rect 14783 2632 14795 2635
rect 14783 2604 14964 2632
rect 14783 2601 14795 2604
rect 14737 2595 14795 2601
rect 14936 2573 14964 2604
rect 15194 2592 15200 2644
rect 15252 2632 15258 2644
rect 17405 2635 17463 2641
rect 15252 2604 15424 2632
rect 15252 2592 15258 2604
rect 14921 2567 14979 2573
rect 14921 2533 14933 2567
rect 14967 2533 14979 2567
rect 15286 2564 15292 2576
rect 15247 2536 15292 2564
rect 14921 2527 14979 2533
rect 15286 2524 15292 2536
rect 15344 2524 15350 2576
rect 15396 2573 15424 2604
rect 17405 2601 17417 2635
rect 17451 2632 17463 2635
rect 17451 2604 17632 2632
rect 17451 2601 17463 2604
rect 17405 2595 17463 2601
rect 15381 2567 15439 2573
rect 15381 2533 15393 2567
rect 15427 2533 15439 2567
rect 15381 2527 15439 2533
rect 16206 2524 16212 2576
rect 16264 2564 16270 2576
rect 16301 2567 16359 2573
rect 16301 2564 16313 2567
rect 16264 2536 16313 2564
rect 16264 2524 16270 2536
rect 16301 2533 16313 2536
rect 16347 2533 16359 2567
rect 16301 2527 16359 2533
rect 16482 2524 16488 2576
rect 16540 2564 16546 2576
rect 16577 2567 16635 2573
rect 16577 2564 16589 2567
rect 16540 2536 16589 2564
rect 16540 2524 16546 2536
rect 16577 2533 16589 2536
rect 16623 2533 16635 2567
rect 16942 2564 16948 2576
rect 16903 2536 16948 2564
rect 16577 2527 16635 2533
rect 16942 2524 16948 2536
rect 17000 2524 17006 2576
rect 17604 2573 17632 2604
rect 17589 2567 17647 2573
rect 17589 2533 17601 2567
rect 17635 2533 17647 2567
rect 17589 2527 17647 2533
rect 18046 2524 18052 2576
rect 18104 2564 18110 2576
rect 18325 2567 18383 2573
rect 18325 2564 18337 2567
rect 18104 2536 18337 2564
rect 18104 2524 18110 2536
rect 18325 2533 18337 2536
rect 18371 2533 18383 2567
rect 18325 2527 18383 2533
rect 14553 2499 14611 2505
rect 14553 2465 14565 2499
rect 14599 2465 14611 2499
rect 14553 2459 14611 2465
rect 16850 2456 16856 2508
rect 16908 2496 16914 2508
rect 17221 2499 17279 2505
rect 17221 2496 17233 2499
rect 16908 2468 17233 2496
rect 16908 2456 16914 2468
rect 17221 2465 17233 2468
rect 17267 2465 17279 2499
rect 17221 2459 17279 2465
rect 17957 2499 18015 2505
rect 17957 2465 17969 2499
rect 18003 2496 18015 2499
rect 18414 2496 18420 2508
rect 18003 2468 18420 2496
rect 18003 2465 18015 2468
rect 17957 2459 18015 2465
rect 18414 2456 18420 2468
rect 18472 2456 18478 2508
rect 6638 2388 6644 2440
rect 6696 2428 6702 2440
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6696 2400 6929 2428
rect 6696 2388 6702 2400
rect 6917 2397 6929 2400
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 10229 2431 10287 2437
rect 10229 2397 10241 2431
rect 10275 2428 10287 2431
rect 11422 2428 11428 2440
rect 10275 2400 11428 2428
rect 10275 2397 10287 2400
rect 10229 2391 10287 2397
rect 11422 2388 11428 2400
rect 11480 2388 11486 2440
rect 11974 2428 11980 2440
rect 11935 2400 11980 2428
rect 11974 2388 11980 2400
rect 12032 2388 12038 2440
rect 12618 2428 12624 2440
rect 12579 2400 12624 2428
rect 12618 2388 12624 2400
rect 12676 2388 12682 2440
rect 15105 2431 15163 2437
rect 15105 2397 15117 2431
rect 15151 2428 15163 2431
rect 16666 2428 16672 2440
rect 15151 2400 16672 2428
rect 15151 2397 15163 2400
rect 15105 2391 15163 2397
rect 16666 2388 16672 2400
rect 16724 2388 16730 2440
rect 17494 2388 17500 2440
rect 17552 2428 17558 2440
rect 17678 2428 17684 2440
rect 17552 2400 17684 2428
rect 17552 2388 17558 2400
rect 17678 2388 17684 2400
rect 17736 2388 17742 2440
rect 6178 2320 6184 2372
rect 6236 2360 6242 2372
rect 6549 2363 6607 2369
rect 6549 2360 6561 2363
rect 6236 2332 6561 2360
rect 6236 2320 6242 2332
rect 6549 2329 6561 2332
rect 6595 2329 6607 2363
rect 6549 2323 6607 2329
rect 7098 2320 7104 2372
rect 7156 2360 7162 2372
rect 7285 2363 7343 2369
rect 7285 2360 7297 2363
rect 7156 2332 7297 2360
rect 7156 2320 7162 2332
rect 7285 2329 7297 2332
rect 7331 2329 7343 2363
rect 7650 2360 7656 2372
rect 7611 2332 7656 2360
rect 7285 2323 7343 2329
rect 7650 2320 7656 2332
rect 7708 2320 7714 2372
rect 8110 2360 8116 2372
rect 8071 2332 8116 2360
rect 8110 2320 8116 2332
rect 8168 2320 8174 2372
rect 8662 2360 8668 2372
rect 8623 2332 8668 2360
rect 8662 2320 8668 2332
rect 8720 2320 8726 2372
rect 11057 2363 11115 2369
rect 11057 2329 11069 2363
rect 11103 2360 11115 2363
rect 15562 2360 15568 2372
rect 11103 2332 15568 2360
rect 11103 2329 11115 2332
rect 11057 2323 11115 2329
rect 15562 2320 15568 2332
rect 15620 2320 15626 2372
rect 15654 2320 15660 2372
rect 15712 2360 15718 2372
rect 16393 2363 16451 2369
rect 16393 2360 16405 2363
rect 15712 2332 16405 2360
rect 15712 2320 15718 2332
rect 16393 2329 16405 2332
rect 16439 2329 16451 2363
rect 17770 2360 17776 2372
rect 17731 2332 17776 2360
rect 16393 2323 16451 2329
rect 17770 2320 17776 2332
rect 17828 2320 17834 2372
rect 17862 2320 17868 2372
rect 17920 2360 17926 2372
rect 18509 2363 18567 2369
rect 18509 2360 18521 2363
rect 17920 2332 18521 2360
rect 17920 2320 17926 2332
rect 18509 2329 18521 2332
rect 18555 2329 18567 2363
rect 18509 2323 18567 2329
rect 8018 2292 8024 2304
rect 5552 2264 8024 2292
rect 3513 2255 3571 2261
rect 8018 2252 8024 2264
rect 8076 2252 8082 2304
rect 9122 2252 9128 2304
rect 9180 2292 9186 2304
rect 11333 2295 11391 2301
rect 11333 2292 11345 2295
rect 9180 2264 11345 2292
rect 9180 2252 9186 2264
rect 11333 2261 11345 2264
rect 11379 2261 11391 2295
rect 11333 2255 11391 2261
rect 13906 2252 13912 2304
rect 13964 2292 13970 2304
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 13964 2264 14289 2292
rect 13964 2252 13970 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 14277 2255 14335 2261
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 16172 2264 16865 2292
rect 16172 2252 16178 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 17678 2252 17684 2304
rect 17736 2292 17742 2304
rect 18049 2295 18107 2301
rect 18049 2292 18061 2295
rect 17736 2264 18061 2292
rect 17736 2252 17742 2264
rect 18049 2261 18061 2264
rect 18095 2261 18107 2295
rect 18049 2255 18107 2261
rect 1104 2202 18860 2224
rect 1104 2150 3947 2202
rect 3999 2150 4011 2202
rect 4063 2150 4075 2202
rect 4127 2150 4139 2202
rect 4191 2150 9878 2202
rect 9930 2150 9942 2202
rect 9994 2150 10006 2202
rect 10058 2150 10070 2202
rect 10122 2150 15808 2202
rect 15860 2150 15872 2202
rect 15924 2150 15936 2202
rect 15988 2150 16000 2202
rect 16052 2150 18860 2202
rect 1104 2128 18860 2150
rect 3418 2048 3424 2100
rect 3476 2088 3482 2100
rect 10686 2088 10692 2100
rect 3476 2060 10692 2088
rect 3476 2048 3482 2060
rect 10686 2048 10692 2060
rect 10744 2048 10750 2100
rect 13170 1708 13176 1760
rect 13228 1748 13234 1760
rect 13906 1748 13912 1760
rect 13228 1720 13912 1748
rect 13228 1708 13234 1720
rect 13906 1708 13912 1720
rect 13964 1708 13970 1760
rect 16758 1096 16764 1148
rect 16816 1136 16822 1148
rect 18138 1136 18144 1148
rect 16816 1108 18144 1136
rect 16816 1096 16822 1108
rect 18138 1096 18144 1108
rect 18196 1096 18202 1148
<< via1 >>
rect 296 15104 348 15156
rect 3240 15104 3292 15156
rect 8208 15104 8260 15156
rect 2688 15036 2740 15088
rect 4252 15036 4304 15088
rect 4988 15036 5040 15088
rect 15016 15036 15068 15088
rect 1584 14968 1636 15020
rect 4528 14968 4580 15020
rect 10876 14968 10928 15020
rect 4712 14900 4764 14952
rect 12716 14900 12768 14952
rect 13268 14900 13320 14952
rect 15292 14900 15344 14952
rect 17224 14900 17276 14952
rect 1952 14832 2004 14884
rect 7656 14832 7708 14884
rect 13544 14832 13596 14884
rect 17684 14832 17736 14884
rect 14004 14764 14056 14816
rect 17040 14764 17092 14816
rect 6912 14662 6964 14714
rect 6976 14662 7028 14714
rect 7040 14662 7092 14714
rect 7104 14662 7156 14714
rect 12843 14662 12895 14714
rect 12907 14662 12959 14714
rect 12971 14662 13023 14714
rect 13035 14662 13087 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 1952 14603 2004 14612
rect 1952 14569 1961 14603
rect 1961 14569 1995 14603
rect 1995 14569 2004 14603
rect 1952 14560 2004 14569
rect 2688 14603 2740 14612
rect 2688 14569 2697 14603
rect 2697 14569 2731 14603
rect 2731 14569 2740 14603
rect 2688 14560 2740 14569
rect 1860 14535 1912 14544
rect 1860 14501 1869 14535
rect 1869 14501 1903 14535
rect 1903 14501 1912 14535
rect 1860 14492 1912 14501
rect 2780 14492 2832 14544
rect 8668 14560 8720 14612
rect 3240 14535 3292 14544
rect 3240 14501 3249 14535
rect 3249 14501 3283 14535
rect 3283 14501 3292 14535
rect 3240 14492 3292 14501
rect 3516 14492 3568 14544
rect 4160 14492 4212 14544
rect 4804 14535 4856 14544
rect 4804 14501 4813 14535
rect 4813 14501 4847 14535
rect 4847 14501 4856 14535
rect 4804 14492 4856 14501
rect 4988 14535 5040 14544
rect 4988 14501 4997 14535
rect 4997 14501 5031 14535
rect 5031 14501 5040 14535
rect 4988 14492 5040 14501
rect 5448 14535 5500 14544
rect 5448 14501 5457 14535
rect 5457 14501 5491 14535
rect 5491 14501 5500 14535
rect 5448 14492 5500 14501
rect 6736 14535 6788 14544
rect 6736 14501 6745 14535
rect 6745 14501 6779 14535
rect 6779 14501 6788 14535
rect 6736 14492 6788 14501
rect 7380 14492 7432 14544
rect 1492 14467 1544 14476
rect 1492 14433 1501 14467
rect 1501 14433 1535 14467
rect 1535 14433 1544 14467
rect 1492 14424 1544 14433
rect 2596 14467 2648 14476
rect 2596 14433 2605 14467
rect 2605 14433 2639 14467
rect 2639 14433 2648 14467
rect 2596 14424 2648 14433
rect 3148 14424 3200 14476
rect 3424 14467 3476 14476
rect 3424 14433 3433 14467
rect 3433 14433 3467 14467
rect 3467 14433 3476 14467
rect 3424 14424 3476 14433
rect 3608 14467 3660 14476
rect 3608 14433 3617 14467
rect 3617 14433 3651 14467
rect 3651 14433 3660 14467
rect 3608 14424 3660 14433
rect 2780 14288 2832 14340
rect 2596 14220 2648 14272
rect 3700 14288 3752 14340
rect 5540 14424 5592 14476
rect 5724 14424 5776 14476
rect 6092 14424 6144 14476
rect 6644 14424 6696 14476
rect 11152 14560 11204 14612
rect 13268 14603 13320 14612
rect 13268 14569 13277 14603
rect 13277 14569 13311 14603
rect 13311 14569 13320 14603
rect 13268 14560 13320 14569
rect 13544 14603 13596 14612
rect 13544 14569 13553 14603
rect 13553 14569 13587 14603
rect 13587 14569 13596 14603
rect 13544 14560 13596 14569
rect 13820 14560 13872 14612
rect 17224 14603 17276 14612
rect 11612 14492 11664 14544
rect 12440 14492 12492 14544
rect 12716 14492 12768 14544
rect 14004 14535 14056 14544
rect 14004 14501 14013 14535
rect 14013 14501 14047 14535
rect 14047 14501 14056 14535
rect 14004 14492 14056 14501
rect 14464 14492 14516 14544
rect 15108 14535 15160 14544
rect 15108 14501 15117 14535
rect 15117 14501 15151 14535
rect 15151 14501 15160 14535
rect 15108 14492 15160 14501
rect 9312 14467 9364 14476
rect 9312 14433 9321 14467
rect 9321 14433 9355 14467
rect 9355 14433 9364 14467
rect 9312 14424 9364 14433
rect 9956 14467 10008 14476
rect 9956 14433 9965 14467
rect 9965 14433 9999 14467
rect 9999 14433 10008 14467
rect 9956 14424 10008 14433
rect 10600 14467 10652 14476
rect 10600 14433 10609 14467
rect 10609 14433 10643 14467
rect 10643 14433 10652 14467
rect 10600 14424 10652 14433
rect 11244 14467 11296 14476
rect 11244 14433 11253 14467
rect 11253 14433 11287 14467
rect 11287 14433 11296 14467
rect 11244 14424 11296 14433
rect 11888 14467 11940 14476
rect 11888 14433 11897 14467
rect 11897 14433 11931 14467
rect 11931 14433 11940 14467
rect 11888 14424 11940 14433
rect 12532 14467 12584 14476
rect 12532 14433 12541 14467
rect 12541 14433 12575 14467
rect 12575 14433 12584 14467
rect 12532 14424 12584 14433
rect 13176 14424 13228 14476
rect 13268 14424 13320 14476
rect 13820 14467 13872 14476
rect 13820 14433 13829 14467
rect 13829 14433 13863 14467
rect 13863 14433 13872 14467
rect 13820 14424 13872 14433
rect 14188 14467 14240 14476
rect 14188 14433 14197 14467
rect 14197 14433 14231 14467
rect 14231 14433 14240 14467
rect 14188 14424 14240 14433
rect 14280 14424 14332 14476
rect 14832 14424 14884 14476
rect 17224 14569 17233 14603
rect 17233 14569 17267 14603
rect 17267 14569 17276 14603
rect 17224 14560 17276 14569
rect 15752 14535 15804 14544
rect 15752 14501 15761 14535
rect 15761 14501 15795 14535
rect 15795 14501 15804 14535
rect 15752 14492 15804 14501
rect 16120 14492 16172 14544
rect 16948 14535 17000 14544
rect 16948 14501 16957 14535
rect 16957 14501 16991 14535
rect 16991 14501 17000 14535
rect 16948 14492 17000 14501
rect 17776 14492 17828 14544
rect 17868 14492 17920 14544
rect 15568 14424 15620 14476
rect 16580 14467 16632 14476
rect 16580 14433 16589 14467
rect 16589 14433 16623 14467
rect 16623 14433 16632 14467
rect 17408 14467 17460 14476
rect 16580 14424 16632 14433
rect 17408 14433 17417 14467
rect 17417 14433 17451 14467
rect 17451 14433 17460 14467
rect 17408 14424 17460 14433
rect 18420 14467 18472 14476
rect 18420 14433 18429 14467
rect 18429 14433 18463 14467
rect 18463 14433 18472 14467
rect 18420 14424 18472 14433
rect 15384 14356 15436 14408
rect 3516 14220 3568 14272
rect 5908 14263 5960 14272
rect 5908 14229 5917 14263
rect 5917 14229 5951 14263
rect 5951 14229 5960 14263
rect 5908 14220 5960 14229
rect 6000 14220 6052 14272
rect 8024 14220 8076 14272
rect 8484 14220 8536 14272
rect 10508 14288 10560 14340
rect 10784 14263 10836 14272
rect 10784 14229 10793 14263
rect 10793 14229 10827 14263
rect 10827 14229 10836 14263
rect 10784 14220 10836 14229
rect 11336 14288 11388 14340
rect 13452 14288 13504 14340
rect 13636 14288 13688 14340
rect 14280 14288 14332 14340
rect 16396 14288 16448 14340
rect 16764 14288 16816 14340
rect 18144 14288 18196 14340
rect 14464 14220 14516 14272
rect 15476 14220 15528 14272
rect 17316 14220 17368 14272
rect 17776 14220 17828 14272
rect 3947 14118 3999 14170
rect 4011 14118 4063 14170
rect 4075 14118 4127 14170
rect 4139 14118 4191 14170
rect 9878 14118 9930 14170
rect 9942 14118 9994 14170
rect 10006 14118 10058 14170
rect 10070 14118 10122 14170
rect 15808 14118 15860 14170
rect 15872 14118 15924 14170
rect 15936 14118 15988 14170
rect 16000 14118 16052 14170
rect 3424 14016 3476 14068
rect 3700 14016 3752 14068
rect 4712 14059 4764 14068
rect 4712 14025 4721 14059
rect 4721 14025 4755 14059
rect 4755 14025 4764 14059
rect 4712 14016 4764 14025
rect 5540 14016 5592 14068
rect 6644 14059 6696 14068
rect 2228 13991 2280 14000
rect 2228 13957 2237 13991
rect 2237 13957 2271 13991
rect 2271 13957 2280 13991
rect 2228 13948 2280 13957
rect 2872 13991 2924 14000
rect 2872 13957 2881 13991
rect 2881 13957 2915 13991
rect 2915 13957 2924 13991
rect 2872 13948 2924 13957
rect 5816 13948 5868 14000
rect 940 13744 992 13796
rect 1492 13744 1544 13796
rect 2872 13812 2924 13864
rect 3424 13855 3476 13864
rect 3424 13821 3433 13855
rect 3433 13821 3467 13855
rect 3467 13821 3476 13855
rect 4344 13880 4396 13932
rect 6644 14025 6653 14059
rect 6653 14025 6687 14059
rect 6687 14025 6696 14059
rect 6644 14016 6696 14025
rect 13176 14016 13228 14068
rect 14188 14016 14240 14068
rect 6736 13948 6788 14000
rect 11152 13948 11204 14000
rect 11796 13948 11848 14000
rect 13268 13991 13320 14000
rect 13268 13957 13277 13991
rect 13277 13957 13311 13991
rect 13311 13957 13320 13991
rect 13268 13948 13320 13957
rect 13452 13991 13504 14000
rect 13452 13957 13461 13991
rect 13461 13957 13495 13991
rect 13495 13957 13504 13991
rect 13452 13948 13504 13957
rect 15016 14016 15068 14068
rect 15384 14016 15436 14068
rect 16580 14059 16632 14068
rect 16580 14025 16589 14059
rect 16589 14025 16623 14059
rect 16623 14025 16632 14059
rect 16580 14016 16632 14025
rect 16948 14016 17000 14068
rect 18328 14016 18380 14068
rect 15752 13948 15804 14000
rect 3424 13812 3476 13821
rect 3792 13855 3844 13864
rect 3792 13821 3801 13855
rect 3801 13821 3835 13855
rect 3835 13821 3844 13855
rect 3792 13812 3844 13821
rect 4620 13812 4672 13864
rect 3240 13744 3292 13796
rect 6000 13855 6052 13864
rect 6000 13821 6009 13855
rect 6009 13821 6043 13855
rect 6043 13821 6052 13855
rect 6000 13812 6052 13821
rect 6184 13812 6236 13864
rect 9496 13812 9548 13864
rect 11704 13812 11756 13864
rect 13636 13855 13688 13864
rect 13636 13821 13645 13855
rect 13645 13821 13679 13855
rect 13679 13821 13688 13855
rect 13636 13812 13688 13821
rect 14832 13812 14884 13864
rect 15568 13812 15620 13864
rect 15752 13855 15804 13864
rect 15752 13821 15761 13855
rect 15761 13821 15795 13855
rect 15795 13821 15804 13855
rect 15752 13812 15804 13821
rect 16212 13812 16264 13864
rect 16396 13855 16448 13864
rect 16396 13821 16405 13855
rect 16405 13821 16439 13855
rect 16439 13821 16448 13855
rect 16396 13812 16448 13821
rect 18420 13855 18472 13864
rect 1676 13676 1728 13728
rect 5908 13676 5960 13728
rect 17040 13744 17092 13796
rect 13820 13676 13872 13728
rect 17500 13676 17552 13728
rect 18420 13821 18429 13855
rect 18429 13821 18463 13855
rect 18463 13821 18472 13855
rect 18420 13812 18472 13821
rect 18972 13812 19024 13864
rect 6912 13574 6964 13626
rect 6976 13574 7028 13626
rect 7040 13574 7092 13626
rect 7104 13574 7156 13626
rect 12843 13574 12895 13626
rect 12907 13574 12959 13626
rect 12971 13574 13023 13626
rect 13035 13574 13087 13626
rect 2596 13472 2648 13524
rect 1860 13447 1912 13456
rect 1860 13413 1869 13447
rect 1869 13413 1903 13447
rect 1903 13413 1912 13447
rect 1860 13404 1912 13413
rect 1492 13379 1544 13388
rect 1492 13345 1501 13379
rect 1501 13345 1535 13379
rect 1535 13345 1544 13379
rect 1492 13336 1544 13345
rect 2136 13379 2188 13388
rect 2136 13345 2145 13379
rect 2145 13345 2179 13379
rect 2179 13345 2188 13379
rect 2136 13336 2188 13345
rect 2596 13379 2648 13388
rect 2596 13345 2605 13379
rect 2605 13345 2639 13379
rect 2639 13345 2648 13379
rect 2596 13336 2648 13345
rect 2688 13379 2740 13388
rect 2688 13345 2706 13379
rect 2706 13345 2740 13379
rect 3148 13472 3200 13524
rect 3332 13515 3384 13524
rect 3332 13481 3341 13515
rect 3341 13481 3375 13515
rect 3375 13481 3384 13515
rect 3332 13472 3384 13481
rect 17040 13515 17092 13524
rect 3884 13404 3936 13456
rect 11060 13404 11112 13456
rect 17040 13481 17049 13515
rect 17049 13481 17083 13515
rect 17083 13481 17092 13515
rect 17040 13472 17092 13481
rect 17500 13472 17552 13524
rect 17868 13472 17920 13524
rect 17684 13404 17736 13456
rect 19616 13404 19668 13456
rect 2688 13336 2740 13345
rect 18420 13379 18472 13388
rect 3884 13311 3936 13320
rect 3884 13277 3893 13311
rect 3893 13277 3927 13311
rect 3927 13277 3936 13311
rect 3884 13268 3936 13277
rect 1676 13243 1728 13252
rect 1676 13209 1685 13243
rect 1685 13209 1719 13243
rect 1719 13209 1728 13243
rect 1676 13200 1728 13209
rect 1952 13175 2004 13184
rect 1952 13141 1961 13175
rect 1961 13141 1995 13175
rect 1995 13141 2004 13175
rect 1952 13132 2004 13141
rect 2228 13132 2280 13184
rect 3240 13200 3292 13252
rect 5724 13268 5776 13320
rect 4344 13243 4396 13252
rect 4344 13209 4353 13243
rect 4353 13209 4387 13243
rect 4387 13209 4396 13243
rect 4344 13200 4396 13209
rect 14556 13200 14608 13252
rect 18420 13345 18429 13379
rect 18429 13345 18463 13379
rect 18463 13345 18472 13379
rect 18420 13336 18472 13345
rect 16948 13200 17000 13252
rect 3424 13132 3476 13184
rect 14188 13132 14240 13184
rect 16396 13132 16448 13184
rect 3947 13030 3999 13082
rect 4011 13030 4063 13082
rect 4075 13030 4127 13082
rect 4139 13030 4191 13082
rect 9878 13030 9930 13082
rect 9942 13030 9994 13082
rect 10006 13030 10058 13082
rect 10070 13030 10122 13082
rect 15808 13030 15860 13082
rect 15872 13030 15924 13082
rect 15936 13030 15988 13082
rect 16000 13030 16052 13082
rect 2688 12928 2740 12980
rect 2964 12971 3016 12980
rect 2964 12937 2973 12971
rect 2973 12937 3007 12971
rect 3007 12937 3016 12971
rect 2964 12928 3016 12937
rect 3240 12928 3292 12980
rect 12072 12928 12124 12980
rect 17408 12928 17460 12980
rect 1584 12860 1636 12912
rect 1492 12767 1544 12776
rect 1492 12733 1501 12767
rect 1501 12733 1535 12767
rect 1535 12733 1544 12767
rect 1492 12724 1544 12733
rect 2044 12724 2096 12776
rect 2596 12792 2648 12844
rect 2872 12792 2924 12844
rect 3792 12792 3844 12844
rect 16856 12792 16908 12844
rect 18420 12767 18472 12776
rect 18420 12733 18429 12767
rect 18429 12733 18463 12767
rect 18463 12733 18472 12767
rect 18420 12724 18472 12733
rect 1584 12656 1636 12708
rect 3056 12656 3108 12708
rect 18052 12699 18104 12708
rect 18052 12665 18061 12699
rect 18061 12665 18095 12699
rect 18095 12665 18104 12699
rect 18052 12656 18104 12665
rect 1768 12588 1820 12640
rect 2136 12631 2188 12640
rect 2136 12597 2145 12631
rect 2145 12597 2179 12631
rect 2179 12597 2188 12631
rect 2136 12588 2188 12597
rect 2872 12588 2924 12640
rect 3240 12631 3292 12640
rect 3240 12597 3249 12631
rect 3249 12597 3283 12631
rect 3283 12597 3292 12631
rect 3240 12588 3292 12597
rect 3792 12631 3844 12640
rect 3792 12597 3801 12631
rect 3801 12597 3835 12631
rect 3835 12597 3844 12631
rect 3792 12588 3844 12597
rect 17500 12588 17552 12640
rect 6912 12486 6964 12538
rect 6976 12486 7028 12538
rect 7040 12486 7092 12538
rect 7104 12486 7156 12538
rect 12843 12486 12895 12538
rect 12907 12486 12959 12538
rect 12971 12486 13023 12538
rect 13035 12486 13087 12538
rect 3056 12427 3108 12436
rect 3056 12393 3065 12427
rect 3065 12393 3099 12427
rect 3099 12393 3108 12427
rect 3056 12384 3108 12393
rect 2688 12359 2740 12368
rect 2688 12325 2697 12359
rect 2697 12325 2731 12359
rect 2731 12325 2740 12359
rect 2688 12316 2740 12325
rect 10876 12316 10928 12368
rect 1400 12248 1452 12300
rect 1860 12291 1912 12300
rect 1860 12257 1869 12291
rect 1869 12257 1903 12291
rect 1903 12257 1912 12291
rect 1860 12248 1912 12257
rect 3424 12248 3476 12300
rect 4620 12248 4672 12300
rect 18052 12291 18104 12300
rect 18052 12257 18061 12291
rect 18061 12257 18095 12291
rect 18095 12257 18104 12291
rect 18052 12248 18104 12257
rect 18420 12291 18472 12300
rect 18420 12257 18429 12291
rect 18429 12257 18463 12291
rect 18463 12257 18472 12291
rect 18420 12248 18472 12257
rect 2412 12112 2464 12164
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 2320 12044 2372 12096
rect 2596 12112 2648 12164
rect 2872 12112 2924 12164
rect 4344 12180 4396 12232
rect 16580 12112 16632 12164
rect 3332 12087 3384 12096
rect 3332 12053 3341 12087
rect 3341 12053 3375 12087
rect 3375 12053 3384 12087
rect 3332 12044 3384 12053
rect 3516 12044 3568 12096
rect 3792 12044 3844 12096
rect 6552 12044 6604 12096
rect 18696 12044 18748 12096
rect 3947 11942 3999 11994
rect 4011 11942 4063 11994
rect 4075 11942 4127 11994
rect 4139 11942 4191 11994
rect 9878 11942 9930 11994
rect 9942 11942 9994 11994
rect 10006 11942 10058 11994
rect 10070 11942 10122 11994
rect 15808 11942 15860 11994
rect 15872 11942 15924 11994
rect 15936 11942 15988 11994
rect 16000 11942 16052 11994
rect 1952 11840 2004 11892
rect 6276 11840 6328 11892
rect 2320 11747 2372 11756
rect 2320 11713 2329 11747
rect 2329 11713 2363 11747
rect 2363 11713 2372 11747
rect 2320 11704 2372 11713
rect 2504 11747 2556 11756
rect 2504 11713 2513 11747
rect 2513 11713 2547 11747
rect 2547 11713 2556 11747
rect 2504 11704 2556 11713
rect 1492 11679 1544 11688
rect 1492 11645 1501 11679
rect 1501 11645 1535 11679
rect 1535 11645 1544 11679
rect 1492 11636 1544 11645
rect 2136 11636 2188 11688
rect 4344 11636 4396 11688
rect 6552 11636 6604 11688
rect 2964 11568 3016 11620
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 1952 11500 2004 11552
rect 2504 11500 2556 11552
rect 4712 11568 4764 11620
rect 15108 11704 15160 11756
rect 7564 11636 7616 11688
rect 8116 11636 8168 11688
rect 17868 11679 17920 11688
rect 17868 11645 17877 11679
rect 17877 11645 17911 11679
rect 17911 11645 17920 11679
rect 17868 11636 17920 11645
rect 8944 11568 8996 11620
rect 18420 11611 18472 11620
rect 18420 11577 18429 11611
rect 18429 11577 18463 11611
rect 18463 11577 18472 11611
rect 18420 11568 18472 11577
rect 4620 11500 4672 11552
rect 7288 11500 7340 11552
rect 7840 11543 7892 11552
rect 7840 11509 7849 11543
rect 7849 11509 7883 11543
rect 7883 11509 7892 11543
rect 7840 11500 7892 11509
rect 17316 11500 17368 11552
rect 18236 11500 18288 11552
rect 18788 11500 18840 11552
rect 6912 11398 6964 11450
rect 6976 11398 7028 11450
rect 7040 11398 7092 11450
rect 7104 11398 7156 11450
rect 12843 11398 12895 11450
rect 12907 11398 12959 11450
rect 12971 11398 13023 11450
rect 13035 11398 13087 11450
rect 4712 11296 4764 11348
rect 5908 11296 5960 11348
rect 6460 11296 6512 11348
rect 17868 11296 17920 11348
rect 18604 11296 18656 11348
rect 1400 11160 1452 11212
rect 2228 11203 2280 11212
rect 2228 11169 2237 11203
rect 2237 11169 2271 11203
rect 2271 11169 2280 11203
rect 2228 11160 2280 11169
rect 2412 11160 2464 11212
rect 2320 11135 2372 11144
rect 2320 11101 2329 11135
rect 2329 11101 2363 11135
rect 2363 11101 2372 11135
rect 2320 11092 2372 11101
rect 2504 11135 2556 11144
rect 2504 11101 2513 11135
rect 2513 11101 2547 11135
rect 2547 11101 2556 11135
rect 2504 11092 2556 11101
rect 3056 11024 3108 11076
rect 1860 10999 1912 11008
rect 1860 10965 1869 10999
rect 1869 10965 1903 10999
rect 1903 10965 1912 10999
rect 1860 10956 1912 10965
rect 2688 10999 2740 11008
rect 2688 10965 2697 10999
rect 2697 10965 2731 10999
rect 2731 10965 2740 10999
rect 2688 10956 2740 10965
rect 4528 11160 4580 11212
rect 4988 11160 5040 11212
rect 3424 11092 3476 11144
rect 6644 11228 6696 11280
rect 7012 11228 7064 11280
rect 7840 11228 7892 11280
rect 11888 11228 11940 11280
rect 11980 11228 12032 11280
rect 3516 11067 3568 11076
rect 3516 11033 3525 11067
rect 3525 11033 3559 11067
rect 3559 11033 3568 11067
rect 3516 11024 3568 11033
rect 4712 11024 4764 11076
rect 3700 10956 3752 11008
rect 5724 10999 5776 11008
rect 5724 10965 5733 10999
rect 5733 10965 5767 10999
rect 5767 10965 5776 10999
rect 5724 10956 5776 10965
rect 5908 11024 5960 11076
rect 6276 11135 6328 11144
rect 6276 11101 6285 11135
rect 6285 11101 6319 11135
rect 6319 11101 6328 11135
rect 6276 11092 6328 11101
rect 7380 11160 7432 11212
rect 11704 11160 11756 11212
rect 13544 11203 13596 11212
rect 6552 11092 6604 11144
rect 11888 11092 11940 11144
rect 13544 11169 13562 11203
rect 13562 11169 13596 11203
rect 13544 11160 13596 11169
rect 18512 11160 18564 11212
rect 6828 10999 6880 11008
rect 6828 10965 6837 10999
rect 6837 10965 6871 10999
rect 6871 10965 6880 10999
rect 6828 10956 6880 10965
rect 9772 10956 9824 11008
rect 10324 10956 10376 11008
rect 12256 11024 12308 11076
rect 11612 10956 11664 11008
rect 11888 10999 11940 11008
rect 11888 10965 11897 10999
rect 11897 10965 11931 10999
rect 11931 10965 11940 10999
rect 11888 10956 11940 10965
rect 16028 11092 16080 11144
rect 16304 11092 16356 11144
rect 18052 11092 18104 11144
rect 14096 11024 14148 11076
rect 17776 11067 17828 11076
rect 14924 10956 14976 11008
rect 16948 10999 17000 11008
rect 16948 10965 16957 10999
rect 16957 10965 16991 10999
rect 16991 10965 17000 10999
rect 16948 10956 17000 10965
rect 17132 10956 17184 11008
rect 17776 11033 17785 11067
rect 17785 11033 17819 11067
rect 17819 11033 17828 11067
rect 17776 11024 17828 11033
rect 3947 10854 3999 10906
rect 4011 10854 4063 10906
rect 4075 10854 4127 10906
rect 4139 10854 4191 10906
rect 9878 10854 9930 10906
rect 9942 10854 9994 10906
rect 10006 10854 10058 10906
rect 10070 10854 10122 10906
rect 15808 10854 15860 10906
rect 15872 10854 15924 10906
rect 15936 10854 15988 10906
rect 16000 10854 16052 10906
rect 2228 10752 2280 10804
rect 2136 10684 2188 10736
rect 11888 10752 11940 10804
rect 13544 10795 13596 10804
rect 13544 10761 13553 10795
rect 13553 10761 13587 10795
rect 13587 10761 13596 10795
rect 13544 10752 13596 10761
rect 6092 10684 6144 10736
rect 6828 10684 6880 10736
rect 1768 10616 1820 10668
rect 2688 10616 2740 10668
rect 4252 10616 4304 10668
rect 2136 10591 2188 10600
rect 2136 10557 2145 10591
rect 2145 10557 2179 10591
rect 2179 10557 2188 10591
rect 2136 10548 2188 10557
rect 3332 10548 3384 10600
rect 1492 10523 1544 10532
rect 1492 10489 1501 10523
rect 1501 10489 1535 10523
rect 1535 10489 1544 10523
rect 1492 10480 1544 10489
rect 3424 10480 3476 10532
rect 3608 10480 3660 10532
rect 4344 10548 4396 10600
rect 5448 10548 5500 10600
rect 5908 10616 5960 10668
rect 7012 10659 7064 10668
rect 7012 10625 7021 10659
rect 7021 10625 7055 10659
rect 7055 10625 7064 10659
rect 7012 10616 7064 10625
rect 7196 10684 7248 10736
rect 7380 10684 7432 10736
rect 6460 10548 6512 10600
rect 7196 10548 7248 10600
rect 7288 10548 7340 10600
rect 10324 10616 10376 10668
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 1768 10412 1820 10464
rect 2596 10455 2648 10464
rect 2596 10421 2605 10455
rect 2605 10421 2639 10455
rect 2639 10421 2648 10455
rect 2596 10412 2648 10421
rect 2964 10412 3016 10464
rect 4896 10412 4948 10464
rect 5724 10412 5776 10464
rect 6000 10412 6052 10464
rect 9772 10480 9824 10532
rect 10692 10548 10744 10600
rect 11704 10548 11756 10600
rect 12256 10616 12308 10668
rect 13268 10659 13320 10668
rect 13268 10625 13277 10659
rect 13277 10625 13311 10659
rect 13311 10625 13320 10659
rect 16764 10684 16816 10736
rect 17224 10684 17276 10736
rect 14924 10659 14976 10668
rect 13268 10616 13320 10625
rect 14924 10625 14933 10659
rect 14933 10625 14967 10659
rect 14967 10625 14976 10659
rect 14924 10616 14976 10625
rect 16488 10616 16540 10668
rect 17776 10616 17828 10668
rect 16672 10548 16724 10600
rect 8760 10455 8812 10464
rect 8760 10421 8769 10455
rect 8769 10421 8803 10455
rect 8803 10421 8812 10455
rect 8760 10412 8812 10421
rect 10140 10412 10192 10464
rect 10416 10412 10468 10464
rect 11244 10455 11296 10464
rect 11244 10421 11253 10455
rect 11253 10421 11287 10455
rect 11287 10421 11296 10455
rect 11244 10412 11296 10421
rect 11888 10480 11940 10532
rect 13360 10480 13412 10532
rect 14004 10480 14056 10532
rect 17684 10480 17736 10532
rect 17868 10523 17920 10532
rect 17868 10489 17877 10523
rect 17877 10489 17911 10523
rect 17911 10489 17920 10523
rect 17868 10480 17920 10489
rect 18144 10480 18196 10532
rect 18420 10523 18472 10532
rect 18420 10489 18429 10523
rect 18429 10489 18463 10523
rect 18463 10489 18472 10523
rect 18420 10480 18472 10489
rect 13176 10412 13228 10464
rect 13728 10412 13780 10464
rect 16580 10412 16632 10464
rect 16948 10455 17000 10464
rect 16948 10421 16957 10455
rect 16957 10421 16991 10455
rect 16991 10421 17000 10455
rect 16948 10412 17000 10421
rect 17592 10412 17644 10464
rect 17776 10412 17828 10464
rect 6912 10310 6964 10362
rect 6976 10310 7028 10362
rect 7040 10310 7092 10362
rect 7104 10310 7156 10362
rect 12843 10310 12895 10362
rect 12907 10310 12959 10362
rect 12971 10310 13023 10362
rect 13035 10310 13087 10362
rect 1860 10251 1912 10260
rect 1860 10217 1869 10251
rect 1869 10217 1903 10251
rect 1903 10217 1912 10251
rect 1860 10208 1912 10217
rect 1952 10251 2004 10260
rect 1952 10217 1961 10251
rect 1961 10217 1995 10251
rect 1995 10217 2004 10251
rect 1952 10208 2004 10217
rect 2320 10208 2372 10260
rect 2872 10251 2924 10260
rect 2872 10217 2881 10251
rect 2881 10217 2915 10251
rect 2915 10217 2924 10251
rect 2872 10208 2924 10217
rect 3424 10251 3476 10260
rect 3424 10217 3433 10251
rect 3433 10217 3467 10251
rect 3467 10217 3476 10251
rect 3424 10208 3476 10217
rect 3516 10208 3568 10260
rect 3700 10251 3752 10260
rect 3700 10217 3709 10251
rect 3709 10217 3743 10251
rect 3743 10217 3752 10251
rect 3700 10208 3752 10217
rect 4896 10251 4948 10260
rect 4896 10217 4905 10251
rect 4905 10217 4939 10251
rect 4939 10217 4948 10251
rect 4896 10208 4948 10217
rect 4620 10140 4672 10192
rect 6368 10208 6420 10260
rect 8208 10208 8260 10260
rect 10876 10251 10928 10260
rect 10876 10217 10885 10251
rect 10885 10217 10919 10251
rect 10919 10217 10928 10251
rect 10876 10208 10928 10217
rect 6000 10140 6052 10192
rect 3700 10072 3752 10124
rect 3884 10072 3936 10124
rect 8760 10140 8812 10192
rect 11612 10208 11664 10260
rect 12072 10208 12124 10260
rect 12348 10251 12400 10260
rect 12348 10217 12357 10251
rect 12357 10217 12391 10251
rect 12391 10217 12400 10251
rect 12348 10208 12400 10217
rect 13544 10208 13596 10260
rect 13728 10251 13780 10260
rect 13728 10217 13737 10251
rect 13737 10217 13771 10251
rect 13771 10217 13780 10251
rect 13728 10208 13780 10217
rect 16488 10208 16540 10260
rect 16672 10208 16724 10260
rect 17592 10251 17644 10260
rect 17592 10217 17601 10251
rect 17601 10217 17635 10251
rect 17635 10217 17644 10251
rect 17592 10208 17644 10217
rect 17684 10251 17736 10260
rect 17684 10217 17693 10251
rect 17693 10217 17727 10251
rect 17727 10217 17736 10251
rect 18052 10251 18104 10260
rect 17684 10208 17736 10217
rect 18052 10217 18061 10251
rect 18061 10217 18095 10251
rect 18095 10217 18104 10251
rect 18052 10208 18104 10217
rect 2964 10047 3016 10056
rect 2964 10013 2973 10047
rect 2973 10013 3007 10047
rect 3007 10013 3016 10047
rect 2964 10004 3016 10013
rect 3792 10004 3844 10056
rect 1400 9911 1452 9920
rect 1400 9877 1409 9911
rect 1409 9877 1443 9911
rect 1443 9877 1452 9911
rect 1400 9868 1452 9877
rect 3056 9868 3108 9920
rect 3240 9911 3292 9920
rect 3240 9877 3249 9911
rect 3249 9877 3283 9911
rect 3283 9877 3292 9911
rect 3240 9868 3292 9877
rect 4344 9868 4396 9920
rect 7288 10072 7340 10124
rect 5908 10047 5960 10056
rect 5908 10013 5917 10047
rect 5917 10013 5951 10047
rect 5951 10013 5960 10047
rect 5908 10004 5960 10013
rect 6644 10047 6696 10056
rect 6644 10013 6653 10047
rect 6653 10013 6687 10047
rect 6687 10013 6696 10047
rect 6644 10004 6696 10013
rect 10692 10072 10744 10124
rect 17960 10140 18012 10192
rect 11612 10115 11664 10124
rect 9772 10047 9824 10056
rect 6368 9936 6420 9988
rect 9772 10013 9781 10047
rect 9781 10013 9815 10047
rect 9815 10013 9824 10047
rect 9772 10004 9824 10013
rect 11612 10081 11621 10115
rect 11621 10081 11655 10115
rect 11655 10081 11664 10115
rect 11612 10072 11664 10081
rect 11888 10072 11940 10124
rect 7196 9868 7248 9920
rect 7380 9868 7432 9920
rect 11704 9936 11756 9988
rect 12256 9936 12308 9988
rect 8852 9868 8904 9920
rect 10324 9911 10376 9920
rect 10324 9877 10333 9911
rect 10333 9877 10367 9911
rect 10367 9877 10376 9911
rect 10324 9868 10376 9877
rect 10876 9868 10928 9920
rect 12532 9868 12584 9920
rect 14924 10072 14976 10124
rect 13268 10004 13320 10056
rect 13176 9936 13228 9988
rect 13820 9936 13872 9988
rect 13912 9868 13964 9920
rect 17592 10072 17644 10124
rect 17132 10047 17184 10056
rect 17132 10013 17141 10047
rect 17141 10013 17175 10047
rect 17175 10013 17184 10047
rect 17132 10004 17184 10013
rect 17316 9936 17368 9988
rect 15384 9868 15436 9920
rect 16120 9868 16172 9920
rect 16764 9911 16816 9920
rect 16764 9877 16773 9911
rect 16773 9877 16807 9911
rect 16807 9877 16816 9911
rect 16764 9868 16816 9877
rect 3947 9766 3999 9818
rect 4011 9766 4063 9818
rect 4075 9766 4127 9818
rect 4139 9766 4191 9818
rect 9878 9766 9930 9818
rect 9942 9766 9994 9818
rect 10006 9766 10058 9818
rect 10070 9766 10122 9818
rect 15808 9766 15860 9818
rect 15872 9766 15924 9818
rect 15936 9766 15988 9818
rect 16000 9766 16052 9818
rect 1584 9664 1636 9716
rect 5448 9707 5500 9716
rect 2136 9460 2188 9512
rect 3516 9596 3568 9648
rect 5448 9673 5457 9707
rect 5457 9673 5491 9707
rect 5491 9673 5500 9707
rect 5448 9664 5500 9673
rect 5724 9664 5776 9716
rect 7196 9664 7248 9716
rect 8668 9664 8720 9716
rect 9128 9707 9180 9716
rect 9128 9673 9137 9707
rect 9137 9673 9171 9707
rect 9171 9673 9180 9707
rect 9128 9664 9180 9673
rect 9772 9664 9824 9716
rect 3332 9528 3384 9580
rect 6000 9596 6052 9648
rect 6644 9596 6696 9648
rect 8208 9596 8260 9648
rect 8300 9596 8352 9648
rect 10140 9596 10192 9648
rect 10232 9596 10284 9648
rect 10692 9664 10744 9716
rect 16396 9664 16448 9716
rect 16580 9664 16632 9716
rect 17776 9664 17828 9716
rect 15660 9639 15712 9648
rect 6552 9528 6604 9580
rect 8852 9528 8904 9580
rect 10416 9571 10468 9580
rect 10416 9537 10425 9571
rect 10425 9537 10459 9571
rect 10459 9537 10468 9571
rect 10416 9528 10468 9537
rect 11612 9528 11664 9580
rect 12072 9571 12124 9580
rect 12072 9537 12081 9571
rect 12081 9537 12115 9571
rect 12115 9537 12124 9571
rect 12072 9528 12124 9537
rect 15660 9605 15669 9639
rect 15669 9605 15703 9639
rect 15703 9605 15712 9639
rect 15660 9596 15712 9605
rect 18052 9596 18104 9648
rect 3792 9460 3844 9512
rect 4068 9503 4120 9512
rect 4068 9469 4077 9503
rect 4077 9469 4111 9503
rect 4111 9469 4120 9503
rect 4068 9460 4120 9469
rect 8208 9460 8260 9512
rect 9404 9460 9456 9512
rect 9864 9460 9916 9512
rect 10324 9503 10376 9512
rect 10324 9469 10333 9503
rect 10333 9469 10367 9503
rect 10367 9469 10376 9503
rect 10324 9460 10376 9469
rect 10968 9460 11020 9512
rect 12624 9460 12676 9512
rect 13268 9528 13320 9580
rect 16488 9571 16540 9580
rect 14372 9460 14424 9512
rect 16488 9537 16497 9571
rect 16497 9537 16531 9571
rect 16531 9537 16540 9571
rect 16488 9528 16540 9537
rect 15384 9503 15436 9512
rect 15384 9469 15393 9503
rect 15393 9469 15427 9503
rect 15427 9469 15436 9503
rect 17408 9528 17460 9580
rect 17592 9571 17644 9580
rect 17592 9537 17601 9571
rect 17601 9537 17635 9571
rect 17635 9537 17644 9571
rect 17592 9528 17644 9537
rect 15384 9460 15436 9469
rect 1492 9435 1544 9444
rect 1492 9401 1501 9435
rect 1501 9401 1535 9435
rect 1535 9401 1544 9435
rect 1492 9392 1544 9401
rect 3976 9392 4028 9444
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 1952 9367 2004 9376
rect 1952 9333 1961 9367
rect 1961 9333 1995 9367
rect 1995 9333 2004 9367
rect 1952 9324 2004 9333
rect 2136 9367 2188 9376
rect 2136 9333 2145 9367
rect 2145 9333 2179 9367
rect 2179 9333 2188 9367
rect 2136 9324 2188 9333
rect 2596 9367 2648 9376
rect 2596 9333 2605 9367
rect 2605 9333 2639 9367
rect 2639 9333 2648 9367
rect 2596 9324 2648 9333
rect 2872 9367 2924 9376
rect 2872 9333 2881 9367
rect 2881 9333 2915 9367
rect 2915 9333 2924 9367
rect 2872 9324 2924 9333
rect 3424 9324 3476 9376
rect 3700 9367 3752 9376
rect 3700 9333 3709 9367
rect 3709 9333 3743 9367
rect 3743 9333 3752 9367
rect 3700 9324 3752 9333
rect 4620 9392 4672 9444
rect 4436 9324 4488 9376
rect 4896 9367 4948 9376
rect 4896 9333 4905 9367
rect 4905 9333 4939 9367
rect 4939 9333 4948 9367
rect 4896 9324 4948 9333
rect 5908 9367 5960 9376
rect 5908 9333 5917 9367
rect 5917 9333 5951 9367
rect 5951 9333 5960 9367
rect 5908 9324 5960 9333
rect 6368 9392 6420 9444
rect 6736 9392 6788 9444
rect 7380 9392 7432 9444
rect 10692 9392 10744 9444
rect 13268 9435 13320 9444
rect 6644 9324 6696 9376
rect 8300 9324 8352 9376
rect 9680 9324 9732 9376
rect 10140 9324 10192 9376
rect 13268 9401 13277 9435
rect 13277 9401 13311 9435
rect 13311 9401 13320 9435
rect 13268 9392 13320 9401
rect 11060 9324 11112 9376
rect 11336 9324 11388 9376
rect 11888 9324 11940 9376
rect 12440 9367 12492 9376
rect 12440 9333 12449 9367
rect 12449 9333 12483 9367
rect 12483 9333 12492 9367
rect 12440 9324 12492 9333
rect 12624 9324 12676 9376
rect 14740 9392 14792 9444
rect 15016 9392 15068 9444
rect 16764 9460 16816 9512
rect 17316 9435 17368 9444
rect 14004 9367 14056 9376
rect 14004 9333 14013 9367
rect 14013 9333 14047 9367
rect 14047 9333 14056 9367
rect 14004 9324 14056 9333
rect 15936 9367 15988 9376
rect 15936 9333 15945 9367
rect 15945 9333 15979 9367
rect 15979 9333 15988 9367
rect 15936 9324 15988 9333
rect 16212 9324 16264 9376
rect 17316 9401 17325 9435
rect 17325 9401 17359 9435
rect 17359 9401 17368 9435
rect 17316 9392 17368 9401
rect 17868 9435 17920 9444
rect 17868 9401 17877 9435
rect 17877 9401 17911 9435
rect 17911 9401 17920 9435
rect 17868 9392 17920 9401
rect 18052 9435 18104 9444
rect 18052 9401 18061 9435
rect 18061 9401 18095 9435
rect 18095 9401 18104 9435
rect 18052 9392 18104 9401
rect 18144 9392 18196 9444
rect 18420 9435 18472 9444
rect 18420 9401 18429 9435
rect 18429 9401 18463 9435
rect 18463 9401 18472 9435
rect 18420 9392 18472 9401
rect 17408 9367 17460 9376
rect 17408 9333 17417 9367
rect 17417 9333 17451 9367
rect 17451 9333 17460 9367
rect 17408 9324 17460 9333
rect 6912 9222 6964 9274
rect 6976 9222 7028 9274
rect 7040 9222 7092 9274
rect 7104 9222 7156 9274
rect 12843 9222 12895 9274
rect 12907 9222 12959 9274
rect 12971 9222 13023 9274
rect 13035 9222 13087 9274
rect 3332 9120 3384 9172
rect 3516 9120 3568 9172
rect 4620 9120 4672 9172
rect 4712 9120 4764 9172
rect 4896 9120 4948 9172
rect 5908 9120 5960 9172
rect 6000 9120 6052 9172
rect 7748 9120 7800 9172
rect 9956 9120 10008 9172
rect 10968 9163 11020 9172
rect 10968 9129 10977 9163
rect 10977 9129 11011 9163
rect 11011 9129 11020 9163
rect 10968 9120 11020 9129
rect 11244 9120 11296 9172
rect 12440 9163 12492 9172
rect 12440 9129 12449 9163
rect 12449 9129 12483 9163
rect 12483 9129 12492 9163
rect 12440 9120 12492 9129
rect 14648 9120 14700 9172
rect 15384 9120 15436 9172
rect 15936 9120 15988 9172
rect 16212 9163 16264 9172
rect 16212 9129 16221 9163
rect 16221 9129 16255 9163
rect 16255 9129 16264 9163
rect 16212 9120 16264 9129
rect 17776 9120 17828 9172
rect 1584 9052 1636 9104
rect 5356 9052 5408 9104
rect 6644 9095 6696 9104
rect 6644 9061 6653 9095
rect 6653 9061 6687 9095
rect 6687 9061 6696 9095
rect 6644 9052 6696 9061
rect 8852 9052 8904 9104
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 1676 8984 1728 9036
rect 2412 8984 2464 9036
rect 1860 8959 1912 8968
rect 1860 8925 1869 8959
rect 1869 8925 1903 8959
rect 1903 8925 1912 8959
rect 1860 8916 1912 8925
rect 3424 8959 3476 8968
rect 3424 8925 3433 8959
rect 3433 8925 3467 8959
rect 3467 8925 3476 8959
rect 3424 8916 3476 8925
rect 3976 8891 4028 8900
rect 3976 8857 3985 8891
rect 3985 8857 4019 8891
rect 4019 8857 4028 8891
rect 3976 8848 4028 8857
rect 6368 8984 6420 9036
rect 7288 9027 7340 9036
rect 7288 8993 7297 9027
rect 7297 8993 7331 9027
rect 7331 8993 7340 9027
rect 7288 8984 7340 8993
rect 7840 8984 7892 9036
rect 9588 9027 9640 9036
rect 9588 8993 9597 9027
rect 9597 8993 9631 9027
rect 9631 8993 9640 9027
rect 9588 8984 9640 8993
rect 10324 8984 10376 9036
rect 10968 8984 11020 9036
rect 12256 9052 12308 9104
rect 12532 9052 12584 9104
rect 13268 9052 13320 9104
rect 15660 9052 15712 9104
rect 11888 8984 11940 9036
rect 6552 8916 6604 8968
rect 8668 8916 8720 8968
rect 9772 8916 9824 8968
rect 3792 8780 3844 8832
rect 11612 8916 11664 8968
rect 16948 8984 17000 9036
rect 10692 8848 10744 8900
rect 12808 8848 12860 8900
rect 13728 8959 13780 8968
rect 13728 8925 13737 8959
rect 13737 8925 13771 8959
rect 13771 8925 13780 8959
rect 13728 8916 13780 8925
rect 14004 8916 14056 8968
rect 16488 8916 16540 8968
rect 16672 8959 16724 8968
rect 16672 8925 16681 8959
rect 16681 8925 16715 8959
rect 16715 8925 16724 8959
rect 16672 8916 16724 8925
rect 17684 8984 17736 9036
rect 18420 9027 18472 9036
rect 16212 8848 16264 8900
rect 17316 8916 17368 8968
rect 17592 8959 17644 8968
rect 17592 8925 17601 8959
rect 17601 8925 17635 8959
rect 17635 8925 17644 8959
rect 17592 8916 17644 8925
rect 8024 8780 8076 8832
rect 8668 8823 8720 8832
rect 8668 8789 8677 8823
rect 8677 8789 8711 8823
rect 8711 8789 8720 8823
rect 8668 8780 8720 8789
rect 9036 8780 9088 8832
rect 9312 8780 9364 8832
rect 9680 8780 9732 8832
rect 10416 8780 10468 8832
rect 11336 8780 11388 8832
rect 11704 8780 11756 8832
rect 12348 8780 12400 8832
rect 13268 8780 13320 8832
rect 13544 8780 13596 8832
rect 13820 8780 13872 8832
rect 14004 8780 14056 8832
rect 14924 8780 14976 8832
rect 16396 8780 16448 8832
rect 18420 8993 18429 9027
rect 18429 8993 18463 9027
rect 18463 8993 18472 9027
rect 18420 8984 18472 8993
rect 18236 8959 18288 8968
rect 18236 8925 18245 8959
rect 18245 8925 18279 8959
rect 18279 8925 18288 8959
rect 18236 8916 18288 8925
rect 18236 8780 18288 8832
rect 3947 8678 3999 8730
rect 4011 8678 4063 8730
rect 4075 8678 4127 8730
rect 4139 8678 4191 8730
rect 9878 8678 9930 8730
rect 9942 8678 9994 8730
rect 10006 8678 10058 8730
rect 10070 8678 10122 8730
rect 15808 8678 15860 8730
rect 15872 8678 15924 8730
rect 15936 8678 15988 8730
rect 16000 8678 16052 8730
rect 2596 8576 2648 8628
rect 3424 8576 3476 8628
rect 6000 8576 6052 8628
rect 6368 8576 6420 8628
rect 13820 8576 13872 8628
rect 16212 8576 16264 8628
rect 16396 8576 16448 8628
rect 16672 8576 16724 8628
rect 2964 8551 3016 8560
rect 2964 8517 2973 8551
rect 2973 8517 3007 8551
rect 3007 8517 3016 8551
rect 2964 8508 3016 8517
rect 6092 8551 6144 8560
rect 6092 8517 6101 8551
rect 6101 8517 6135 8551
rect 6135 8517 6144 8551
rect 6092 8508 6144 8517
rect 8024 8551 8076 8560
rect 1860 8372 1912 8424
rect 3608 8372 3660 8424
rect 2964 8304 3016 8356
rect 5448 8440 5500 8492
rect 8024 8517 8033 8551
rect 8033 8517 8067 8551
rect 8067 8517 8076 8551
rect 8024 8508 8076 8517
rect 8668 8508 8720 8560
rect 9956 8551 10008 8560
rect 7840 8483 7892 8492
rect 7840 8449 7849 8483
rect 7849 8449 7883 8483
rect 7883 8449 7892 8483
rect 7840 8440 7892 8449
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 9956 8517 9965 8551
rect 9965 8517 9999 8551
rect 9999 8517 10008 8551
rect 9956 8508 10008 8517
rect 13452 8508 13504 8560
rect 13636 8508 13688 8560
rect 13728 8483 13780 8492
rect 7288 8372 7340 8424
rect 9312 8372 9364 8424
rect 11704 8415 11756 8424
rect 11704 8381 11713 8415
rect 11713 8381 11747 8415
rect 11747 8381 11756 8415
rect 11704 8372 11756 8381
rect 13728 8449 13737 8483
rect 13737 8449 13771 8483
rect 13771 8449 13780 8483
rect 13728 8440 13780 8449
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 16948 8508 17000 8560
rect 15844 8440 15896 8492
rect 16212 8440 16264 8492
rect 17592 8483 17644 8492
rect 17592 8449 17601 8483
rect 17601 8449 17635 8483
rect 17635 8449 17644 8483
rect 17592 8440 17644 8449
rect 1584 8236 1636 8288
rect 6552 8304 6604 8356
rect 7564 8347 7616 8356
rect 7564 8313 7582 8347
rect 7582 8313 7616 8347
rect 7564 8304 7616 8313
rect 7748 8304 7800 8356
rect 3608 8279 3660 8288
rect 3608 8245 3617 8279
rect 3617 8245 3651 8279
rect 3651 8245 3660 8279
rect 3608 8236 3660 8245
rect 5172 8279 5224 8288
rect 5172 8245 5181 8279
rect 5181 8245 5215 8279
rect 5215 8245 5224 8279
rect 5172 8236 5224 8245
rect 5632 8279 5684 8288
rect 5632 8245 5641 8279
rect 5641 8245 5675 8279
rect 5675 8245 5684 8279
rect 5632 8236 5684 8245
rect 6276 8236 6328 8288
rect 8208 8236 8260 8288
rect 8300 8236 8352 8288
rect 10232 8304 10284 8356
rect 15752 8372 15804 8424
rect 18144 8440 18196 8492
rect 18328 8415 18380 8424
rect 15660 8304 15712 8356
rect 16764 8347 16816 8356
rect 16764 8313 16773 8347
rect 16773 8313 16807 8347
rect 16807 8313 16816 8347
rect 16764 8304 16816 8313
rect 11796 8236 11848 8288
rect 11980 8236 12032 8288
rect 12716 8236 12768 8288
rect 13176 8279 13228 8288
rect 13176 8245 13185 8279
rect 13185 8245 13219 8279
rect 13219 8245 13228 8279
rect 13176 8236 13228 8245
rect 13820 8236 13872 8288
rect 15752 8236 15804 8288
rect 15844 8236 15896 8288
rect 16672 8236 16724 8288
rect 16948 8304 17000 8356
rect 17776 8304 17828 8356
rect 18328 8381 18337 8415
rect 18337 8381 18371 8415
rect 18371 8381 18380 8415
rect 18328 8372 18380 8381
rect 18512 8347 18564 8356
rect 18512 8313 18521 8347
rect 18521 8313 18555 8347
rect 18555 8313 18564 8347
rect 18512 8304 18564 8313
rect 18052 8279 18104 8288
rect 18052 8245 18061 8279
rect 18061 8245 18095 8279
rect 18095 8245 18104 8279
rect 18052 8236 18104 8245
rect 6912 8134 6964 8186
rect 6976 8134 7028 8186
rect 7040 8134 7092 8186
rect 7104 8134 7156 8186
rect 12843 8134 12895 8186
rect 12907 8134 12959 8186
rect 12971 8134 13023 8186
rect 13035 8134 13087 8186
rect 1860 8075 1912 8084
rect 1860 8041 1869 8075
rect 1869 8041 1903 8075
rect 1903 8041 1912 8075
rect 1860 8032 1912 8041
rect 3424 8075 3476 8084
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 4252 8075 4304 8084
rect 4252 8041 4261 8075
rect 4261 8041 4295 8075
rect 4295 8041 4304 8075
rect 4252 8032 4304 8041
rect 5080 8032 5132 8084
rect 5264 8032 5316 8084
rect 5356 8032 5408 8084
rect 5632 8032 5684 8084
rect 6552 8075 6604 8084
rect 6552 8041 6561 8075
rect 6561 8041 6595 8075
rect 6595 8041 6604 8075
rect 6552 8032 6604 8041
rect 6644 8032 6696 8084
rect 2872 7964 2924 8016
rect 5816 7964 5868 8016
rect 7380 8032 7432 8084
rect 9128 8032 9180 8084
rect 9312 8032 9364 8084
rect 16304 8075 16356 8084
rect 2136 7896 2188 7948
rect 3424 7896 3476 7948
rect 3700 7896 3752 7948
rect 5356 7896 5408 7948
rect 5632 7896 5684 7948
rect 6368 7896 6420 7948
rect 8300 7964 8352 8016
rect 7748 7896 7800 7948
rect 8116 7896 8168 7948
rect 11980 7964 12032 8016
rect 12716 7964 12768 8016
rect 12992 8007 13044 8016
rect 12992 7973 13001 8007
rect 13001 7973 13035 8007
rect 13035 7973 13044 8007
rect 12992 7964 13044 7973
rect 8944 7896 8996 7948
rect 9404 7896 9456 7948
rect 13084 7896 13136 7948
rect 2964 7828 3016 7880
rect 3516 7828 3568 7880
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5307 7871
rect 5307 7837 5316 7871
rect 5264 7828 5316 7837
rect 5448 7871 5500 7880
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 6276 7871 6328 7880
rect 6276 7837 6285 7871
rect 6285 7837 6319 7871
rect 6319 7837 6328 7871
rect 7104 7871 7156 7880
rect 6276 7828 6328 7837
rect 7104 7837 7113 7871
rect 7113 7837 7147 7871
rect 7147 7837 7156 7871
rect 7104 7828 7156 7837
rect 7564 7828 7616 7880
rect 8392 7828 8444 7880
rect 8668 7828 8720 7880
rect 12348 7871 12400 7880
rect 12348 7837 12357 7871
rect 12357 7837 12391 7871
rect 12391 7837 12400 7871
rect 12348 7828 12400 7837
rect 7288 7760 7340 7812
rect 12808 7803 12860 7812
rect 1492 7735 1544 7744
rect 1492 7701 1501 7735
rect 1501 7701 1535 7735
rect 1535 7701 1544 7735
rect 1492 7692 1544 7701
rect 2412 7692 2464 7744
rect 4620 7692 4672 7744
rect 7748 7692 7800 7744
rect 11060 7692 11112 7744
rect 12808 7769 12817 7803
rect 12817 7769 12851 7803
rect 12851 7769 12860 7803
rect 12808 7760 12860 7769
rect 13728 7964 13780 8016
rect 13820 7896 13872 7948
rect 14096 7964 14148 8016
rect 15384 7964 15436 8016
rect 14648 7896 14700 7948
rect 15660 7896 15712 7948
rect 16304 8041 16313 8075
rect 16313 8041 16347 8075
rect 16347 8041 16356 8075
rect 16304 8032 16356 8041
rect 16672 8032 16724 8084
rect 16948 8075 17000 8084
rect 16948 8041 16957 8075
rect 16957 8041 16991 8075
rect 16991 8041 17000 8075
rect 16948 8032 17000 8041
rect 17408 8032 17460 8084
rect 17960 8032 18012 8084
rect 18696 8032 18748 8084
rect 17316 7964 17368 8016
rect 18236 7964 18288 8016
rect 17132 7828 17184 7880
rect 17776 7896 17828 7948
rect 17684 7871 17736 7880
rect 14648 7760 14700 7812
rect 17684 7837 17693 7871
rect 17693 7837 17727 7871
rect 17727 7837 17736 7871
rect 17684 7828 17736 7837
rect 18512 7803 18564 7812
rect 18512 7769 18521 7803
rect 18521 7769 18555 7803
rect 18555 7769 18564 7803
rect 18512 7760 18564 7769
rect 11704 7692 11756 7744
rect 13544 7692 13596 7744
rect 14372 7692 14424 7744
rect 16304 7692 16356 7744
rect 16488 7735 16540 7744
rect 16488 7701 16497 7735
rect 16497 7701 16531 7735
rect 16531 7701 16540 7735
rect 16488 7692 16540 7701
rect 16764 7692 16816 7744
rect 18420 7692 18472 7744
rect 3947 7590 3999 7642
rect 4011 7590 4063 7642
rect 4075 7590 4127 7642
rect 4139 7590 4191 7642
rect 9878 7590 9930 7642
rect 9942 7590 9994 7642
rect 10006 7590 10058 7642
rect 10070 7590 10122 7642
rect 15808 7590 15860 7642
rect 15872 7590 15924 7642
rect 15936 7590 15988 7642
rect 16000 7590 16052 7642
rect 2044 7488 2096 7540
rect 3332 7488 3384 7540
rect 5080 7531 5132 7540
rect 5080 7497 5089 7531
rect 5089 7497 5123 7531
rect 5123 7497 5132 7531
rect 5080 7488 5132 7497
rect 5264 7488 5316 7540
rect 6644 7488 6696 7540
rect 11888 7531 11940 7540
rect 2872 7463 2924 7472
rect 2872 7429 2881 7463
rect 2881 7429 2915 7463
rect 2915 7429 2924 7463
rect 2872 7420 2924 7429
rect 1584 7352 1636 7404
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 2964 7352 3016 7404
rect 3424 7420 3476 7472
rect 4252 7420 4304 7472
rect 5816 7420 5868 7472
rect 2412 7327 2464 7336
rect 2412 7293 2421 7327
rect 2421 7293 2455 7327
rect 2455 7293 2464 7327
rect 2412 7284 2464 7293
rect 3608 7352 3660 7404
rect 5356 7395 5408 7404
rect 5356 7361 5365 7395
rect 5365 7361 5399 7395
rect 5399 7361 5408 7395
rect 5356 7352 5408 7361
rect 4620 7327 4672 7336
rect 4620 7293 4629 7327
rect 4629 7293 4663 7327
rect 4663 7293 4672 7327
rect 4620 7284 4672 7293
rect 5172 7284 5224 7336
rect 5540 7284 5592 7336
rect 6644 7352 6696 7404
rect 7104 7395 7156 7404
rect 7104 7361 7113 7395
rect 7113 7361 7147 7395
rect 7147 7361 7156 7395
rect 7104 7352 7156 7361
rect 8392 7395 8444 7404
rect 8392 7361 8401 7395
rect 8401 7361 8435 7395
rect 8435 7361 8444 7395
rect 8392 7352 8444 7361
rect 3240 7148 3292 7200
rect 5632 7216 5684 7268
rect 6368 7216 6420 7268
rect 8576 7284 8628 7336
rect 9312 7284 9364 7336
rect 10140 7463 10192 7472
rect 10140 7429 10149 7463
rect 10149 7429 10183 7463
rect 10183 7429 10192 7463
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 12348 7488 12400 7540
rect 10140 7420 10192 7429
rect 12164 7463 12216 7472
rect 12164 7429 12173 7463
rect 12173 7429 12207 7463
rect 12207 7429 12216 7463
rect 12164 7420 12216 7429
rect 6644 7148 6696 7200
rect 7380 7191 7432 7200
rect 7380 7157 7389 7191
rect 7389 7157 7423 7191
rect 7423 7157 7432 7191
rect 7380 7148 7432 7157
rect 7656 7148 7708 7200
rect 8116 7191 8168 7200
rect 8116 7157 8125 7191
rect 8125 7157 8159 7191
rect 8159 7157 8168 7191
rect 8116 7148 8168 7157
rect 8208 7191 8260 7200
rect 8208 7157 8217 7191
rect 8217 7157 8251 7191
rect 8251 7157 8260 7191
rect 8760 7216 8812 7268
rect 10968 7284 11020 7336
rect 11704 7327 11756 7336
rect 11704 7293 11713 7327
rect 11713 7293 11747 7327
rect 11747 7293 11756 7327
rect 11704 7284 11756 7293
rect 12992 7488 13044 7540
rect 13268 7488 13320 7540
rect 15200 7488 15252 7540
rect 15384 7488 15436 7540
rect 17960 7488 18012 7540
rect 12716 7420 12768 7472
rect 13084 7352 13136 7404
rect 13544 7395 13596 7404
rect 12624 7327 12676 7336
rect 12624 7293 12633 7327
rect 12633 7293 12667 7327
rect 12667 7293 12676 7327
rect 12624 7284 12676 7293
rect 13176 7284 13228 7336
rect 13544 7361 13553 7395
rect 13553 7361 13587 7395
rect 13587 7361 13596 7395
rect 13544 7352 13596 7361
rect 13820 7420 13872 7472
rect 18328 7420 18380 7472
rect 11980 7216 12032 7268
rect 8208 7148 8260 7157
rect 12072 7148 12124 7200
rect 12808 7216 12860 7268
rect 14004 7216 14056 7268
rect 14372 7284 14424 7336
rect 15384 7284 15436 7336
rect 18144 7395 18196 7404
rect 18144 7361 18153 7395
rect 18153 7361 18187 7395
rect 18187 7361 18196 7395
rect 18144 7352 18196 7361
rect 15660 7284 15712 7336
rect 15844 7284 15896 7336
rect 16488 7284 16540 7336
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 17408 7284 17460 7336
rect 18052 7284 18104 7336
rect 13636 7148 13688 7200
rect 15384 7148 15436 7200
rect 17224 7216 17276 7268
rect 17500 7216 17552 7268
rect 18512 7259 18564 7268
rect 18512 7225 18521 7259
rect 18521 7225 18555 7259
rect 18555 7225 18564 7259
rect 18512 7216 18564 7225
rect 16304 7191 16356 7200
rect 16304 7157 16313 7191
rect 16313 7157 16347 7191
rect 16347 7157 16356 7191
rect 17132 7191 17184 7200
rect 16304 7148 16356 7157
rect 17132 7157 17141 7191
rect 17141 7157 17175 7191
rect 17175 7157 17184 7191
rect 17132 7148 17184 7157
rect 17776 7191 17828 7200
rect 17776 7157 17785 7191
rect 17785 7157 17819 7191
rect 17819 7157 17828 7191
rect 17776 7148 17828 7157
rect 6912 7046 6964 7098
rect 6976 7046 7028 7098
rect 7040 7046 7092 7098
rect 7104 7046 7156 7098
rect 12843 7046 12895 7098
rect 12907 7046 12959 7098
rect 12971 7046 13023 7098
rect 13035 7046 13087 7098
rect 2504 6876 2556 6928
rect 2780 6876 2832 6928
rect 1768 6851 1820 6860
rect 1768 6817 1777 6851
rect 1777 6817 1811 6851
rect 1811 6817 1820 6851
rect 1768 6808 1820 6817
rect 2964 6876 3016 6928
rect 6276 6944 6328 6996
rect 7748 6987 7800 6996
rect 7748 6953 7757 6987
rect 7757 6953 7791 6987
rect 7791 6953 7800 6987
rect 7748 6944 7800 6953
rect 8208 6944 8260 6996
rect 8300 6944 8352 6996
rect 11244 6944 11296 6996
rect 11980 6987 12032 6996
rect 11980 6953 11989 6987
rect 11989 6953 12023 6987
rect 12023 6953 12032 6987
rect 11980 6944 12032 6953
rect 12348 6944 12400 6996
rect 13636 6987 13688 6996
rect 13636 6953 13645 6987
rect 13645 6953 13679 6987
rect 13679 6953 13688 6987
rect 13636 6944 13688 6953
rect 1492 6647 1544 6656
rect 1492 6613 1501 6647
rect 1501 6613 1535 6647
rect 1535 6613 1544 6647
rect 1492 6604 1544 6613
rect 3516 6808 3568 6860
rect 7380 6876 7432 6928
rect 7656 6919 7708 6928
rect 7656 6885 7665 6919
rect 7665 6885 7699 6919
rect 7699 6885 7708 6919
rect 7656 6876 7708 6885
rect 11060 6876 11112 6928
rect 6920 6808 6972 6860
rect 7564 6808 7616 6860
rect 8208 6808 8260 6860
rect 3608 6672 3660 6724
rect 2504 6604 2556 6656
rect 4252 6740 4304 6792
rect 6828 6740 6880 6792
rect 8300 6740 8352 6792
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 11888 6808 11940 6860
rect 12072 6783 12124 6792
rect 10140 6672 10192 6724
rect 12072 6749 12081 6783
rect 12081 6749 12115 6783
rect 12115 6749 12124 6783
rect 12072 6740 12124 6749
rect 13268 6876 13320 6928
rect 15016 6944 15068 6996
rect 15384 6944 15436 6996
rect 16120 6944 16172 6996
rect 16304 6944 16356 6996
rect 16580 6944 16632 6996
rect 16948 6944 17000 6996
rect 17132 6944 17184 6996
rect 13820 6876 13872 6928
rect 17316 6876 17368 6928
rect 12808 6740 12860 6792
rect 13084 6740 13136 6792
rect 14280 6808 14332 6860
rect 15384 6808 15436 6860
rect 15752 6808 15804 6860
rect 16580 6808 16632 6860
rect 16672 6808 16724 6860
rect 18328 6851 18380 6860
rect 14372 6783 14424 6792
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 5264 6604 5316 6656
rect 7472 6604 7524 6656
rect 11336 6604 11388 6656
rect 11520 6647 11572 6656
rect 11520 6613 11529 6647
rect 11529 6613 11563 6647
rect 11563 6613 11572 6647
rect 11520 6604 11572 6613
rect 11980 6604 12032 6656
rect 16948 6740 17000 6792
rect 16488 6672 16540 6724
rect 17132 6740 17184 6792
rect 18328 6817 18337 6851
rect 18337 6817 18371 6851
rect 18371 6817 18380 6851
rect 18328 6808 18380 6817
rect 17224 6715 17276 6724
rect 17224 6681 17233 6715
rect 17233 6681 17267 6715
rect 17267 6681 17276 6715
rect 17224 6672 17276 6681
rect 18512 6715 18564 6724
rect 18512 6681 18521 6715
rect 18521 6681 18555 6715
rect 18555 6681 18564 6715
rect 18512 6672 18564 6681
rect 16396 6604 16448 6656
rect 16672 6604 16724 6656
rect 18052 6647 18104 6656
rect 18052 6613 18061 6647
rect 18061 6613 18095 6647
rect 18095 6613 18104 6647
rect 18052 6604 18104 6613
rect 3947 6502 3999 6554
rect 4011 6502 4063 6554
rect 4075 6502 4127 6554
rect 4139 6502 4191 6554
rect 9878 6502 9930 6554
rect 9942 6502 9994 6554
rect 10006 6502 10058 6554
rect 10070 6502 10122 6554
rect 15808 6502 15860 6554
rect 15872 6502 15924 6554
rect 15936 6502 15988 6554
rect 16000 6502 16052 6554
rect 3516 6443 3568 6452
rect 3516 6409 3525 6443
rect 3525 6409 3559 6443
rect 3559 6409 3568 6443
rect 3516 6400 3568 6409
rect 3608 6400 3660 6452
rect 7840 6400 7892 6452
rect 8116 6400 8168 6452
rect 4896 6332 4948 6384
rect 5816 6332 5868 6384
rect 7656 6332 7708 6384
rect 3424 6307 3476 6316
rect 3424 6273 3433 6307
rect 3433 6273 3467 6307
rect 3467 6273 3476 6307
rect 3424 6264 3476 6273
rect 1952 6239 2004 6248
rect 1952 6205 1961 6239
rect 1961 6205 1995 6239
rect 1995 6205 2004 6239
rect 1952 6196 2004 6205
rect 4988 6264 5040 6316
rect 10784 6400 10836 6452
rect 8392 6332 8444 6384
rect 10692 6375 10744 6384
rect 10692 6341 10701 6375
rect 10701 6341 10735 6375
rect 10735 6341 10744 6375
rect 10692 6332 10744 6341
rect 1492 6103 1544 6112
rect 1492 6069 1501 6103
rect 1501 6069 1535 6103
rect 1535 6069 1544 6103
rect 1492 6060 1544 6069
rect 3332 6060 3384 6112
rect 3424 6060 3476 6112
rect 4252 6060 4304 6112
rect 5540 6196 5592 6248
rect 5816 6239 5868 6248
rect 5816 6205 5825 6239
rect 5825 6205 5859 6239
rect 5859 6205 5868 6239
rect 5816 6196 5868 6205
rect 6828 6239 6880 6248
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 6920 6239 6972 6248
rect 6920 6205 6929 6239
rect 6929 6205 6963 6239
rect 6963 6205 6972 6239
rect 8760 6264 8812 6316
rect 6920 6196 6972 6205
rect 9128 6196 9180 6248
rect 10324 6239 10376 6248
rect 10324 6205 10342 6239
rect 10342 6205 10376 6239
rect 10324 6196 10376 6205
rect 10784 6196 10836 6248
rect 17500 6443 17552 6452
rect 17500 6409 17509 6443
rect 17509 6409 17543 6443
rect 17543 6409 17552 6443
rect 17500 6400 17552 6409
rect 11336 6196 11388 6248
rect 13176 6332 13228 6384
rect 16856 6332 16908 6384
rect 17408 6332 17460 6384
rect 15660 6264 15712 6316
rect 16120 6307 16172 6316
rect 16120 6273 16129 6307
rect 16129 6273 16163 6307
rect 16163 6273 16172 6307
rect 16120 6264 16172 6273
rect 16672 6307 16724 6316
rect 16672 6273 16681 6307
rect 16681 6273 16715 6307
rect 16715 6273 16724 6307
rect 16672 6264 16724 6273
rect 13176 6239 13228 6248
rect 5264 6128 5316 6180
rect 13176 6205 13185 6239
rect 13185 6205 13219 6239
rect 13219 6205 13228 6239
rect 13176 6196 13228 6205
rect 15200 6196 15252 6248
rect 16028 6196 16080 6248
rect 16580 6196 16632 6248
rect 17684 6196 17736 6248
rect 18052 6196 18104 6248
rect 11888 6128 11940 6180
rect 5448 6103 5500 6112
rect 5448 6069 5457 6103
rect 5457 6069 5491 6103
rect 5491 6069 5500 6103
rect 5448 6060 5500 6069
rect 6000 6060 6052 6112
rect 6460 6103 6512 6112
rect 6460 6069 6469 6103
rect 6469 6069 6503 6103
rect 6503 6069 6512 6103
rect 6460 6060 6512 6069
rect 7840 6060 7892 6112
rect 12992 6128 13044 6180
rect 12348 6060 12400 6112
rect 17224 6128 17276 6180
rect 14648 6060 14700 6112
rect 15844 6060 15896 6112
rect 16120 6060 16172 6112
rect 16396 6060 16448 6112
rect 16580 6060 16632 6112
rect 18512 6171 18564 6180
rect 18512 6137 18521 6171
rect 18521 6137 18555 6171
rect 18555 6137 18564 6171
rect 18512 6128 18564 6137
rect 18236 6060 18288 6112
rect 6912 5958 6964 6010
rect 6976 5958 7028 6010
rect 7040 5958 7092 6010
rect 7104 5958 7156 6010
rect 12843 5958 12895 6010
rect 12907 5958 12959 6010
rect 12971 5958 13023 6010
rect 13035 5958 13087 6010
rect 1952 5856 2004 5908
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 5448 5856 5500 5908
rect 6000 5856 6052 5908
rect 7288 5856 7340 5908
rect 10784 5856 10836 5908
rect 10968 5856 11020 5908
rect 11336 5856 11388 5908
rect 11520 5856 11572 5908
rect 15660 5856 15712 5908
rect 15844 5899 15896 5908
rect 15844 5865 15853 5899
rect 15853 5865 15887 5899
rect 15887 5865 15896 5899
rect 15844 5856 15896 5865
rect 16028 5856 16080 5908
rect 18052 5899 18104 5908
rect 2596 5788 2648 5840
rect 2780 5831 2832 5840
rect 2780 5797 2789 5831
rect 2789 5797 2823 5831
rect 2823 5797 2832 5831
rect 2780 5788 2832 5797
rect 6460 5788 6512 5840
rect 17316 5788 17368 5840
rect 2872 5720 2924 5772
rect 3332 5720 3384 5772
rect 3424 5695 3476 5704
rect 3424 5661 3433 5695
rect 3433 5661 3467 5695
rect 3467 5661 3476 5695
rect 3424 5652 3476 5661
rect 5816 5720 5868 5772
rect 6092 5720 6144 5772
rect 6736 5720 6788 5772
rect 7932 5720 7984 5772
rect 8852 5720 8904 5772
rect 9128 5763 9180 5772
rect 9128 5729 9137 5763
rect 9137 5729 9171 5763
rect 9171 5729 9180 5763
rect 9128 5720 9180 5729
rect 12256 5720 12308 5772
rect 13268 5763 13320 5772
rect 13268 5729 13277 5763
rect 13277 5729 13311 5763
rect 13311 5729 13320 5763
rect 13268 5720 13320 5729
rect 13912 5720 13964 5772
rect 14648 5763 14700 5772
rect 14648 5729 14682 5763
rect 14682 5729 14700 5763
rect 14648 5720 14700 5729
rect 15660 5720 15712 5772
rect 16028 5720 16080 5772
rect 16580 5720 16632 5772
rect 4988 5652 5040 5704
rect 5356 5652 5408 5704
rect 11520 5652 11572 5704
rect 11980 5695 12032 5704
rect 11980 5661 11989 5695
rect 11989 5661 12023 5695
rect 12023 5661 12032 5695
rect 11980 5652 12032 5661
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 1584 5516 1636 5568
rect 2964 5559 3016 5568
rect 2964 5525 2973 5559
rect 2973 5525 3007 5559
rect 3007 5525 3016 5559
rect 2964 5516 3016 5525
rect 4252 5516 4304 5568
rect 4712 5559 4764 5568
rect 4712 5525 4721 5559
rect 4721 5525 4755 5559
rect 4755 5525 4764 5559
rect 4712 5516 4764 5525
rect 4804 5516 4856 5568
rect 6000 5584 6052 5636
rect 7932 5584 7984 5636
rect 5540 5516 5592 5568
rect 6276 5516 6328 5568
rect 7380 5516 7432 5568
rect 7656 5516 7708 5568
rect 12072 5584 12124 5636
rect 12348 5584 12400 5636
rect 12440 5584 12492 5636
rect 13176 5652 13228 5704
rect 14372 5695 14424 5704
rect 14372 5661 14381 5695
rect 14381 5661 14415 5695
rect 14415 5661 14424 5695
rect 14372 5652 14424 5661
rect 15384 5584 15436 5636
rect 16488 5652 16540 5704
rect 17408 5720 17460 5772
rect 18052 5865 18061 5899
rect 18061 5865 18095 5899
rect 18095 5865 18104 5899
rect 18052 5856 18104 5865
rect 18236 5788 18288 5840
rect 9312 5559 9364 5568
rect 9312 5525 9321 5559
rect 9321 5525 9355 5559
rect 9355 5525 9364 5559
rect 9588 5559 9640 5568
rect 9312 5516 9364 5525
rect 9588 5525 9597 5559
rect 9597 5525 9631 5559
rect 9631 5525 9640 5559
rect 9588 5516 9640 5525
rect 10324 5516 10376 5568
rect 11612 5516 11664 5568
rect 13912 5516 13964 5568
rect 17224 5695 17276 5704
rect 17224 5661 17233 5695
rect 17233 5661 17267 5695
rect 17267 5661 17276 5695
rect 17224 5652 17276 5661
rect 18512 5627 18564 5636
rect 18512 5593 18521 5627
rect 18521 5593 18555 5627
rect 18555 5593 18564 5627
rect 18512 5584 18564 5593
rect 16764 5516 16816 5568
rect 17960 5516 18012 5568
rect 3947 5414 3999 5466
rect 4011 5414 4063 5466
rect 4075 5414 4127 5466
rect 4139 5414 4191 5466
rect 9878 5414 9930 5466
rect 9942 5414 9994 5466
rect 10006 5414 10058 5466
rect 10070 5414 10122 5466
rect 15808 5414 15860 5466
rect 15872 5414 15924 5466
rect 15936 5414 15988 5466
rect 16000 5414 16052 5466
rect 2872 5355 2924 5364
rect 2872 5321 2881 5355
rect 2881 5321 2915 5355
rect 2915 5321 2924 5355
rect 2872 5312 2924 5321
rect 3424 5312 3476 5364
rect 4804 5244 4856 5296
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 2964 5176 3016 5228
rect 3516 5219 3568 5228
rect 3516 5185 3525 5219
rect 3525 5185 3559 5219
rect 3559 5185 3568 5219
rect 3516 5176 3568 5185
rect 4988 5312 5040 5364
rect 5264 5312 5316 5364
rect 9312 5312 9364 5364
rect 11244 5355 11296 5364
rect 11244 5321 11253 5355
rect 11253 5321 11287 5355
rect 11287 5321 11296 5355
rect 11244 5312 11296 5321
rect 11336 5312 11388 5364
rect 14648 5312 14700 5364
rect 15108 5312 15160 5364
rect 15384 5312 15436 5364
rect 15660 5355 15712 5364
rect 15660 5321 15669 5355
rect 15669 5321 15703 5355
rect 15703 5321 15712 5355
rect 15660 5312 15712 5321
rect 16120 5312 16172 5364
rect 16304 5312 16356 5364
rect 11888 5244 11940 5296
rect 16396 5244 16448 5296
rect 9312 5176 9364 5228
rect 1952 5083 2004 5092
rect 1952 5049 1961 5083
rect 1961 5049 1995 5083
rect 1995 5049 2004 5083
rect 1952 5040 2004 5049
rect 4712 5108 4764 5160
rect 6276 5151 6328 5160
rect 6276 5117 6285 5151
rect 6285 5117 6319 5151
rect 6319 5117 6328 5151
rect 6276 5108 6328 5117
rect 7748 5108 7800 5160
rect 2872 5040 2924 5092
rect 3700 5040 3752 5092
rect 4988 5040 5040 5092
rect 5448 5040 5500 5092
rect 7380 5040 7432 5092
rect 8576 5108 8628 5160
rect 10600 5176 10652 5228
rect 13268 5176 13320 5228
rect 14004 5219 14056 5228
rect 14004 5185 14013 5219
rect 14013 5185 14047 5219
rect 14047 5185 14056 5219
rect 14004 5176 14056 5185
rect 10968 5151 11020 5160
rect 8760 5040 8812 5092
rect 10968 5117 10977 5151
rect 10977 5117 11011 5151
rect 11011 5117 11020 5151
rect 10968 5108 11020 5117
rect 12532 5108 12584 5160
rect 13820 5151 13872 5160
rect 13820 5117 13829 5151
rect 13829 5117 13863 5151
rect 13863 5117 13872 5151
rect 13820 5108 13872 5117
rect 14096 5108 14148 5160
rect 14648 5108 14700 5160
rect 15292 5108 15344 5160
rect 15660 5108 15712 5160
rect 10784 5040 10836 5092
rect 1860 5015 1912 5024
rect 1860 4981 1869 5015
rect 1869 4981 1903 5015
rect 1903 4981 1912 5015
rect 1860 4972 1912 4981
rect 2136 5015 2188 5024
rect 2136 4981 2145 5015
rect 2145 4981 2179 5015
rect 2179 4981 2188 5015
rect 2136 4972 2188 4981
rect 4160 5015 4212 5024
rect 4160 4981 4169 5015
rect 4169 4981 4203 5015
rect 4203 4981 4212 5015
rect 4160 4972 4212 4981
rect 6092 4972 6144 5024
rect 6184 4972 6236 5024
rect 6552 4972 6604 5024
rect 8668 4972 8720 5024
rect 11060 4972 11112 5024
rect 15200 5040 15252 5092
rect 15752 5040 15804 5092
rect 16304 5176 16356 5228
rect 16488 5176 16540 5228
rect 17224 5176 17276 5228
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 16672 5108 16724 5160
rect 17132 5108 17184 5160
rect 17868 5151 17920 5160
rect 17868 5117 17877 5151
rect 17877 5117 17911 5151
rect 17911 5117 17920 5151
rect 17868 5108 17920 5117
rect 18604 5108 18656 5160
rect 16764 5040 16816 5092
rect 16856 5040 16908 5092
rect 12716 4972 12768 5024
rect 13820 4972 13872 5024
rect 14004 4972 14056 5024
rect 15108 5015 15160 5024
rect 15108 4981 15117 5015
rect 15117 4981 15151 5015
rect 15151 4981 15160 5015
rect 15108 4972 15160 4981
rect 16120 4972 16172 5024
rect 18236 4972 18288 5024
rect 6912 4870 6964 4922
rect 6976 4870 7028 4922
rect 7040 4870 7092 4922
rect 7104 4870 7156 4922
rect 12843 4870 12895 4922
rect 12907 4870 12959 4922
rect 12971 4870 13023 4922
rect 13035 4870 13087 4922
rect 1952 4768 2004 4820
rect 2872 4811 2924 4820
rect 2872 4777 2881 4811
rect 2881 4777 2915 4811
rect 2915 4777 2924 4811
rect 2872 4768 2924 4777
rect 3792 4768 3844 4820
rect 4160 4811 4212 4820
rect 4160 4777 4169 4811
rect 4169 4777 4203 4811
rect 4203 4777 4212 4811
rect 4160 4768 4212 4777
rect 4528 4811 4580 4820
rect 4528 4777 4537 4811
rect 4537 4777 4571 4811
rect 4571 4777 4580 4811
rect 4528 4768 4580 4777
rect 4988 4811 5040 4820
rect 4988 4777 4997 4811
rect 4997 4777 5031 4811
rect 5031 4777 5040 4811
rect 4988 4768 5040 4777
rect 5080 4768 5132 4820
rect 2136 4700 2188 4752
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 6552 4700 6604 4752
rect 3792 4632 3844 4684
rect 4712 4632 4764 4684
rect 3148 4428 3200 4480
rect 6000 4632 6052 4684
rect 9496 4768 9548 4820
rect 9588 4768 9640 4820
rect 10784 4700 10836 4752
rect 11244 4700 11296 4752
rect 11612 4700 11664 4752
rect 12532 4768 12584 4820
rect 12716 4768 12768 4820
rect 13176 4700 13228 4752
rect 13360 4768 13412 4820
rect 14648 4700 14700 4752
rect 5172 4564 5224 4616
rect 6276 4607 6328 4616
rect 5540 4496 5592 4548
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 5816 4539 5868 4548
rect 5816 4505 5825 4539
rect 5825 4505 5859 4539
rect 5859 4505 5868 4539
rect 5816 4496 5868 4505
rect 6092 4496 6144 4548
rect 6552 4564 6604 4616
rect 10600 4564 10652 4616
rect 13820 4632 13872 4684
rect 7564 4496 7616 4548
rect 10416 4428 10468 4480
rect 10784 4428 10836 4480
rect 10968 4428 11020 4480
rect 11520 4428 11572 4480
rect 12440 4564 12492 4616
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 14464 4632 14516 4684
rect 15108 4632 15160 4684
rect 15752 4632 15804 4684
rect 16304 4632 16356 4684
rect 16580 4768 16632 4820
rect 17040 4811 17092 4820
rect 17040 4777 17049 4811
rect 17049 4777 17083 4811
rect 17083 4777 17092 4811
rect 17040 4768 17092 4777
rect 18788 4768 18840 4820
rect 16488 4700 16540 4752
rect 17316 4700 17368 4752
rect 17960 4743 18012 4752
rect 17960 4709 17969 4743
rect 17969 4709 18003 4743
rect 18003 4709 18012 4743
rect 17960 4700 18012 4709
rect 18052 4700 18104 4752
rect 16948 4632 17000 4684
rect 18144 4675 18196 4684
rect 18144 4641 18153 4675
rect 18153 4641 18187 4675
rect 18187 4641 18196 4675
rect 18144 4632 18196 4641
rect 13912 4496 13964 4548
rect 15292 4496 15344 4548
rect 15752 4496 15804 4548
rect 17224 4607 17276 4616
rect 17224 4573 17233 4607
rect 17233 4573 17267 4607
rect 17267 4573 17276 4607
rect 17224 4564 17276 4573
rect 17040 4496 17092 4548
rect 18512 4539 18564 4548
rect 18512 4505 18521 4539
rect 18521 4505 18555 4539
rect 18555 4505 18564 4539
rect 18512 4496 18564 4505
rect 11888 4428 11940 4480
rect 13452 4428 13504 4480
rect 14280 4428 14332 4480
rect 15200 4428 15252 4480
rect 15384 4471 15436 4480
rect 15384 4437 15393 4471
rect 15393 4437 15427 4471
rect 15427 4437 15436 4471
rect 15384 4428 15436 4437
rect 16580 4471 16632 4480
rect 16580 4437 16589 4471
rect 16589 4437 16623 4471
rect 16623 4437 16632 4471
rect 16580 4428 16632 4437
rect 17960 4428 18012 4480
rect 3947 4326 3999 4378
rect 4011 4326 4063 4378
rect 4075 4326 4127 4378
rect 4139 4326 4191 4378
rect 9878 4326 9930 4378
rect 9942 4326 9994 4378
rect 10006 4326 10058 4378
rect 10070 4326 10122 4378
rect 15808 4326 15860 4378
rect 15872 4326 15924 4378
rect 15936 4326 15988 4378
rect 16000 4326 16052 4378
rect 2688 4224 2740 4276
rect 3608 4224 3660 4276
rect 4528 4224 4580 4276
rect 2504 4020 2556 4072
rect 5448 4224 5500 4276
rect 6276 4224 6328 4276
rect 6552 4224 6604 4276
rect 8760 4267 8812 4276
rect 8760 4233 8769 4267
rect 8769 4233 8803 4267
rect 8803 4233 8812 4267
rect 8760 4224 8812 4233
rect 10600 4224 10652 4276
rect 11152 4224 11204 4276
rect 5172 4156 5224 4208
rect 7380 4131 7432 4140
rect 7380 4097 7389 4131
rect 7389 4097 7423 4131
rect 7423 4097 7432 4131
rect 7380 4088 7432 4097
rect 9404 4088 9456 4140
rect 12348 4224 12400 4276
rect 15108 4224 15160 4276
rect 15568 4199 15620 4208
rect 15568 4165 15577 4199
rect 15577 4165 15611 4199
rect 15611 4165 15620 4199
rect 15568 4156 15620 4165
rect 16120 4224 16172 4276
rect 16948 4224 17000 4276
rect 15936 4156 15988 4208
rect 1952 3995 2004 4004
rect 1952 3961 1961 3995
rect 1961 3961 1995 3995
rect 1995 3961 2004 3995
rect 1952 3952 2004 3961
rect 5172 4020 5224 4072
rect 6736 4020 6788 4072
rect 8852 4063 8904 4072
rect 1492 3927 1544 3936
rect 1492 3893 1501 3927
rect 1501 3893 1535 3927
rect 1535 3893 1544 3927
rect 1492 3884 1544 3893
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 2228 3927 2280 3936
rect 2228 3893 2237 3927
rect 2237 3893 2271 3927
rect 2271 3893 2280 3927
rect 2228 3884 2280 3893
rect 2780 3927 2832 3936
rect 2780 3893 2789 3927
rect 2789 3893 2823 3927
rect 2823 3893 2832 3927
rect 4620 3952 4672 4004
rect 2780 3884 2832 3893
rect 3608 3884 3660 3936
rect 3792 3884 3844 3936
rect 8024 3952 8076 4004
rect 8852 4029 8861 4063
rect 8861 4029 8895 4063
rect 8895 4029 8904 4063
rect 8852 4020 8904 4029
rect 9496 4063 9548 4072
rect 9496 4029 9505 4063
rect 9505 4029 9539 4063
rect 9539 4029 9548 4063
rect 9496 4020 9548 4029
rect 10324 4020 10376 4072
rect 11520 4063 11572 4072
rect 10416 3952 10468 4004
rect 11520 4029 11529 4063
rect 11529 4029 11563 4063
rect 11563 4029 11572 4063
rect 11520 4020 11572 4029
rect 11704 4088 11756 4140
rect 12716 4088 12768 4140
rect 14832 4131 14884 4140
rect 11980 4020 12032 4072
rect 14832 4097 14841 4131
rect 14841 4097 14875 4131
rect 14875 4097 14884 4131
rect 14832 4088 14884 4097
rect 15384 4088 15436 4140
rect 15660 4088 15712 4140
rect 17316 4088 17368 4140
rect 18052 4088 18104 4140
rect 14004 4020 14056 4072
rect 15752 4063 15804 4072
rect 15752 4029 15761 4063
rect 15761 4029 15795 4063
rect 15795 4029 15804 4063
rect 15752 4020 15804 4029
rect 15936 4063 15988 4072
rect 15936 4029 15945 4063
rect 15945 4029 15979 4063
rect 15979 4029 15988 4063
rect 15936 4020 15988 4029
rect 16764 4020 16816 4072
rect 16948 4063 17000 4072
rect 16948 4029 16957 4063
rect 16957 4029 16991 4063
rect 16991 4029 17000 4063
rect 16948 4020 17000 4029
rect 17132 4020 17184 4072
rect 12440 3995 12492 4004
rect 12440 3961 12449 3995
rect 12449 3961 12483 3995
rect 12483 3961 12492 3995
rect 12440 3952 12492 3961
rect 13636 3952 13688 4004
rect 4804 3884 4856 3936
rect 6000 3884 6052 3936
rect 7748 3884 7800 3936
rect 8116 3884 8168 3936
rect 10232 3884 10284 3936
rect 10600 3884 10652 3936
rect 11336 3884 11388 3936
rect 11612 3884 11664 3936
rect 11888 3927 11940 3936
rect 11888 3893 11897 3927
rect 11897 3893 11931 3927
rect 11931 3893 11940 3927
rect 11888 3884 11940 3893
rect 13176 3884 13228 3936
rect 13360 3927 13412 3936
rect 13360 3893 13369 3927
rect 13369 3893 13403 3927
rect 13403 3893 13412 3927
rect 13360 3884 13412 3893
rect 14280 3995 14332 4004
rect 14280 3961 14289 3995
rect 14289 3961 14323 3995
rect 14323 3961 14332 3995
rect 14280 3952 14332 3961
rect 15200 3952 15252 4004
rect 18236 4020 18288 4072
rect 15016 3884 15068 3936
rect 18144 3995 18196 4004
rect 17132 3927 17184 3936
rect 17132 3893 17141 3927
rect 17141 3893 17175 3927
rect 17175 3893 17184 3927
rect 17132 3884 17184 3893
rect 17316 3884 17368 3936
rect 18144 3961 18153 3995
rect 18153 3961 18187 3995
rect 18187 3961 18196 3995
rect 18144 3952 18196 3961
rect 18512 3995 18564 4004
rect 18512 3961 18521 3995
rect 18521 3961 18555 3995
rect 18555 3961 18564 3995
rect 18512 3952 18564 3961
rect 19156 3884 19208 3936
rect 6912 3782 6964 3834
rect 6976 3782 7028 3834
rect 7040 3782 7092 3834
rect 7104 3782 7156 3834
rect 12843 3782 12895 3834
rect 12907 3782 12959 3834
rect 12971 3782 13023 3834
rect 13035 3782 13087 3834
rect 1952 3680 2004 3732
rect 3608 3680 3660 3732
rect 8024 3723 8076 3732
rect 1952 3587 2004 3596
rect 1952 3553 1961 3587
rect 1961 3553 1995 3587
rect 1995 3553 2004 3587
rect 1952 3544 2004 3553
rect 2688 3587 2740 3596
rect 2688 3553 2697 3587
rect 2697 3553 2731 3587
rect 2731 3553 2740 3587
rect 2688 3544 2740 3553
rect 2872 3476 2924 3528
rect 3148 3544 3200 3596
rect 5264 3544 5316 3596
rect 6184 3544 6236 3596
rect 6552 3612 6604 3664
rect 7472 3544 7524 3596
rect 8024 3689 8033 3723
rect 8033 3689 8067 3723
rect 8067 3689 8076 3723
rect 8024 3680 8076 3689
rect 8852 3680 8904 3732
rect 7932 3612 7984 3664
rect 8208 3544 8260 3596
rect 5172 3519 5224 3528
rect 5172 3485 5181 3519
rect 5181 3485 5215 3519
rect 5215 3485 5224 3519
rect 5172 3476 5224 3485
rect 4988 3408 5040 3460
rect 1400 3340 1452 3392
rect 1860 3383 1912 3392
rect 1860 3349 1869 3383
rect 1869 3349 1903 3383
rect 1903 3349 1912 3383
rect 1860 3340 1912 3349
rect 2228 3383 2280 3392
rect 2228 3349 2237 3383
rect 2237 3349 2271 3383
rect 2271 3349 2280 3383
rect 2228 3340 2280 3349
rect 3332 3383 3384 3392
rect 3332 3349 3341 3383
rect 3341 3349 3375 3383
rect 3375 3349 3384 3383
rect 3700 3383 3752 3392
rect 3332 3340 3384 3349
rect 3700 3349 3709 3383
rect 3709 3349 3743 3383
rect 3743 3349 3752 3383
rect 3700 3340 3752 3349
rect 4804 3340 4856 3392
rect 6552 3451 6604 3460
rect 6552 3417 6561 3451
rect 6561 3417 6595 3451
rect 6595 3417 6604 3451
rect 6552 3408 6604 3417
rect 7840 3476 7892 3528
rect 10600 3612 10652 3664
rect 10784 3544 10836 3596
rect 12348 3612 12400 3664
rect 12532 3612 12584 3664
rect 13912 3680 13964 3732
rect 15660 3680 15712 3732
rect 16948 3680 17000 3732
rect 17132 3680 17184 3732
rect 17040 3612 17092 3664
rect 17960 3655 18012 3664
rect 17960 3621 17969 3655
rect 17969 3621 18003 3655
rect 18003 3621 18012 3655
rect 17960 3612 18012 3621
rect 10968 3544 11020 3596
rect 11612 3587 11664 3596
rect 11612 3553 11621 3587
rect 11621 3553 11655 3587
rect 11655 3553 11664 3587
rect 11612 3544 11664 3553
rect 11704 3587 11756 3596
rect 11704 3553 11713 3587
rect 11713 3553 11747 3587
rect 11747 3553 11756 3587
rect 11704 3544 11756 3553
rect 11888 3544 11940 3596
rect 11060 3476 11112 3528
rect 11980 3519 12032 3528
rect 7748 3408 7800 3460
rect 11428 3451 11480 3460
rect 7380 3340 7432 3392
rect 8300 3340 8352 3392
rect 9680 3340 9732 3392
rect 9772 3340 9824 3392
rect 10416 3383 10468 3392
rect 10416 3349 10425 3383
rect 10425 3349 10459 3383
rect 10459 3349 10468 3383
rect 10416 3340 10468 3349
rect 11060 3383 11112 3392
rect 11060 3349 11069 3383
rect 11069 3349 11103 3383
rect 11103 3349 11112 3383
rect 11060 3340 11112 3349
rect 11428 3417 11437 3451
rect 11437 3417 11471 3451
rect 11471 3417 11480 3451
rect 11428 3408 11480 3417
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 12440 3476 12492 3528
rect 13360 3544 13412 3596
rect 13912 3587 13964 3596
rect 13912 3553 13921 3587
rect 13921 3553 13955 3587
rect 13955 3553 13964 3587
rect 13912 3544 13964 3553
rect 12072 3408 12124 3460
rect 12164 3408 12216 3460
rect 13820 3476 13872 3528
rect 14464 3587 14516 3596
rect 14464 3553 14508 3587
rect 14508 3553 14516 3587
rect 14740 3587 14792 3596
rect 14464 3544 14516 3553
rect 14740 3553 14749 3587
rect 14749 3553 14783 3587
rect 14783 3553 14792 3587
rect 14740 3544 14792 3553
rect 15016 3587 15068 3596
rect 15016 3553 15025 3587
rect 15025 3553 15059 3587
rect 15059 3553 15068 3587
rect 15016 3544 15068 3553
rect 15200 3476 15252 3528
rect 13636 3408 13688 3460
rect 15660 3544 15712 3596
rect 16304 3544 16356 3596
rect 16396 3544 16448 3596
rect 15568 3408 15620 3460
rect 11612 3340 11664 3392
rect 11980 3340 12032 3392
rect 13268 3340 13320 3392
rect 13728 3383 13780 3392
rect 13728 3349 13737 3383
rect 13737 3349 13771 3383
rect 13771 3349 13780 3383
rect 13728 3340 13780 3349
rect 19616 3544 19668 3596
rect 17224 3408 17276 3460
rect 18604 3476 18656 3528
rect 18144 3451 18196 3460
rect 18144 3417 18153 3451
rect 18153 3417 18187 3451
rect 18187 3417 18196 3451
rect 18144 3408 18196 3417
rect 16396 3383 16448 3392
rect 16396 3349 16405 3383
rect 16405 3349 16439 3383
rect 16439 3349 16448 3383
rect 16396 3340 16448 3349
rect 16672 3383 16724 3392
rect 16672 3349 16681 3383
rect 16681 3349 16715 3383
rect 16715 3349 16724 3383
rect 16672 3340 16724 3349
rect 17592 3340 17644 3392
rect 17868 3340 17920 3392
rect 3947 3238 3999 3290
rect 4011 3238 4063 3290
rect 4075 3238 4127 3290
rect 4139 3238 4191 3290
rect 9878 3238 9930 3290
rect 9942 3238 9994 3290
rect 10006 3238 10058 3290
rect 10070 3238 10122 3290
rect 15808 3238 15860 3290
rect 15872 3238 15924 3290
rect 15936 3238 15988 3290
rect 16000 3238 16052 3290
rect 1952 3136 2004 3188
rect 2964 3136 3016 3188
rect 3700 3136 3752 3188
rect 4620 3179 4672 3188
rect 4620 3145 4629 3179
rect 4629 3145 4663 3179
rect 4663 3145 4672 3179
rect 4620 3136 4672 3145
rect 6184 3136 6236 3188
rect 8024 3136 8076 3188
rect 1676 3068 1728 3120
rect 4160 3068 4212 3120
rect 2780 3000 2832 3052
rect 3056 3000 3108 3052
rect 2044 2932 2096 2984
rect 2136 2932 2188 2984
rect 1768 2907 1820 2916
rect 1768 2873 1777 2907
rect 1777 2873 1811 2907
rect 1811 2873 1820 2907
rect 1768 2864 1820 2873
rect 2320 2907 2372 2916
rect 2320 2873 2329 2907
rect 2329 2873 2363 2907
rect 2363 2873 2372 2907
rect 2320 2864 2372 2873
rect 2596 2932 2648 2984
rect 2964 2975 3016 2984
rect 2964 2941 2973 2975
rect 2973 2941 3007 2975
rect 3007 2941 3016 2975
rect 2964 2932 3016 2941
rect 3240 2975 3292 2984
rect 3240 2941 3249 2975
rect 3249 2941 3283 2975
rect 3283 2941 3292 2975
rect 3240 2932 3292 2941
rect 3700 3000 3752 3052
rect 5080 3068 5132 3120
rect 7472 3068 7524 3120
rect 8484 3068 8536 3120
rect 10416 3136 10468 3188
rect 9680 3068 9732 3120
rect 10140 3068 10192 3120
rect 10232 3068 10284 3120
rect 12532 3136 12584 3188
rect 12992 3136 13044 3188
rect 13820 3136 13872 3188
rect 6828 3000 6880 3052
rect 3792 2975 3844 2984
rect 3792 2941 3801 2975
rect 3801 2941 3835 2975
rect 3835 2941 3844 2975
rect 3792 2932 3844 2941
rect 4068 2975 4120 2984
rect 4068 2941 4077 2975
rect 4077 2941 4111 2975
rect 4111 2941 4120 2975
rect 4068 2932 4120 2941
rect 4344 2975 4396 2984
rect 4344 2941 4353 2975
rect 4353 2941 4387 2975
rect 4387 2941 4396 2975
rect 4344 2932 4396 2941
rect 4620 2932 4672 2984
rect 7288 3000 7340 3052
rect 7932 3000 7984 3052
rect 4252 2864 4304 2916
rect 7748 2932 7800 2984
rect 9404 2932 9456 2984
rect 9772 2932 9824 2984
rect 10416 3000 10468 3052
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 13728 3000 13780 3052
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 10600 2932 10652 2984
rect 10784 2975 10836 2984
rect 10784 2941 10793 2975
rect 10793 2941 10827 2975
rect 10827 2941 10836 2975
rect 10784 2932 10836 2941
rect 10876 2975 10928 2984
rect 10876 2941 10885 2975
rect 10885 2941 10919 2975
rect 10919 2941 10928 2975
rect 11060 2975 11112 2984
rect 10876 2932 10928 2941
rect 11060 2941 11069 2975
rect 11069 2941 11103 2975
rect 11103 2941 11112 2975
rect 11060 2932 11112 2941
rect 1308 2796 1360 2848
rect 2228 2839 2280 2848
rect 2228 2805 2237 2839
rect 2237 2805 2271 2839
rect 2271 2805 2280 2839
rect 2228 2796 2280 2805
rect 2504 2839 2556 2848
rect 2504 2805 2513 2839
rect 2513 2805 2547 2839
rect 2547 2805 2556 2839
rect 2504 2796 2556 2805
rect 3056 2839 3108 2848
rect 3056 2805 3065 2839
rect 3065 2805 3099 2839
rect 3099 2805 3108 2839
rect 3056 2796 3108 2805
rect 3148 2796 3200 2848
rect 3608 2839 3660 2848
rect 3608 2805 3617 2839
rect 3617 2805 3651 2839
rect 3651 2805 3660 2839
rect 3608 2796 3660 2805
rect 3884 2839 3936 2848
rect 3884 2805 3893 2839
rect 3893 2805 3927 2839
rect 3927 2805 3936 2839
rect 3884 2796 3936 2805
rect 4528 2839 4580 2848
rect 4528 2805 4537 2839
rect 4537 2805 4571 2839
rect 4571 2805 4580 2839
rect 4528 2796 4580 2805
rect 7840 2796 7892 2848
rect 8116 2839 8168 2848
rect 8116 2805 8125 2839
rect 8125 2805 8159 2839
rect 8159 2805 8168 2839
rect 8116 2796 8168 2805
rect 9680 2907 9732 2916
rect 9312 2839 9364 2848
rect 9312 2805 9321 2839
rect 9321 2805 9355 2839
rect 9355 2805 9364 2839
rect 9312 2796 9364 2805
rect 9680 2873 9689 2907
rect 9689 2873 9723 2907
rect 9723 2873 9732 2907
rect 9680 2864 9732 2873
rect 9772 2796 9824 2848
rect 11612 2864 11664 2916
rect 10600 2796 10652 2848
rect 12440 2907 12492 2916
rect 12440 2873 12449 2907
rect 12449 2873 12483 2907
rect 12483 2873 12492 2907
rect 12440 2864 12492 2873
rect 12808 2975 12860 2984
rect 12808 2941 12852 2975
rect 12852 2941 12860 2975
rect 12808 2932 12860 2941
rect 13268 2907 13320 2916
rect 13268 2873 13277 2907
rect 13277 2873 13311 2907
rect 13311 2873 13320 2907
rect 13268 2864 13320 2873
rect 15660 3136 15712 3188
rect 16488 3136 16540 3188
rect 16856 3136 16908 3188
rect 17132 3136 17184 3188
rect 17684 3136 17736 3188
rect 14740 3068 14792 3120
rect 16672 3068 16724 3120
rect 15476 3000 15528 3052
rect 15752 3043 15804 3052
rect 15752 3009 15761 3043
rect 15761 3009 15795 3043
rect 15795 3009 15804 3043
rect 15752 3000 15804 3009
rect 16396 3000 16448 3052
rect 16580 2975 16632 2984
rect 16580 2941 16589 2975
rect 16589 2941 16623 2975
rect 16623 2941 16632 2975
rect 16580 2932 16632 2941
rect 17132 2975 17184 2984
rect 17132 2941 17141 2975
rect 17141 2941 17175 2975
rect 17175 2941 17184 2975
rect 17132 2932 17184 2941
rect 17224 2932 17276 2984
rect 17776 3000 17828 3052
rect 14556 2864 14608 2916
rect 16488 2864 16540 2916
rect 16764 2907 16816 2916
rect 16764 2873 16773 2907
rect 16773 2873 16807 2907
rect 16807 2873 16816 2907
rect 16764 2864 16816 2873
rect 17776 2907 17828 2916
rect 17776 2873 17785 2907
rect 17785 2873 17819 2907
rect 17819 2873 17828 2907
rect 17776 2864 17828 2873
rect 17408 2796 17460 2848
rect 6912 2694 6964 2746
rect 6976 2694 7028 2746
rect 7040 2694 7092 2746
rect 7104 2694 7156 2746
rect 12843 2694 12895 2746
rect 12907 2694 12959 2746
rect 12971 2694 13023 2746
rect 13035 2694 13087 2746
rect 1584 2567 1636 2576
rect 1584 2533 1593 2567
rect 1593 2533 1627 2567
rect 1627 2533 1636 2567
rect 1584 2524 1636 2533
rect 3056 2592 3108 2644
rect 4160 2592 4212 2644
rect 5724 2592 5776 2644
rect 2596 2567 2648 2576
rect 2596 2533 2605 2567
rect 2605 2533 2639 2567
rect 2639 2533 2648 2567
rect 2596 2524 2648 2533
rect 3148 2524 3200 2576
rect 3608 2524 3660 2576
rect 3884 2524 3936 2576
rect 4436 2567 4488 2576
rect 4436 2533 4445 2567
rect 4445 2533 4479 2567
rect 4479 2533 4488 2567
rect 4436 2524 4488 2533
rect 4528 2524 4580 2576
rect 4988 2524 5040 2576
rect 6644 2524 6696 2576
rect 9772 2592 9824 2644
rect 7472 2567 7524 2576
rect 7472 2533 7481 2567
rect 7481 2533 7515 2567
rect 7515 2533 7524 2567
rect 7472 2524 7524 2533
rect 8116 2524 8168 2576
rect 8300 2567 8352 2576
rect 8300 2533 8309 2567
rect 8309 2533 8343 2567
rect 8343 2533 8352 2567
rect 8300 2524 8352 2533
rect 9220 2567 9272 2576
rect 9220 2533 9229 2567
rect 9229 2533 9263 2567
rect 9263 2533 9272 2567
rect 9220 2524 9272 2533
rect 10140 2567 10192 2576
rect 10140 2533 10149 2567
rect 10149 2533 10183 2567
rect 10183 2533 10192 2567
rect 10140 2524 10192 2533
rect 10508 2567 10560 2576
rect 10508 2533 10517 2567
rect 10517 2533 10551 2567
rect 10551 2533 10560 2567
rect 10508 2524 10560 2533
rect 10968 2592 11020 2644
rect 12440 2592 12492 2644
rect 11336 2524 11388 2576
rect 12072 2567 12124 2576
rect 12072 2533 12081 2567
rect 12081 2533 12115 2567
rect 12115 2533 12124 2567
rect 12072 2524 12124 2533
rect 13176 2567 13228 2576
rect 13176 2533 13185 2567
rect 13185 2533 13219 2567
rect 13219 2533 13228 2567
rect 13176 2524 13228 2533
rect 13452 2524 13504 2576
rect 14188 2567 14240 2576
rect 14188 2533 14197 2567
rect 14197 2533 14231 2567
rect 14231 2533 14240 2567
rect 14188 2524 14240 2533
rect 3424 2456 3476 2508
rect 3700 2499 3752 2508
rect 3700 2465 3709 2499
rect 3709 2465 3743 2499
rect 3743 2465 3752 2499
rect 3700 2456 3752 2465
rect 4252 2456 4304 2508
rect 1124 2388 1176 2440
rect 204 2320 256 2372
rect 2688 2363 2740 2372
rect 2688 2329 2697 2363
rect 2697 2329 2731 2363
rect 2731 2329 2740 2363
rect 2688 2320 2740 2329
rect 3148 2363 3200 2372
rect 3148 2329 3157 2363
rect 3157 2329 3191 2363
rect 3191 2329 3200 2363
rect 3148 2320 3200 2329
rect 3608 2320 3660 2372
rect 4252 2363 4304 2372
rect 4252 2329 4261 2363
rect 4261 2329 4295 2363
rect 4295 2329 4304 2363
rect 4252 2320 4304 2329
rect 5172 2320 5224 2372
rect 664 2252 716 2304
rect 2872 2252 2924 2304
rect 5632 2456 5684 2508
rect 7288 2456 7340 2508
rect 9312 2456 9364 2508
rect 15200 2592 15252 2644
rect 15292 2567 15344 2576
rect 15292 2533 15301 2567
rect 15301 2533 15335 2567
rect 15335 2533 15344 2567
rect 15292 2524 15344 2533
rect 16212 2524 16264 2576
rect 16488 2524 16540 2576
rect 16948 2567 17000 2576
rect 16948 2533 16957 2567
rect 16957 2533 16991 2567
rect 16991 2533 17000 2567
rect 16948 2524 17000 2533
rect 18052 2524 18104 2576
rect 16856 2456 16908 2508
rect 18420 2456 18472 2508
rect 6644 2388 6696 2440
rect 11428 2388 11480 2440
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 16672 2388 16724 2440
rect 17500 2388 17552 2440
rect 17684 2388 17736 2440
rect 6184 2320 6236 2372
rect 7104 2320 7156 2372
rect 7656 2363 7708 2372
rect 7656 2329 7665 2363
rect 7665 2329 7699 2363
rect 7699 2329 7708 2363
rect 7656 2320 7708 2329
rect 8116 2363 8168 2372
rect 8116 2329 8125 2363
rect 8125 2329 8159 2363
rect 8159 2329 8168 2363
rect 8116 2320 8168 2329
rect 8668 2363 8720 2372
rect 8668 2329 8677 2363
rect 8677 2329 8711 2363
rect 8711 2329 8720 2363
rect 8668 2320 8720 2329
rect 15568 2320 15620 2372
rect 15660 2320 15712 2372
rect 17776 2363 17828 2372
rect 17776 2329 17785 2363
rect 17785 2329 17819 2363
rect 17819 2329 17828 2363
rect 17776 2320 17828 2329
rect 17868 2320 17920 2372
rect 8024 2252 8076 2304
rect 9128 2252 9180 2304
rect 13912 2252 13964 2304
rect 16120 2252 16172 2304
rect 17684 2252 17736 2304
rect 3947 2150 3999 2202
rect 4011 2150 4063 2202
rect 4075 2150 4127 2202
rect 4139 2150 4191 2202
rect 9878 2150 9930 2202
rect 9942 2150 9994 2202
rect 10006 2150 10058 2202
rect 10070 2150 10122 2202
rect 15808 2150 15860 2202
rect 15872 2150 15924 2202
rect 15936 2150 15988 2202
rect 16000 2150 16052 2202
rect 3424 2048 3476 2100
rect 10692 2048 10744 2100
rect 13176 1708 13228 1760
rect 13912 1708 13964 1760
rect 16764 1096 16816 1148
rect 18144 1096 18196 1148
<< metal2 >>
rect 294 16400 350 17200
rect 938 16400 994 17200
rect 1582 16400 1638 17200
rect 2226 16400 2282 17200
rect 2870 16400 2926 17200
rect 3146 16416 3202 16425
rect 308 15162 336 16400
rect 296 15156 348 15162
rect 296 15098 348 15104
rect 952 13802 980 16400
rect 1596 15178 1624 16400
rect 1596 15150 1716 15178
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1596 14618 1624 14962
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1490 14512 1546 14521
rect 1490 14447 1492 14456
rect 1544 14447 1546 14456
rect 1492 14418 1544 14424
rect 940 13796 992 13802
rect 940 13738 992 13744
rect 1492 13796 1544 13802
rect 1492 13738 1544 13744
rect 1504 13394 1532 13738
rect 1688 13734 1716 15150
rect 1952 14884 2004 14890
rect 1952 14826 2004 14832
rect 1858 14784 1914 14793
rect 1858 14719 1914 14728
rect 1872 14550 1900 14719
rect 1964 14618 1992 14826
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1860 14544 1912 14550
rect 1860 14486 1912 14492
rect 2240 14006 2268 16400
rect 2594 16008 2650 16017
rect 2594 15943 2650 15952
rect 2608 14482 2636 15943
rect 2778 15600 2834 15609
rect 2778 15535 2834 15544
rect 2688 15088 2740 15094
rect 2688 15030 2740 15036
rect 2700 14618 2728 15030
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2792 14550 2820 15535
rect 2780 14544 2832 14550
rect 2780 14486 2832 14492
rect 2596 14476 2648 14482
rect 2596 14418 2648 14424
rect 2608 14278 2636 14418
rect 2780 14340 2832 14346
rect 2780 14282 2832 14288
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 2792 14090 2820 14282
rect 2700 14062 2820 14090
rect 2228 14000 2280 14006
rect 2228 13942 2280 13948
rect 2594 13968 2650 13977
rect 2594 13903 2650 13912
rect 1676 13728 1728 13734
rect 1676 13670 1728 13676
rect 1858 13560 1914 13569
rect 2608 13530 2636 13903
rect 2700 13818 2728 14062
rect 2884 14006 2912 16400
rect 3514 16400 3570 17200
rect 3790 16824 3846 16833
rect 3790 16759 3846 16768
rect 3146 16351 3202 16360
rect 2962 15192 3018 15201
rect 2962 15127 3018 15136
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 2872 13864 2924 13870
rect 2700 13790 2820 13818
rect 2872 13806 2924 13812
rect 1858 13495 1914 13504
rect 2596 13524 2648 13530
rect 1872 13462 1900 13495
rect 2596 13466 2648 13472
rect 1860 13456 1912 13462
rect 1860 13398 1912 13404
rect 2608 13394 2636 13466
rect 1492 13388 1544 13394
rect 1492 13330 1544 13336
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 1504 13161 1532 13330
rect 2148 13297 2176 13330
rect 2134 13288 2190 13297
rect 1676 13252 1728 13258
rect 2134 13223 2190 13232
rect 1676 13194 1728 13200
rect 1490 13152 1546 13161
rect 1490 13087 1546 13096
rect 1584 12912 1636 12918
rect 1584 12854 1636 12860
rect 1492 12776 1544 12782
rect 1596 12753 1624 12854
rect 1492 12718 1544 12724
rect 1582 12744 1638 12753
rect 1504 12345 1532 12718
rect 1582 12679 1584 12688
rect 1636 12679 1638 12688
rect 1584 12650 1636 12656
rect 1490 12336 1546 12345
rect 1400 12300 1452 12306
rect 1490 12271 1546 12280
rect 1400 12242 1452 12248
rect 1412 11393 1440 12242
rect 1490 11792 1546 11801
rect 1490 11727 1546 11736
rect 1504 11694 1532 11727
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1398 11384 1454 11393
rect 1398 11319 1454 11328
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1412 10577 1440 11154
rect 1504 10985 1532 11630
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1490 10976 1546 10985
rect 1490 10911 1546 10920
rect 1596 10713 1624 11494
rect 1688 10985 1716 13194
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 1964 12753 1992 13126
rect 2044 12776 2096 12782
rect 1950 12744 2006 12753
rect 2044 12718 2096 12724
rect 1950 12679 2006 12688
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1674 10976 1730 10985
rect 1674 10911 1730 10920
rect 1780 10826 1808 12582
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1872 11937 1900 12242
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1858 11928 1914 11937
rect 1964 11898 1992 12038
rect 1858 11863 1914 11872
rect 1952 11892 2004 11898
rect 1952 11834 2004 11840
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1688 10798 1808 10826
rect 1582 10704 1638 10713
rect 1582 10639 1638 10648
rect 1398 10568 1454 10577
rect 1398 10503 1454 10512
rect 1492 10532 1544 10538
rect 1492 10474 1544 10480
rect 1504 10169 1532 10474
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1490 10160 1546 10169
rect 1490 10095 1546 10104
rect 1400 9920 1452 9926
rect 1400 9862 1452 9868
rect 1412 9042 1440 9862
rect 1596 9722 1624 10406
rect 1688 10248 1716 10798
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 1780 10470 1808 10610
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1872 10266 1900 10950
rect 1964 10266 1992 11494
rect 1860 10260 1912 10266
rect 1688 10220 1808 10248
rect 1584 9716 1636 9722
rect 1584 9658 1636 9664
rect 1492 9444 1544 9450
rect 1492 9386 1544 9392
rect 1504 9353 1532 9386
rect 1584 9376 1636 9382
rect 1490 9344 1546 9353
rect 1584 9318 1636 9324
rect 1490 9279 1546 9288
rect 1596 9110 1624 9318
rect 1584 9104 1636 9110
rect 1584 9046 1636 9052
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1412 8945 1440 8978
rect 1398 8936 1454 8945
rect 1688 8922 1716 8978
rect 1398 8871 1454 8880
rect 1596 8894 1716 8922
rect 1596 8294 1624 8894
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 1492 7744 1544 7750
rect 1490 7712 1492 7721
rect 1544 7712 1546 7721
rect 1490 7647 1546 7656
rect 1596 7410 1624 8230
rect 1780 7857 1808 10220
rect 1860 10202 1912 10208
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 2056 10146 2084 12718
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 2148 11694 2176 12582
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2240 11370 2268 13126
rect 2700 12986 2728 13330
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2608 12170 2636 12786
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2412 12164 2464 12170
rect 2412 12106 2464 12112
rect 2596 12164 2648 12170
rect 2596 12106 2648 12112
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2332 11762 2360 12038
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2148 11342 2268 11370
rect 2148 10742 2176 11342
rect 2424 11218 2452 12106
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2516 11558 2544 11698
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2240 10810 2268 11154
rect 2516 11150 2544 11494
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2136 10736 2188 10742
rect 2136 10678 2188 10684
rect 2148 10606 2176 10678
rect 2136 10600 2188 10606
rect 2136 10542 2188 10548
rect 2332 10266 2360 11086
rect 2502 10976 2558 10985
rect 2502 10911 2558 10920
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2056 10118 2452 10146
rect 2134 9616 2190 9625
rect 2134 9551 2190 9560
rect 2148 9518 2176 9551
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 1952 9376 2004 9382
rect 1950 9344 1952 9353
rect 2136 9376 2188 9382
rect 2004 9344 2006 9353
rect 2136 9318 2188 9324
rect 1950 9279 2006 9288
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1872 8430 1900 8910
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1858 8120 1914 8129
rect 1858 8055 1860 8064
rect 1912 8055 1914 8064
rect 1860 8026 1912 8032
rect 2148 7954 2176 9318
rect 2424 9042 2452 10118
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 1766 7848 1822 7857
rect 1766 7783 1822 7792
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1400 7336 1452 7342
rect 1398 7304 1400 7313
rect 1452 7304 1454 7313
rect 1398 7239 1454 7248
rect 1766 6896 1822 6905
rect 1766 6831 1768 6840
rect 1820 6831 1822 6840
rect 1768 6802 1820 6808
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1504 6497 1532 6598
rect 1490 6488 1546 6497
rect 1490 6423 1546 6432
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1492 6112 1544 6118
rect 1490 6080 1492 6089
rect 1544 6080 1546 6089
rect 1490 6015 1546 6024
rect 1964 5914 1992 6190
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 1492 5568 1544 5574
rect 1490 5536 1492 5545
rect 1584 5568 1636 5574
rect 1544 5536 1546 5545
rect 1584 5510 1636 5516
rect 1490 5471 1546 5480
rect 1400 5160 1452 5166
rect 1398 5128 1400 5137
rect 1452 5128 1454 5137
rect 1398 5063 1454 5072
rect 1398 4720 1454 4729
rect 1398 4655 1400 4664
rect 1452 4655 1454 4664
rect 1400 4626 1452 4632
rect 1492 3936 1544 3942
rect 1492 3878 1544 3884
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 1308 2848 1360 2854
rect 1308 2790 1360 2796
rect 1124 2440 1176 2446
rect 1124 2382 1176 2388
rect 204 2372 256 2378
rect 204 2314 256 2320
rect 216 800 244 2314
rect 664 2304 716 2310
rect 664 2246 716 2252
rect 676 800 704 2246
rect 1136 800 1164 2382
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1320 649 1348 2790
rect 1412 1465 1440 3334
rect 1504 2689 1532 3878
rect 1490 2680 1546 2689
rect 1490 2615 1546 2624
rect 1596 2582 1624 5510
rect 1952 5092 2004 5098
rect 1952 5034 2004 5040
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1872 4321 1900 4966
rect 1964 4826 1992 5034
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1858 4312 1914 4321
rect 1858 4247 1914 4256
rect 1952 4004 2004 4010
rect 1952 3946 2004 3952
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1872 3505 1900 3878
rect 1964 3738 1992 3946
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1858 3496 1914 3505
rect 1858 3431 1914 3440
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1676 3120 1728 3126
rect 1676 3062 1728 3068
rect 1584 2576 1636 2582
rect 1584 2518 1636 2524
rect 1398 1456 1454 1465
rect 1398 1391 1454 1400
rect 1688 800 1716 3062
rect 1768 2916 1820 2922
rect 1768 2858 1820 2864
rect 1780 1057 1808 2858
rect 1872 2281 1900 3334
rect 1964 3194 1992 3538
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 2056 2990 2084 7482
rect 2424 7342 2452 7686
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2516 6934 2544 10911
rect 2608 10470 2636 12106
rect 2700 11098 2728 12310
rect 2792 11200 2820 13790
rect 2884 13705 2912 13806
rect 2870 13696 2926 13705
rect 2870 13631 2926 13640
rect 2976 12986 3004 15127
rect 3160 14482 3188 16351
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 3252 14550 3280 15098
rect 3330 14784 3386 14793
rect 3330 14719 3386 14728
rect 3240 14544 3292 14550
rect 3240 14486 3292 14492
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 3160 13530 3188 14418
rect 3238 13832 3294 13841
rect 3238 13767 3240 13776
rect 3292 13767 3294 13776
rect 3240 13738 3292 13744
rect 3344 13530 3372 14719
rect 3528 14550 3556 16400
rect 3516 14544 3568 14550
rect 3516 14486 3568 14492
rect 3606 14512 3662 14521
rect 3424 14476 3476 14482
rect 3606 14447 3608 14456
rect 3424 14418 3476 14424
rect 3660 14447 3662 14456
rect 3608 14418 3660 14424
rect 3436 14074 3464 14418
rect 3700 14340 3752 14346
rect 3700 14282 3752 14288
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 3252 12986 3280 13194
rect 3436 13190 3464 13806
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2884 12646 2912 12786
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 3068 12442 3096 12650
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 2884 11608 2912 12106
rect 3252 11937 3280 12582
rect 3528 12322 3556 14214
rect 3712 14074 3740 14282
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 3804 13870 3832 16759
rect 4158 16400 4214 17200
rect 4802 16400 4858 17200
rect 5446 16400 5502 17200
rect 6090 16400 6146 17200
rect 6734 16400 6790 17200
rect 7378 16400 7434 17200
rect 8022 16400 8078 17200
rect 8666 16400 8722 17200
rect 9310 16400 9366 17200
rect 9954 16400 10010 17200
rect 10598 16400 10654 17200
rect 11242 16400 11298 17200
rect 11886 16400 11942 17200
rect 12530 16400 12586 17200
rect 13174 16400 13230 17200
rect 13818 16400 13874 17200
rect 14462 16400 14518 17200
rect 15106 16400 15162 17200
rect 15750 16400 15806 17200
rect 16394 16400 16450 17200
rect 17038 16400 17094 17200
rect 17406 16824 17462 16833
rect 17406 16759 17462 16768
rect 4172 14550 4200 16400
rect 4252 15088 4304 15094
rect 4252 15030 4304 15036
rect 4160 14544 4212 14550
rect 4160 14486 4212 14492
rect 3921 14172 4217 14192
rect 3977 14170 4001 14172
rect 4057 14170 4081 14172
rect 4137 14170 4161 14172
rect 3999 14118 4001 14170
rect 4063 14118 4075 14170
rect 4137 14118 4139 14170
rect 3977 14116 4001 14118
rect 4057 14116 4081 14118
rect 4137 14116 4161 14118
rect 3921 14096 4217 14116
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 3884 13456 3936 13462
rect 3884 13398 3936 13404
rect 3896 13326 3924 13398
rect 3884 13320 3936 13326
rect 3882 13288 3884 13297
rect 3936 13288 3938 13297
rect 3882 13223 3938 13232
rect 3921 13084 4217 13104
rect 3977 13082 4001 13084
rect 4057 13082 4081 13084
rect 4137 13082 4161 13084
rect 3999 13030 4001 13082
rect 4063 13030 4075 13082
rect 4137 13030 4139 13082
rect 3977 13028 4001 13030
rect 4057 13028 4081 13030
rect 4137 13028 4161 13030
rect 3921 13008 4217 13028
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3804 12646 3832 12786
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 3804 12434 3832 12582
rect 3436 12306 3556 12322
rect 3424 12300 3556 12306
rect 3476 12294 3556 12300
rect 3424 12242 3476 12248
rect 3528 12102 3556 12294
rect 3712 12406 3832 12434
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3238 11928 3294 11937
rect 3238 11863 3294 11872
rect 3344 11801 3372 12038
rect 3330 11792 3386 11801
rect 3330 11727 3386 11736
rect 2964 11620 3016 11626
rect 2884 11580 2964 11608
rect 2964 11562 3016 11568
rect 2792 11172 3188 11200
rect 2700 11070 2820 11098
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2700 10674 2728 10950
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2792 10554 2820 11070
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 2700 10526 2820 10554
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2608 8634 2636 9318
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2700 7562 2728 10526
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2884 9382 2912 10202
rect 2976 10062 3004 10406
rect 3068 10169 3096 11018
rect 3054 10160 3110 10169
rect 3054 10095 3110 10104
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2964 8560 3016 8566
rect 2962 8528 2964 8537
rect 3016 8528 3018 8537
rect 2962 8463 3018 8472
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 2872 8016 2924 8022
rect 2872 7958 2924 7964
rect 2608 7534 2728 7562
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2504 6656 2556 6662
rect 2424 6616 2504 6644
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2148 4758 2176 4966
rect 2136 4752 2188 4758
rect 2136 4694 2188 4700
rect 2228 3936 2280 3942
rect 2226 3904 2228 3913
rect 2280 3904 2282 3913
rect 2226 3839 2282 3848
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2240 3097 2268 3334
rect 2226 3088 2282 3097
rect 2226 3023 2282 3032
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 2136 2984 2188 2990
rect 2424 2938 2452 6616
rect 2504 6598 2556 6604
rect 2608 5846 2636 7534
rect 2884 7478 2912 7958
rect 2976 7886 3004 8298
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2976 6934 3004 7346
rect 2780 6928 2832 6934
rect 2780 6870 2832 6876
rect 2964 6928 3016 6934
rect 2964 6870 3016 6876
rect 2792 5846 2820 6870
rect 2596 5840 2648 5846
rect 2596 5782 2648 5788
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2884 5370 2912 5714
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2594 5264 2650 5273
rect 2976 5234 3004 5510
rect 2594 5199 2650 5208
rect 2964 5228 3016 5234
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2136 2926 2188 2932
rect 1858 2272 1914 2281
rect 1858 2207 1914 2216
rect 1766 1048 1822 1057
rect 1766 983 1822 992
rect 2148 800 2176 2926
rect 2332 2922 2452 2938
rect 2320 2916 2452 2922
rect 2372 2910 2452 2916
rect 2320 2858 2372 2864
rect 2516 2854 2544 4014
rect 2608 2990 2636 5199
rect 2964 5170 3016 5176
rect 2872 5092 2924 5098
rect 2872 5034 2924 5040
rect 2884 4826 2912 5034
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 2700 3602 2728 4218
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2688 3596 2740 3602
rect 2688 3538 2740 3544
rect 2792 3058 2820 3878
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 2228 2848 2280 2854
rect 2228 2790 2280 2796
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 2240 1873 2268 2790
rect 2608 2582 2636 2926
rect 2596 2576 2648 2582
rect 2596 2518 2648 2524
rect 2688 2372 2740 2378
rect 2688 2314 2740 2320
rect 2226 1864 2282 1873
rect 2226 1799 2282 1808
rect 2700 800 2728 2314
rect 2884 2310 2912 3470
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 2976 2990 3004 3130
rect 3068 3058 3096 9862
rect 3160 6361 3188 11172
rect 3424 11144 3476 11150
rect 3344 11104 3424 11132
rect 3344 10606 3372 11104
rect 3424 11086 3476 11092
rect 3516 11076 3568 11082
rect 3516 11018 3568 11024
rect 3332 10600 3384 10606
rect 3528 10577 3556 11018
rect 3712 11014 3740 12406
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 3332 10542 3384 10548
rect 3514 10568 3570 10577
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3252 9761 3280 9862
rect 3238 9752 3294 9761
rect 3238 9687 3294 9696
rect 3252 9625 3280 9687
rect 3238 9616 3294 9625
rect 3344 9586 3372 10542
rect 3424 10532 3476 10538
rect 3514 10503 3570 10512
rect 3608 10532 3660 10538
rect 3424 10474 3476 10480
rect 3608 10474 3660 10480
rect 3436 10266 3464 10474
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3528 9654 3556 10202
rect 3516 9648 3568 9654
rect 3516 9590 3568 9596
rect 3238 9551 3294 9560
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3344 9178 3372 9522
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3514 9344 3570 9353
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3436 9081 3464 9318
rect 3514 9279 3570 9288
rect 3528 9178 3556 9279
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3422 9072 3478 9081
rect 3422 9007 3478 9016
rect 3436 8974 3464 9007
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3436 8090 3464 8570
rect 3620 8430 3648 10474
rect 3712 10266 3740 10950
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3712 9382 3740 10066
rect 3804 10062 3832 12038
rect 3921 11996 4217 12016
rect 3977 11994 4001 11996
rect 4057 11994 4081 11996
rect 4137 11994 4161 11996
rect 3999 11942 4001 11994
rect 4063 11942 4075 11994
rect 4137 11942 4139 11994
rect 3977 11940 4001 11942
rect 4057 11940 4081 11942
rect 4137 11940 4161 11942
rect 3921 11920 4217 11940
rect 3921 10908 4217 10928
rect 3977 10906 4001 10908
rect 4057 10906 4081 10908
rect 4137 10906 4161 10908
rect 3999 10854 4001 10906
rect 4063 10854 4075 10906
rect 4137 10854 4139 10906
rect 3977 10852 4001 10854
rect 4057 10852 4081 10854
rect 4137 10852 4161 10854
rect 3921 10832 4217 10852
rect 4264 10674 4292 15030
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4344 13932 4396 13938
rect 4344 13874 4396 13880
rect 4356 13258 4384 13874
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4356 11694 4384 12174
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3896 9908 3924 10066
rect 3804 9880 3924 9908
rect 3804 9518 3832 9880
rect 3921 9820 4217 9840
rect 3977 9818 4001 9820
rect 4057 9818 4081 9820
rect 4137 9818 4161 9820
rect 3999 9766 4001 9818
rect 4063 9766 4075 9818
rect 4137 9766 4139 9818
rect 3977 9764 4001 9766
rect 4057 9764 4081 9766
rect 4137 9764 4161 9766
rect 3921 9744 4217 9764
rect 3792 9512 3844 9518
rect 4068 9512 4120 9518
rect 3792 9454 3844 9460
rect 4066 9480 4068 9489
rect 4120 9480 4122 9489
rect 3976 9444 4028 9450
rect 4066 9415 4122 9424
rect 3976 9386 4028 9392
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3988 8945 4016 9386
rect 3974 8936 4030 8945
rect 3974 8871 3976 8880
rect 4028 8871 4030 8880
rect 3976 8842 4028 8848
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3424 8084 3476 8090
rect 3344 8044 3424 8072
rect 3344 7546 3372 8044
rect 3424 8026 3476 8032
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3436 7478 3464 7890
rect 3516 7880 3568 7886
rect 3620 7834 3648 8230
rect 3700 7948 3752 7954
rect 3700 7890 3752 7896
rect 3568 7828 3648 7834
rect 3516 7822 3648 7828
rect 3528 7806 3648 7822
rect 3424 7472 3476 7478
rect 3424 7414 3476 7420
rect 3620 7410 3648 7806
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3146 6352 3202 6361
rect 3146 6287 3202 6296
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3160 3602 3188 4422
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 3252 2990 3280 7142
rect 3516 6860 3568 6866
rect 3516 6802 3568 6808
rect 3528 6458 3556 6802
rect 3608 6724 3660 6730
rect 3608 6666 3660 6672
rect 3620 6458 3648 6666
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3436 6118 3464 6258
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3344 5778 3372 6054
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3436 5370 3464 5646
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3528 5234 3556 6394
rect 3606 5808 3662 5817
rect 3606 5743 3662 5752
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3620 4282 3648 5743
rect 3712 5098 3740 7890
rect 3700 5092 3752 5098
rect 3700 5034 3752 5040
rect 3804 4826 3832 8774
rect 3921 8732 4217 8752
rect 3977 8730 4001 8732
rect 4057 8730 4081 8732
rect 4137 8730 4161 8732
rect 3999 8678 4001 8730
rect 4063 8678 4075 8730
rect 4137 8678 4139 8730
rect 3977 8676 4001 8678
rect 4057 8676 4081 8678
rect 4137 8676 4161 8678
rect 3921 8656 4217 8676
rect 4264 8090 4292 10610
rect 4356 10606 4384 11630
rect 4540 11218 4568 14962
rect 4712 14952 4764 14958
rect 4712 14894 4764 14900
rect 4724 14074 4752 14894
rect 4816 14550 4844 16400
rect 4988 15088 5040 15094
rect 4988 15030 5040 15036
rect 5000 14550 5028 15030
rect 5460 14550 5488 16400
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 4988 14544 5040 14550
rect 4988 14486 5040 14492
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 6104 14482 6132 16400
rect 6748 14550 6776 16400
rect 6886 14716 7182 14736
rect 6942 14714 6966 14716
rect 7022 14714 7046 14716
rect 7102 14714 7126 14716
rect 6964 14662 6966 14714
rect 7028 14662 7040 14714
rect 7102 14662 7104 14714
rect 6942 14660 6966 14662
rect 7022 14660 7046 14662
rect 7102 14660 7126 14662
rect 6886 14640 7182 14660
rect 7392 14550 7420 16400
rect 7656 14884 7708 14890
rect 7656 14826 7708 14832
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 7380 14544 7432 14550
rect 7380 14486 7432 14492
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 5552 14074 5580 14418
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 4620 13864 4672 13870
rect 4618 13832 4620 13841
rect 4672 13832 4674 13841
rect 4618 13767 4674 13776
rect 4724 13705 4752 14010
rect 4710 13696 4766 13705
rect 4710 13631 4766 13640
rect 5736 13326 5764 14418
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 5816 14000 5868 14006
rect 5816 13942 5868 13948
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 4710 12744 4766 12753
rect 4710 12679 4766 12688
rect 4724 12434 4752 12679
rect 5828 12434 5856 13942
rect 5920 13734 5948 14214
rect 6012 13870 6040 14214
rect 6656 14074 6684 14418
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6736 14000 6788 14006
rect 6736 13942 6788 13948
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 4724 12406 4844 12434
rect 5828 12406 5948 12434
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4632 11558 4660 12242
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4632 10198 4660 11494
rect 4724 11354 4752 11562
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 3921 7644 4217 7664
rect 3977 7642 4001 7644
rect 4057 7642 4081 7644
rect 4137 7642 4161 7644
rect 3999 7590 4001 7642
rect 4063 7590 4075 7642
rect 4137 7590 4139 7642
rect 3977 7588 4001 7590
rect 4057 7588 4081 7590
rect 4137 7588 4161 7590
rect 3921 7568 4217 7588
rect 4264 7478 4292 8026
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 3921 6556 4217 6576
rect 3977 6554 4001 6556
rect 4057 6554 4081 6556
rect 4137 6554 4161 6556
rect 3999 6502 4001 6554
rect 4063 6502 4075 6554
rect 4137 6502 4139 6554
rect 3977 6500 4001 6502
rect 4057 6500 4081 6502
rect 4137 6500 4161 6502
rect 3921 6480 4217 6500
rect 4264 6118 4292 6734
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4250 5944 4306 5953
rect 4250 5879 4252 5888
rect 4304 5879 4306 5888
rect 4252 5850 4304 5856
rect 4250 5672 4306 5681
rect 4250 5607 4306 5616
rect 4264 5574 4292 5607
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 3921 5468 4217 5488
rect 3977 5466 4001 5468
rect 4057 5466 4081 5468
rect 4137 5466 4161 5468
rect 3999 5414 4001 5466
rect 4063 5414 4075 5466
rect 4137 5414 4139 5466
rect 3977 5412 4001 5414
rect 4057 5412 4081 5414
rect 4137 5412 4161 5414
rect 3921 5392 4217 5412
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4172 4826 4200 4966
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 3804 4690 3832 4762
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 3921 4380 4217 4400
rect 3977 4378 4001 4380
rect 4057 4378 4081 4380
rect 4137 4378 4161 4380
rect 3999 4326 4001 4378
rect 4063 4326 4075 4378
rect 4137 4326 4139 4378
rect 3977 4324 4001 4326
rect 4057 4324 4081 4326
rect 4137 4324 4161 4326
rect 3921 4304 4217 4324
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3620 3738 3648 3878
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 3068 2650 3096 2790
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3160 2582 3188 2790
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 3148 2372 3200 2378
rect 3148 2314 3200 2320
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 3160 800 3188 2314
rect 1306 640 1362 649
rect 1306 575 1362 584
rect 1674 0 1730 800
rect 2134 0 2190 800
rect 2686 0 2742 800
rect 3146 0 3202 800
rect 3344 241 3372 3334
rect 3712 3194 3740 3334
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3608 2848 3660 2854
rect 3608 2790 3660 2796
rect 3620 2582 3648 2790
rect 3608 2576 3660 2582
rect 3608 2518 3660 2524
rect 3712 2514 3740 2994
rect 3804 2990 3832 3878
rect 3921 3292 4217 3312
rect 3977 3290 4001 3292
rect 4057 3290 4081 3292
rect 4137 3290 4161 3292
rect 3999 3238 4001 3290
rect 4063 3238 4075 3290
rect 4137 3238 4139 3290
rect 3977 3236 4001 3238
rect 4057 3236 4081 3238
rect 4137 3236 4161 3238
rect 3921 3216 4217 3236
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 3792 2984 3844 2990
rect 4068 2984 4120 2990
rect 3792 2926 3844 2932
rect 4066 2952 4068 2961
rect 4120 2952 4122 2961
rect 4066 2887 4122 2896
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3896 2582 3924 2790
rect 4172 2650 4200 3062
rect 4356 2990 4384 9862
rect 4620 9444 4672 9450
rect 4620 9386 4672 9392
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 3884 2576 3936 2582
rect 3884 2518 3936 2524
rect 4264 2514 4292 2858
rect 4448 2582 4476 9318
rect 4632 9178 4660 9386
rect 4724 9178 4752 11018
rect 4816 9625 4844 12406
rect 5920 11354 5948 12406
rect 5908 11348 5960 11354
rect 5908 11290 5960 11296
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4908 10266 4936 10406
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 4802 9616 4858 9625
rect 4802 9551 4858 9560
rect 4894 9480 4950 9489
rect 4894 9415 4950 9424
rect 4908 9382 4936 9415
rect 4896 9376 4948 9382
rect 4816 9336 4896 9364
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4526 8936 4582 8945
rect 4526 8871 4582 8880
rect 4540 4826 4568 8871
rect 4632 8809 4660 9114
rect 4618 8800 4674 8809
rect 4674 8758 4752 8786
rect 4618 8735 4674 8744
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4632 7342 4660 7686
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4724 5658 4752 8758
rect 4816 6474 4844 9336
rect 4896 9318 4948 9324
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4908 7154 4936 9114
rect 5000 7721 5028 11154
rect 5908 11076 5960 11082
rect 5828 11036 5908 11064
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5538 10704 5594 10713
rect 5538 10639 5594 10648
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5460 9722 5488 10542
rect 5448 9716 5500 9722
rect 5448 9658 5500 9664
rect 5262 9616 5318 9625
rect 5262 9551 5318 9560
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4986 7712 5042 7721
rect 4986 7647 5042 7656
rect 5092 7546 5120 8026
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5184 7342 5212 8230
rect 5276 8090 5304 9551
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5368 8090 5396 9046
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5276 7546 5304 7822
rect 5368 7585 5396 7890
rect 5460 7886 5488 8434
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5354 7576 5410 7585
rect 5264 7540 5316 7546
rect 5354 7511 5410 7520
rect 5264 7482 5316 7488
rect 5368 7410 5396 7511
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5552 7342 5580 10639
rect 5736 10470 5764 10950
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5644 8090 5672 8230
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5644 7274 5672 7890
rect 5632 7268 5684 7274
rect 5632 7210 5684 7216
rect 4908 7126 5212 7154
rect 4816 6446 5120 6474
rect 4896 6384 4948 6390
rect 4894 6352 4896 6361
rect 4948 6352 4950 6361
rect 4894 6287 4950 6296
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 5000 5710 5028 6258
rect 4632 5630 4752 5658
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4540 4282 4568 4762
rect 4632 4672 4660 5630
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4724 5166 4752 5510
rect 4816 5302 4844 5510
rect 5000 5370 5028 5646
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 5000 4826 5028 5034
rect 5092 4826 5120 6446
rect 5184 6066 5212 7126
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5276 6186 5304 6598
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5264 6180 5316 6186
rect 5264 6122 5316 6128
rect 5448 6112 5500 6118
rect 5184 6038 5304 6066
rect 5448 6054 5500 6060
rect 5276 5370 5304 6038
rect 5354 5944 5410 5953
rect 5460 5914 5488 6054
rect 5354 5879 5410 5888
rect 5448 5908 5500 5914
rect 5368 5710 5396 5879
rect 5448 5850 5500 5856
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5552 5574 5580 6190
rect 5736 5681 5764 9658
rect 5828 8401 5856 11036
rect 5908 11018 5960 11024
rect 6092 10736 6144 10742
rect 6092 10678 6144 10684
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5920 10062 5948 10610
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6012 10198 6040 10406
rect 6000 10192 6052 10198
rect 6000 10134 6052 10140
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 5908 9376 5960 9382
rect 6012 9353 6040 9590
rect 5908 9318 5960 9324
rect 5998 9344 6054 9353
rect 5920 9178 5948 9318
rect 5998 9279 6054 9288
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 6012 8634 6040 9114
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6104 8566 6132 10678
rect 6092 8560 6144 8566
rect 6092 8502 6144 8508
rect 5814 8392 5870 8401
rect 5870 8350 5948 8378
rect 5814 8327 5870 8336
rect 5816 8016 5868 8022
rect 5816 7958 5868 7964
rect 5828 7478 5856 7958
rect 5816 7472 5868 7478
rect 5816 7414 5868 7420
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 5828 6254 5856 6326
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5920 5817 5948 8350
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 6012 5914 6040 6054
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 5906 5808 5962 5817
rect 5816 5772 5868 5778
rect 5906 5743 5962 5752
rect 5816 5714 5868 5720
rect 5722 5672 5778 5681
rect 5722 5607 5778 5616
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 4712 4684 4764 4690
rect 4632 4644 4712 4672
rect 4712 4626 4764 4632
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4632 3194 4660 3946
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4816 3398 4844 3878
rect 4988 3460 5040 3466
rect 4988 3402 5040 3408
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 4540 2582 4568 2790
rect 4436 2576 4488 2582
rect 4436 2518 4488 2524
rect 4528 2576 4580 2582
rect 4528 2518 4580 2524
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 4252 2508 4304 2514
rect 4252 2450 4304 2456
rect 3436 2106 3464 2450
rect 3608 2372 3660 2378
rect 3608 2314 3660 2320
rect 4252 2372 4304 2378
rect 4252 2314 4304 2320
rect 3424 2100 3476 2106
rect 3424 2042 3476 2048
rect 3620 800 3648 2314
rect 3921 2204 4217 2224
rect 3977 2202 4001 2204
rect 4057 2202 4081 2204
rect 4137 2202 4161 2204
rect 3999 2150 4001 2202
rect 4063 2150 4075 2202
rect 4137 2150 4139 2202
rect 3977 2148 4001 2150
rect 4057 2148 4081 2150
rect 4137 2148 4161 2150
rect 3921 2128 4217 2148
rect 4264 1170 4292 2314
rect 4172 1142 4292 1170
rect 4172 800 4200 1142
rect 4632 800 4660 2926
rect 5000 2582 5028 3402
rect 5092 3126 5120 4762
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5184 4214 5212 4558
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5184 3534 5212 4014
rect 5276 3602 5304 5306
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5460 4570 5488 5034
rect 5460 4554 5580 4570
rect 5828 4554 5856 5714
rect 6012 5642 6040 5850
rect 6104 5778 6132 8502
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 6196 5114 6224 13806
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6288 11150 6316 11834
rect 6564 11694 6592 12038
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6288 8294 6316 11086
rect 6472 10606 6500 11290
rect 6564 11150 6592 11630
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6380 9994 6408 10202
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6564 9586 6592 11086
rect 6656 10062 6684 11222
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6656 9654 6684 9998
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6368 9444 6420 9450
rect 6420 9404 6500 9432
rect 6368 9386 6420 9392
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6380 8634 6408 8978
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6380 7954 6408 8570
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6288 7002 6316 7822
rect 6368 7268 6420 7274
rect 6368 7210 6420 7216
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6288 5166 6316 5510
rect 6380 5273 6408 7210
rect 6472 7018 6500 9404
rect 6564 8974 6592 9522
rect 6748 9450 6776 13942
rect 6886 13628 7182 13648
rect 6942 13626 6966 13628
rect 7022 13626 7046 13628
rect 7102 13626 7126 13628
rect 6964 13574 6966 13626
rect 7028 13574 7040 13626
rect 7102 13574 7104 13626
rect 6942 13572 6966 13574
rect 7022 13572 7046 13574
rect 7102 13572 7126 13574
rect 6886 13552 7182 13572
rect 6886 12540 7182 12560
rect 6942 12538 6966 12540
rect 7022 12538 7046 12540
rect 7102 12538 7126 12540
rect 6964 12486 6966 12538
rect 7028 12486 7040 12538
rect 7102 12486 7104 12538
rect 6942 12484 6966 12486
rect 7022 12484 7046 12486
rect 7102 12484 7126 12486
rect 6886 12464 7182 12484
rect 7564 11688 7616 11694
rect 7484 11636 7564 11642
rect 7484 11630 7616 11636
rect 7484 11614 7604 11630
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 6886 11452 7182 11472
rect 6942 11450 6966 11452
rect 7022 11450 7046 11452
rect 7102 11450 7126 11452
rect 6964 11398 6966 11450
rect 7028 11398 7040 11450
rect 7102 11398 7104 11450
rect 6942 11396 6966 11398
rect 7022 11396 7046 11398
rect 7102 11396 7126 11398
rect 6886 11376 7182 11396
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6840 10742 6868 10950
rect 6828 10736 6880 10742
rect 6828 10678 6880 10684
rect 7024 10674 7052 11222
rect 7300 11200 7328 11494
rect 7380 11212 7432 11218
rect 7300 11172 7380 11200
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 7208 10606 7236 10678
rect 7300 10606 7328 11172
rect 7380 11154 7432 11160
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 6886 10364 7182 10384
rect 6942 10362 6966 10364
rect 7022 10362 7046 10364
rect 7102 10362 7126 10364
rect 6964 10310 6966 10362
rect 7028 10310 7040 10362
rect 7102 10310 7104 10362
rect 6942 10308 6966 10310
rect 7022 10308 7046 10310
rect 7102 10308 7126 10310
rect 6886 10288 7182 10308
rect 7300 10130 7328 10542
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7208 9722 7236 9862
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6644 9376 6696 9382
rect 6642 9344 6644 9353
rect 6696 9344 6698 9353
rect 6642 9279 6698 9288
rect 6656 9110 6684 9279
rect 6886 9276 7182 9296
rect 6942 9274 6966 9276
rect 7022 9274 7046 9276
rect 7102 9274 7126 9276
rect 6964 9222 6966 9274
rect 7028 9222 7040 9274
rect 7102 9222 7104 9274
rect 6942 9220 6966 9222
rect 7022 9220 7046 9222
rect 7102 9220 7126 9222
rect 6886 9200 7182 9220
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6564 8090 6592 8298
rect 6656 8090 6684 9046
rect 7300 9042 7328 10066
rect 7392 9926 7420 10678
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7380 9444 7432 9450
rect 7380 9386 7432 9392
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 6886 8188 7182 8208
rect 6942 8186 6966 8188
rect 7022 8186 7046 8188
rect 7102 8186 7126 8188
rect 6964 8134 6966 8186
rect 7028 8134 7040 8186
rect 7102 8134 7104 8186
rect 6942 8132 6966 8134
rect 7022 8132 7046 8134
rect 7102 8132 7126 8134
rect 6886 8112 7182 8132
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6656 7546 6684 8026
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 7116 7410 7144 7822
rect 7300 7818 7328 8366
rect 7392 8090 7420 9386
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 6656 7206 6684 7346
rect 7392 7206 7420 8026
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 6886 7100 7182 7120
rect 6942 7098 6966 7100
rect 7022 7098 7046 7100
rect 7102 7098 7126 7100
rect 6964 7046 6966 7098
rect 7028 7046 7040 7098
rect 7102 7046 7104 7098
rect 6942 7044 6966 7046
rect 7022 7044 7046 7046
rect 7102 7044 7126 7046
rect 6886 7024 7182 7044
rect 6472 6990 6684 7018
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 6472 5846 6500 6054
rect 6460 5840 6512 5846
rect 6460 5782 6512 5788
rect 6366 5264 6422 5273
rect 6366 5199 6422 5208
rect 5920 5086 6224 5114
rect 6276 5160 6328 5166
rect 6276 5102 6328 5108
rect 5460 4548 5592 4554
rect 5460 4542 5540 4548
rect 5460 4282 5488 4542
rect 5540 4490 5592 4496
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 5920 2774 5948 5086
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6184 5024 6236 5030
rect 6552 5024 6604 5030
rect 6184 4966 6236 4972
rect 6288 4984 6552 5012
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6012 3942 6040 4626
rect 6104 4554 6132 4966
rect 6092 4548 6144 4554
rect 6092 4490 6144 4496
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 6196 3602 6224 4966
rect 6288 4622 6316 4984
rect 6552 4966 6604 4972
rect 6552 4752 6604 4758
rect 6552 4694 6604 4700
rect 6564 4622 6592 4694
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6288 4282 6316 4558
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6564 3670 6592 4218
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6196 3194 6224 3538
rect 6564 3466 6592 3606
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 5736 2746 5948 2774
rect 5736 2650 5764 2746
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 6656 2582 6684 6990
rect 7392 6934 7420 7142
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6840 6254 6868 6734
rect 6932 6254 6960 6802
rect 7484 6746 7512 11614
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7576 7886 7604 8298
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7668 7732 7696 14826
rect 8036 14498 8064 16400
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8036 14470 8156 14498
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 8036 12434 8064 14214
rect 7944 12406 8064 12434
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7852 11286 7880 11494
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 7746 9208 7802 9217
rect 7746 9143 7748 9152
rect 7800 9143 7802 9152
rect 7748 9114 7800 9120
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7852 8498 7880 8978
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 7760 7954 7788 8298
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7576 7704 7696 7732
rect 7748 7744 7800 7750
rect 7576 6866 7604 7704
rect 7748 7686 7800 7692
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7668 6934 7696 7142
rect 7760 7002 7788 7686
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7484 6718 7604 6746
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6886 6012 7182 6032
rect 6942 6010 6966 6012
rect 7022 6010 7046 6012
rect 7102 6010 7126 6012
rect 6964 5958 6966 6010
rect 7028 5958 7040 6010
rect 7102 5958 7104 6010
rect 6942 5956 6966 5958
rect 7022 5956 7046 5958
rect 7102 5956 7126 5958
rect 6886 5936 7182 5956
rect 7286 5944 7342 5953
rect 7286 5879 7288 5888
rect 7340 5879 7342 5888
rect 7288 5850 7340 5856
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6748 4078 6776 5714
rect 7378 5672 7434 5681
rect 7378 5607 7434 5616
rect 7392 5574 7420 5607
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7380 5092 7432 5098
rect 7380 5034 7432 5040
rect 6886 4924 7182 4944
rect 6942 4922 6966 4924
rect 7022 4922 7046 4924
rect 7102 4922 7126 4924
rect 6964 4870 6966 4922
rect 7028 4870 7040 4922
rect 7102 4870 7104 4922
rect 6942 4868 6966 4870
rect 7022 4868 7046 4870
rect 7102 4868 7126 4870
rect 6886 4848 7182 4868
rect 7392 4146 7420 5034
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6748 3040 6776 4014
rect 6886 3836 7182 3856
rect 6942 3834 6966 3836
rect 7022 3834 7046 3836
rect 7102 3834 7126 3836
rect 6964 3782 6966 3834
rect 7028 3782 7040 3834
rect 7102 3782 7104 3834
rect 6942 3780 6966 3782
rect 7022 3780 7046 3782
rect 7102 3780 7126 3782
rect 6886 3760 7182 3780
rect 7392 3398 7420 4082
rect 7484 3602 7512 6598
rect 7576 4554 7604 6718
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7668 5574 7696 6326
rect 7852 6118 7880 6394
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7944 5778 7972 12406
rect 8128 11694 8156 14470
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8220 10266 8248 15098
rect 8680 14618 8708 16400
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 9324 14482 9352 16400
rect 9968 14482 9996 16400
rect 10612 14482 10640 16400
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10508 14340 10560 14346
rect 10508 14282 10560 14288
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8220 9654 8248 10202
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8220 9353 8248 9454
rect 8312 9382 8340 9590
rect 8300 9376 8352 9382
rect 8206 9344 8262 9353
rect 8300 9318 8352 9324
rect 8206 9279 8262 9288
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 8566 8064 8774
rect 8024 8560 8076 8566
rect 8076 8520 8156 8548
rect 8024 8502 8076 8508
rect 8128 7954 8156 8520
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8220 7834 8248 8230
rect 8312 8022 8340 8230
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8392 7880 8444 7886
rect 8220 7806 8340 7834
rect 8392 7822 8444 7828
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8128 6458 8156 7142
rect 8220 7002 8248 7142
rect 8312 7002 8340 7806
rect 8404 7449 8432 7822
rect 8390 7440 8446 7449
rect 8390 7375 8392 7384
rect 8444 7375 8446 7384
rect 8392 7346 8444 7352
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8220 6361 8248 6802
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8206 6352 8262 6361
rect 8206 6287 8262 6296
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 7746 5672 7802 5681
rect 7746 5607 7802 5616
rect 7932 5636 7984 5642
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7760 5166 7788 5607
rect 7932 5578 7984 5584
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7760 3466 7788 3878
rect 7944 3670 7972 5578
rect 8024 4004 8076 4010
rect 8024 3946 8076 3952
rect 8036 3738 8064 3946
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 7932 3664 7984 3670
rect 7932 3606 7984 3612
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 6828 3052 6880 3058
rect 6748 3012 6828 3040
rect 6828 2994 6880 3000
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 6886 2748 7182 2768
rect 6942 2746 6966 2748
rect 7022 2746 7046 2748
rect 7102 2746 7126 2748
rect 6964 2694 6966 2746
rect 7028 2694 7040 2746
rect 7102 2694 7104 2746
rect 6942 2692 6966 2694
rect 7022 2692 7046 2694
rect 7102 2692 7126 2694
rect 6886 2672 7182 2692
rect 4988 2576 5040 2582
rect 4988 2518 5040 2524
rect 6644 2576 6696 2582
rect 6644 2518 6696 2524
rect 7300 2514 7328 2994
rect 7484 2582 7512 3062
rect 7760 2990 7788 3402
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7852 2854 7880 3470
rect 7944 3058 7972 3606
rect 8036 3194 8064 3674
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8128 3074 8156 3878
rect 8312 3618 8340 6734
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 8404 5681 8432 6326
rect 8390 5672 8446 5681
rect 8390 5607 8446 5616
rect 8220 3602 8340 3618
rect 8208 3596 8340 3602
rect 8260 3590 8340 3596
rect 8208 3538 8260 3544
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 8036 3046 8156 3074
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7472 2576 7524 2582
rect 7472 2518 7524 2524
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 5172 2372 5224 2378
rect 5172 2314 5224 2320
rect 5184 800 5212 2314
rect 5644 800 5672 2450
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6184 2372 6236 2378
rect 6184 2314 6236 2320
rect 6196 800 6224 2314
rect 6656 800 6684 2382
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 7656 2372 7708 2378
rect 7656 2314 7708 2320
rect 7116 800 7144 2314
rect 7668 800 7696 2314
rect 8036 2310 8064 3046
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8128 2582 8156 2790
rect 8312 2582 8340 3334
rect 8496 3126 8524 14214
rect 9852 14172 10148 14192
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 9930 14118 9932 14170
rect 9994 14118 10006 14170
rect 10068 14118 10070 14170
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 9852 14096 10148 14116
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9508 12434 9536 13806
rect 9852 13084 10148 13104
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 9930 13030 9932 13082
rect 9994 13030 10006 13082
rect 10068 13030 10070 13082
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 9852 13008 10148 13028
rect 9232 12406 9536 12434
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8772 10198 8800 10406
rect 8760 10192 8812 10198
rect 8666 10160 8722 10169
rect 8760 10134 8812 10140
rect 8666 10095 8722 10104
rect 8680 9722 8708 10095
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8668 9716 8720 9722
rect 8588 9676 8668 9704
rect 8588 7732 8616 9676
rect 8668 9658 8720 9664
rect 8864 9586 8892 9862
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8864 9110 8892 9522
rect 8852 9104 8904 9110
rect 8666 9072 8722 9081
rect 8852 9046 8904 9052
rect 8666 9007 8722 9016
rect 8680 8974 8708 9007
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8680 8566 8708 8774
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8680 7886 8708 8502
rect 8956 7954 8984 11562
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9048 8498 9076 8774
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9140 8090 9168 9658
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8668 7880 8720 7886
rect 8720 7840 8800 7868
rect 8668 7822 8720 7828
rect 8588 7704 8708 7732
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8588 5166 8616 7278
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8680 5030 8708 7704
rect 8772 7274 8800 7840
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 8772 6798 8800 7210
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 8772 6322 8800 6734
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 9140 6254 9168 6734
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 8852 5772 8904 5778
rect 9128 5772 9180 5778
rect 8904 5732 9128 5760
rect 8852 5714 8904 5720
rect 9128 5714 9180 5720
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8772 4282 8800 5034
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8864 4078 8892 5714
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8864 3738 8892 4014
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 8484 3120 8536 3126
rect 8484 3062 8536 3068
rect 9232 2582 9260 12406
rect 9852 11996 10148 12016
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 9930 11942 9932 11994
rect 9994 11942 10006 11994
rect 10068 11942 10070 11994
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 9852 11920 10148 11940
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 9784 10538 9812 10950
rect 9852 10908 10148 10928
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 9930 10854 9932 10906
rect 9994 10854 10006 10906
rect 10068 10854 10070 10906
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 9852 10832 10148 10852
rect 10336 10674 10364 10950
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9784 10062 9812 10474
rect 10140 10464 10192 10470
rect 10416 10464 10468 10470
rect 10192 10424 10272 10452
rect 10140 10406 10192 10412
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9852 9820 10148 9840
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 9930 9766 9932 9818
rect 9994 9766 10006 9818
rect 10068 9766 10070 9818
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 9852 9744 10148 9764
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9324 9574 9628 9602
rect 9324 9353 9352 9574
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9310 9344 9366 9353
rect 9310 9279 9366 9288
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9324 8430 9352 8774
rect 9416 8650 9444 9454
rect 9600 9364 9628 9574
rect 9680 9376 9732 9382
rect 9600 9336 9680 9364
rect 9680 9318 9732 9324
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9600 8945 9628 8978
rect 9784 8974 9812 9658
rect 10244 9654 10272 10424
rect 10416 10406 10468 10412
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 9876 9353 9904 9454
rect 10152 9382 10180 9590
rect 10140 9376 10192 9382
rect 9862 9344 9918 9353
rect 10140 9318 10192 9324
rect 9862 9279 9918 9288
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 9772 8968 9824 8974
rect 9586 8936 9642 8945
rect 9772 8910 9824 8916
rect 9586 8871 9642 8880
rect 9680 8832 9732 8838
rect 9968 8820 9996 9114
rect 9784 8792 9996 8820
rect 9784 8786 9812 8792
rect 9732 8780 9812 8786
rect 9680 8774 9812 8780
rect 9692 8758 9812 8774
rect 9852 8732 10148 8752
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 9930 8678 9932 8730
rect 9994 8678 10006 8730
rect 10068 8678 10070 8730
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 9852 8656 10148 8676
rect 9416 8622 9628 8650
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9402 8392 9458 8401
rect 9402 8327 9458 8336
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9324 7585 9352 8026
rect 9416 7954 9444 8327
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9310 7576 9366 7585
rect 9310 7511 9366 7520
rect 9310 7440 9366 7449
rect 9310 7375 9366 7384
rect 9324 7342 9352 7375
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9600 5794 9628 8622
rect 9956 8560 10008 8566
rect 9954 8528 9956 8537
rect 10008 8528 10010 8537
rect 10244 8514 10272 9590
rect 10336 9518 10364 9862
rect 10428 9586 10456 10406
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10414 9480 10470 9489
rect 10414 9415 10470 9424
rect 10324 9036 10376 9042
rect 10428 9024 10456 9415
rect 10376 8996 10456 9024
rect 10324 8978 10376 8984
rect 10428 8838 10456 8996
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10244 8486 10364 8514
rect 9954 8463 10010 8472
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 9852 7644 10148 7664
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 9930 7590 9932 7642
rect 9994 7590 10006 7642
rect 10068 7590 10070 7642
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 9852 7568 10148 7588
rect 10140 7472 10192 7478
rect 10244 7460 10272 8298
rect 10192 7432 10272 7460
rect 10140 7414 10192 7420
rect 10152 6730 10180 7414
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 9852 6556 10148 6576
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 9930 6502 9932 6554
rect 9994 6502 10006 6554
rect 10068 6502 10070 6554
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 9852 6480 10148 6500
rect 10336 6254 10364 8486
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 9508 5766 9628 5794
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9324 5370 9352 5510
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9324 5234 9352 5306
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9508 4826 9536 5766
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 9600 4826 9628 5510
rect 9852 5468 10148 5488
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 9930 5414 9932 5466
rect 9994 5414 10006 5466
rect 10068 5414 10070 5466
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 9852 5392 10148 5412
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9416 2990 9444 4082
rect 9496 4072 9548 4078
rect 9600 4060 9628 4762
rect 9852 4380 10148 4400
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 9930 4326 9932 4378
rect 9994 4326 10006 4378
rect 10068 4326 10070 4378
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 9852 4304 10148 4324
rect 10336 4078 10364 5510
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 9548 4032 9628 4060
rect 10324 4072 10376 4078
rect 9496 4014 9548 4020
rect 10324 4014 10376 4020
rect 10428 4010 10456 4422
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9692 3126 9720 3334
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9784 2990 9812 3334
rect 9852 3292 10148 3312
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 9930 3238 9932 3290
rect 9994 3238 10006 3290
rect 10068 3238 10070 3290
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 9852 3216 10148 3236
rect 10244 3126 10272 3878
rect 10428 3398 10456 3946
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 9220 2576 9272 2582
rect 9220 2518 9272 2524
rect 9324 2514 9352 2790
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 8116 2372 8168 2378
rect 8116 2314 8168 2320
rect 8668 2372 8720 2378
rect 8668 2314 8720 2320
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 8128 800 8156 2314
rect 8680 800 8708 2314
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9140 800 9168 2246
rect 9692 800 9720 2858
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9784 2650 9812 2790
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 10152 2582 10180 3062
rect 10428 3058 10456 3130
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10230 2816 10286 2825
rect 10230 2751 10286 2760
rect 10140 2576 10192 2582
rect 10140 2518 10192 2524
rect 9852 2204 10148 2224
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 9930 2150 9932 2202
rect 9994 2150 10006 2202
rect 10068 2150 10070 2202
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 9852 2128 10148 2148
rect 10244 1034 10272 2751
rect 10520 2582 10548 14282
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10704 10130 10732 10542
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10704 9722 10732 10066
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10704 8906 10732 9386
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 10796 7834 10824 14214
rect 10888 12374 10916 14962
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 11164 14006 11192 14554
rect 11256 14482 11284 16400
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11336 14340 11388 14346
rect 11336 14282 11388 14288
rect 11152 14000 11204 14006
rect 11152 13942 11204 13948
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 11072 12434 11100 13398
rect 11348 12434 11376 14282
rect 11624 12434 11652 14486
rect 11900 14482 11928 16400
rect 12440 14544 12492 14550
rect 12440 14486 12492 14492
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11072 12406 11192 12434
rect 11348 12406 11468 12434
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10888 10266 10916 12310
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10888 9926 10916 10202
rect 11058 10024 11114 10033
rect 11058 9959 11114 9968
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10980 9178 11008 9454
rect 11072 9382 11100 9959
rect 11060 9376 11112 9382
rect 11058 9344 11060 9353
rect 11112 9344 11114 9353
rect 11058 9279 11114 9288
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10980 8537 11008 8978
rect 10966 8528 11022 8537
rect 10966 8463 11022 8472
rect 10796 7806 10916 7834
rect 10782 6760 10838 6769
rect 10782 6695 10838 6704
rect 10796 6458 10824 6695
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10612 4622 10640 5170
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 10612 3942 10640 4218
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10600 3664 10652 3670
rect 10600 3606 10652 3612
rect 10612 3505 10640 3606
rect 10598 3496 10654 3505
rect 10598 3431 10654 3440
rect 10598 3360 10654 3369
rect 10598 3295 10654 3304
rect 10612 2990 10640 3295
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 10508 2576 10560 2582
rect 10508 2518 10560 2524
rect 10152 1006 10272 1034
rect 10152 800 10180 1006
rect 10612 800 10640 2790
rect 10704 2106 10732 6326
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10796 5914 10824 6190
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10796 5098 10824 5850
rect 10784 5092 10836 5098
rect 10784 5034 10836 5040
rect 10796 4758 10824 5034
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10796 3602 10824 4422
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10796 2990 10824 3538
rect 10888 3233 10916 7806
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10980 5914 11008 7278
rect 11072 6934 11100 7686
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10980 4486 11008 5102
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10874 3224 10930 3233
rect 10874 3159 10930 3168
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10888 2825 10916 2926
rect 10874 2816 10930 2825
rect 10874 2751 10930 2760
rect 10980 2650 11008 3538
rect 11072 3534 11100 4966
rect 11164 4282 11192 12406
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11256 9178 11284 10406
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11348 8838 11376 9318
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11256 5522 11284 6938
rect 11334 6896 11390 6905
rect 11334 6831 11390 6840
rect 11348 6662 11376 6831
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11336 6248 11388 6254
rect 11336 6190 11388 6196
rect 11348 5914 11376 6190
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11256 5494 11376 5522
rect 11348 5370 11376 5494
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11256 4758 11284 5306
rect 11440 4842 11468 12406
rect 11532 12406 11652 12434
rect 11532 6746 11560 12406
rect 11716 11370 11744 13806
rect 11624 11342 11744 11370
rect 11624 11014 11652 11342
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11624 10266 11652 10950
rect 11716 10606 11744 11154
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11612 10260 11664 10266
rect 11808 10248 11836 13942
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12084 12434 12112 12922
rect 12084 12406 12204 12434
rect 11888 11280 11940 11286
rect 11888 11222 11940 11228
rect 11980 11280 12032 11286
rect 11980 11222 12032 11228
rect 11900 11150 11928 11222
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11888 11008 11940 11014
rect 11992 10996 12020 11222
rect 11940 10968 12020 10996
rect 11888 10950 11940 10956
rect 11900 10810 11928 10950
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11900 10538 11928 10746
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 12072 10260 12124 10266
rect 11808 10220 12020 10248
rect 11612 10202 11664 10208
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11624 9586 11652 10066
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11716 9466 11744 9930
rect 11624 9438 11744 9466
rect 11624 8974 11652 9438
rect 11900 9382 11928 10066
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11716 8430 11744 8774
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11716 7342 11744 7686
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11532 6718 11744 6746
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11532 5914 11560 6598
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11520 5704 11572 5710
rect 11572 5664 11652 5692
rect 11520 5646 11572 5652
rect 11624 5574 11652 5664
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11440 4814 11652 4842
rect 11624 4758 11652 4814
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11612 4752 11664 4758
rect 11612 4694 11664 4700
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11532 4078 11560 4422
rect 11716 4146 11744 6718
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 11072 2990 11100 3334
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 11348 2582 11376 3878
rect 11624 3602 11652 3878
rect 11612 3596 11664 3602
rect 11532 3556 11612 3584
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 11336 2576 11388 2582
rect 11336 2518 11388 2524
rect 11440 2446 11468 3402
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 11532 2292 11560 3556
rect 11612 3538 11664 3544
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11624 2922 11652 3334
rect 11612 2916 11664 2922
rect 11612 2858 11664 2864
rect 11716 2774 11744 3538
rect 11808 3058 11836 8230
rect 11900 7546 11928 8978
rect 11992 8294 12020 10220
rect 12072 10202 12124 10208
rect 12084 9586 12112 10202
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11980 8016 12032 8022
rect 11978 7984 11980 7993
rect 12032 7984 12034 7993
rect 11978 7919 12034 7928
rect 11888 7540 11940 7546
rect 11940 7500 12112 7528
rect 11888 7482 11940 7488
rect 12084 7290 12112 7500
rect 12176 7478 12204 12406
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 12268 10674 12296 11018
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12268 9994 12296 10610
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12256 9988 12308 9994
rect 12256 9930 12308 9936
rect 12360 9674 12388 10202
rect 12268 9646 12388 9674
rect 12268 9110 12296 9646
rect 12452 9466 12480 14486
rect 12544 14482 12572 16400
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12728 14550 12756 14894
rect 12817 14716 13113 14736
rect 12873 14714 12897 14716
rect 12953 14714 12977 14716
rect 13033 14714 13057 14716
rect 12895 14662 12897 14714
rect 12959 14662 12971 14714
rect 13033 14662 13035 14714
rect 12873 14660 12897 14662
rect 12953 14660 12977 14662
rect 13033 14660 13057 14662
rect 12817 14640 13113 14660
rect 12716 14544 12768 14550
rect 12716 14486 12768 14492
rect 13188 14482 13216 16400
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13280 14618 13308 14894
rect 13544 14884 13596 14890
rect 13544 14826 13596 14832
rect 13556 14618 13584 14826
rect 13832 14618 13860 16400
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 14016 14550 14044 14758
rect 14476 14550 14504 16400
rect 15016 15088 15068 15094
rect 15016 15030 15068 15036
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 14464 14544 14516 14550
rect 14464 14486 14516 14492
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14832 14476 14884 14482
rect 14832 14418 14884 14424
rect 13188 14074 13216 14418
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13280 14006 13308 14418
rect 13452 14340 13504 14346
rect 13452 14282 13504 14288
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13464 14006 13492 14282
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13648 13870 13676 14282
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 12817 13628 13113 13648
rect 12873 13626 12897 13628
rect 12953 13626 12977 13628
rect 13033 13626 13057 13628
rect 12895 13574 12897 13626
rect 12959 13574 12971 13626
rect 13033 13574 13035 13626
rect 12873 13572 12897 13574
rect 12953 13572 12977 13574
rect 13033 13572 13057 13574
rect 12817 13552 13113 13572
rect 12817 12540 13113 12560
rect 12873 12538 12897 12540
rect 12953 12538 12977 12540
rect 13033 12538 13057 12540
rect 12895 12486 12897 12538
rect 12959 12486 12971 12538
rect 13033 12486 13035 12538
rect 12873 12484 12897 12486
rect 12953 12484 12977 12486
rect 13033 12484 13057 12486
rect 12817 12464 13113 12484
rect 12817 11452 13113 11472
rect 12873 11450 12897 11452
rect 12953 11450 12977 11452
rect 13033 11450 13057 11452
rect 12895 11398 12897 11450
rect 12959 11398 12971 11450
rect 13033 11398 13035 11450
rect 12873 11396 12897 11398
rect 12953 11396 12977 11398
rect 13033 11396 13057 11398
rect 12817 11376 13113 11396
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13556 10810 13584 11154
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 12817 10364 13113 10384
rect 12873 10362 12897 10364
rect 12953 10362 12977 10364
rect 13033 10362 13057 10364
rect 12895 10310 12897 10362
rect 12959 10310 12971 10362
rect 13033 10310 13035 10362
rect 12873 10308 12897 10310
rect 12953 10308 12977 10310
rect 13033 10308 13057 10310
rect 12817 10288 13113 10308
rect 13188 9994 13216 10406
rect 13280 10062 13308 10610
rect 13360 10532 13412 10538
rect 13360 10474 13412 10480
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13176 9988 13228 9994
rect 13176 9930 13228 9936
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12360 9438 12480 9466
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 12360 9058 12388 9438
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12452 9178 12480 9318
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12544 9110 12572 9862
rect 13280 9586 13308 9998
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12636 9382 12664 9454
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12817 9276 13113 9296
rect 12873 9274 12897 9276
rect 12953 9274 12977 9276
rect 13033 9274 13057 9276
rect 12895 9222 12897 9274
rect 12959 9222 12971 9274
rect 13033 9222 13035 9274
rect 12873 9220 12897 9222
rect 12953 9220 12977 9222
rect 13033 9220 13057 9222
rect 12817 9200 13113 9220
rect 13280 9110 13308 9386
rect 12532 9104 12584 9110
rect 12360 9030 12480 9058
rect 12532 9046 12584 9052
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12360 7886 12388 8774
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12346 7576 12402 7585
rect 12346 7511 12348 7520
rect 12400 7511 12402 7520
rect 12348 7482 12400 7488
rect 12164 7472 12216 7478
rect 12216 7432 12296 7460
rect 12164 7414 12216 7420
rect 12268 7392 12296 7432
rect 12268 7364 12388 7392
rect 12360 7313 12388 7364
rect 12346 7304 12402 7313
rect 11980 7268 12032 7274
rect 12084 7262 12296 7290
rect 11980 7210 12032 7216
rect 11992 7002 12020 7210
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11900 6186 11928 6802
rect 12084 6798 12112 7142
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11888 6180 11940 6186
rect 11888 6122 11940 6128
rect 11992 5710 12020 6598
rect 12070 5808 12126 5817
rect 12268 5778 12296 7262
rect 12346 7239 12402 7248
rect 12360 7002 12388 7239
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12452 6882 12480 9030
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12820 8378 12848 8842
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 12636 8350 12848 8378
rect 12636 7342 12664 8350
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 12728 8022 12756 8230
rect 12817 8188 13113 8208
rect 12873 8186 12897 8188
rect 12953 8186 12977 8188
rect 13033 8186 13057 8188
rect 12895 8134 12897 8186
rect 12959 8134 12971 8186
rect 13033 8134 13035 8186
rect 12873 8132 12897 8134
rect 12953 8132 12977 8134
rect 13033 8132 13057 8134
rect 12817 8112 13113 8132
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12992 8016 13044 8022
rect 12992 7958 13044 7964
rect 12728 7478 12756 7958
rect 12806 7848 12862 7857
rect 12806 7783 12808 7792
rect 12860 7783 12862 7792
rect 12808 7754 12860 7760
rect 12716 7472 12768 7478
rect 12716 7414 12768 7420
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12728 6882 12756 7414
rect 12820 7274 12848 7754
rect 13004 7546 13032 7958
rect 13084 7948 13136 7954
rect 13084 7890 13136 7896
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 13096 7410 13124 7890
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 13188 7342 13216 8230
rect 13280 7546 13308 8774
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 12817 7100 13113 7120
rect 12873 7098 12897 7100
rect 12953 7098 12977 7100
rect 13033 7098 13057 7100
rect 12895 7046 12897 7098
rect 12959 7046 12971 7098
rect 13033 7046 13035 7098
rect 12873 7044 12897 7046
rect 12953 7044 12977 7046
rect 13033 7044 13057 7046
rect 12817 7024 13113 7044
rect 13268 6928 13320 6934
rect 12452 6854 12664 6882
rect 12728 6854 12848 6882
rect 13372 6905 13400 10474
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13556 8838 13584 10202
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13648 8566 13676 13806
rect 13832 13734 13860 14418
rect 14200 14074 14228 14418
rect 14292 14346 14320 14418
rect 14280 14340 14332 14346
rect 14280 14282 14332 14288
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14096 11076 14148 11082
rect 14096 11018 14148 11024
rect 14004 10532 14056 10538
rect 14004 10474 14056 10480
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10266 13768 10406
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13464 7154 13492 8502
rect 13740 8498 13768 8910
rect 13832 8838 13860 9930
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13924 9489 13952 9862
rect 13910 9480 13966 9489
rect 13910 9415 13966 9424
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13740 8022 13768 8434
rect 13832 8294 13860 8570
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13556 7410 13584 7686
rect 13832 7585 13860 7890
rect 13818 7576 13874 7585
rect 13818 7511 13874 7520
rect 13820 7472 13872 7478
rect 13726 7440 13782 7449
rect 13544 7404 13596 7410
rect 13820 7414 13872 7420
rect 13726 7375 13782 7384
rect 13544 7346 13596 7352
rect 13636 7200 13688 7206
rect 13464 7126 13584 7154
rect 13636 7142 13688 7148
rect 13268 6870 13320 6876
rect 13358 6896 13414 6905
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12070 5743 12126 5752
rect 12256 5772 12308 5778
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 12084 5642 12112 5743
rect 12256 5714 12308 5720
rect 12360 5642 12388 6054
rect 12072 5636 12124 5642
rect 12072 5578 12124 5584
rect 12348 5636 12400 5642
rect 12348 5578 12400 5584
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 11888 5296 11940 5302
rect 11888 5238 11940 5244
rect 11900 4486 11928 5238
rect 12452 4622 12480 5578
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12544 4826 12572 5102
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11900 3602 11928 3878
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11992 3534 12020 4014
rect 12360 3670 12388 4218
rect 12440 4004 12492 4010
rect 12440 3946 12492 3952
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 12452 3534 12480 3946
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11164 2264 11560 2292
rect 11624 2746 11744 2774
rect 10692 2100 10744 2106
rect 10692 2042 10744 2048
rect 11164 800 11192 2264
rect 11624 800 11652 2746
rect 11992 2446 12020 3334
rect 12084 2582 12112 3402
rect 12072 2576 12124 2582
rect 12072 2518 12124 2524
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 12176 800 12204 3402
rect 12544 3194 12572 3606
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12440 2916 12492 2922
rect 12440 2858 12492 2864
rect 12452 2650 12480 2858
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12636 2446 12664 6854
rect 12820 6798 12848 6854
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13096 6644 13124 6734
rect 13004 6616 13124 6644
rect 13004 6186 13032 6616
rect 13174 6488 13230 6497
rect 13174 6423 13230 6432
rect 13188 6390 13216 6423
rect 13176 6384 13228 6390
rect 13176 6326 13228 6332
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 12817 6012 13113 6032
rect 12873 6010 12897 6012
rect 12953 6010 12977 6012
rect 13033 6010 13057 6012
rect 12895 5958 12897 6010
rect 12959 5958 12971 6010
rect 13033 5958 13035 6010
rect 12873 5956 12897 5958
rect 12953 5956 12977 5958
rect 13033 5956 13057 5958
rect 12817 5936 13113 5956
rect 13188 5710 13216 6190
rect 13280 5778 13308 6870
rect 13358 6831 13414 6840
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13280 5234 13308 5714
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12728 4826 12756 4966
rect 12817 4924 13113 4944
rect 12873 4922 12897 4924
rect 12953 4922 12977 4924
rect 13033 4922 13057 4924
rect 12895 4870 12897 4922
rect 12959 4870 12971 4922
rect 13033 4870 13035 4922
rect 12873 4868 12897 4870
rect 12953 4868 12977 4870
rect 13033 4868 13057 4870
rect 12817 4848 13113 4868
rect 12716 4820 12768 4826
rect 13360 4820 13412 4826
rect 12716 4762 12768 4768
rect 13280 4780 13360 4808
rect 13176 4752 13228 4758
rect 13280 4740 13308 4780
rect 13360 4762 13412 4768
rect 13228 4712 13308 4740
rect 13450 4720 13506 4729
rect 13176 4694 13228 4700
rect 13450 4655 13506 4664
rect 13464 4486 13492 4655
rect 13556 4622 13584 7126
rect 13648 7002 13676 7142
rect 13740 7041 13768 7375
rect 13726 7032 13782 7041
rect 13636 6996 13688 7002
rect 13726 6967 13782 6976
rect 13636 6938 13688 6944
rect 13832 6934 13860 7414
rect 13820 6928 13872 6934
rect 13726 6896 13782 6905
rect 13820 6870 13872 6876
rect 13726 6831 13782 6840
rect 13740 6225 13768 6831
rect 13726 6216 13782 6225
rect 13726 6151 13782 6160
rect 13924 5778 13952 9415
rect 14016 9382 14044 10474
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14016 8974 14044 9318
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 14004 8832 14056 8838
rect 14004 8774 14056 8780
rect 14016 7993 14044 8774
rect 14108 8022 14136 11018
rect 14096 8016 14148 8022
rect 14002 7984 14058 7993
rect 14096 7958 14148 7964
rect 14002 7919 14058 7928
rect 14016 7698 14044 7919
rect 14016 7670 14136 7698
rect 14004 7268 14056 7274
rect 14004 7210 14056 7216
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 13924 5574 13952 5714
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 14016 5234 14044 7210
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 14108 5166 14136 7670
rect 13820 5160 13872 5166
rect 13818 5128 13820 5137
rect 14096 5160 14148 5166
rect 13872 5128 13874 5137
rect 14096 5102 14148 5108
rect 13818 5063 13874 5072
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 13832 4690 13860 4966
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13912 4548 13964 4554
rect 13912 4490 13964 4496
rect 13452 4480 13504 4486
rect 13452 4422 13504 4428
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12728 1442 12756 4082
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 12817 3836 13113 3856
rect 12873 3834 12897 3836
rect 12953 3834 12977 3836
rect 13033 3834 13057 3836
rect 12895 3782 12897 3834
rect 12959 3782 12971 3834
rect 13033 3782 13035 3834
rect 12873 3780 12897 3782
rect 12953 3780 12977 3782
rect 13033 3780 13057 3782
rect 12817 3760 13113 3780
rect 12806 3496 12862 3505
rect 12806 3431 12862 3440
rect 12820 2990 12848 3431
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13004 3097 13032 3130
rect 12990 3088 13046 3097
rect 12990 3023 13046 3032
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 12817 2748 13113 2768
rect 12873 2746 12897 2748
rect 12953 2746 12977 2748
rect 13033 2746 13057 2748
rect 12895 2694 12897 2746
rect 12959 2694 12971 2746
rect 13033 2694 13035 2746
rect 12873 2692 12897 2694
rect 12953 2692 12977 2694
rect 13033 2692 13057 2694
rect 12817 2672 13113 2692
rect 13188 2582 13216 3878
rect 13372 3602 13400 3878
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13648 3466 13676 3946
rect 13924 3738 13952 4490
rect 14016 4078 14044 4966
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13280 2922 13308 3334
rect 13450 3088 13506 3097
rect 13740 3058 13768 3334
rect 13832 3194 13860 3470
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13450 3023 13506 3032
rect 13728 3052 13780 3058
rect 13268 2916 13320 2922
rect 13268 2858 13320 2864
rect 13464 2582 13492 3023
rect 13728 2994 13780 3000
rect 13832 2938 13860 3130
rect 13648 2910 13860 2938
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 13452 2576 13504 2582
rect 13452 2518 13504 2524
rect 13176 1760 13228 1766
rect 13176 1702 13228 1708
rect 12636 1414 12756 1442
rect 12636 800 12664 1414
rect 13188 800 13216 1702
rect 13648 800 13676 2910
rect 13924 2310 13952 3538
rect 14016 2774 14044 4014
rect 14016 2746 14136 2774
rect 13912 2304 13964 2310
rect 13912 2246 13964 2252
rect 13924 1766 13952 2246
rect 13912 1760 13964 1766
rect 13912 1702 13964 1708
rect 14108 800 14136 2746
rect 14200 2582 14228 13126
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14384 7750 14412 9454
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 14278 7440 14334 7449
rect 14278 7375 14334 7384
rect 14292 6866 14320 7375
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14292 6497 14320 6802
rect 14384 6798 14412 7278
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14278 6488 14334 6497
rect 14278 6423 14334 6432
rect 14384 5710 14412 6734
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14476 4690 14504 14214
rect 14844 13870 14872 14418
rect 15028 14074 15056 15030
rect 15120 14550 15148 16400
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15108 14544 15160 14550
rect 15108 14486 15160 14492
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14292 4010 14320 4422
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14476 3369 14504 3538
rect 14462 3360 14518 3369
rect 14462 3295 14518 3304
rect 14278 3224 14334 3233
rect 14278 3159 14334 3168
rect 14292 3058 14320 3159
rect 14476 3097 14504 3295
rect 14462 3088 14518 3097
rect 14280 3052 14332 3058
rect 14462 3023 14518 3032
rect 14280 2994 14332 3000
rect 14568 2922 14596 13194
rect 14740 9444 14792 9450
rect 14740 9386 14792 9392
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14660 8498 14688 9114
rect 14752 8945 14780 9386
rect 14738 8936 14794 8945
rect 14738 8871 14794 8880
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14660 7954 14688 8434
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14660 6225 14688 7754
rect 14646 6216 14702 6225
rect 14646 6151 14702 6160
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14660 5778 14688 6054
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14646 5672 14702 5681
rect 14646 5607 14702 5616
rect 14660 5370 14688 5607
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 14646 5264 14702 5273
rect 14646 5199 14702 5208
rect 14660 5166 14688 5199
rect 14648 5160 14700 5166
rect 14752 5137 14780 8871
rect 14648 5102 14700 5108
rect 14738 5128 14794 5137
rect 14738 5063 14794 5072
rect 14648 4752 14700 4758
rect 14648 4694 14700 4700
rect 14556 2916 14608 2922
rect 14556 2858 14608 2864
rect 14188 2576 14240 2582
rect 14188 2518 14240 2524
rect 14660 800 14688 4694
rect 14844 4146 14872 13806
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14936 10674 14964 10950
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14936 10130 14964 10610
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 14752 3126 14780 3538
rect 14740 3120 14792 3126
rect 14740 3062 14792 3068
rect 14936 2961 14964 8774
rect 15028 7002 15056 9386
rect 15016 6996 15068 7002
rect 15016 6938 15068 6944
rect 15120 5370 15148 11698
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15212 6254 15240 7482
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15198 6080 15254 6089
rect 15198 6015 15254 6024
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15212 5250 15240 6015
rect 15120 5222 15240 5250
rect 15120 5030 15148 5222
rect 15304 5166 15332 14894
rect 15764 14550 15792 16400
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15396 14074 15424 14350
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15396 9518 15424 9862
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15396 9178 15424 9454
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15384 8016 15436 8022
rect 15384 7958 15436 7964
rect 15396 7546 15424 7958
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15396 7342 15424 7482
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15396 7002 15424 7142
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15396 5642 15424 6802
rect 15384 5636 15436 5642
rect 15384 5578 15436 5584
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 15200 5092 15252 5098
rect 15200 5034 15252 5040
rect 15108 5024 15160 5030
rect 15108 4966 15160 4972
rect 15212 4808 15240 5034
rect 15028 4780 15240 4808
rect 15028 4026 15056 4780
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15120 4282 15148 4626
rect 15396 4593 15424 5306
rect 15382 4584 15438 4593
rect 15292 4548 15344 4554
rect 15382 4519 15438 4528
rect 15292 4490 15344 4496
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15108 4276 15160 4282
rect 15108 4218 15160 4224
rect 15028 3998 15148 4026
rect 15212 4010 15240 4422
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 15028 3602 15056 3878
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 14922 2952 14978 2961
rect 14922 2887 14978 2896
rect 15120 800 15148 3998
rect 15200 4004 15252 4010
rect 15200 3946 15252 3952
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15212 2650 15240 3470
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15304 2582 15332 4490
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15396 4146 15424 4422
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15488 3058 15516 14214
rect 15580 13870 15608 14418
rect 15782 14172 16078 14192
rect 15838 14170 15862 14172
rect 15918 14170 15942 14172
rect 15998 14170 16022 14172
rect 15860 14118 15862 14170
rect 15924 14118 15936 14170
rect 15998 14118 16000 14170
rect 15838 14116 15862 14118
rect 15918 14116 15942 14118
rect 15998 14116 16022 14118
rect 15782 14096 16078 14116
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15764 13870 15792 13942
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15580 4214 15608 13806
rect 15782 13084 16078 13104
rect 15838 13082 15862 13084
rect 15918 13082 15942 13084
rect 15998 13082 16022 13084
rect 15860 13030 15862 13082
rect 15924 13030 15936 13082
rect 15998 13030 16000 13082
rect 15838 13028 15862 13030
rect 15918 13028 15942 13030
rect 15998 13028 16022 13030
rect 15782 13008 16078 13028
rect 15782 11996 16078 12016
rect 15838 11994 15862 11996
rect 15918 11994 15942 11996
rect 15998 11994 16022 11996
rect 15860 11942 15862 11994
rect 15924 11942 15936 11994
rect 15998 11942 16000 11994
rect 15838 11940 15862 11942
rect 15918 11940 15942 11942
rect 15998 11940 16022 11942
rect 15782 11920 16078 11940
rect 16132 11642 16160 14486
rect 16408 14346 16436 16400
rect 16578 16008 16634 16017
rect 16578 15943 16634 15952
rect 16592 14482 16620 15943
rect 16946 15600 17002 15609
rect 16946 15535 17002 15544
rect 16960 14550 16988 15535
rect 17052 14822 17080 16400
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17040 14816 17092 14822
rect 17040 14758 17092 14764
rect 17236 14618 17264 14894
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 16948 14544 17000 14550
rect 16948 14486 17000 14492
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16396 14340 16448 14346
rect 16396 14282 16448 14288
rect 16592 14074 16620 14418
rect 16764 14340 16816 14346
rect 16764 14282 16816 14288
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16040 11614 16160 11642
rect 16040 11150 16068 11614
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15782 10908 16078 10928
rect 15838 10906 15862 10908
rect 15918 10906 15942 10908
rect 15998 10906 16022 10908
rect 15860 10854 15862 10906
rect 15924 10854 15936 10906
rect 15998 10854 16000 10906
rect 15838 10852 15862 10854
rect 15918 10852 15942 10854
rect 15998 10852 16022 10854
rect 15782 10832 16078 10852
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 15782 9820 16078 9840
rect 15838 9818 15862 9820
rect 15918 9818 15942 9820
rect 15998 9818 16022 9820
rect 15860 9766 15862 9818
rect 15924 9766 15936 9818
rect 15998 9766 16000 9818
rect 15838 9764 15862 9766
rect 15918 9764 15942 9766
rect 15998 9764 16022 9766
rect 15782 9744 16078 9764
rect 16132 9704 16160 9862
rect 16040 9676 16160 9704
rect 15660 9648 15712 9654
rect 15658 9616 15660 9625
rect 15712 9616 15714 9625
rect 15658 9551 15714 9560
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15948 9178 15976 9318
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15660 9104 15712 9110
rect 16040 9081 16068 9676
rect 16224 9466 16252 13806
rect 16408 13190 16436 13806
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 16132 9438 16252 9466
rect 15660 9046 15712 9052
rect 16026 9072 16082 9081
rect 15672 8514 15700 9046
rect 16026 9007 16082 9016
rect 15782 8732 16078 8752
rect 15838 8730 15862 8732
rect 15918 8730 15942 8732
rect 15998 8730 16022 8732
rect 15860 8678 15862 8730
rect 15924 8678 15936 8730
rect 15998 8678 16000 8730
rect 15838 8676 15862 8678
rect 15918 8676 15942 8678
rect 15998 8676 16022 8678
rect 15782 8656 16078 8676
rect 15672 8498 15884 8514
rect 15672 8492 15896 8498
rect 15672 8486 15844 8492
rect 15844 8434 15896 8440
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15660 8356 15712 8362
rect 15660 8298 15712 8304
rect 15672 8129 15700 8298
rect 15764 8294 15792 8366
rect 15856 8294 15884 8434
rect 15752 8288 15804 8294
rect 15752 8230 15804 8236
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15658 8120 15714 8129
rect 15658 8055 15714 8064
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15672 7342 15700 7890
rect 15782 7644 16078 7664
rect 15838 7642 15862 7644
rect 15918 7642 15942 7644
rect 15998 7642 16022 7644
rect 15860 7590 15862 7642
rect 15924 7590 15936 7642
rect 15998 7590 16000 7642
rect 15838 7588 15862 7590
rect 15918 7588 15942 7590
rect 15998 7588 16022 7590
rect 15782 7568 16078 7588
rect 16132 7562 16160 9438
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16224 9178 16252 9318
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16212 8900 16264 8906
rect 16212 8842 16264 8848
rect 16224 8634 16252 8842
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16316 8514 16344 11086
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16500 10266 16528 10610
rect 16592 10470 16620 12106
rect 16776 10742 16804 14282
rect 16960 14074 16988 14486
rect 17420 14482 17448 16759
rect 17498 16416 17554 16425
rect 17682 16400 17738 17200
rect 18326 16400 18382 17200
rect 18970 16400 19026 17200
rect 19614 16400 19670 17200
rect 17498 16351 17554 16360
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 17040 13796 17092 13802
rect 17040 13738 17092 13744
rect 17052 13530 17080 13738
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16948 13252 17000 13258
rect 16948 13194 17000 13200
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16764 10736 16816 10742
rect 16764 10678 16816 10684
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16868 10554 16896 12786
rect 16960 11014 16988 13194
rect 17328 11558 17356 14214
rect 17420 12986 17448 14418
rect 17512 13734 17540 16351
rect 17696 14890 17724 16400
rect 17774 15192 17830 15201
rect 17774 15127 17830 15136
rect 17684 14884 17736 14890
rect 17684 14826 17736 14832
rect 17788 14550 17816 15127
rect 17866 14784 17922 14793
rect 17866 14719 17922 14728
rect 17880 14550 17908 14719
rect 17776 14544 17828 14550
rect 17696 14504 17776 14532
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17512 13530 17540 13670
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17696 13462 17724 14504
rect 17776 14486 17828 14492
rect 17868 14544 17920 14550
rect 17868 14486 17920 14492
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17684 13456 17736 13462
rect 17684 13398 17736 13404
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17512 12434 17540 12582
rect 17788 12434 17816 14214
rect 17880 13530 17908 14486
rect 18144 14340 18196 14346
rect 18144 14282 18196 14288
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 18052 12708 18104 12714
rect 18052 12650 18104 12656
rect 18064 12617 18092 12650
rect 18050 12608 18106 12617
rect 18050 12543 18106 12552
rect 18156 12434 18184 14282
rect 18340 14074 18368 16400
rect 18420 14476 18472 14482
rect 18420 14418 18472 14424
rect 18432 14249 18460 14418
rect 18418 14240 18474 14249
rect 18418 14175 18474 14184
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18984 13870 19012 16400
rect 18420 13864 18472 13870
rect 18418 13832 18420 13841
rect 18972 13864 19024 13870
rect 18472 13832 18474 13841
rect 18972 13806 19024 13812
rect 18418 13767 18474 13776
rect 19628 13462 19656 16400
rect 19616 13456 19668 13462
rect 18418 13424 18474 13433
rect 19616 13398 19668 13404
rect 18418 13359 18420 13368
rect 18472 13359 18474 13368
rect 18420 13330 18472 13336
rect 18418 13016 18474 13025
rect 18418 12951 18474 12960
rect 18432 12782 18460 12951
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 17420 12406 17540 12434
rect 17604 12406 17816 12434
rect 17972 12406 18184 12434
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16684 10266 16712 10542
rect 16868 10526 17080 10554
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 16408 8838 16436 9658
rect 16500 9586 16528 10202
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 16488 8968 16540 8974
rect 16592 8956 16620 9658
rect 16684 9330 16712 10202
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16776 9518 16804 9862
rect 16854 9616 16910 9625
rect 16854 9551 16910 9560
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16684 9302 16804 9330
rect 16540 8928 16620 8956
rect 16672 8968 16724 8974
rect 16488 8910 16540 8916
rect 16672 8910 16724 8916
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16408 8634 16436 8774
rect 16684 8634 16712 8910
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16212 8492 16264 8498
rect 16316 8486 16528 8514
rect 16212 8434 16264 8440
rect 16224 8106 16252 8434
rect 16302 8120 16358 8129
rect 16224 8078 16302 8106
rect 16302 8055 16304 8064
rect 16356 8055 16358 8064
rect 16304 8026 16356 8032
rect 16500 7750 16528 8486
rect 16776 8362 16804 9302
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16684 8090 16712 8230
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16304 7744 16356 7750
rect 16488 7744 16540 7750
rect 16356 7704 16436 7732
rect 16304 7686 16356 7692
rect 16132 7534 16252 7562
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15672 6322 15700 7278
rect 15750 6896 15806 6905
rect 15750 6831 15752 6840
rect 15804 6831 15806 6840
rect 15752 6802 15804 6808
rect 15856 6769 15884 7278
rect 16120 6996 16172 7002
rect 16120 6938 16172 6944
rect 15842 6760 15898 6769
rect 15842 6695 15898 6704
rect 15782 6556 16078 6576
rect 15838 6554 15862 6556
rect 15918 6554 15942 6556
rect 15998 6554 16022 6556
rect 15860 6502 15862 6554
rect 15924 6502 15936 6554
rect 15998 6502 16000 6554
rect 15838 6500 15862 6502
rect 15918 6500 15942 6502
rect 15998 6500 16022 6502
rect 15782 6480 16078 6500
rect 16132 6322 16160 6938
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15856 5914 15884 6054
rect 16040 5914 16068 6190
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 15672 5778 15700 5850
rect 16040 5778 16068 5850
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 15672 5370 15700 5714
rect 15782 5468 16078 5488
rect 15838 5466 15862 5468
rect 15918 5466 15942 5468
rect 15998 5466 16022 5468
rect 15860 5414 15862 5466
rect 15924 5414 15936 5466
rect 15998 5414 16000 5466
rect 15838 5412 15862 5414
rect 15918 5412 15942 5414
rect 15998 5412 16022 5414
rect 15782 5392 16078 5412
rect 16132 5370 16160 6054
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15672 4264 15700 5102
rect 15752 5092 15804 5098
rect 15752 5034 15804 5040
rect 15764 4690 15792 5034
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15750 4584 15806 4593
rect 15750 4519 15752 4528
rect 15804 4519 15806 4528
rect 15752 4490 15804 4496
rect 15782 4380 16078 4400
rect 15838 4378 15862 4380
rect 15918 4378 15942 4380
rect 15998 4378 16022 4380
rect 15860 4326 15862 4378
rect 15924 4326 15936 4378
rect 15998 4326 16000 4378
rect 15838 4324 15862 4326
rect 15918 4324 15942 4326
rect 15998 4324 16022 4326
rect 15782 4304 16078 4324
rect 16132 4282 16160 4966
rect 16120 4276 16172 4282
rect 15672 4236 15792 4264
rect 15568 4208 15620 4214
rect 15568 4150 15620 4156
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15672 3738 15700 4082
rect 15764 4078 15792 4236
rect 16120 4218 16172 4224
rect 15936 4208 15988 4214
rect 15936 4150 15988 4156
rect 15948 4078 15976 4150
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 15580 2378 15608 3402
rect 15672 3194 15700 3538
rect 15782 3292 16078 3312
rect 15838 3290 15862 3292
rect 15918 3290 15942 3292
rect 15998 3290 16022 3292
rect 15860 3238 15862 3290
rect 15924 3238 15936 3290
rect 15998 3238 16000 3290
rect 15838 3236 15862 3238
rect 15918 3236 15942 3238
rect 15998 3236 16022 3238
rect 15782 3216 16078 3236
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15750 3088 15806 3097
rect 15750 3023 15752 3032
rect 15804 3023 15806 3032
rect 15752 2994 15804 3000
rect 16224 2582 16252 7534
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16316 7002 16344 7142
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16408 6746 16436 7704
rect 16488 7686 16540 7692
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16500 7342 16528 7686
rect 16488 7336 16540 7342
rect 16672 7336 16724 7342
rect 16488 7278 16540 7284
rect 16670 7304 16672 7313
rect 16724 7304 16726 7313
rect 16670 7239 16726 7248
rect 16580 6996 16632 7002
rect 16580 6938 16632 6944
rect 16592 6866 16620 6938
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16316 6718 16436 6746
rect 16488 6724 16540 6730
rect 16316 5370 16344 6718
rect 16488 6666 16540 6672
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 16408 6118 16436 6598
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16408 5817 16436 6054
rect 16394 5808 16450 5817
rect 16394 5743 16450 5752
rect 16500 5710 16528 6666
rect 16684 6662 16712 6802
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16670 6352 16726 6361
rect 16670 6287 16672 6296
rect 16724 6287 16726 6296
rect 16672 6258 16724 6264
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16592 6118 16620 6190
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16316 5234 16344 5306
rect 16396 5296 16448 5302
rect 16396 5238 16448 5244
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16316 3602 16344 4626
rect 16408 3602 16436 5238
rect 16500 5234 16528 5646
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16592 4826 16620 5714
rect 16776 5681 16804 7686
rect 16868 6390 16896 9551
rect 16960 9042 16988 10406
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16948 8560 17000 8566
rect 16948 8502 17000 8508
rect 16960 8362 16988 8502
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 16960 8090 16988 8298
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 17052 7460 17080 10526
rect 17144 10062 17172 10950
rect 17224 10736 17276 10742
rect 17224 10678 17276 10684
rect 17132 10056 17184 10062
rect 17132 9998 17184 10004
rect 17144 7886 17172 9998
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 16960 7432 17080 7460
rect 16960 7002 16988 7432
rect 17236 7392 17264 10678
rect 17328 9994 17356 11494
rect 17316 9988 17368 9994
rect 17316 9930 17368 9936
rect 17314 9616 17370 9625
rect 17420 9586 17448 12406
rect 17604 10554 17632 12406
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17880 11354 17908 11630
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17776 11076 17828 11082
rect 17776 11018 17828 11024
rect 17788 10674 17816 11018
rect 17776 10668 17828 10674
rect 17776 10610 17828 10616
rect 17512 10526 17632 10554
rect 17684 10532 17736 10538
rect 17314 9551 17370 9560
rect 17408 9580 17460 9586
rect 17328 9450 17356 9551
rect 17408 9522 17460 9528
rect 17316 9444 17368 9450
rect 17316 9386 17368 9392
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17328 8022 17356 8910
rect 17420 8090 17448 9318
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17316 8016 17368 8022
rect 17316 7958 17368 7964
rect 17052 7364 17264 7392
rect 16948 6996 17000 7002
rect 16948 6938 17000 6944
rect 17052 6882 17080 7364
rect 17328 7324 17356 7958
rect 17512 7449 17540 10526
rect 17684 10474 17736 10480
rect 17868 10532 17920 10538
rect 17868 10474 17920 10480
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 17604 10266 17632 10406
rect 17696 10266 17724 10474
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17604 9586 17632 10066
rect 17788 9722 17816 10406
rect 17880 10033 17908 10474
rect 17972 10198 18000 12406
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 18064 12209 18092 12242
rect 18050 12200 18106 12209
rect 18050 12135 18106 12144
rect 18432 11801 18460 12242
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18418 11792 18474 11801
rect 18418 11727 18474 11736
rect 18420 11620 18472 11626
rect 18420 11562 18472 11568
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 18064 10266 18092 11086
rect 18144 10532 18196 10538
rect 18144 10474 18196 10480
rect 18156 10441 18184 10474
rect 18142 10432 18198 10441
rect 18142 10367 18198 10376
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 17866 10024 17922 10033
rect 17866 9959 17922 9968
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17592 9580 17644 9586
rect 17644 9540 17724 9568
rect 17592 9522 17644 9528
rect 17696 9042 17724 9540
rect 17788 9178 17816 9658
rect 18064 9654 18092 9685
rect 18052 9648 18104 9654
rect 18050 9616 18052 9625
rect 18104 9616 18106 9625
rect 18050 9551 18106 9560
rect 18248 9568 18276 11494
rect 18432 11257 18460 11562
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 18418 11248 18474 11257
rect 18418 11183 18474 11192
rect 18512 11212 18564 11218
rect 18512 11154 18564 11160
rect 18524 10849 18552 11154
rect 18510 10840 18566 10849
rect 18510 10775 18566 10784
rect 18420 10532 18472 10538
rect 18420 10474 18472 10480
rect 18432 10033 18460 10474
rect 18418 10024 18474 10033
rect 18418 9959 18474 9968
rect 17866 9480 17922 9489
rect 18064 9450 18092 9551
rect 18248 9540 18368 9568
rect 17866 9415 17868 9424
rect 17920 9415 17922 9424
rect 18052 9444 18104 9450
rect 17868 9386 17920 9392
rect 18052 9386 18104 9392
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17604 8498 17632 8910
rect 18156 8498 18184 9386
rect 18236 8968 18288 8974
rect 18234 8936 18236 8945
rect 18288 8936 18290 8945
rect 18234 8871 18290 8880
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 17604 7868 17632 8434
rect 17776 8356 17828 8362
rect 17776 8298 17828 8304
rect 17788 7954 17816 8298
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17684 7880 17736 7886
rect 17604 7840 17684 7868
rect 17684 7822 17736 7828
rect 17972 7546 18000 8026
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17498 7440 17554 7449
rect 17498 7375 17554 7384
rect 18064 7342 18092 8230
rect 18248 8022 18276 8774
rect 18340 8430 18368 9540
rect 18420 9444 18472 9450
rect 18420 9386 18472 9392
rect 18432 9217 18460 9386
rect 18418 9208 18474 9217
rect 18418 9143 18474 9152
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18432 8809 18460 8978
rect 18418 8800 18474 8809
rect 18418 8735 18474 8744
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18524 8265 18552 8298
rect 18510 8256 18566 8265
rect 18510 8191 18566 8200
rect 18236 8016 18288 8022
rect 18236 7958 18288 7964
rect 18510 7848 18566 7857
rect 18510 7783 18512 7792
rect 18564 7783 18566 7792
rect 18512 7754 18564 7760
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18328 7472 18380 7478
rect 18142 7440 18198 7449
rect 18328 7414 18380 7420
rect 18142 7375 18144 7384
rect 18196 7375 18198 7384
rect 18144 7346 18196 7352
rect 17408 7336 17460 7342
rect 17328 7296 17408 7324
rect 17408 7278 17460 7284
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 17224 7268 17276 7274
rect 17224 7210 17276 7216
rect 17500 7268 17552 7274
rect 17500 7210 17552 7216
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 17144 7002 17172 7142
rect 17132 6996 17184 7002
rect 17132 6938 17184 6944
rect 16960 6854 17080 6882
rect 16960 6798 16988 6854
rect 16948 6792 17000 6798
rect 17132 6792 17184 6798
rect 16948 6734 17000 6740
rect 17130 6760 17132 6769
rect 17184 6760 17186 6769
rect 17236 6730 17264 7210
rect 17316 6928 17368 6934
rect 17316 6870 17368 6876
rect 17130 6695 17186 6704
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 16856 6384 16908 6390
rect 16856 6326 16908 6332
rect 17224 6180 17276 6186
rect 17224 6122 17276 6128
rect 17236 5710 17264 6122
rect 17328 5846 17356 6870
rect 17512 6458 17540 7210
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 17682 7032 17738 7041
rect 17682 6967 17738 6976
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17408 6384 17460 6390
rect 17408 6326 17460 6332
rect 17316 5840 17368 5846
rect 17316 5782 17368 5788
rect 17224 5704 17276 5710
rect 16762 5672 16818 5681
rect 16818 5630 16988 5658
rect 17224 5646 17276 5652
rect 16762 5607 16818 5616
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16776 5352 16804 5510
rect 16684 5324 16804 5352
rect 16684 5166 16712 5324
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 16854 5128 16910 5137
rect 16764 5092 16816 5098
rect 16854 5063 16856 5072
rect 16764 5034 16816 5040
rect 16908 5063 16910 5072
rect 16856 5034 16908 5040
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16488 4752 16540 4758
rect 16488 4694 16540 4700
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16408 3058 16436 3334
rect 16500 3194 16528 4694
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16592 2990 16620 4422
rect 16776 4078 16804 5034
rect 16960 4690 16988 5630
rect 17236 5234 17264 5646
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17132 5160 17184 5166
rect 17132 5102 17184 5108
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 17052 4729 17080 4762
rect 17038 4720 17094 4729
rect 16948 4684 17000 4690
rect 17038 4655 17094 4664
rect 16948 4626 17000 4632
rect 17040 4548 17092 4554
rect 17040 4490 17092 4496
rect 16948 4276 17000 4282
rect 16948 4218 17000 4224
rect 16960 4078 16988 4218
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16684 3126 16712 3334
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16672 3120 16724 3126
rect 16672 3062 16724 3068
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 16764 2916 16816 2922
rect 16764 2858 16816 2864
rect 16500 2582 16528 2858
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 16488 2576 16540 2582
rect 16488 2518 16540 2524
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 15568 2372 15620 2378
rect 15568 2314 15620 2320
rect 15660 2372 15712 2378
rect 15660 2314 15712 2320
rect 15672 800 15700 2314
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 15782 2204 16078 2224
rect 15838 2202 15862 2204
rect 15918 2202 15942 2204
rect 15998 2202 16022 2204
rect 15860 2150 15862 2202
rect 15924 2150 15936 2202
rect 15998 2150 16000 2202
rect 15838 2148 15862 2150
rect 15918 2148 15942 2150
rect 15998 2148 16022 2150
rect 15782 2128 16078 2148
rect 16132 800 16160 2246
rect 16684 800 16712 2382
rect 16776 1154 16804 2858
rect 16868 2514 16896 3130
rect 16960 2582 16988 3674
rect 17052 3670 17080 4490
rect 17144 4078 17172 5102
rect 17236 4622 17264 5170
rect 17328 4758 17356 5782
rect 17420 5778 17448 6326
rect 17696 6254 17724 6967
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 17316 4752 17368 4758
rect 17316 4694 17368 4700
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17132 4072 17184 4078
rect 17184 4032 17264 4060
rect 17132 4014 17184 4020
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 17144 3738 17172 3878
rect 17132 3732 17184 3738
rect 17132 3674 17184 3680
rect 17040 3664 17092 3670
rect 17040 3606 17092 3612
rect 17236 3584 17264 4032
rect 17328 3942 17356 4082
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17144 3556 17264 3584
rect 17144 3194 17172 3556
rect 17224 3460 17276 3466
rect 17224 3402 17276 3408
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17236 2990 17264 3402
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17132 2984 17184 2990
rect 17132 2926 17184 2932
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 16948 2576 17000 2582
rect 16948 2518 17000 2524
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 16764 1148 16816 1154
rect 16764 1090 16816 1096
rect 17144 800 17172 2926
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 17420 1873 17448 2790
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 17406 1864 17462 1873
rect 17406 1799 17462 1808
rect 17512 1465 17540 2382
rect 17498 1456 17554 1465
rect 17498 1391 17554 1400
rect 17604 800 17632 3334
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17696 2446 17724 3130
rect 17788 3058 17816 7142
rect 18340 6866 18368 7414
rect 18328 6860 18380 6866
rect 18328 6802 18380 6808
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 18064 6254 18092 6598
rect 18052 6248 18104 6254
rect 18052 6190 18104 6196
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17866 5264 17922 5273
rect 17866 5199 17922 5208
rect 17880 5166 17908 5199
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17972 4758 18000 5510
rect 18064 4758 18092 5850
rect 18248 5846 18276 6054
rect 18236 5840 18288 5846
rect 18236 5782 18288 5788
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18142 4856 18198 4865
rect 18142 4791 18198 4800
rect 17960 4752 18012 4758
rect 17960 4694 18012 4700
rect 18052 4752 18104 4758
rect 18052 4694 18104 4700
rect 18156 4690 18184 4791
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17972 3670 18000 4422
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 17960 3664 18012 3670
rect 17960 3606 18012 3612
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17776 2916 17828 2922
rect 17776 2858 17828 2864
rect 17788 2689 17816 2858
rect 17774 2680 17830 2689
rect 17774 2615 17830 2624
rect 17880 2553 17908 3334
rect 18064 2582 18092 4082
rect 18248 4078 18276 4966
rect 18236 4072 18288 4078
rect 18142 4040 18198 4049
rect 18236 4014 18288 4020
rect 18142 3975 18144 3984
rect 18196 3975 18198 3984
rect 18144 3946 18196 3952
rect 18144 3460 18196 3466
rect 18144 3402 18196 3408
rect 18156 3233 18184 3402
rect 18142 3224 18198 3233
rect 18142 3159 18198 3168
rect 18052 2576 18104 2582
rect 17866 2544 17922 2553
rect 18052 2518 18104 2524
rect 18432 2514 18460 7686
rect 18512 7268 18564 7274
rect 18512 7210 18564 7216
rect 18524 7041 18552 7210
rect 18510 7032 18566 7041
rect 18510 6967 18566 6976
rect 18512 6724 18564 6730
rect 18512 6666 18564 6672
rect 18524 6633 18552 6666
rect 18510 6624 18566 6633
rect 18510 6559 18566 6568
rect 18510 6216 18566 6225
rect 18510 6151 18512 6160
rect 18564 6151 18566 6160
rect 18512 6122 18564 6128
rect 18510 5672 18566 5681
rect 18510 5607 18512 5616
rect 18564 5607 18566 5616
rect 18512 5578 18564 5584
rect 18510 5264 18566 5273
rect 18510 5199 18512 5208
rect 18564 5199 18566 5208
rect 18512 5170 18564 5176
rect 18616 5166 18644 11290
rect 18708 8090 18736 12038
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18800 4826 18828 11494
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18512 4548 18564 4554
rect 18512 4490 18564 4496
rect 18524 4457 18552 4490
rect 18510 4448 18566 4457
rect 18510 4383 18566 4392
rect 18512 4004 18564 4010
rect 18512 3946 18564 3952
rect 18524 3641 18552 3946
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 18510 3632 18566 3641
rect 18510 3567 18566 3576
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 17866 2479 17922 2488
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 17776 2372 17828 2378
rect 17776 2314 17828 2320
rect 17868 2372 17920 2378
rect 17868 2314 17920 2320
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 3330 232 3386 241
rect 3330 167 3386 176
rect 3606 0 3662 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5170 0 5226 800
rect 5630 0 5686 800
rect 6182 0 6238 800
rect 6642 0 6698 800
rect 7102 0 7158 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9126 0 9182 800
rect 9678 0 9734 800
rect 10138 0 10194 800
rect 10598 0 10654 800
rect 11150 0 11206 800
rect 11610 0 11666 800
rect 12162 0 12218 800
rect 12622 0 12678 800
rect 13174 0 13230 800
rect 13634 0 13690 800
rect 14094 0 14150 800
rect 14646 0 14702 800
rect 15106 0 15162 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16670 0 16726 800
rect 17130 0 17186 800
rect 17590 0 17646 800
rect 17696 649 17724 2246
rect 17788 1057 17816 2314
rect 17774 1048 17830 1057
rect 17774 983 17830 992
rect 17682 640 17738 649
rect 17682 575 17738 584
rect 17880 241 17908 2314
rect 18144 1148 18196 1154
rect 18144 1090 18196 1096
rect 18156 800 18184 1090
rect 18616 800 18644 3470
rect 19168 800 19196 3878
rect 19616 3596 19668 3602
rect 19616 3538 19668 3544
rect 19628 800 19656 3538
rect 17866 232 17922 241
rect 17866 167 17922 176
rect 18142 0 18198 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19614 0 19670 800
<< via2 >>
rect 1490 14476 1546 14512
rect 1490 14456 1492 14476
rect 1492 14456 1544 14476
rect 1544 14456 1546 14476
rect 1858 14728 1914 14784
rect 2594 15952 2650 16008
rect 2778 15544 2834 15600
rect 2594 13912 2650 13968
rect 1858 13504 1914 13560
rect 3146 16360 3202 16416
rect 3790 16768 3846 16824
rect 2962 15136 3018 15192
rect 2134 13232 2190 13288
rect 1490 13096 1546 13152
rect 1582 12708 1638 12744
rect 1582 12688 1584 12708
rect 1584 12688 1636 12708
rect 1636 12688 1638 12708
rect 1490 12280 1546 12336
rect 1490 11736 1546 11792
rect 1398 11328 1454 11384
rect 1490 10920 1546 10976
rect 1950 12688 2006 12744
rect 1674 10920 1730 10976
rect 1858 11872 1914 11928
rect 1582 10648 1638 10704
rect 1398 10512 1454 10568
rect 1490 10104 1546 10160
rect 1490 9288 1546 9344
rect 1398 8880 1454 8936
rect 1490 7692 1492 7712
rect 1492 7692 1544 7712
rect 1544 7692 1546 7712
rect 1490 7656 1546 7692
rect 2502 10920 2558 10976
rect 2134 9560 2190 9616
rect 1950 9324 1952 9344
rect 1952 9324 2004 9344
rect 2004 9324 2006 9344
rect 1950 9288 2006 9324
rect 1858 8084 1914 8120
rect 1858 8064 1860 8084
rect 1860 8064 1912 8084
rect 1912 8064 1914 8084
rect 1766 7792 1822 7848
rect 1398 7284 1400 7304
rect 1400 7284 1452 7304
rect 1452 7284 1454 7304
rect 1398 7248 1454 7284
rect 1766 6860 1822 6896
rect 1766 6840 1768 6860
rect 1768 6840 1820 6860
rect 1820 6840 1822 6860
rect 1490 6432 1546 6488
rect 1490 6060 1492 6080
rect 1492 6060 1544 6080
rect 1544 6060 1546 6080
rect 1490 6024 1546 6060
rect 1490 5516 1492 5536
rect 1492 5516 1544 5536
rect 1544 5516 1546 5536
rect 1490 5480 1546 5516
rect 1398 5108 1400 5128
rect 1400 5108 1452 5128
rect 1452 5108 1454 5128
rect 1398 5072 1454 5108
rect 1398 4684 1454 4720
rect 1398 4664 1400 4684
rect 1400 4664 1452 4684
rect 1452 4664 1454 4684
rect 1490 2624 1546 2680
rect 1858 4256 1914 4312
rect 1858 3440 1914 3496
rect 1398 1400 1454 1456
rect 2870 13640 2926 13696
rect 3330 14728 3386 14784
rect 3238 13796 3294 13832
rect 3238 13776 3240 13796
rect 3240 13776 3292 13796
rect 3292 13776 3294 13796
rect 3606 14476 3662 14512
rect 3606 14456 3608 14476
rect 3608 14456 3660 14476
rect 3660 14456 3662 14476
rect 17406 16768 17462 16824
rect 3921 14170 3977 14172
rect 4001 14170 4057 14172
rect 4081 14170 4137 14172
rect 4161 14170 4217 14172
rect 3921 14118 3947 14170
rect 3947 14118 3977 14170
rect 4001 14118 4011 14170
rect 4011 14118 4057 14170
rect 4081 14118 4127 14170
rect 4127 14118 4137 14170
rect 4161 14118 4191 14170
rect 4191 14118 4217 14170
rect 3921 14116 3977 14118
rect 4001 14116 4057 14118
rect 4081 14116 4137 14118
rect 4161 14116 4217 14118
rect 3882 13268 3884 13288
rect 3884 13268 3936 13288
rect 3936 13268 3938 13288
rect 3882 13232 3938 13268
rect 3921 13082 3977 13084
rect 4001 13082 4057 13084
rect 4081 13082 4137 13084
rect 4161 13082 4217 13084
rect 3921 13030 3947 13082
rect 3947 13030 3977 13082
rect 4001 13030 4011 13082
rect 4011 13030 4057 13082
rect 4081 13030 4127 13082
rect 4127 13030 4137 13082
rect 4161 13030 4191 13082
rect 4191 13030 4217 13082
rect 3921 13028 3977 13030
rect 4001 13028 4057 13030
rect 4081 13028 4137 13030
rect 4161 13028 4217 13030
rect 3238 11872 3294 11928
rect 3330 11736 3386 11792
rect 3054 10104 3110 10160
rect 2962 8508 2964 8528
rect 2964 8508 3016 8528
rect 3016 8508 3018 8528
rect 2962 8472 3018 8508
rect 2226 3884 2228 3904
rect 2228 3884 2280 3904
rect 2280 3884 2282 3904
rect 2226 3848 2282 3884
rect 2226 3032 2282 3088
rect 2594 5208 2650 5264
rect 1858 2216 1914 2272
rect 1766 992 1822 1048
rect 2226 1808 2282 1864
rect 3238 9696 3294 9752
rect 3238 9560 3294 9616
rect 3514 10512 3570 10568
rect 3514 9288 3570 9344
rect 3422 9016 3478 9072
rect 3921 11994 3977 11996
rect 4001 11994 4057 11996
rect 4081 11994 4137 11996
rect 4161 11994 4217 11996
rect 3921 11942 3947 11994
rect 3947 11942 3977 11994
rect 4001 11942 4011 11994
rect 4011 11942 4057 11994
rect 4081 11942 4127 11994
rect 4127 11942 4137 11994
rect 4161 11942 4191 11994
rect 4191 11942 4217 11994
rect 3921 11940 3977 11942
rect 4001 11940 4057 11942
rect 4081 11940 4137 11942
rect 4161 11940 4217 11942
rect 3921 10906 3977 10908
rect 4001 10906 4057 10908
rect 4081 10906 4137 10908
rect 4161 10906 4217 10908
rect 3921 10854 3947 10906
rect 3947 10854 3977 10906
rect 4001 10854 4011 10906
rect 4011 10854 4057 10906
rect 4081 10854 4127 10906
rect 4127 10854 4137 10906
rect 4161 10854 4191 10906
rect 4191 10854 4217 10906
rect 3921 10852 3977 10854
rect 4001 10852 4057 10854
rect 4081 10852 4137 10854
rect 4161 10852 4217 10854
rect 3921 9818 3977 9820
rect 4001 9818 4057 9820
rect 4081 9818 4137 9820
rect 4161 9818 4217 9820
rect 3921 9766 3947 9818
rect 3947 9766 3977 9818
rect 4001 9766 4011 9818
rect 4011 9766 4057 9818
rect 4081 9766 4127 9818
rect 4127 9766 4137 9818
rect 4161 9766 4191 9818
rect 4191 9766 4217 9818
rect 3921 9764 3977 9766
rect 4001 9764 4057 9766
rect 4081 9764 4137 9766
rect 4161 9764 4217 9766
rect 4066 9460 4068 9480
rect 4068 9460 4120 9480
rect 4120 9460 4122 9480
rect 4066 9424 4122 9460
rect 3974 8900 4030 8936
rect 3974 8880 3976 8900
rect 3976 8880 4028 8900
rect 4028 8880 4030 8900
rect 3146 6296 3202 6352
rect 3606 5752 3662 5808
rect 3921 8730 3977 8732
rect 4001 8730 4057 8732
rect 4081 8730 4137 8732
rect 4161 8730 4217 8732
rect 3921 8678 3947 8730
rect 3947 8678 3977 8730
rect 4001 8678 4011 8730
rect 4011 8678 4057 8730
rect 4081 8678 4127 8730
rect 4127 8678 4137 8730
rect 4161 8678 4191 8730
rect 4191 8678 4217 8730
rect 3921 8676 3977 8678
rect 4001 8676 4057 8678
rect 4081 8676 4137 8678
rect 4161 8676 4217 8678
rect 6886 14714 6942 14716
rect 6966 14714 7022 14716
rect 7046 14714 7102 14716
rect 7126 14714 7182 14716
rect 6886 14662 6912 14714
rect 6912 14662 6942 14714
rect 6966 14662 6976 14714
rect 6976 14662 7022 14714
rect 7046 14662 7092 14714
rect 7092 14662 7102 14714
rect 7126 14662 7156 14714
rect 7156 14662 7182 14714
rect 6886 14660 6942 14662
rect 6966 14660 7022 14662
rect 7046 14660 7102 14662
rect 7126 14660 7182 14662
rect 4618 13812 4620 13832
rect 4620 13812 4672 13832
rect 4672 13812 4674 13832
rect 4618 13776 4674 13812
rect 4710 13640 4766 13696
rect 4710 12688 4766 12744
rect 3921 7642 3977 7644
rect 4001 7642 4057 7644
rect 4081 7642 4137 7644
rect 4161 7642 4217 7644
rect 3921 7590 3947 7642
rect 3947 7590 3977 7642
rect 4001 7590 4011 7642
rect 4011 7590 4057 7642
rect 4081 7590 4127 7642
rect 4127 7590 4137 7642
rect 4161 7590 4191 7642
rect 4191 7590 4217 7642
rect 3921 7588 3977 7590
rect 4001 7588 4057 7590
rect 4081 7588 4137 7590
rect 4161 7588 4217 7590
rect 3921 6554 3977 6556
rect 4001 6554 4057 6556
rect 4081 6554 4137 6556
rect 4161 6554 4217 6556
rect 3921 6502 3947 6554
rect 3947 6502 3977 6554
rect 4001 6502 4011 6554
rect 4011 6502 4057 6554
rect 4081 6502 4127 6554
rect 4127 6502 4137 6554
rect 4161 6502 4191 6554
rect 4191 6502 4217 6554
rect 3921 6500 3977 6502
rect 4001 6500 4057 6502
rect 4081 6500 4137 6502
rect 4161 6500 4217 6502
rect 4250 5908 4306 5944
rect 4250 5888 4252 5908
rect 4252 5888 4304 5908
rect 4304 5888 4306 5908
rect 4250 5616 4306 5672
rect 3921 5466 3977 5468
rect 4001 5466 4057 5468
rect 4081 5466 4137 5468
rect 4161 5466 4217 5468
rect 3921 5414 3947 5466
rect 3947 5414 3977 5466
rect 4001 5414 4011 5466
rect 4011 5414 4057 5466
rect 4081 5414 4127 5466
rect 4127 5414 4137 5466
rect 4161 5414 4191 5466
rect 4191 5414 4217 5466
rect 3921 5412 3977 5414
rect 4001 5412 4057 5414
rect 4081 5412 4137 5414
rect 4161 5412 4217 5414
rect 3921 4378 3977 4380
rect 4001 4378 4057 4380
rect 4081 4378 4137 4380
rect 4161 4378 4217 4380
rect 3921 4326 3947 4378
rect 3947 4326 3977 4378
rect 4001 4326 4011 4378
rect 4011 4326 4057 4378
rect 4081 4326 4127 4378
rect 4127 4326 4137 4378
rect 4161 4326 4191 4378
rect 4191 4326 4217 4378
rect 3921 4324 3977 4326
rect 4001 4324 4057 4326
rect 4081 4324 4137 4326
rect 4161 4324 4217 4326
rect 1306 584 1362 640
rect 3921 3290 3977 3292
rect 4001 3290 4057 3292
rect 4081 3290 4137 3292
rect 4161 3290 4217 3292
rect 3921 3238 3947 3290
rect 3947 3238 3977 3290
rect 4001 3238 4011 3290
rect 4011 3238 4057 3290
rect 4081 3238 4127 3290
rect 4127 3238 4137 3290
rect 4161 3238 4191 3290
rect 4191 3238 4217 3290
rect 3921 3236 3977 3238
rect 4001 3236 4057 3238
rect 4081 3236 4137 3238
rect 4161 3236 4217 3238
rect 4066 2932 4068 2952
rect 4068 2932 4120 2952
rect 4120 2932 4122 2952
rect 4066 2896 4122 2932
rect 4802 9560 4858 9616
rect 4894 9424 4950 9480
rect 4526 8880 4582 8936
rect 4618 8744 4674 8800
rect 5538 10648 5594 10704
rect 5262 9560 5318 9616
rect 4986 7656 5042 7712
rect 5354 7520 5410 7576
rect 4894 6332 4896 6352
rect 4896 6332 4948 6352
rect 4948 6332 4950 6352
rect 4894 6296 4950 6332
rect 5354 5888 5410 5944
rect 5998 9288 6054 9344
rect 5814 8336 5870 8392
rect 5906 5752 5962 5808
rect 5722 5616 5778 5672
rect 3921 2202 3977 2204
rect 4001 2202 4057 2204
rect 4081 2202 4137 2204
rect 4161 2202 4217 2204
rect 3921 2150 3947 2202
rect 3947 2150 3977 2202
rect 4001 2150 4011 2202
rect 4011 2150 4057 2202
rect 4081 2150 4127 2202
rect 4127 2150 4137 2202
rect 4161 2150 4191 2202
rect 4191 2150 4217 2202
rect 3921 2148 3977 2150
rect 4001 2148 4057 2150
rect 4081 2148 4137 2150
rect 4161 2148 4217 2150
rect 6886 13626 6942 13628
rect 6966 13626 7022 13628
rect 7046 13626 7102 13628
rect 7126 13626 7182 13628
rect 6886 13574 6912 13626
rect 6912 13574 6942 13626
rect 6966 13574 6976 13626
rect 6976 13574 7022 13626
rect 7046 13574 7092 13626
rect 7092 13574 7102 13626
rect 7126 13574 7156 13626
rect 7156 13574 7182 13626
rect 6886 13572 6942 13574
rect 6966 13572 7022 13574
rect 7046 13572 7102 13574
rect 7126 13572 7182 13574
rect 6886 12538 6942 12540
rect 6966 12538 7022 12540
rect 7046 12538 7102 12540
rect 7126 12538 7182 12540
rect 6886 12486 6912 12538
rect 6912 12486 6942 12538
rect 6966 12486 6976 12538
rect 6976 12486 7022 12538
rect 7046 12486 7092 12538
rect 7092 12486 7102 12538
rect 7126 12486 7156 12538
rect 7156 12486 7182 12538
rect 6886 12484 6942 12486
rect 6966 12484 7022 12486
rect 7046 12484 7102 12486
rect 7126 12484 7182 12486
rect 6886 11450 6942 11452
rect 6966 11450 7022 11452
rect 7046 11450 7102 11452
rect 7126 11450 7182 11452
rect 6886 11398 6912 11450
rect 6912 11398 6942 11450
rect 6966 11398 6976 11450
rect 6976 11398 7022 11450
rect 7046 11398 7092 11450
rect 7092 11398 7102 11450
rect 7126 11398 7156 11450
rect 7156 11398 7182 11450
rect 6886 11396 6942 11398
rect 6966 11396 7022 11398
rect 7046 11396 7102 11398
rect 7126 11396 7182 11398
rect 6886 10362 6942 10364
rect 6966 10362 7022 10364
rect 7046 10362 7102 10364
rect 7126 10362 7182 10364
rect 6886 10310 6912 10362
rect 6912 10310 6942 10362
rect 6966 10310 6976 10362
rect 6976 10310 7022 10362
rect 7046 10310 7092 10362
rect 7092 10310 7102 10362
rect 7126 10310 7156 10362
rect 7156 10310 7182 10362
rect 6886 10308 6942 10310
rect 6966 10308 7022 10310
rect 7046 10308 7102 10310
rect 7126 10308 7182 10310
rect 6642 9324 6644 9344
rect 6644 9324 6696 9344
rect 6696 9324 6698 9344
rect 6642 9288 6698 9324
rect 6886 9274 6942 9276
rect 6966 9274 7022 9276
rect 7046 9274 7102 9276
rect 7126 9274 7182 9276
rect 6886 9222 6912 9274
rect 6912 9222 6942 9274
rect 6966 9222 6976 9274
rect 6976 9222 7022 9274
rect 7046 9222 7092 9274
rect 7092 9222 7102 9274
rect 7126 9222 7156 9274
rect 7156 9222 7182 9274
rect 6886 9220 6942 9222
rect 6966 9220 7022 9222
rect 7046 9220 7102 9222
rect 7126 9220 7182 9222
rect 6886 8186 6942 8188
rect 6966 8186 7022 8188
rect 7046 8186 7102 8188
rect 7126 8186 7182 8188
rect 6886 8134 6912 8186
rect 6912 8134 6942 8186
rect 6966 8134 6976 8186
rect 6976 8134 7022 8186
rect 7046 8134 7092 8186
rect 7092 8134 7102 8186
rect 7126 8134 7156 8186
rect 7156 8134 7182 8186
rect 6886 8132 6942 8134
rect 6966 8132 7022 8134
rect 7046 8132 7102 8134
rect 7126 8132 7182 8134
rect 6886 7098 6942 7100
rect 6966 7098 7022 7100
rect 7046 7098 7102 7100
rect 7126 7098 7182 7100
rect 6886 7046 6912 7098
rect 6912 7046 6942 7098
rect 6966 7046 6976 7098
rect 6976 7046 7022 7098
rect 7046 7046 7092 7098
rect 7092 7046 7102 7098
rect 7126 7046 7156 7098
rect 7156 7046 7182 7098
rect 6886 7044 6942 7046
rect 6966 7044 7022 7046
rect 7046 7044 7102 7046
rect 7126 7044 7182 7046
rect 6366 5208 6422 5264
rect 7746 9172 7802 9208
rect 7746 9152 7748 9172
rect 7748 9152 7800 9172
rect 7800 9152 7802 9172
rect 6886 6010 6942 6012
rect 6966 6010 7022 6012
rect 7046 6010 7102 6012
rect 7126 6010 7182 6012
rect 6886 5958 6912 6010
rect 6912 5958 6942 6010
rect 6966 5958 6976 6010
rect 6976 5958 7022 6010
rect 7046 5958 7092 6010
rect 7092 5958 7102 6010
rect 7126 5958 7156 6010
rect 7156 5958 7182 6010
rect 6886 5956 6942 5958
rect 6966 5956 7022 5958
rect 7046 5956 7102 5958
rect 7126 5956 7182 5958
rect 7286 5908 7342 5944
rect 7286 5888 7288 5908
rect 7288 5888 7340 5908
rect 7340 5888 7342 5908
rect 7378 5616 7434 5672
rect 6886 4922 6942 4924
rect 6966 4922 7022 4924
rect 7046 4922 7102 4924
rect 7126 4922 7182 4924
rect 6886 4870 6912 4922
rect 6912 4870 6942 4922
rect 6966 4870 6976 4922
rect 6976 4870 7022 4922
rect 7046 4870 7092 4922
rect 7092 4870 7102 4922
rect 7126 4870 7156 4922
rect 7156 4870 7182 4922
rect 6886 4868 6942 4870
rect 6966 4868 7022 4870
rect 7046 4868 7102 4870
rect 7126 4868 7182 4870
rect 6886 3834 6942 3836
rect 6966 3834 7022 3836
rect 7046 3834 7102 3836
rect 7126 3834 7182 3836
rect 6886 3782 6912 3834
rect 6912 3782 6942 3834
rect 6966 3782 6976 3834
rect 6976 3782 7022 3834
rect 7046 3782 7092 3834
rect 7092 3782 7102 3834
rect 7126 3782 7156 3834
rect 7156 3782 7182 3834
rect 6886 3780 6942 3782
rect 6966 3780 7022 3782
rect 7046 3780 7102 3782
rect 7126 3780 7182 3782
rect 8206 9288 8262 9344
rect 8390 7404 8446 7440
rect 8390 7384 8392 7404
rect 8392 7384 8444 7404
rect 8444 7384 8446 7404
rect 8206 6296 8262 6352
rect 7746 5616 7802 5672
rect 6886 2746 6942 2748
rect 6966 2746 7022 2748
rect 7046 2746 7102 2748
rect 7126 2746 7182 2748
rect 6886 2694 6912 2746
rect 6912 2694 6942 2746
rect 6966 2694 6976 2746
rect 6976 2694 7022 2746
rect 7046 2694 7092 2746
rect 7092 2694 7102 2746
rect 7126 2694 7156 2746
rect 7156 2694 7182 2746
rect 6886 2692 6942 2694
rect 6966 2692 7022 2694
rect 7046 2692 7102 2694
rect 7126 2692 7182 2694
rect 8390 5616 8446 5672
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9878 14170
rect 9878 14118 9908 14170
rect 9932 14118 9942 14170
rect 9942 14118 9988 14170
rect 10012 14118 10058 14170
rect 10058 14118 10068 14170
rect 10092 14118 10122 14170
rect 10122 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9878 13082
rect 9878 13030 9908 13082
rect 9932 13030 9942 13082
rect 9942 13030 9988 13082
rect 10012 13030 10058 13082
rect 10058 13030 10068 13082
rect 10092 13030 10122 13082
rect 10122 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 8666 10104 8722 10160
rect 8666 9016 8722 9072
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9878 11994
rect 9878 11942 9908 11994
rect 9932 11942 9942 11994
rect 9942 11942 9988 11994
rect 10012 11942 10058 11994
rect 10058 11942 10068 11994
rect 10092 11942 10122 11994
rect 10122 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9878 10906
rect 9878 10854 9908 10906
rect 9932 10854 9942 10906
rect 9942 10854 9988 10906
rect 10012 10854 10058 10906
rect 10058 10854 10068 10906
rect 10092 10854 10122 10906
rect 10122 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9878 9818
rect 9878 9766 9908 9818
rect 9932 9766 9942 9818
rect 9942 9766 9988 9818
rect 10012 9766 10058 9818
rect 10058 9766 10068 9818
rect 10092 9766 10122 9818
rect 10122 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 9310 9288 9366 9344
rect 9862 9288 9918 9344
rect 9586 8880 9642 8936
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9878 8730
rect 9878 8678 9908 8730
rect 9932 8678 9942 8730
rect 9942 8678 9988 8730
rect 10012 8678 10058 8730
rect 10058 8678 10068 8730
rect 10092 8678 10122 8730
rect 10122 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 9402 8336 9458 8392
rect 9310 7520 9366 7576
rect 9310 7384 9366 7440
rect 9954 8508 9956 8528
rect 9956 8508 10008 8528
rect 10008 8508 10010 8528
rect 9954 8472 10010 8508
rect 10414 9424 10470 9480
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9878 7642
rect 9878 7590 9908 7642
rect 9932 7590 9942 7642
rect 9942 7590 9988 7642
rect 10012 7590 10058 7642
rect 10058 7590 10068 7642
rect 10092 7590 10122 7642
rect 10122 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9878 6554
rect 9878 6502 9908 6554
rect 9932 6502 9942 6554
rect 9942 6502 9988 6554
rect 10012 6502 10058 6554
rect 10058 6502 10068 6554
rect 10092 6502 10122 6554
rect 10122 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9878 5466
rect 9878 5414 9908 5466
rect 9932 5414 9942 5466
rect 9942 5414 9988 5466
rect 10012 5414 10058 5466
rect 10058 5414 10068 5466
rect 10092 5414 10122 5466
rect 10122 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9878 4378
rect 9878 4326 9908 4378
rect 9932 4326 9942 4378
rect 9942 4326 9988 4378
rect 10012 4326 10058 4378
rect 10058 4326 10068 4378
rect 10092 4326 10122 4378
rect 10122 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9878 3290
rect 9878 3238 9908 3290
rect 9932 3238 9942 3290
rect 9942 3238 9988 3290
rect 10012 3238 10058 3290
rect 10058 3238 10068 3290
rect 10092 3238 10122 3290
rect 10122 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 10230 2760 10286 2816
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9878 2202
rect 9878 2150 9908 2202
rect 9932 2150 9942 2202
rect 9942 2150 9988 2202
rect 10012 2150 10058 2202
rect 10058 2150 10068 2202
rect 10092 2150 10122 2202
rect 10122 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 11058 9968 11114 10024
rect 11058 9324 11060 9344
rect 11060 9324 11112 9344
rect 11112 9324 11114 9344
rect 11058 9288 11114 9324
rect 10966 8472 11022 8528
rect 10782 6704 10838 6760
rect 10598 3440 10654 3496
rect 10598 3304 10654 3360
rect 10874 3168 10930 3224
rect 10874 2760 10930 2816
rect 11334 6840 11390 6896
rect 11978 7964 11980 7984
rect 11980 7964 12032 7984
rect 12032 7964 12034 7984
rect 11978 7928 12034 7964
rect 12817 14714 12873 14716
rect 12897 14714 12953 14716
rect 12977 14714 13033 14716
rect 13057 14714 13113 14716
rect 12817 14662 12843 14714
rect 12843 14662 12873 14714
rect 12897 14662 12907 14714
rect 12907 14662 12953 14714
rect 12977 14662 13023 14714
rect 13023 14662 13033 14714
rect 13057 14662 13087 14714
rect 13087 14662 13113 14714
rect 12817 14660 12873 14662
rect 12897 14660 12953 14662
rect 12977 14660 13033 14662
rect 13057 14660 13113 14662
rect 12817 13626 12873 13628
rect 12897 13626 12953 13628
rect 12977 13626 13033 13628
rect 13057 13626 13113 13628
rect 12817 13574 12843 13626
rect 12843 13574 12873 13626
rect 12897 13574 12907 13626
rect 12907 13574 12953 13626
rect 12977 13574 13023 13626
rect 13023 13574 13033 13626
rect 13057 13574 13087 13626
rect 13087 13574 13113 13626
rect 12817 13572 12873 13574
rect 12897 13572 12953 13574
rect 12977 13572 13033 13574
rect 13057 13572 13113 13574
rect 12817 12538 12873 12540
rect 12897 12538 12953 12540
rect 12977 12538 13033 12540
rect 13057 12538 13113 12540
rect 12817 12486 12843 12538
rect 12843 12486 12873 12538
rect 12897 12486 12907 12538
rect 12907 12486 12953 12538
rect 12977 12486 13023 12538
rect 13023 12486 13033 12538
rect 13057 12486 13087 12538
rect 13087 12486 13113 12538
rect 12817 12484 12873 12486
rect 12897 12484 12953 12486
rect 12977 12484 13033 12486
rect 13057 12484 13113 12486
rect 12817 11450 12873 11452
rect 12897 11450 12953 11452
rect 12977 11450 13033 11452
rect 13057 11450 13113 11452
rect 12817 11398 12843 11450
rect 12843 11398 12873 11450
rect 12897 11398 12907 11450
rect 12907 11398 12953 11450
rect 12977 11398 13023 11450
rect 13023 11398 13033 11450
rect 13057 11398 13087 11450
rect 13087 11398 13113 11450
rect 12817 11396 12873 11398
rect 12897 11396 12953 11398
rect 12977 11396 13033 11398
rect 13057 11396 13113 11398
rect 12817 10362 12873 10364
rect 12897 10362 12953 10364
rect 12977 10362 13033 10364
rect 13057 10362 13113 10364
rect 12817 10310 12843 10362
rect 12843 10310 12873 10362
rect 12897 10310 12907 10362
rect 12907 10310 12953 10362
rect 12977 10310 13023 10362
rect 13023 10310 13033 10362
rect 13057 10310 13087 10362
rect 13087 10310 13113 10362
rect 12817 10308 12873 10310
rect 12897 10308 12953 10310
rect 12977 10308 13033 10310
rect 13057 10308 13113 10310
rect 12817 9274 12873 9276
rect 12897 9274 12953 9276
rect 12977 9274 13033 9276
rect 13057 9274 13113 9276
rect 12817 9222 12843 9274
rect 12843 9222 12873 9274
rect 12897 9222 12907 9274
rect 12907 9222 12953 9274
rect 12977 9222 13023 9274
rect 13023 9222 13033 9274
rect 13057 9222 13087 9274
rect 13087 9222 13113 9274
rect 12817 9220 12873 9222
rect 12897 9220 12953 9222
rect 12977 9220 13033 9222
rect 13057 9220 13113 9222
rect 12346 7540 12402 7576
rect 12346 7520 12348 7540
rect 12348 7520 12400 7540
rect 12400 7520 12402 7540
rect 12070 5752 12126 5808
rect 12346 7248 12402 7304
rect 12817 8186 12873 8188
rect 12897 8186 12953 8188
rect 12977 8186 13033 8188
rect 13057 8186 13113 8188
rect 12817 8134 12843 8186
rect 12843 8134 12873 8186
rect 12897 8134 12907 8186
rect 12907 8134 12953 8186
rect 12977 8134 13023 8186
rect 13023 8134 13033 8186
rect 13057 8134 13087 8186
rect 13087 8134 13113 8186
rect 12817 8132 12873 8134
rect 12897 8132 12953 8134
rect 12977 8132 13033 8134
rect 13057 8132 13113 8134
rect 12806 7812 12862 7848
rect 12806 7792 12808 7812
rect 12808 7792 12860 7812
rect 12860 7792 12862 7812
rect 12817 7098 12873 7100
rect 12897 7098 12953 7100
rect 12977 7098 13033 7100
rect 13057 7098 13113 7100
rect 12817 7046 12843 7098
rect 12843 7046 12873 7098
rect 12897 7046 12907 7098
rect 12907 7046 12953 7098
rect 12977 7046 13023 7098
rect 13023 7046 13033 7098
rect 13057 7046 13087 7098
rect 13087 7046 13113 7098
rect 12817 7044 12873 7046
rect 12897 7044 12953 7046
rect 12977 7044 13033 7046
rect 13057 7044 13113 7046
rect 13910 9424 13966 9480
rect 13818 7520 13874 7576
rect 13726 7384 13782 7440
rect 13174 6432 13230 6488
rect 12817 6010 12873 6012
rect 12897 6010 12953 6012
rect 12977 6010 13033 6012
rect 13057 6010 13113 6012
rect 12817 5958 12843 6010
rect 12843 5958 12873 6010
rect 12897 5958 12907 6010
rect 12907 5958 12953 6010
rect 12977 5958 13023 6010
rect 13023 5958 13033 6010
rect 13057 5958 13087 6010
rect 13087 5958 13113 6010
rect 12817 5956 12873 5958
rect 12897 5956 12953 5958
rect 12977 5956 13033 5958
rect 13057 5956 13113 5958
rect 13358 6840 13414 6896
rect 12817 4922 12873 4924
rect 12897 4922 12953 4924
rect 12977 4922 13033 4924
rect 13057 4922 13113 4924
rect 12817 4870 12843 4922
rect 12843 4870 12873 4922
rect 12897 4870 12907 4922
rect 12907 4870 12953 4922
rect 12977 4870 13023 4922
rect 13023 4870 13033 4922
rect 13057 4870 13087 4922
rect 13087 4870 13113 4922
rect 12817 4868 12873 4870
rect 12897 4868 12953 4870
rect 12977 4868 13033 4870
rect 13057 4868 13113 4870
rect 13450 4664 13506 4720
rect 13726 6976 13782 7032
rect 13726 6840 13782 6896
rect 13726 6160 13782 6216
rect 14002 7928 14058 7984
rect 13818 5108 13820 5128
rect 13820 5108 13872 5128
rect 13872 5108 13874 5128
rect 13818 5072 13874 5108
rect 12817 3834 12873 3836
rect 12897 3834 12953 3836
rect 12977 3834 13033 3836
rect 13057 3834 13113 3836
rect 12817 3782 12843 3834
rect 12843 3782 12873 3834
rect 12897 3782 12907 3834
rect 12907 3782 12953 3834
rect 12977 3782 13023 3834
rect 13023 3782 13033 3834
rect 13057 3782 13087 3834
rect 13087 3782 13113 3834
rect 12817 3780 12873 3782
rect 12897 3780 12953 3782
rect 12977 3780 13033 3782
rect 13057 3780 13113 3782
rect 12806 3440 12862 3496
rect 12990 3032 13046 3088
rect 12817 2746 12873 2748
rect 12897 2746 12953 2748
rect 12977 2746 13033 2748
rect 13057 2746 13113 2748
rect 12817 2694 12843 2746
rect 12843 2694 12873 2746
rect 12897 2694 12907 2746
rect 12907 2694 12953 2746
rect 12977 2694 13023 2746
rect 13023 2694 13033 2746
rect 13057 2694 13087 2746
rect 13087 2694 13113 2746
rect 12817 2692 12873 2694
rect 12897 2692 12953 2694
rect 12977 2692 13033 2694
rect 13057 2692 13113 2694
rect 13450 3032 13506 3088
rect 14278 7384 14334 7440
rect 14278 6432 14334 6488
rect 14462 3304 14518 3360
rect 14278 3168 14334 3224
rect 14462 3032 14518 3088
rect 14738 8880 14794 8936
rect 14646 6160 14702 6216
rect 14646 5616 14702 5672
rect 14646 5208 14702 5264
rect 14738 5072 14794 5128
rect 15198 6024 15254 6080
rect 15382 4528 15438 4584
rect 14922 2896 14978 2952
rect 15782 14170 15838 14172
rect 15862 14170 15918 14172
rect 15942 14170 15998 14172
rect 16022 14170 16078 14172
rect 15782 14118 15808 14170
rect 15808 14118 15838 14170
rect 15862 14118 15872 14170
rect 15872 14118 15918 14170
rect 15942 14118 15988 14170
rect 15988 14118 15998 14170
rect 16022 14118 16052 14170
rect 16052 14118 16078 14170
rect 15782 14116 15838 14118
rect 15862 14116 15918 14118
rect 15942 14116 15998 14118
rect 16022 14116 16078 14118
rect 15782 13082 15838 13084
rect 15862 13082 15918 13084
rect 15942 13082 15998 13084
rect 16022 13082 16078 13084
rect 15782 13030 15808 13082
rect 15808 13030 15838 13082
rect 15862 13030 15872 13082
rect 15872 13030 15918 13082
rect 15942 13030 15988 13082
rect 15988 13030 15998 13082
rect 16022 13030 16052 13082
rect 16052 13030 16078 13082
rect 15782 13028 15838 13030
rect 15862 13028 15918 13030
rect 15942 13028 15998 13030
rect 16022 13028 16078 13030
rect 15782 11994 15838 11996
rect 15862 11994 15918 11996
rect 15942 11994 15998 11996
rect 16022 11994 16078 11996
rect 15782 11942 15808 11994
rect 15808 11942 15838 11994
rect 15862 11942 15872 11994
rect 15872 11942 15918 11994
rect 15942 11942 15988 11994
rect 15988 11942 15998 11994
rect 16022 11942 16052 11994
rect 16052 11942 16078 11994
rect 15782 11940 15838 11942
rect 15862 11940 15918 11942
rect 15942 11940 15998 11942
rect 16022 11940 16078 11942
rect 16578 15952 16634 16008
rect 16946 15544 17002 15600
rect 15782 10906 15838 10908
rect 15862 10906 15918 10908
rect 15942 10906 15998 10908
rect 16022 10906 16078 10908
rect 15782 10854 15808 10906
rect 15808 10854 15838 10906
rect 15862 10854 15872 10906
rect 15872 10854 15918 10906
rect 15942 10854 15988 10906
rect 15988 10854 15998 10906
rect 16022 10854 16052 10906
rect 16052 10854 16078 10906
rect 15782 10852 15838 10854
rect 15862 10852 15918 10854
rect 15942 10852 15998 10854
rect 16022 10852 16078 10854
rect 15782 9818 15838 9820
rect 15862 9818 15918 9820
rect 15942 9818 15998 9820
rect 16022 9818 16078 9820
rect 15782 9766 15808 9818
rect 15808 9766 15838 9818
rect 15862 9766 15872 9818
rect 15872 9766 15918 9818
rect 15942 9766 15988 9818
rect 15988 9766 15998 9818
rect 16022 9766 16052 9818
rect 16052 9766 16078 9818
rect 15782 9764 15838 9766
rect 15862 9764 15918 9766
rect 15942 9764 15998 9766
rect 16022 9764 16078 9766
rect 15658 9596 15660 9616
rect 15660 9596 15712 9616
rect 15712 9596 15714 9616
rect 15658 9560 15714 9596
rect 16026 9016 16082 9072
rect 15782 8730 15838 8732
rect 15862 8730 15918 8732
rect 15942 8730 15998 8732
rect 16022 8730 16078 8732
rect 15782 8678 15808 8730
rect 15808 8678 15838 8730
rect 15862 8678 15872 8730
rect 15872 8678 15918 8730
rect 15942 8678 15988 8730
rect 15988 8678 15998 8730
rect 16022 8678 16052 8730
rect 16052 8678 16078 8730
rect 15782 8676 15838 8678
rect 15862 8676 15918 8678
rect 15942 8676 15998 8678
rect 16022 8676 16078 8678
rect 15658 8064 15714 8120
rect 15782 7642 15838 7644
rect 15862 7642 15918 7644
rect 15942 7642 15998 7644
rect 16022 7642 16078 7644
rect 15782 7590 15808 7642
rect 15808 7590 15838 7642
rect 15862 7590 15872 7642
rect 15872 7590 15918 7642
rect 15942 7590 15988 7642
rect 15988 7590 15998 7642
rect 16022 7590 16052 7642
rect 16052 7590 16078 7642
rect 15782 7588 15838 7590
rect 15862 7588 15918 7590
rect 15942 7588 15998 7590
rect 16022 7588 16078 7590
rect 17498 16360 17554 16416
rect 17774 15136 17830 15192
rect 17866 14728 17922 14784
rect 18050 12552 18106 12608
rect 18418 14184 18474 14240
rect 18418 13812 18420 13832
rect 18420 13812 18472 13832
rect 18472 13812 18474 13832
rect 18418 13776 18474 13812
rect 18418 13388 18474 13424
rect 18418 13368 18420 13388
rect 18420 13368 18472 13388
rect 18472 13368 18474 13388
rect 18418 12960 18474 13016
rect 16854 9560 16910 9616
rect 16302 8084 16358 8120
rect 16302 8064 16304 8084
rect 16304 8064 16356 8084
rect 16356 8064 16358 8084
rect 15750 6860 15806 6896
rect 15750 6840 15752 6860
rect 15752 6840 15804 6860
rect 15804 6840 15806 6860
rect 15842 6704 15898 6760
rect 15782 6554 15838 6556
rect 15862 6554 15918 6556
rect 15942 6554 15998 6556
rect 16022 6554 16078 6556
rect 15782 6502 15808 6554
rect 15808 6502 15838 6554
rect 15862 6502 15872 6554
rect 15872 6502 15918 6554
rect 15942 6502 15988 6554
rect 15988 6502 15998 6554
rect 16022 6502 16052 6554
rect 16052 6502 16078 6554
rect 15782 6500 15838 6502
rect 15862 6500 15918 6502
rect 15942 6500 15998 6502
rect 16022 6500 16078 6502
rect 15782 5466 15838 5468
rect 15862 5466 15918 5468
rect 15942 5466 15998 5468
rect 16022 5466 16078 5468
rect 15782 5414 15808 5466
rect 15808 5414 15838 5466
rect 15862 5414 15872 5466
rect 15872 5414 15918 5466
rect 15942 5414 15988 5466
rect 15988 5414 15998 5466
rect 16022 5414 16052 5466
rect 16052 5414 16078 5466
rect 15782 5412 15838 5414
rect 15862 5412 15918 5414
rect 15942 5412 15998 5414
rect 16022 5412 16078 5414
rect 15750 4548 15806 4584
rect 15750 4528 15752 4548
rect 15752 4528 15804 4548
rect 15804 4528 15806 4548
rect 15782 4378 15838 4380
rect 15862 4378 15918 4380
rect 15942 4378 15998 4380
rect 16022 4378 16078 4380
rect 15782 4326 15808 4378
rect 15808 4326 15838 4378
rect 15862 4326 15872 4378
rect 15872 4326 15918 4378
rect 15942 4326 15988 4378
rect 15988 4326 15998 4378
rect 16022 4326 16052 4378
rect 16052 4326 16078 4378
rect 15782 4324 15838 4326
rect 15862 4324 15918 4326
rect 15942 4324 15998 4326
rect 16022 4324 16078 4326
rect 15782 3290 15838 3292
rect 15862 3290 15918 3292
rect 15942 3290 15998 3292
rect 16022 3290 16078 3292
rect 15782 3238 15808 3290
rect 15808 3238 15838 3290
rect 15862 3238 15872 3290
rect 15872 3238 15918 3290
rect 15942 3238 15988 3290
rect 15988 3238 15998 3290
rect 16022 3238 16052 3290
rect 16052 3238 16078 3290
rect 15782 3236 15838 3238
rect 15862 3236 15918 3238
rect 15942 3236 15998 3238
rect 16022 3236 16078 3238
rect 15750 3052 15806 3088
rect 15750 3032 15752 3052
rect 15752 3032 15804 3052
rect 15804 3032 15806 3052
rect 16670 7284 16672 7304
rect 16672 7284 16724 7304
rect 16724 7284 16726 7304
rect 16670 7248 16726 7284
rect 16394 5752 16450 5808
rect 16670 6316 16726 6352
rect 16670 6296 16672 6316
rect 16672 6296 16724 6316
rect 16724 6296 16726 6316
rect 17314 9560 17370 9616
rect 18050 12144 18106 12200
rect 18418 11736 18474 11792
rect 18142 10376 18198 10432
rect 17866 9968 17922 10024
rect 18050 9596 18052 9616
rect 18052 9596 18104 9616
rect 18104 9596 18106 9616
rect 18050 9560 18106 9596
rect 18418 11192 18474 11248
rect 18510 10784 18566 10840
rect 18418 9968 18474 10024
rect 17866 9444 17922 9480
rect 17866 9424 17868 9444
rect 17868 9424 17920 9444
rect 17920 9424 17922 9444
rect 18234 8916 18236 8936
rect 18236 8916 18288 8936
rect 18288 8916 18290 8936
rect 18234 8880 18290 8916
rect 17498 7384 17554 7440
rect 18418 9152 18474 9208
rect 18418 8744 18474 8800
rect 18510 8200 18566 8256
rect 18510 7812 18566 7848
rect 18510 7792 18512 7812
rect 18512 7792 18564 7812
rect 18564 7792 18566 7812
rect 18142 7404 18198 7440
rect 18142 7384 18144 7404
rect 18144 7384 18196 7404
rect 18196 7384 18198 7404
rect 17130 6740 17132 6760
rect 17132 6740 17184 6760
rect 17184 6740 17186 6760
rect 17130 6704 17186 6740
rect 17682 6976 17738 7032
rect 16762 5616 16818 5672
rect 16854 5092 16910 5128
rect 16854 5072 16856 5092
rect 16856 5072 16908 5092
rect 16908 5072 16910 5092
rect 17038 4664 17094 4720
rect 15782 2202 15838 2204
rect 15862 2202 15918 2204
rect 15942 2202 15998 2204
rect 16022 2202 16078 2204
rect 15782 2150 15808 2202
rect 15808 2150 15838 2202
rect 15862 2150 15872 2202
rect 15872 2150 15918 2202
rect 15942 2150 15988 2202
rect 15988 2150 15998 2202
rect 16022 2150 16052 2202
rect 16052 2150 16078 2202
rect 15782 2148 15838 2150
rect 15862 2148 15918 2150
rect 15942 2148 15998 2150
rect 16022 2148 16078 2150
rect 17406 1808 17462 1864
rect 17498 1400 17554 1456
rect 17866 5208 17922 5264
rect 18142 4800 18198 4856
rect 17774 2624 17830 2680
rect 18142 4004 18198 4040
rect 18142 3984 18144 4004
rect 18144 3984 18196 4004
rect 18196 3984 18198 4004
rect 18142 3168 18198 3224
rect 17866 2488 17922 2544
rect 18510 6976 18566 7032
rect 18510 6568 18566 6624
rect 18510 6180 18566 6216
rect 18510 6160 18512 6180
rect 18512 6160 18564 6180
rect 18564 6160 18566 6180
rect 18510 5636 18566 5672
rect 18510 5616 18512 5636
rect 18512 5616 18564 5636
rect 18564 5616 18566 5636
rect 18510 5228 18566 5264
rect 18510 5208 18512 5228
rect 18512 5208 18564 5228
rect 18564 5208 18566 5228
rect 18510 4392 18566 4448
rect 18510 3576 18566 3632
rect 3330 176 3386 232
rect 17774 992 17830 1048
rect 17682 584 17738 640
rect 17866 176 17922 232
<< metal3 >>
rect 0 16826 800 16856
rect 3785 16826 3851 16829
rect 0 16824 3851 16826
rect 0 16768 3790 16824
rect 3846 16768 3851 16824
rect 0 16766 3851 16768
rect 0 16736 800 16766
rect 3785 16763 3851 16766
rect 17401 16826 17467 16829
rect 19200 16826 20000 16856
rect 17401 16824 20000 16826
rect 17401 16768 17406 16824
rect 17462 16768 20000 16824
rect 17401 16766 20000 16768
rect 17401 16763 17467 16766
rect 19200 16736 20000 16766
rect 0 16418 800 16448
rect 3141 16418 3207 16421
rect 0 16416 3207 16418
rect 0 16360 3146 16416
rect 3202 16360 3207 16416
rect 0 16358 3207 16360
rect 0 16328 800 16358
rect 3141 16355 3207 16358
rect 17493 16418 17559 16421
rect 19200 16418 20000 16448
rect 17493 16416 20000 16418
rect 17493 16360 17498 16416
rect 17554 16360 20000 16416
rect 17493 16358 20000 16360
rect 17493 16355 17559 16358
rect 19200 16328 20000 16358
rect 0 16010 800 16040
rect 2589 16010 2655 16013
rect 0 16008 2655 16010
rect 0 15952 2594 16008
rect 2650 15952 2655 16008
rect 0 15950 2655 15952
rect 0 15920 800 15950
rect 2589 15947 2655 15950
rect 16573 16010 16639 16013
rect 19200 16010 20000 16040
rect 16573 16008 20000 16010
rect 16573 15952 16578 16008
rect 16634 15952 20000 16008
rect 16573 15950 20000 15952
rect 16573 15947 16639 15950
rect 19200 15920 20000 15950
rect 0 15602 800 15632
rect 2773 15602 2839 15605
rect 0 15600 2839 15602
rect 0 15544 2778 15600
rect 2834 15544 2839 15600
rect 0 15542 2839 15544
rect 0 15512 800 15542
rect 2773 15539 2839 15542
rect 16941 15602 17007 15605
rect 19200 15602 20000 15632
rect 16941 15600 20000 15602
rect 16941 15544 16946 15600
rect 17002 15544 20000 15600
rect 16941 15542 20000 15544
rect 16941 15539 17007 15542
rect 19200 15512 20000 15542
rect 0 15194 800 15224
rect 2957 15194 3023 15197
rect 0 15192 3023 15194
rect 0 15136 2962 15192
rect 3018 15136 3023 15192
rect 0 15134 3023 15136
rect 0 15104 800 15134
rect 2957 15131 3023 15134
rect 17769 15194 17835 15197
rect 19200 15194 20000 15224
rect 17769 15192 20000 15194
rect 17769 15136 17774 15192
rect 17830 15136 20000 15192
rect 17769 15134 20000 15136
rect 17769 15131 17835 15134
rect 19200 15104 20000 15134
rect 0 14786 800 14816
rect 1853 14786 1919 14789
rect 3325 14786 3391 14789
rect 0 14784 3391 14786
rect 0 14728 1858 14784
rect 1914 14728 3330 14784
rect 3386 14728 3391 14784
rect 0 14726 3391 14728
rect 0 14696 800 14726
rect 1853 14723 1919 14726
rect 3325 14723 3391 14726
rect 17861 14786 17927 14789
rect 19200 14786 20000 14816
rect 17861 14784 20000 14786
rect 17861 14728 17866 14784
rect 17922 14728 20000 14784
rect 17861 14726 20000 14728
rect 17861 14723 17927 14726
rect 6874 14720 7194 14721
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7194 14720
rect 6874 14655 7194 14656
rect 12805 14720 13125 14721
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 19200 14696 20000 14726
rect 12805 14655 13125 14656
rect 1485 14514 1551 14517
rect 3601 14514 3667 14517
rect 1485 14512 3667 14514
rect 1485 14456 1490 14512
rect 1546 14456 3606 14512
rect 3662 14456 3667 14512
rect 1485 14454 3667 14456
rect 1485 14451 1551 14454
rect 3601 14451 3667 14454
rect 0 14378 800 14408
rect 1488 14378 1548 14451
rect 0 14318 1548 14378
rect 0 14288 800 14318
rect 18413 14242 18479 14245
rect 19200 14242 20000 14272
rect 18413 14240 20000 14242
rect 18413 14184 18418 14240
rect 18474 14184 20000 14240
rect 18413 14182 20000 14184
rect 18413 14179 18479 14182
rect 3909 14176 4229 14177
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 14111 4229 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 15770 14176 16090 14177
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 19200 14152 20000 14182
rect 15770 14111 16090 14112
rect 0 13970 800 14000
rect 2589 13970 2655 13973
rect 0 13968 2655 13970
rect 0 13912 2594 13968
rect 2650 13912 2655 13968
rect 0 13910 2655 13912
rect 0 13880 800 13910
rect 2589 13907 2655 13910
rect 3233 13834 3299 13837
rect 4613 13834 4679 13837
rect 3233 13832 4679 13834
rect 3233 13776 3238 13832
rect 3294 13776 4618 13832
rect 4674 13776 4679 13832
rect 3233 13774 4679 13776
rect 3233 13771 3299 13774
rect 4613 13771 4679 13774
rect 18413 13834 18479 13837
rect 19200 13834 20000 13864
rect 18413 13832 20000 13834
rect 18413 13776 18418 13832
rect 18474 13776 20000 13832
rect 18413 13774 20000 13776
rect 18413 13771 18479 13774
rect 19200 13744 20000 13774
rect 2865 13698 2931 13701
rect 4705 13698 4771 13701
rect 2865 13696 4771 13698
rect 2865 13640 2870 13696
rect 2926 13640 4710 13696
rect 4766 13640 4771 13696
rect 2865 13638 4771 13640
rect 2865 13635 2931 13638
rect 4705 13635 4771 13638
rect 6874 13632 7194 13633
rect 0 13562 800 13592
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7194 13632
rect 6874 13567 7194 13568
rect 12805 13632 13125 13633
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 13567 13125 13568
rect 1853 13562 1919 13565
rect 0 13560 1919 13562
rect 0 13504 1858 13560
rect 1914 13504 1919 13560
rect 0 13502 1919 13504
rect 0 13472 800 13502
rect 1853 13499 1919 13502
rect 18413 13426 18479 13429
rect 19200 13426 20000 13456
rect 18413 13424 20000 13426
rect 18413 13368 18418 13424
rect 18474 13368 20000 13424
rect 18413 13366 20000 13368
rect 18413 13363 18479 13366
rect 19200 13336 20000 13366
rect 2129 13290 2195 13293
rect 3877 13290 3943 13293
rect 2129 13288 3943 13290
rect 2129 13232 2134 13288
rect 2190 13232 3882 13288
rect 3938 13232 3943 13288
rect 2129 13230 3943 13232
rect 2129 13227 2195 13230
rect 3877 13227 3943 13230
rect 0 13154 800 13184
rect 1485 13154 1551 13157
rect 0 13152 1551 13154
rect 0 13096 1490 13152
rect 1546 13096 1551 13152
rect 0 13094 1551 13096
rect 0 13064 800 13094
rect 1485 13091 1551 13094
rect 3909 13088 4229 13089
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 13023 4229 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 15770 13088 16090 13089
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 13023 16090 13024
rect 18413 13018 18479 13021
rect 19200 13018 20000 13048
rect 18413 13016 20000 13018
rect 18413 12960 18418 13016
rect 18474 12960 20000 13016
rect 18413 12958 20000 12960
rect 18413 12955 18479 12958
rect 19200 12928 20000 12958
rect 0 12746 800 12776
rect 1577 12746 1643 12749
rect 0 12744 1643 12746
rect 0 12688 1582 12744
rect 1638 12688 1643 12744
rect 0 12686 1643 12688
rect 0 12656 800 12686
rect 1577 12683 1643 12686
rect 1945 12746 2011 12749
rect 4705 12746 4771 12749
rect 1945 12744 4771 12746
rect 1945 12688 1950 12744
rect 2006 12688 4710 12744
rect 4766 12688 4771 12744
rect 1945 12686 4771 12688
rect 1945 12683 2011 12686
rect 4705 12683 4771 12686
rect 18045 12610 18111 12613
rect 19200 12610 20000 12640
rect 18045 12608 20000 12610
rect 18045 12552 18050 12608
rect 18106 12552 20000 12608
rect 18045 12550 20000 12552
rect 18045 12547 18111 12550
rect 6874 12544 7194 12545
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7194 12544
rect 6874 12479 7194 12480
rect 12805 12544 13125 12545
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 19200 12520 20000 12550
rect 12805 12479 13125 12480
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 18045 12202 18111 12205
rect 19200 12202 20000 12232
rect 18045 12200 20000 12202
rect 18045 12144 18050 12200
rect 18106 12144 20000 12200
rect 18045 12142 20000 12144
rect 18045 12139 18111 12142
rect 19200 12112 20000 12142
rect 3909 12000 4229 12001
rect 0 11930 800 11960
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 11935 4229 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 15770 12000 16090 12001
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 11935 16090 11936
rect 1853 11930 1919 11933
rect 3233 11930 3299 11933
rect 0 11928 3299 11930
rect 0 11872 1858 11928
rect 1914 11872 3238 11928
rect 3294 11872 3299 11928
rect 0 11870 3299 11872
rect 0 11840 800 11870
rect 1853 11867 1919 11870
rect 3233 11867 3299 11870
rect 1485 11794 1551 11797
rect 3325 11794 3391 11797
rect 1485 11792 3391 11794
rect 1485 11736 1490 11792
rect 1546 11736 3330 11792
rect 3386 11736 3391 11792
rect 1485 11734 3391 11736
rect 1485 11731 1551 11734
rect 3325 11731 3391 11734
rect 18413 11794 18479 11797
rect 19200 11794 20000 11824
rect 18413 11792 20000 11794
rect 18413 11736 18418 11792
rect 18474 11736 20000 11792
rect 18413 11734 20000 11736
rect 18413 11731 18479 11734
rect 19200 11704 20000 11734
rect 6874 11456 7194 11457
rect 0 11386 800 11416
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7194 11456
rect 6874 11391 7194 11392
rect 12805 11456 13125 11457
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 11391 13125 11392
rect 1393 11386 1459 11389
rect 0 11384 1459 11386
rect 0 11328 1398 11384
rect 1454 11328 1459 11384
rect 0 11326 1459 11328
rect 0 11296 800 11326
rect 1393 11323 1459 11326
rect 18413 11250 18479 11253
rect 19200 11250 20000 11280
rect 18413 11248 20000 11250
rect 18413 11192 18418 11248
rect 18474 11192 20000 11248
rect 18413 11190 20000 11192
rect 18413 11187 18479 11190
rect 19200 11160 20000 11190
rect 0 10978 800 11008
rect 1485 10978 1551 10981
rect 0 10976 1551 10978
rect 0 10920 1490 10976
rect 1546 10920 1551 10976
rect 0 10918 1551 10920
rect 0 10888 800 10918
rect 1485 10915 1551 10918
rect 1669 10978 1735 10981
rect 2497 10978 2563 10981
rect 1669 10976 2563 10978
rect 1669 10920 1674 10976
rect 1730 10920 2502 10976
rect 2558 10920 2563 10976
rect 1669 10918 2563 10920
rect 1669 10915 1735 10918
rect 2497 10915 2563 10918
rect 3909 10912 4229 10913
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 10847 4229 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 15770 10912 16090 10913
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 10847 16090 10848
rect 18505 10842 18571 10845
rect 19200 10842 20000 10872
rect 18505 10840 20000 10842
rect 18505 10784 18510 10840
rect 18566 10784 20000 10840
rect 18505 10782 20000 10784
rect 18505 10779 18571 10782
rect 19200 10752 20000 10782
rect 1577 10706 1643 10709
rect 5533 10706 5599 10709
rect 1577 10704 5599 10706
rect 1577 10648 1582 10704
rect 1638 10648 5538 10704
rect 5594 10648 5599 10704
rect 1577 10646 5599 10648
rect 1577 10643 1643 10646
rect 5533 10643 5599 10646
rect 0 10570 800 10600
rect 1393 10570 1459 10573
rect 3509 10570 3575 10573
rect 0 10568 3575 10570
rect 0 10512 1398 10568
rect 1454 10512 3514 10568
rect 3570 10512 3575 10568
rect 0 10510 3575 10512
rect 0 10480 800 10510
rect 1393 10507 1459 10510
rect 3509 10507 3575 10510
rect 18137 10434 18203 10437
rect 19200 10434 20000 10464
rect 18137 10432 20000 10434
rect 18137 10376 18142 10432
rect 18198 10376 20000 10432
rect 18137 10374 20000 10376
rect 18137 10371 18203 10374
rect 6874 10368 7194 10369
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7194 10368
rect 6874 10303 7194 10304
rect 12805 10368 13125 10369
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 19200 10344 20000 10374
rect 12805 10303 13125 10304
rect 0 10162 800 10192
rect 1485 10162 1551 10165
rect 0 10160 1551 10162
rect 0 10104 1490 10160
rect 1546 10104 1551 10160
rect 0 10102 1551 10104
rect 0 10072 800 10102
rect 1485 10099 1551 10102
rect 3049 10162 3115 10165
rect 8661 10162 8727 10165
rect 3049 10160 8727 10162
rect 3049 10104 3054 10160
rect 3110 10104 8666 10160
rect 8722 10104 8727 10160
rect 3049 10102 8727 10104
rect 3049 10099 3115 10102
rect 8661 10099 8727 10102
rect 11053 10026 11119 10029
rect 17861 10026 17927 10029
rect 11053 10024 17927 10026
rect 11053 9968 11058 10024
rect 11114 9968 17866 10024
rect 17922 9968 17927 10024
rect 11053 9966 17927 9968
rect 11053 9963 11119 9966
rect 17861 9963 17927 9966
rect 18413 10026 18479 10029
rect 19200 10026 20000 10056
rect 18413 10024 20000 10026
rect 18413 9968 18418 10024
rect 18474 9968 20000 10024
rect 18413 9966 20000 9968
rect 18413 9963 18479 9966
rect 19200 9936 20000 9966
rect 3909 9824 4229 9825
rect 0 9754 800 9784
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 9759 4229 9760
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 15770 9824 16090 9825
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 15770 9759 16090 9760
rect 3233 9754 3299 9757
rect 0 9752 3299 9754
rect 0 9696 3238 9752
rect 3294 9696 3299 9752
rect 0 9694 3299 9696
rect 0 9664 800 9694
rect 3233 9691 3299 9694
rect 2129 9618 2195 9621
rect 3233 9618 3299 9621
rect 2129 9616 3299 9618
rect 2129 9560 2134 9616
rect 2190 9560 3238 9616
rect 3294 9560 3299 9616
rect 2129 9558 3299 9560
rect 2129 9555 2195 9558
rect 3233 9555 3299 9558
rect 4797 9618 4863 9621
rect 5257 9618 5323 9621
rect 15653 9618 15719 9621
rect 16849 9618 16915 9621
rect 17309 9618 17375 9621
rect 4797 9616 17375 9618
rect 4797 9560 4802 9616
rect 4858 9560 5262 9616
rect 5318 9560 15658 9616
rect 15714 9560 16854 9616
rect 16910 9560 17314 9616
rect 17370 9560 17375 9616
rect 4797 9558 17375 9560
rect 4797 9555 4863 9558
rect 5257 9555 5323 9558
rect 15653 9555 15719 9558
rect 16849 9555 16915 9558
rect 17309 9555 17375 9558
rect 18045 9618 18111 9621
rect 19200 9618 20000 9648
rect 18045 9616 20000 9618
rect 18045 9560 18050 9616
rect 18106 9560 20000 9616
rect 18045 9558 20000 9560
rect 18045 9555 18111 9558
rect 19200 9528 20000 9558
rect 4061 9482 4127 9485
rect 4889 9482 4955 9485
rect 10409 9482 10475 9485
rect 4061 9480 10475 9482
rect 4061 9424 4066 9480
rect 4122 9424 4894 9480
rect 4950 9424 10414 9480
rect 10470 9424 10475 9480
rect 4061 9422 10475 9424
rect 4061 9419 4127 9422
rect 4889 9419 4955 9422
rect 10409 9419 10475 9422
rect 13905 9482 13971 9485
rect 17861 9482 17927 9485
rect 13905 9480 17927 9482
rect 13905 9424 13910 9480
rect 13966 9424 17866 9480
rect 17922 9424 17927 9480
rect 13905 9422 17927 9424
rect 13905 9419 13971 9422
rect 17861 9419 17927 9422
rect 0 9346 800 9376
rect 1485 9346 1551 9349
rect 0 9344 1551 9346
rect 0 9288 1490 9344
rect 1546 9288 1551 9344
rect 0 9286 1551 9288
rect 0 9256 800 9286
rect 1485 9283 1551 9286
rect 1945 9346 2011 9349
rect 3509 9346 3575 9349
rect 1945 9344 3575 9346
rect 1945 9288 1950 9344
rect 2006 9288 3514 9344
rect 3570 9288 3575 9344
rect 1945 9286 3575 9288
rect 1945 9283 2011 9286
rect 3509 9283 3575 9286
rect 5993 9346 6059 9349
rect 6637 9346 6703 9349
rect 5993 9344 6703 9346
rect 5993 9288 5998 9344
rect 6054 9288 6642 9344
rect 6698 9288 6703 9344
rect 5993 9286 6703 9288
rect 5993 9283 6059 9286
rect 6637 9283 6703 9286
rect 8201 9346 8267 9349
rect 9305 9346 9371 9349
rect 8201 9344 9371 9346
rect 8201 9288 8206 9344
rect 8262 9288 9310 9344
rect 9366 9288 9371 9344
rect 8201 9286 9371 9288
rect 8201 9283 8267 9286
rect 9305 9283 9371 9286
rect 9857 9346 9923 9349
rect 11053 9346 11119 9349
rect 9857 9344 11119 9346
rect 9857 9288 9862 9344
rect 9918 9288 11058 9344
rect 11114 9288 11119 9344
rect 9857 9286 11119 9288
rect 9857 9283 9923 9286
rect 11053 9283 11119 9286
rect 6874 9280 7194 9281
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7194 9280
rect 6874 9215 7194 9216
rect 12805 9280 13125 9281
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 9215 13125 9216
rect 7741 9210 7807 9213
rect 18413 9210 18479 9213
rect 19200 9210 20000 9240
rect 7741 9208 12634 9210
rect 7741 9152 7746 9208
rect 7802 9152 12634 9208
rect 7741 9150 12634 9152
rect 7741 9147 7807 9150
rect 3417 9074 3483 9077
rect 8661 9074 8727 9077
rect 3417 9072 8727 9074
rect 3417 9016 3422 9072
rect 3478 9016 8666 9072
rect 8722 9016 8727 9072
rect 3417 9014 8727 9016
rect 12574 9074 12634 9150
rect 18413 9208 20000 9210
rect 18413 9152 18418 9208
rect 18474 9152 20000 9208
rect 18413 9150 20000 9152
rect 18413 9147 18479 9150
rect 19200 9120 20000 9150
rect 16021 9074 16087 9077
rect 12574 9072 16087 9074
rect 12574 9016 16026 9072
rect 16082 9016 16087 9072
rect 12574 9014 16087 9016
rect 3417 9011 3483 9014
rect 8661 9011 8727 9014
rect 16021 9011 16087 9014
rect 0 8938 800 8968
rect 1393 8938 1459 8941
rect 0 8936 1459 8938
rect 0 8880 1398 8936
rect 1454 8880 1459 8936
rect 0 8878 1459 8880
rect 0 8848 800 8878
rect 1393 8875 1459 8878
rect 3969 8938 4035 8941
rect 4521 8938 4587 8941
rect 9581 8938 9647 8941
rect 3969 8936 9647 8938
rect 3969 8880 3974 8936
rect 4030 8880 4526 8936
rect 4582 8880 9586 8936
rect 9642 8880 9647 8936
rect 3969 8878 9647 8880
rect 3969 8875 4035 8878
rect 4521 8875 4587 8878
rect 9581 8875 9647 8878
rect 14733 8938 14799 8941
rect 18229 8938 18295 8941
rect 14733 8936 18295 8938
rect 14733 8880 14738 8936
rect 14794 8880 18234 8936
rect 18290 8880 18295 8936
rect 14733 8878 18295 8880
rect 14733 8875 14799 8878
rect 18229 8875 18295 8878
rect 4613 8802 4679 8805
rect 18413 8802 18479 8805
rect 19200 8802 20000 8832
rect 4613 8800 9690 8802
rect 4613 8744 4618 8800
rect 4674 8744 9690 8800
rect 4613 8742 9690 8744
rect 4613 8739 4679 8742
rect 3909 8736 4229 8737
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 8671 4229 8672
rect 0 8530 800 8560
rect 2957 8530 3023 8533
rect 0 8528 3023 8530
rect 0 8472 2962 8528
rect 3018 8472 3023 8528
rect 0 8470 3023 8472
rect 9630 8530 9690 8742
rect 18413 8800 20000 8802
rect 18413 8744 18418 8800
rect 18474 8744 20000 8800
rect 18413 8742 20000 8744
rect 18413 8739 18479 8742
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 15770 8736 16090 8737
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 19200 8712 20000 8742
rect 15770 8671 16090 8672
rect 9949 8530 10015 8533
rect 10961 8530 11027 8533
rect 9630 8528 11027 8530
rect 9630 8472 9954 8528
rect 10010 8472 10966 8528
rect 11022 8472 11027 8528
rect 9630 8470 11027 8472
rect 0 8440 800 8470
rect 2957 8467 3023 8470
rect 9949 8467 10015 8470
rect 10961 8467 11027 8470
rect 5809 8394 5875 8397
rect 9397 8394 9463 8397
rect 5809 8392 9463 8394
rect 5809 8336 5814 8392
rect 5870 8336 9402 8392
rect 9458 8336 9463 8392
rect 5809 8334 9463 8336
rect 5809 8331 5875 8334
rect 9397 8331 9463 8334
rect 18505 8258 18571 8261
rect 19200 8258 20000 8288
rect 18505 8256 20000 8258
rect 18505 8200 18510 8256
rect 18566 8200 20000 8256
rect 18505 8198 20000 8200
rect 18505 8195 18571 8198
rect 6874 8192 7194 8193
rect 0 8122 800 8152
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7194 8192
rect 6874 8127 7194 8128
rect 12805 8192 13125 8193
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 19200 8168 20000 8198
rect 12805 8127 13125 8128
rect 1853 8122 1919 8125
rect 0 8120 1919 8122
rect 0 8064 1858 8120
rect 1914 8064 1919 8120
rect 0 8062 1919 8064
rect 0 8032 800 8062
rect 1853 8059 1919 8062
rect 15653 8122 15719 8125
rect 16297 8122 16363 8125
rect 15653 8120 16363 8122
rect 15653 8064 15658 8120
rect 15714 8064 16302 8120
rect 16358 8064 16363 8120
rect 15653 8062 16363 8064
rect 15653 8059 15719 8062
rect 16297 8059 16363 8062
rect 11973 7986 12039 7989
rect 13997 7986 14063 7989
rect 11973 7984 14063 7986
rect 11973 7928 11978 7984
rect 12034 7928 14002 7984
rect 14058 7928 14063 7984
rect 11973 7926 14063 7928
rect 11973 7923 12039 7926
rect 13997 7923 14063 7926
rect 1761 7850 1827 7853
rect 12801 7850 12867 7853
rect 1761 7848 12867 7850
rect 1761 7792 1766 7848
rect 1822 7792 12806 7848
rect 12862 7792 12867 7848
rect 1761 7790 12867 7792
rect 1761 7787 1827 7790
rect 12801 7787 12867 7790
rect 18505 7850 18571 7853
rect 19200 7850 20000 7880
rect 18505 7848 20000 7850
rect 18505 7792 18510 7848
rect 18566 7792 20000 7848
rect 18505 7790 20000 7792
rect 18505 7787 18571 7790
rect 19200 7760 20000 7790
rect 0 7714 800 7744
rect 1485 7714 1551 7717
rect 0 7712 1551 7714
rect 0 7656 1490 7712
rect 1546 7656 1551 7712
rect 0 7654 1551 7656
rect 0 7624 800 7654
rect 1485 7651 1551 7654
rect 4981 7714 5047 7717
rect 4981 7712 9690 7714
rect 4981 7656 4986 7712
rect 5042 7656 9690 7712
rect 4981 7654 9690 7656
rect 4981 7651 5047 7654
rect 3909 7648 4229 7649
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 7583 4229 7584
rect 5349 7578 5415 7581
rect 9305 7578 9371 7581
rect 5349 7576 9371 7578
rect 5349 7520 5354 7576
rect 5410 7520 9310 7576
rect 9366 7520 9371 7576
rect 5349 7518 9371 7520
rect 5349 7515 5415 7518
rect 9305 7515 9371 7518
rect 8385 7442 8451 7445
rect 9305 7442 9371 7445
rect 8385 7440 9371 7442
rect 8385 7384 8390 7440
rect 8446 7384 9310 7440
rect 9366 7384 9371 7440
rect 8385 7382 9371 7384
rect 9630 7442 9690 7654
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 15770 7648 16090 7649
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 7583 16090 7584
rect 12341 7578 12407 7581
rect 13813 7578 13879 7581
rect 12341 7576 13879 7578
rect 12341 7520 12346 7576
rect 12402 7520 13818 7576
rect 13874 7520 13879 7576
rect 12341 7518 13879 7520
rect 12341 7515 12407 7518
rect 13813 7515 13879 7518
rect 13721 7442 13787 7445
rect 9630 7440 13787 7442
rect 9630 7384 13726 7440
rect 13782 7384 13787 7440
rect 9630 7382 13787 7384
rect 8385 7379 8451 7382
rect 9305 7379 9371 7382
rect 13721 7379 13787 7382
rect 14273 7442 14339 7445
rect 17493 7442 17559 7445
rect 14273 7440 17559 7442
rect 14273 7384 14278 7440
rect 14334 7384 17498 7440
rect 17554 7384 17559 7440
rect 14273 7382 17559 7384
rect 14273 7379 14339 7382
rect 17493 7379 17559 7382
rect 18137 7442 18203 7445
rect 19200 7442 20000 7472
rect 18137 7440 20000 7442
rect 18137 7384 18142 7440
rect 18198 7384 20000 7440
rect 18137 7382 20000 7384
rect 18137 7379 18203 7382
rect 19200 7352 20000 7382
rect 0 7306 800 7336
rect 1393 7306 1459 7309
rect 0 7304 1459 7306
rect 0 7248 1398 7304
rect 1454 7248 1459 7304
rect 0 7246 1459 7248
rect 0 7216 800 7246
rect 1393 7243 1459 7246
rect 12341 7306 12407 7309
rect 16665 7306 16731 7309
rect 12341 7304 16731 7306
rect 12341 7248 12346 7304
rect 12402 7248 16670 7304
rect 16726 7248 16731 7304
rect 12341 7246 16731 7248
rect 12341 7243 12407 7246
rect 16665 7243 16731 7246
rect 6874 7104 7194 7105
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7194 7104
rect 6874 7039 7194 7040
rect 12805 7104 13125 7105
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 7039 13125 7040
rect 13721 7034 13787 7037
rect 17677 7034 17743 7037
rect 13721 7032 17743 7034
rect 13721 6976 13726 7032
rect 13782 6976 17682 7032
rect 17738 6976 17743 7032
rect 13721 6974 17743 6976
rect 13721 6971 13787 6974
rect 17677 6971 17743 6974
rect 18505 7034 18571 7037
rect 19200 7034 20000 7064
rect 18505 7032 20000 7034
rect 18505 6976 18510 7032
rect 18566 6976 20000 7032
rect 18505 6974 20000 6976
rect 18505 6971 18571 6974
rect 19200 6944 20000 6974
rect 0 6898 800 6928
rect 1761 6898 1827 6901
rect 0 6896 1827 6898
rect 0 6840 1766 6896
rect 1822 6840 1827 6896
rect 0 6838 1827 6840
rect 0 6808 800 6838
rect 1761 6835 1827 6838
rect 11329 6898 11395 6901
rect 13353 6898 13419 6901
rect 11329 6896 13419 6898
rect 11329 6840 11334 6896
rect 11390 6840 13358 6896
rect 13414 6840 13419 6896
rect 11329 6838 13419 6840
rect 11329 6835 11395 6838
rect 13353 6835 13419 6838
rect 13721 6898 13787 6901
rect 15745 6898 15811 6901
rect 13721 6896 15811 6898
rect 13721 6840 13726 6896
rect 13782 6840 15750 6896
rect 15806 6840 15811 6896
rect 13721 6838 15811 6840
rect 13721 6835 13787 6838
rect 15745 6835 15811 6838
rect 10777 6762 10843 6765
rect 15837 6762 15903 6765
rect 17125 6762 17191 6765
rect 10777 6760 17191 6762
rect 10777 6704 10782 6760
rect 10838 6704 15842 6760
rect 15898 6704 17130 6760
rect 17186 6704 17191 6760
rect 10777 6702 17191 6704
rect 10777 6699 10843 6702
rect 15837 6699 15903 6702
rect 17125 6699 17191 6702
rect 18505 6626 18571 6629
rect 19200 6626 20000 6656
rect 18505 6624 20000 6626
rect 18505 6568 18510 6624
rect 18566 6568 20000 6624
rect 18505 6566 20000 6568
rect 18505 6563 18571 6566
rect 3909 6560 4229 6561
rect 0 6490 800 6520
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 6495 4229 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 15770 6560 16090 6561
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 19200 6536 20000 6566
rect 15770 6495 16090 6496
rect 1485 6490 1551 6493
rect 0 6488 1551 6490
rect 0 6432 1490 6488
rect 1546 6432 1551 6488
rect 0 6430 1551 6432
rect 0 6400 800 6430
rect 1485 6427 1551 6430
rect 13169 6490 13235 6493
rect 14273 6490 14339 6493
rect 13169 6488 14339 6490
rect 13169 6432 13174 6488
rect 13230 6432 14278 6488
rect 14334 6432 14339 6488
rect 13169 6430 14339 6432
rect 13169 6427 13235 6430
rect 14273 6427 14339 6430
rect 3141 6354 3207 6357
rect 4889 6354 4955 6357
rect 3141 6352 4955 6354
rect 3141 6296 3146 6352
rect 3202 6296 4894 6352
rect 4950 6296 4955 6352
rect 3141 6294 4955 6296
rect 3141 6291 3207 6294
rect 4889 6291 4955 6294
rect 8201 6354 8267 6357
rect 16665 6354 16731 6357
rect 8201 6352 16731 6354
rect 8201 6296 8206 6352
rect 8262 6296 16670 6352
rect 16726 6296 16731 6352
rect 8201 6294 16731 6296
rect 8201 6291 8267 6294
rect 16665 6291 16731 6294
rect 13721 6218 13787 6221
rect 8250 6216 13787 6218
rect 8250 6160 13726 6216
rect 13782 6160 13787 6216
rect 8250 6158 13787 6160
rect 0 6082 800 6112
rect 1485 6082 1551 6085
rect 0 6080 1551 6082
rect 0 6024 1490 6080
rect 1546 6024 1551 6080
rect 0 6022 1551 6024
rect 0 5992 800 6022
rect 1485 6019 1551 6022
rect 6874 6016 7194 6017
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7194 6016
rect 6874 5951 7194 5952
rect 4245 5946 4311 5949
rect 5349 5946 5415 5949
rect 4245 5944 5415 5946
rect 4245 5888 4250 5944
rect 4306 5888 5354 5944
rect 5410 5888 5415 5944
rect 4245 5886 5415 5888
rect 4245 5883 4311 5886
rect 5349 5883 5415 5886
rect 7281 5946 7347 5949
rect 8250 5946 8310 6158
rect 13721 6155 13787 6158
rect 14641 6218 14707 6221
rect 18505 6218 18571 6221
rect 19200 6218 20000 6248
rect 14641 6216 15256 6218
rect 14641 6160 14646 6216
rect 14702 6160 15256 6216
rect 14641 6158 15256 6160
rect 14641 6155 14707 6158
rect 15196 6085 15256 6158
rect 18505 6216 20000 6218
rect 18505 6160 18510 6216
rect 18566 6160 20000 6216
rect 18505 6158 20000 6160
rect 18505 6155 18571 6158
rect 19200 6128 20000 6158
rect 15193 6080 15259 6085
rect 15193 6024 15198 6080
rect 15254 6024 15259 6080
rect 15193 6019 15259 6024
rect 12805 6016 13125 6017
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 5951 13125 5952
rect 7281 5944 8310 5946
rect 7281 5888 7286 5944
rect 7342 5888 8310 5944
rect 7281 5886 8310 5888
rect 7281 5883 7347 5886
rect 3601 5810 3667 5813
rect 5901 5810 5967 5813
rect 3601 5808 5967 5810
rect 3601 5752 3606 5808
rect 3662 5752 5906 5808
rect 5962 5752 5967 5808
rect 3601 5750 5967 5752
rect 3601 5747 3667 5750
rect 5901 5747 5967 5750
rect 12065 5810 12131 5813
rect 16389 5810 16455 5813
rect 12065 5808 16455 5810
rect 12065 5752 12070 5808
rect 12126 5752 16394 5808
rect 16450 5752 16455 5808
rect 12065 5750 16455 5752
rect 12065 5747 12131 5750
rect 16389 5747 16455 5750
rect 4245 5674 4311 5677
rect 5717 5674 5783 5677
rect 4245 5672 5783 5674
rect 4245 5616 4250 5672
rect 4306 5616 5722 5672
rect 5778 5616 5783 5672
rect 4245 5614 5783 5616
rect 4245 5611 4311 5614
rect 5717 5611 5783 5614
rect 7373 5674 7439 5677
rect 7741 5674 7807 5677
rect 8385 5674 8451 5677
rect 7373 5672 8451 5674
rect 7373 5616 7378 5672
rect 7434 5616 7746 5672
rect 7802 5616 8390 5672
rect 8446 5616 8451 5672
rect 7373 5614 8451 5616
rect 7373 5611 7439 5614
rect 7741 5611 7807 5614
rect 8385 5611 8451 5614
rect 14641 5674 14707 5677
rect 16757 5674 16823 5677
rect 14641 5672 16823 5674
rect 14641 5616 14646 5672
rect 14702 5616 16762 5672
rect 16818 5616 16823 5672
rect 14641 5614 16823 5616
rect 14641 5611 14707 5614
rect 16757 5611 16823 5614
rect 18505 5674 18571 5677
rect 19200 5674 20000 5704
rect 18505 5672 20000 5674
rect 18505 5616 18510 5672
rect 18566 5616 20000 5672
rect 18505 5614 20000 5616
rect 18505 5611 18571 5614
rect 19200 5584 20000 5614
rect 0 5538 800 5568
rect 1485 5538 1551 5541
rect 0 5536 1551 5538
rect 0 5480 1490 5536
rect 1546 5480 1551 5536
rect 0 5478 1551 5480
rect 0 5448 800 5478
rect 1485 5475 1551 5478
rect 3909 5472 4229 5473
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 5407 4229 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 15770 5472 16090 5473
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 5407 16090 5408
rect 2589 5266 2655 5269
rect 6361 5266 6427 5269
rect 2589 5264 6427 5266
rect 2589 5208 2594 5264
rect 2650 5208 6366 5264
rect 6422 5208 6427 5264
rect 2589 5206 6427 5208
rect 2589 5203 2655 5206
rect 6361 5203 6427 5206
rect 14641 5266 14707 5269
rect 17861 5266 17927 5269
rect 14641 5264 17927 5266
rect 14641 5208 14646 5264
rect 14702 5208 17866 5264
rect 17922 5208 17927 5264
rect 14641 5206 17927 5208
rect 14641 5203 14707 5206
rect 17861 5203 17927 5206
rect 18505 5266 18571 5269
rect 19200 5266 20000 5296
rect 18505 5264 20000 5266
rect 18505 5208 18510 5264
rect 18566 5208 20000 5264
rect 18505 5206 20000 5208
rect 18505 5203 18571 5206
rect 19200 5176 20000 5206
rect 0 5130 800 5160
rect 1393 5130 1459 5133
rect 0 5128 1459 5130
rect 0 5072 1398 5128
rect 1454 5072 1459 5128
rect 0 5070 1459 5072
rect 0 5040 800 5070
rect 1393 5067 1459 5070
rect 13813 5130 13879 5133
rect 14733 5130 14799 5133
rect 16849 5130 16915 5133
rect 13813 5128 16915 5130
rect 13813 5072 13818 5128
rect 13874 5072 14738 5128
rect 14794 5072 16854 5128
rect 16910 5072 16915 5128
rect 13813 5070 16915 5072
rect 13813 5067 13879 5070
rect 14733 5067 14799 5070
rect 16849 5067 16915 5070
rect 6874 4928 7194 4929
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7194 4928
rect 6874 4863 7194 4864
rect 12805 4928 13125 4929
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 4863 13125 4864
rect 18137 4858 18203 4861
rect 19200 4858 20000 4888
rect 18137 4856 20000 4858
rect 18137 4800 18142 4856
rect 18198 4800 20000 4856
rect 18137 4798 20000 4800
rect 18137 4795 18203 4798
rect 19200 4768 20000 4798
rect 0 4722 800 4752
rect 1393 4722 1459 4725
rect 0 4720 1459 4722
rect 0 4664 1398 4720
rect 1454 4664 1459 4720
rect 0 4662 1459 4664
rect 0 4632 800 4662
rect 1393 4659 1459 4662
rect 13445 4722 13511 4725
rect 17033 4722 17099 4725
rect 13445 4720 17099 4722
rect 13445 4664 13450 4720
rect 13506 4664 17038 4720
rect 17094 4664 17099 4720
rect 13445 4662 17099 4664
rect 13445 4659 13511 4662
rect 17033 4659 17099 4662
rect 15377 4586 15443 4589
rect 15745 4586 15811 4589
rect 15377 4584 15811 4586
rect 15377 4528 15382 4584
rect 15438 4528 15750 4584
rect 15806 4528 15811 4584
rect 15377 4526 15811 4528
rect 15377 4523 15443 4526
rect 15745 4523 15811 4526
rect 18505 4450 18571 4453
rect 19200 4450 20000 4480
rect 18505 4448 20000 4450
rect 18505 4392 18510 4448
rect 18566 4392 20000 4448
rect 18505 4390 20000 4392
rect 18505 4387 18571 4390
rect 3909 4384 4229 4385
rect 0 4314 800 4344
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 4319 4229 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 15770 4384 16090 4385
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 19200 4360 20000 4390
rect 15770 4319 16090 4320
rect 1853 4314 1919 4317
rect 0 4312 1919 4314
rect 0 4256 1858 4312
rect 1914 4256 1919 4312
rect 0 4254 1919 4256
rect 0 4224 800 4254
rect 1853 4251 1919 4254
rect 18137 4042 18203 4045
rect 19200 4042 20000 4072
rect 18137 4040 20000 4042
rect 18137 3984 18142 4040
rect 18198 3984 20000 4040
rect 18137 3982 20000 3984
rect 18137 3979 18203 3982
rect 19200 3952 20000 3982
rect 0 3906 800 3936
rect 2221 3906 2287 3909
rect 0 3904 2287 3906
rect 0 3848 2226 3904
rect 2282 3848 2287 3904
rect 0 3846 2287 3848
rect 0 3816 800 3846
rect 2221 3843 2287 3846
rect 6874 3840 7194 3841
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7194 3840
rect 6874 3775 7194 3776
rect 12805 3840 13125 3841
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 3775 13125 3776
rect 18505 3634 18571 3637
rect 19200 3634 20000 3664
rect 18505 3632 20000 3634
rect 18505 3576 18510 3632
rect 18566 3576 20000 3632
rect 18505 3574 20000 3576
rect 18505 3571 18571 3574
rect 19200 3544 20000 3574
rect 0 3498 800 3528
rect 1853 3498 1919 3501
rect 0 3496 1919 3498
rect 0 3440 1858 3496
rect 1914 3440 1919 3496
rect 0 3438 1919 3440
rect 0 3408 800 3438
rect 1853 3435 1919 3438
rect 10593 3498 10659 3501
rect 12801 3498 12867 3501
rect 10593 3496 12867 3498
rect 10593 3440 10598 3496
rect 10654 3440 12806 3496
rect 12862 3440 12867 3496
rect 10593 3438 12867 3440
rect 10593 3435 10659 3438
rect 12801 3435 12867 3438
rect 10593 3362 10659 3365
rect 14457 3362 14523 3365
rect 10593 3360 14523 3362
rect 10593 3304 10598 3360
rect 10654 3304 14462 3360
rect 14518 3304 14523 3360
rect 10593 3302 14523 3304
rect 10593 3299 10659 3302
rect 14457 3299 14523 3302
rect 3909 3296 4229 3297
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 3231 4229 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 15770 3296 16090 3297
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 3231 16090 3232
rect 10869 3226 10935 3229
rect 14273 3226 14339 3229
rect 10869 3224 14339 3226
rect 10869 3168 10874 3224
rect 10930 3168 14278 3224
rect 14334 3168 14339 3224
rect 10869 3166 14339 3168
rect 10869 3163 10935 3166
rect 14273 3163 14339 3166
rect 18137 3226 18203 3229
rect 19200 3226 20000 3256
rect 18137 3224 20000 3226
rect 18137 3168 18142 3224
rect 18198 3168 20000 3224
rect 18137 3166 20000 3168
rect 18137 3163 18203 3166
rect 19200 3136 20000 3166
rect 0 3090 800 3120
rect 2221 3090 2287 3093
rect 0 3088 2287 3090
rect 0 3032 2226 3088
rect 2282 3032 2287 3088
rect 0 3030 2287 3032
rect 0 3000 800 3030
rect 2221 3027 2287 3030
rect 12985 3090 13051 3093
rect 13445 3090 13511 3093
rect 12985 3088 13511 3090
rect 12985 3032 12990 3088
rect 13046 3032 13450 3088
rect 13506 3032 13511 3088
rect 12985 3030 13511 3032
rect 12985 3027 13051 3030
rect 13445 3027 13511 3030
rect 14457 3090 14523 3093
rect 15745 3090 15811 3093
rect 14457 3088 15811 3090
rect 14457 3032 14462 3088
rect 14518 3032 15750 3088
rect 15806 3032 15811 3088
rect 14457 3030 15811 3032
rect 14457 3027 14523 3030
rect 15745 3027 15811 3030
rect 4061 2954 4127 2957
rect 14917 2954 14983 2957
rect 4061 2952 14983 2954
rect 4061 2896 4066 2952
rect 4122 2896 14922 2952
rect 14978 2896 14983 2952
rect 4061 2894 14983 2896
rect 4061 2891 4127 2894
rect 14917 2891 14983 2894
rect 10225 2818 10291 2821
rect 10869 2818 10935 2821
rect 10225 2816 10935 2818
rect 10225 2760 10230 2816
rect 10286 2760 10874 2816
rect 10930 2760 10935 2816
rect 10225 2758 10935 2760
rect 10225 2755 10291 2758
rect 10869 2755 10935 2758
rect 6874 2752 7194 2753
rect 0 2682 800 2712
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7194 2752
rect 6874 2687 7194 2688
rect 12805 2752 13125 2753
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2687 13125 2688
rect 1485 2682 1551 2685
rect 0 2680 1551 2682
rect 0 2624 1490 2680
rect 1546 2624 1551 2680
rect 0 2622 1551 2624
rect 0 2592 800 2622
rect 1485 2619 1551 2622
rect 17769 2682 17835 2685
rect 19200 2682 20000 2712
rect 17769 2680 20000 2682
rect 17769 2624 17774 2680
rect 17830 2624 20000 2680
rect 17769 2622 20000 2624
rect 17769 2619 17835 2622
rect 19200 2592 20000 2622
rect 17861 2546 17927 2549
rect 17861 2544 18154 2546
rect 17861 2488 17866 2544
rect 17922 2488 18154 2544
rect 17861 2486 18154 2488
rect 17861 2483 17927 2486
rect 0 2274 800 2304
rect 1853 2274 1919 2277
rect 0 2272 1919 2274
rect 0 2216 1858 2272
rect 1914 2216 1919 2272
rect 0 2214 1919 2216
rect 18094 2274 18154 2486
rect 19200 2274 20000 2304
rect 18094 2214 20000 2274
rect 0 2184 800 2214
rect 1853 2211 1919 2214
rect 3909 2208 4229 2209
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2143 4229 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 15770 2208 16090 2209
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 19200 2184 20000 2214
rect 15770 2143 16090 2144
rect 0 1866 800 1896
rect 2221 1866 2287 1869
rect 0 1864 2287 1866
rect 0 1808 2226 1864
rect 2282 1808 2287 1864
rect 0 1806 2287 1808
rect 0 1776 800 1806
rect 2221 1803 2287 1806
rect 17401 1866 17467 1869
rect 19200 1866 20000 1896
rect 17401 1864 20000 1866
rect 17401 1808 17406 1864
rect 17462 1808 20000 1864
rect 17401 1806 20000 1808
rect 17401 1803 17467 1806
rect 19200 1776 20000 1806
rect 0 1458 800 1488
rect 1393 1458 1459 1461
rect 0 1456 1459 1458
rect 0 1400 1398 1456
rect 1454 1400 1459 1456
rect 0 1398 1459 1400
rect 0 1368 800 1398
rect 1393 1395 1459 1398
rect 17493 1458 17559 1461
rect 19200 1458 20000 1488
rect 17493 1456 20000 1458
rect 17493 1400 17498 1456
rect 17554 1400 20000 1456
rect 17493 1398 20000 1400
rect 17493 1395 17559 1398
rect 19200 1368 20000 1398
rect 0 1050 800 1080
rect 1761 1050 1827 1053
rect 0 1048 1827 1050
rect 0 992 1766 1048
rect 1822 992 1827 1048
rect 0 990 1827 992
rect 0 960 800 990
rect 1761 987 1827 990
rect 17769 1050 17835 1053
rect 19200 1050 20000 1080
rect 17769 1048 20000 1050
rect 17769 992 17774 1048
rect 17830 992 20000 1048
rect 17769 990 20000 992
rect 17769 987 17835 990
rect 19200 960 20000 990
rect 0 642 800 672
rect 1301 642 1367 645
rect 0 640 1367 642
rect 0 584 1306 640
rect 1362 584 1367 640
rect 0 582 1367 584
rect 0 552 800 582
rect 1301 579 1367 582
rect 17677 642 17743 645
rect 19200 642 20000 672
rect 17677 640 20000 642
rect 17677 584 17682 640
rect 17738 584 20000 640
rect 17677 582 20000 584
rect 17677 579 17743 582
rect 19200 552 20000 582
rect 0 234 800 264
rect 3325 234 3391 237
rect 0 232 3391 234
rect 0 176 3330 232
rect 3386 176 3391 232
rect 0 174 3391 176
rect 0 144 800 174
rect 3325 171 3391 174
rect 17861 234 17927 237
rect 19200 234 20000 264
rect 17861 232 20000 234
rect 17861 176 17866 232
rect 17922 176 20000 232
rect 17861 174 20000 176
rect 17861 171 17927 174
rect 19200 144 20000 174
<< via3 >>
rect 6882 14716 6946 14720
rect 6882 14660 6886 14716
rect 6886 14660 6942 14716
rect 6942 14660 6946 14716
rect 6882 14656 6946 14660
rect 6962 14716 7026 14720
rect 6962 14660 6966 14716
rect 6966 14660 7022 14716
rect 7022 14660 7026 14716
rect 6962 14656 7026 14660
rect 7042 14716 7106 14720
rect 7042 14660 7046 14716
rect 7046 14660 7102 14716
rect 7102 14660 7106 14716
rect 7042 14656 7106 14660
rect 7122 14716 7186 14720
rect 7122 14660 7126 14716
rect 7126 14660 7182 14716
rect 7182 14660 7186 14716
rect 7122 14656 7186 14660
rect 12813 14716 12877 14720
rect 12813 14660 12817 14716
rect 12817 14660 12873 14716
rect 12873 14660 12877 14716
rect 12813 14656 12877 14660
rect 12893 14716 12957 14720
rect 12893 14660 12897 14716
rect 12897 14660 12953 14716
rect 12953 14660 12957 14716
rect 12893 14656 12957 14660
rect 12973 14716 13037 14720
rect 12973 14660 12977 14716
rect 12977 14660 13033 14716
rect 13033 14660 13037 14716
rect 12973 14656 13037 14660
rect 13053 14716 13117 14720
rect 13053 14660 13057 14716
rect 13057 14660 13113 14716
rect 13113 14660 13117 14716
rect 13053 14656 13117 14660
rect 3917 14172 3981 14176
rect 3917 14116 3921 14172
rect 3921 14116 3977 14172
rect 3977 14116 3981 14172
rect 3917 14112 3981 14116
rect 3997 14172 4061 14176
rect 3997 14116 4001 14172
rect 4001 14116 4057 14172
rect 4057 14116 4061 14172
rect 3997 14112 4061 14116
rect 4077 14172 4141 14176
rect 4077 14116 4081 14172
rect 4081 14116 4137 14172
rect 4137 14116 4141 14172
rect 4077 14112 4141 14116
rect 4157 14172 4221 14176
rect 4157 14116 4161 14172
rect 4161 14116 4217 14172
rect 4217 14116 4221 14172
rect 4157 14112 4221 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 15778 14172 15842 14176
rect 15778 14116 15782 14172
rect 15782 14116 15838 14172
rect 15838 14116 15842 14172
rect 15778 14112 15842 14116
rect 15858 14172 15922 14176
rect 15858 14116 15862 14172
rect 15862 14116 15918 14172
rect 15918 14116 15922 14172
rect 15858 14112 15922 14116
rect 15938 14172 16002 14176
rect 15938 14116 15942 14172
rect 15942 14116 15998 14172
rect 15998 14116 16002 14172
rect 15938 14112 16002 14116
rect 16018 14172 16082 14176
rect 16018 14116 16022 14172
rect 16022 14116 16078 14172
rect 16078 14116 16082 14172
rect 16018 14112 16082 14116
rect 6882 13628 6946 13632
rect 6882 13572 6886 13628
rect 6886 13572 6942 13628
rect 6942 13572 6946 13628
rect 6882 13568 6946 13572
rect 6962 13628 7026 13632
rect 6962 13572 6966 13628
rect 6966 13572 7022 13628
rect 7022 13572 7026 13628
rect 6962 13568 7026 13572
rect 7042 13628 7106 13632
rect 7042 13572 7046 13628
rect 7046 13572 7102 13628
rect 7102 13572 7106 13628
rect 7042 13568 7106 13572
rect 7122 13628 7186 13632
rect 7122 13572 7126 13628
rect 7126 13572 7182 13628
rect 7182 13572 7186 13628
rect 7122 13568 7186 13572
rect 12813 13628 12877 13632
rect 12813 13572 12817 13628
rect 12817 13572 12873 13628
rect 12873 13572 12877 13628
rect 12813 13568 12877 13572
rect 12893 13628 12957 13632
rect 12893 13572 12897 13628
rect 12897 13572 12953 13628
rect 12953 13572 12957 13628
rect 12893 13568 12957 13572
rect 12973 13628 13037 13632
rect 12973 13572 12977 13628
rect 12977 13572 13033 13628
rect 13033 13572 13037 13628
rect 12973 13568 13037 13572
rect 13053 13628 13117 13632
rect 13053 13572 13057 13628
rect 13057 13572 13113 13628
rect 13113 13572 13117 13628
rect 13053 13568 13117 13572
rect 3917 13084 3981 13088
rect 3917 13028 3921 13084
rect 3921 13028 3977 13084
rect 3977 13028 3981 13084
rect 3917 13024 3981 13028
rect 3997 13084 4061 13088
rect 3997 13028 4001 13084
rect 4001 13028 4057 13084
rect 4057 13028 4061 13084
rect 3997 13024 4061 13028
rect 4077 13084 4141 13088
rect 4077 13028 4081 13084
rect 4081 13028 4137 13084
rect 4137 13028 4141 13084
rect 4077 13024 4141 13028
rect 4157 13084 4221 13088
rect 4157 13028 4161 13084
rect 4161 13028 4217 13084
rect 4217 13028 4221 13084
rect 4157 13024 4221 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 15778 13084 15842 13088
rect 15778 13028 15782 13084
rect 15782 13028 15838 13084
rect 15838 13028 15842 13084
rect 15778 13024 15842 13028
rect 15858 13084 15922 13088
rect 15858 13028 15862 13084
rect 15862 13028 15918 13084
rect 15918 13028 15922 13084
rect 15858 13024 15922 13028
rect 15938 13084 16002 13088
rect 15938 13028 15942 13084
rect 15942 13028 15998 13084
rect 15998 13028 16002 13084
rect 15938 13024 16002 13028
rect 16018 13084 16082 13088
rect 16018 13028 16022 13084
rect 16022 13028 16078 13084
rect 16078 13028 16082 13084
rect 16018 13024 16082 13028
rect 6882 12540 6946 12544
rect 6882 12484 6886 12540
rect 6886 12484 6942 12540
rect 6942 12484 6946 12540
rect 6882 12480 6946 12484
rect 6962 12540 7026 12544
rect 6962 12484 6966 12540
rect 6966 12484 7022 12540
rect 7022 12484 7026 12540
rect 6962 12480 7026 12484
rect 7042 12540 7106 12544
rect 7042 12484 7046 12540
rect 7046 12484 7102 12540
rect 7102 12484 7106 12540
rect 7042 12480 7106 12484
rect 7122 12540 7186 12544
rect 7122 12484 7126 12540
rect 7126 12484 7182 12540
rect 7182 12484 7186 12540
rect 7122 12480 7186 12484
rect 12813 12540 12877 12544
rect 12813 12484 12817 12540
rect 12817 12484 12873 12540
rect 12873 12484 12877 12540
rect 12813 12480 12877 12484
rect 12893 12540 12957 12544
rect 12893 12484 12897 12540
rect 12897 12484 12953 12540
rect 12953 12484 12957 12540
rect 12893 12480 12957 12484
rect 12973 12540 13037 12544
rect 12973 12484 12977 12540
rect 12977 12484 13033 12540
rect 13033 12484 13037 12540
rect 12973 12480 13037 12484
rect 13053 12540 13117 12544
rect 13053 12484 13057 12540
rect 13057 12484 13113 12540
rect 13113 12484 13117 12540
rect 13053 12480 13117 12484
rect 3917 11996 3981 12000
rect 3917 11940 3921 11996
rect 3921 11940 3977 11996
rect 3977 11940 3981 11996
rect 3917 11936 3981 11940
rect 3997 11996 4061 12000
rect 3997 11940 4001 11996
rect 4001 11940 4057 11996
rect 4057 11940 4061 11996
rect 3997 11936 4061 11940
rect 4077 11996 4141 12000
rect 4077 11940 4081 11996
rect 4081 11940 4137 11996
rect 4137 11940 4141 11996
rect 4077 11936 4141 11940
rect 4157 11996 4221 12000
rect 4157 11940 4161 11996
rect 4161 11940 4217 11996
rect 4217 11940 4221 11996
rect 4157 11936 4221 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 15778 11996 15842 12000
rect 15778 11940 15782 11996
rect 15782 11940 15838 11996
rect 15838 11940 15842 11996
rect 15778 11936 15842 11940
rect 15858 11996 15922 12000
rect 15858 11940 15862 11996
rect 15862 11940 15918 11996
rect 15918 11940 15922 11996
rect 15858 11936 15922 11940
rect 15938 11996 16002 12000
rect 15938 11940 15942 11996
rect 15942 11940 15998 11996
rect 15998 11940 16002 11996
rect 15938 11936 16002 11940
rect 16018 11996 16082 12000
rect 16018 11940 16022 11996
rect 16022 11940 16078 11996
rect 16078 11940 16082 11996
rect 16018 11936 16082 11940
rect 6882 11452 6946 11456
rect 6882 11396 6886 11452
rect 6886 11396 6942 11452
rect 6942 11396 6946 11452
rect 6882 11392 6946 11396
rect 6962 11452 7026 11456
rect 6962 11396 6966 11452
rect 6966 11396 7022 11452
rect 7022 11396 7026 11452
rect 6962 11392 7026 11396
rect 7042 11452 7106 11456
rect 7042 11396 7046 11452
rect 7046 11396 7102 11452
rect 7102 11396 7106 11452
rect 7042 11392 7106 11396
rect 7122 11452 7186 11456
rect 7122 11396 7126 11452
rect 7126 11396 7182 11452
rect 7182 11396 7186 11452
rect 7122 11392 7186 11396
rect 12813 11452 12877 11456
rect 12813 11396 12817 11452
rect 12817 11396 12873 11452
rect 12873 11396 12877 11452
rect 12813 11392 12877 11396
rect 12893 11452 12957 11456
rect 12893 11396 12897 11452
rect 12897 11396 12953 11452
rect 12953 11396 12957 11452
rect 12893 11392 12957 11396
rect 12973 11452 13037 11456
rect 12973 11396 12977 11452
rect 12977 11396 13033 11452
rect 13033 11396 13037 11452
rect 12973 11392 13037 11396
rect 13053 11452 13117 11456
rect 13053 11396 13057 11452
rect 13057 11396 13113 11452
rect 13113 11396 13117 11452
rect 13053 11392 13117 11396
rect 3917 10908 3981 10912
rect 3917 10852 3921 10908
rect 3921 10852 3977 10908
rect 3977 10852 3981 10908
rect 3917 10848 3981 10852
rect 3997 10908 4061 10912
rect 3997 10852 4001 10908
rect 4001 10852 4057 10908
rect 4057 10852 4061 10908
rect 3997 10848 4061 10852
rect 4077 10908 4141 10912
rect 4077 10852 4081 10908
rect 4081 10852 4137 10908
rect 4137 10852 4141 10908
rect 4077 10848 4141 10852
rect 4157 10908 4221 10912
rect 4157 10852 4161 10908
rect 4161 10852 4217 10908
rect 4217 10852 4221 10908
rect 4157 10848 4221 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 15778 10908 15842 10912
rect 15778 10852 15782 10908
rect 15782 10852 15838 10908
rect 15838 10852 15842 10908
rect 15778 10848 15842 10852
rect 15858 10908 15922 10912
rect 15858 10852 15862 10908
rect 15862 10852 15918 10908
rect 15918 10852 15922 10908
rect 15858 10848 15922 10852
rect 15938 10908 16002 10912
rect 15938 10852 15942 10908
rect 15942 10852 15998 10908
rect 15998 10852 16002 10908
rect 15938 10848 16002 10852
rect 16018 10908 16082 10912
rect 16018 10852 16022 10908
rect 16022 10852 16078 10908
rect 16078 10852 16082 10908
rect 16018 10848 16082 10852
rect 6882 10364 6946 10368
rect 6882 10308 6886 10364
rect 6886 10308 6942 10364
rect 6942 10308 6946 10364
rect 6882 10304 6946 10308
rect 6962 10364 7026 10368
rect 6962 10308 6966 10364
rect 6966 10308 7022 10364
rect 7022 10308 7026 10364
rect 6962 10304 7026 10308
rect 7042 10364 7106 10368
rect 7042 10308 7046 10364
rect 7046 10308 7102 10364
rect 7102 10308 7106 10364
rect 7042 10304 7106 10308
rect 7122 10364 7186 10368
rect 7122 10308 7126 10364
rect 7126 10308 7182 10364
rect 7182 10308 7186 10364
rect 7122 10304 7186 10308
rect 12813 10364 12877 10368
rect 12813 10308 12817 10364
rect 12817 10308 12873 10364
rect 12873 10308 12877 10364
rect 12813 10304 12877 10308
rect 12893 10364 12957 10368
rect 12893 10308 12897 10364
rect 12897 10308 12953 10364
rect 12953 10308 12957 10364
rect 12893 10304 12957 10308
rect 12973 10364 13037 10368
rect 12973 10308 12977 10364
rect 12977 10308 13033 10364
rect 13033 10308 13037 10364
rect 12973 10304 13037 10308
rect 13053 10364 13117 10368
rect 13053 10308 13057 10364
rect 13057 10308 13113 10364
rect 13113 10308 13117 10364
rect 13053 10304 13117 10308
rect 3917 9820 3981 9824
rect 3917 9764 3921 9820
rect 3921 9764 3977 9820
rect 3977 9764 3981 9820
rect 3917 9760 3981 9764
rect 3997 9820 4061 9824
rect 3997 9764 4001 9820
rect 4001 9764 4057 9820
rect 4057 9764 4061 9820
rect 3997 9760 4061 9764
rect 4077 9820 4141 9824
rect 4077 9764 4081 9820
rect 4081 9764 4137 9820
rect 4137 9764 4141 9820
rect 4077 9760 4141 9764
rect 4157 9820 4221 9824
rect 4157 9764 4161 9820
rect 4161 9764 4217 9820
rect 4217 9764 4221 9820
rect 4157 9760 4221 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 15778 9820 15842 9824
rect 15778 9764 15782 9820
rect 15782 9764 15838 9820
rect 15838 9764 15842 9820
rect 15778 9760 15842 9764
rect 15858 9820 15922 9824
rect 15858 9764 15862 9820
rect 15862 9764 15918 9820
rect 15918 9764 15922 9820
rect 15858 9760 15922 9764
rect 15938 9820 16002 9824
rect 15938 9764 15942 9820
rect 15942 9764 15998 9820
rect 15998 9764 16002 9820
rect 15938 9760 16002 9764
rect 16018 9820 16082 9824
rect 16018 9764 16022 9820
rect 16022 9764 16078 9820
rect 16078 9764 16082 9820
rect 16018 9760 16082 9764
rect 6882 9276 6946 9280
rect 6882 9220 6886 9276
rect 6886 9220 6942 9276
rect 6942 9220 6946 9276
rect 6882 9216 6946 9220
rect 6962 9276 7026 9280
rect 6962 9220 6966 9276
rect 6966 9220 7022 9276
rect 7022 9220 7026 9276
rect 6962 9216 7026 9220
rect 7042 9276 7106 9280
rect 7042 9220 7046 9276
rect 7046 9220 7102 9276
rect 7102 9220 7106 9276
rect 7042 9216 7106 9220
rect 7122 9276 7186 9280
rect 7122 9220 7126 9276
rect 7126 9220 7182 9276
rect 7182 9220 7186 9276
rect 7122 9216 7186 9220
rect 12813 9276 12877 9280
rect 12813 9220 12817 9276
rect 12817 9220 12873 9276
rect 12873 9220 12877 9276
rect 12813 9216 12877 9220
rect 12893 9276 12957 9280
rect 12893 9220 12897 9276
rect 12897 9220 12953 9276
rect 12953 9220 12957 9276
rect 12893 9216 12957 9220
rect 12973 9276 13037 9280
rect 12973 9220 12977 9276
rect 12977 9220 13033 9276
rect 13033 9220 13037 9276
rect 12973 9216 13037 9220
rect 13053 9276 13117 9280
rect 13053 9220 13057 9276
rect 13057 9220 13113 9276
rect 13113 9220 13117 9276
rect 13053 9216 13117 9220
rect 3917 8732 3981 8736
rect 3917 8676 3921 8732
rect 3921 8676 3977 8732
rect 3977 8676 3981 8732
rect 3917 8672 3981 8676
rect 3997 8732 4061 8736
rect 3997 8676 4001 8732
rect 4001 8676 4057 8732
rect 4057 8676 4061 8732
rect 3997 8672 4061 8676
rect 4077 8732 4141 8736
rect 4077 8676 4081 8732
rect 4081 8676 4137 8732
rect 4137 8676 4141 8732
rect 4077 8672 4141 8676
rect 4157 8732 4221 8736
rect 4157 8676 4161 8732
rect 4161 8676 4217 8732
rect 4217 8676 4221 8732
rect 4157 8672 4221 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 15778 8732 15842 8736
rect 15778 8676 15782 8732
rect 15782 8676 15838 8732
rect 15838 8676 15842 8732
rect 15778 8672 15842 8676
rect 15858 8732 15922 8736
rect 15858 8676 15862 8732
rect 15862 8676 15918 8732
rect 15918 8676 15922 8732
rect 15858 8672 15922 8676
rect 15938 8732 16002 8736
rect 15938 8676 15942 8732
rect 15942 8676 15998 8732
rect 15998 8676 16002 8732
rect 15938 8672 16002 8676
rect 16018 8732 16082 8736
rect 16018 8676 16022 8732
rect 16022 8676 16078 8732
rect 16078 8676 16082 8732
rect 16018 8672 16082 8676
rect 6882 8188 6946 8192
rect 6882 8132 6886 8188
rect 6886 8132 6942 8188
rect 6942 8132 6946 8188
rect 6882 8128 6946 8132
rect 6962 8188 7026 8192
rect 6962 8132 6966 8188
rect 6966 8132 7022 8188
rect 7022 8132 7026 8188
rect 6962 8128 7026 8132
rect 7042 8188 7106 8192
rect 7042 8132 7046 8188
rect 7046 8132 7102 8188
rect 7102 8132 7106 8188
rect 7042 8128 7106 8132
rect 7122 8188 7186 8192
rect 7122 8132 7126 8188
rect 7126 8132 7182 8188
rect 7182 8132 7186 8188
rect 7122 8128 7186 8132
rect 12813 8188 12877 8192
rect 12813 8132 12817 8188
rect 12817 8132 12873 8188
rect 12873 8132 12877 8188
rect 12813 8128 12877 8132
rect 12893 8188 12957 8192
rect 12893 8132 12897 8188
rect 12897 8132 12953 8188
rect 12953 8132 12957 8188
rect 12893 8128 12957 8132
rect 12973 8188 13037 8192
rect 12973 8132 12977 8188
rect 12977 8132 13033 8188
rect 13033 8132 13037 8188
rect 12973 8128 13037 8132
rect 13053 8188 13117 8192
rect 13053 8132 13057 8188
rect 13057 8132 13113 8188
rect 13113 8132 13117 8188
rect 13053 8128 13117 8132
rect 3917 7644 3981 7648
rect 3917 7588 3921 7644
rect 3921 7588 3977 7644
rect 3977 7588 3981 7644
rect 3917 7584 3981 7588
rect 3997 7644 4061 7648
rect 3997 7588 4001 7644
rect 4001 7588 4057 7644
rect 4057 7588 4061 7644
rect 3997 7584 4061 7588
rect 4077 7644 4141 7648
rect 4077 7588 4081 7644
rect 4081 7588 4137 7644
rect 4137 7588 4141 7644
rect 4077 7584 4141 7588
rect 4157 7644 4221 7648
rect 4157 7588 4161 7644
rect 4161 7588 4217 7644
rect 4217 7588 4221 7644
rect 4157 7584 4221 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 15778 7644 15842 7648
rect 15778 7588 15782 7644
rect 15782 7588 15838 7644
rect 15838 7588 15842 7644
rect 15778 7584 15842 7588
rect 15858 7644 15922 7648
rect 15858 7588 15862 7644
rect 15862 7588 15918 7644
rect 15918 7588 15922 7644
rect 15858 7584 15922 7588
rect 15938 7644 16002 7648
rect 15938 7588 15942 7644
rect 15942 7588 15998 7644
rect 15998 7588 16002 7644
rect 15938 7584 16002 7588
rect 16018 7644 16082 7648
rect 16018 7588 16022 7644
rect 16022 7588 16078 7644
rect 16078 7588 16082 7644
rect 16018 7584 16082 7588
rect 6882 7100 6946 7104
rect 6882 7044 6886 7100
rect 6886 7044 6942 7100
rect 6942 7044 6946 7100
rect 6882 7040 6946 7044
rect 6962 7100 7026 7104
rect 6962 7044 6966 7100
rect 6966 7044 7022 7100
rect 7022 7044 7026 7100
rect 6962 7040 7026 7044
rect 7042 7100 7106 7104
rect 7042 7044 7046 7100
rect 7046 7044 7102 7100
rect 7102 7044 7106 7100
rect 7042 7040 7106 7044
rect 7122 7100 7186 7104
rect 7122 7044 7126 7100
rect 7126 7044 7182 7100
rect 7182 7044 7186 7100
rect 7122 7040 7186 7044
rect 12813 7100 12877 7104
rect 12813 7044 12817 7100
rect 12817 7044 12873 7100
rect 12873 7044 12877 7100
rect 12813 7040 12877 7044
rect 12893 7100 12957 7104
rect 12893 7044 12897 7100
rect 12897 7044 12953 7100
rect 12953 7044 12957 7100
rect 12893 7040 12957 7044
rect 12973 7100 13037 7104
rect 12973 7044 12977 7100
rect 12977 7044 13033 7100
rect 13033 7044 13037 7100
rect 12973 7040 13037 7044
rect 13053 7100 13117 7104
rect 13053 7044 13057 7100
rect 13057 7044 13113 7100
rect 13113 7044 13117 7100
rect 13053 7040 13117 7044
rect 3917 6556 3981 6560
rect 3917 6500 3921 6556
rect 3921 6500 3977 6556
rect 3977 6500 3981 6556
rect 3917 6496 3981 6500
rect 3997 6556 4061 6560
rect 3997 6500 4001 6556
rect 4001 6500 4057 6556
rect 4057 6500 4061 6556
rect 3997 6496 4061 6500
rect 4077 6556 4141 6560
rect 4077 6500 4081 6556
rect 4081 6500 4137 6556
rect 4137 6500 4141 6556
rect 4077 6496 4141 6500
rect 4157 6556 4221 6560
rect 4157 6500 4161 6556
rect 4161 6500 4217 6556
rect 4217 6500 4221 6556
rect 4157 6496 4221 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 15778 6556 15842 6560
rect 15778 6500 15782 6556
rect 15782 6500 15838 6556
rect 15838 6500 15842 6556
rect 15778 6496 15842 6500
rect 15858 6556 15922 6560
rect 15858 6500 15862 6556
rect 15862 6500 15918 6556
rect 15918 6500 15922 6556
rect 15858 6496 15922 6500
rect 15938 6556 16002 6560
rect 15938 6500 15942 6556
rect 15942 6500 15998 6556
rect 15998 6500 16002 6556
rect 15938 6496 16002 6500
rect 16018 6556 16082 6560
rect 16018 6500 16022 6556
rect 16022 6500 16078 6556
rect 16078 6500 16082 6556
rect 16018 6496 16082 6500
rect 6882 6012 6946 6016
rect 6882 5956 6886 6012
rect 6886 5956 6942 6012
rect 6942 5956 6946 6012
rect 6882 5952 6946 5956
rect 6962 6012 7026 6016
rect 6962 5956 6966 6012
rect 6966 5956 7022 6012
rect 7022 5956 7026 6012
rect 6962 5952 7026 5956
rect 7042 6012 7106 6016
rect 7042 5956 7046 6012
rect 7046 5956 7102 6012
rect 7102 5956 7106 6012
rect 7042 5952 7106 5956
rect 7122 6012 7186 6016
rect 7122 5956 7126 6012
rect 7126 5956 7182 6012
rect 7182 5956 7186 6012
rect 7122 5952 7186 5956
rect 12813 6012 12877 6016
rect 12813 5956 12817 6012
rect 12817 5956 12873 6012
rect 12873 5956 12877 6012
rect 12813 5952 12877 5956
rect 12893 6012 12957 6016
rect 12893 5956 12897 6012
rect 12897 5956 12953 6012
rect 12953 5956 12957 6012
rect 12893 5952 12957 5956
rect 12973 6012 13037 6016
rect 12973 5956 12977 6012
rect 12977 5956 13033 6012
rect 13033 5956 13037 6012
rect 12973 5952 13037 5956
rect 13053 6012 13117 6016
rect 13053 5956 13057 6012
rect 13057 5956 13113 6012
rect 13113 5956 13117 6012
rect 13053 5952 13117 5956
rect 3917 5468 3981 5472
rect 3917 5412 3921 5468
rect 3921 5412 3977 5468
rect 3977 5412 3981 5468
rect 3917 5408 3981 5412
rect 3997 5468 4061 5472
rect 3997 5412 4001 5468
rect 4001 5412 4057 5468
rect 4057 5412 4061 5468
rect 3997 5408 4061 5412
rect 4077 5468 4141 5472
rect 4077 5412 4081 5468
rect 4081 5412 4137 5468
rect 4137 5412 4141 5468
rect 4077 5408 4141 5412
rect 4157 5468 4221 5472
rect 4157 5412 4161 5468
rect 4161 5412 4217 5468
rect 4217 5412 4221 5468
rect 4157 5408 4221 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 15778 5468 15842 5472
rect 15778 5412 15782 5468
rect 15782 5412 15838 5468
rect 15838 5412 15842 5468
rect 15778 5408 15842 5412
rect 15858 5468 15922 5472
rect 15858 5412 15862 5468
rect 15862 5412 15918 5468
rect 15918 5412 15922 5468
rect 15858 5408 15922 5412
rect 15938 5468 16002 5472
rect 15938 5412 15942 5468
rect 15942 5412 15998 5468
rect 15998 5412 16002 5468
rect 15938 5408 16002 5412
rect 16018 5468 16082 5472
rect 16018 5412 16022 5468
rect 16022 5412 16078 5468
rect 16078 5412 16082 5468
rect 16018 5408 16082 5412
rect 6882 4924 6946 4928
rect 6882 4868 6886 4924
rect 6886 4868 6942 4924
rect 6942 4868 6946 4924
rect 6882 4864 6946 4868
rect 6962 4924 7026 4928
rect 6962 4868 6966 4924
rect 6966 4868 7022 4924
rect 7022 4868 7026 4924
rect 6962 4864 7026 4868
rect 7042 4924 7106 4928
rect 7042 4868 7046 4924
rect 7046 4868 7102 4924
rect 7102 4868 7106 4924
rect 7042 4864 7106 4868
rect 7122 4924 7186 4928
rect 7122 4868 7126 4924
rect 7126 4868 7182 4924
rect 7182 4868 7186 4924
rect 7122 4864 7186 4868
rect 12813 4924 12877 4928
rect 12813 4868 12817 4924
rect 12817 4868 12873 4924
rect 12873 4868 12877 4924
rect 12813 4864 12877 4868
rect 12893 4924 12957 4928
rect 12893 4868 12897 4924
rect 12897 4868 12953 4924
rect 12953 4868 12957 4924
rect 12893 4864 12957 4868
rect 12973 4924 13037 4928
rect 12973 4868 12977 4924
rect 12977 4868 13033 4924
rect 13033 4868 13037 4924
rect 12973 4864 13037 4868
rect 13053 4924 13117 4928
rect 13053 4868 13057 4924
rect 13057 4868 13113 4924
rect 13113 4868 13117 4924
rect 13053 4864 13117 4868
rect 3917 4380 3981 4384
rect 3917 4324 3921 4380
rect 3921 4324 3977 4380
rect 3977 4324 3981 4380
rect 3917 4320 3981 4324
rect 3997 4380 4061 4384
rect 3997 4324 4001 4380
rect 4001 4324 4057 4380
rect 4057 4324 4061 4380
rect 3997 4320 4061 4324
rect 4077 4380 4141 4384
rect 4077 4324 4081 4380
rect 4081 4324 4137 4380
rect 4137 4324 4141 4380
rect 4077 4320 4141 4324
rect 4157 4380 4221 4384
rect 4157 4324 4161 4380
rect 4161 4324 4217 4380
rect 4217 4324 4221 4380
rect 4157 4320 4221 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 15778 4380 15842 4384
rect 15778 4324 15782 4380
rect 15782 4324 15838 4380
rect 15838 4324 15842 4380
rect 15778 4320 15842 4324
rect 15858 4380 15922 4384
rect 15858 4324 15862 4380
rect 15862 4324 15918 4380
rect 15918 4324 15922 4380
rect 15858 4320 15922 4324
rect 15938 4380 16002 4384
rect 15938 4324 15942 4380
rect 15942 4324 15998 4380
rect 15998 4324 16002 4380
rect 15938 4320 16002 4324
rect 16018 4380 16082 4384
rect 16018 4324 16022 4380
rect 16022 4324 16078 4380
rect 16078 4324 16082 4380
rect 16018 4320 16082 4324
rect 6882 3836 6946 3840
rect 6882 3780 6886 3836
rect 6886 3780 6942 3836
rect 6942 3780 6946 3836
rect 6882 3776 6946 3780
rect 6962 3836 7026 3840
rect 6962 3780 6966 3836
rect 6966 3780 7022 3836
rect 7022 3780 7026 3836
rect 6962 3776 7026 3780
rect 7042 3836 7106 3840
rect 7042 3780 7046 3836
rect 7046 3780 7102 3836
rect 7102 3780 7106 3836
rect 7042 3776 7106 3780
rect 7122 3836 7186 3840
rect 7122 3780 7126 3836
rect 7126 3780 7182 3836
rect 7182 3780 7186 3836
rect 7122 3776 7186 3780
rect 12813 3836 12877 3840
rect 12813 3780 12817 3836
rect 12817 3780 12873 3836
rect 12873 3780 12877 3836
rect 12813 3776 12877 3780
rect 12893 3836 12957 3840
rect 12893 3780 12897 3836
rect 12897 3780 12953 3836
rect 12953 3780 12957 3836
rect 12893 3776 12957 3780
rect 12973 3836 13037 3840
rect 12973 3780 12977 3836
rect 12977 3780 13033 3836
rect 13033 3780 13037 3836
rect 12973 3776 13037 3780
rect 13053 3836 13117 3840
rect 13053 3780 13057 3836
rect 13057 3780 13113 3836
rect 13113 3780 13117 3836
rect 13053 3776 13117 3780
rect 3917 3292 3981 3296
rect 3917 3236 3921 3292
rect 3921 3236 3977 3292
rect 3977 3236 3981 3292
rect 3917 3232 3981 3236
rect 3997 3292 4061 3296
rect 3997 3236 4001 3292
rect 4001 3236 4057 3292
rect 4057 3236 4061 3292
rect 3997 3232 4061 3236
rect 4077 3292 4141 3296
rect 4077 3236 4081 3292
rect 4081 3236 4137 3292
rect 4137 3236 4141 3292
rect 4077 3232 4141 3236
rect 4157 3292 4221 3296
rect 4157 3236 4161 3292
rect 4161 3236 4217 3292
rect 4217 3236 4221 3292
rect 4157 3232 4221 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 15778 3292 15842 3296
rect 15778 3236 15782 3292
rect 15782 3236 15838 3292
rect 15838 3236 15842 3292
rect 15778 3232 15842 3236
rect 15858 3292 15922 3296
rect 15858 3236 15862 3292
rect 15862 3236 15918 3292
rect 15918 3236 15922 3292
rect 15858 3232 15922 3236
rect 15938 3292 16002 3296
rect 15938 3236 15942 3292
rect 15942 3236 15998 3292
rect 15998 3236 16002 3292
rect 15938 3232 16002 3236
rect 16018 3292 16082 3296
rect 16018 3236 16022 3292
rect 16022 3236 16078 3292
rect 16078 3236 16082 3292
rect 16018 3232 16082 3236
rect 6882 2748 6946 2752
rect 6882 2692 6886 2748
rect 6886 2692 6942 2748
rect 6942 2692 6946 2748
rect 6882 2688 6946 2692
rect 6962 2748 7026 2752
rect 6962 2692 6966 2748
rect 6966 2692 7022 2748
rect 7022 2692 7026 2748
rect 6962 2688 7026 2692
rect 7042 2748 7106 2752
rect 7042 2692 7046 2748
rect 7046 2692 7102 2748
rect 7102 2692 7106 2748
rect 7042 2688 7106 2692
rect 7122 2748 7186 2752
rect 7122 2692 7126 2748
rect 7126 2692 7182 2748
rect 7182 2692 7186 2748
rect 7122 2688 7186 2692
rect 12813 2748 12877 2752
rect 12813 2692 12817 2748
rect 12817 2692 12873 2748
rect 12873 2692 12877 2748
rect 12813 2688 12877 2692
rect 12893 2748 12957 2752
rect 12893 2692 12897 2748
rect 12897 2692 12953 2748
rect 12953 2692 12957 2748
rect 12893 2688 12957 2692
rect 12973 2748 13037 2752
rect 12973 2692 12977 2748
rect 12977 2692 13033 2748
rect 13033 2692 13037 2748
rect 12973 2688 13037 2692
rect 13053 2748 13117 2752
rect 13053 2692 13057 2748
rect 13057 2692 13113 2748
rect 13113 2692 13117 2748
rect 13053 2688 13117 2692
rect 3917 2204 3981 2208
rect 3917 2148 3921 2204
rect 3921 2148 3977 2204
rect 3977 2148 3981 2204
rect 3917 2144 3981 2148
rect 3997 2204 4061 2208
rect 3997 2148 4001 2204
rect 4001 2148 4057 2204
rect 4057 2148 4061 2204
rect 3997 2144 4061 2148
rect 4077 2204 4141 2208
rect 4077 2148 4081 2204
rect 4081 2148 4137 2204
rect 4137 2148 4141 2204
rect 4077 2144 4141 2148
rect 4157 2204 4221 2208
rect 4157 2148 4161 2204
rect 4161 2148 4217 2204
rect 4217 2148 4221 2204
rect 4157 2144 4221 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 15778 2204 15842 2208
rect 15778 2148 15782 2204
rect 15782 2148 15838 2204
rect 15838 2148 15842 2204
rect 15778 2144 15842 2148
rect 15858 2204 15922 2208
rect 15858 2148 15862 2204
rect 15862 2148 15918 2204
rect 15918 2148 15922 2204
rect 15858 2144 15922 2148
rect 15938 2204 16002 2208
rect 15938 2148 15942 2204
rect 15942 2148 15998 2204
rect 15998 2148 16002 2204
rect 15938 2144 16002 2148
rect 16018 2204 16082 2208
rect 16018 2148 16022 2204
rect 16022 2148 16078 2204
rect 16078 2148 16082 2204
rect 16018 2144 16082 2148
<< metal4 >>
rect 3909 14176 4229 14736
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 13088 4229 14112
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 12000 4229 13024
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 10912 4229 11936
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 9824 4229 10848
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 8736 4229 9760
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 7648 4229 8672
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 6560 4229 7584
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 5472 4229 6496
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 4384 4229 5408
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 3296 4229 4320
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 2208 4229 3232
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2128 4229 2144
rect 6874 14720 7195 14736
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7195 14720
rect 6874 13632 7195 14656
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7195 13632
rect 6874 12544 7195 13568
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7195 12544
rect 6874 11456 7195 12480
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7195 11456
rect 6874 10368 7195 11392
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7195 10368
rect 6874 9280 7195 10304
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7195 9280
rect 6874 8192 7195 9216
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7195 8192
rect 6874 7104 7195 8128
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7195 7104
rect 6874 6016 7195 7040
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7195 6016
rect 6874 4928 7195 5952
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7195 4928
rect 6874 3840 7195 4864
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7195 3840
rect 6874 2752 7195 3776
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7195 2752
rect 6874 2128 7195 2688
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12805 14720 13125 14736
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 13632 13125 14656
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 12544 13125 13568
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 11456 13125 12480
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 10368 13125 11392
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 12805 9280 13125 10304
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 8192 13125 9216
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 7104 13125 8128
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 6016 13125 7040
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 4928 13125 5952
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 3840 13125 4864
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 2752 13125 3776
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2128 13125 2688
rect 15770 14176 16091 14736
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16091 14176
rect 15770 13088 16091 14112
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16091 13088
rect 15770 12000 16091 13024
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16091 12000
rect 15770 10912 16091 11936
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16091 10912
rect 15770 9824 16091 10848
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16091 9824
rect 15770 8736 16091 9760
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16091 8736
rect 15770 7648 16091 8672
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16091 7648
rect 15770 6560 16091 7584
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16091 6560
rect 15770 5472 16091 6496
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16091 5472
rect 15770 4384 16091 5408
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16091 4384
rect 15770 3296 16091 4320
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16091 3296
rect 15770 2208 16091 3232
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16091 2208
rect 15770 2128 16091 2144
use sky130_fd_sc_hd__clkbuf_2  output75 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 1748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output65
timestamp 1624635492
transform -1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output86
timestamp 1624635492
transform -1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output70
timestamp 1624635492
transform -1 0 2116 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output88
timestamp 1624635492
transform -1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output71
timestamp 1624635492
transform -1 0 2484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__18__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 2668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output66
timestamp 1624635492
transform -1 0 3036 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _86_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2760 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _18_
timestamp 1624635492
transform 1 0 2484 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3036 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output67
timestamp 1624635492
transform -1 0 3496 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3312 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3036 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output68
timestamp 1624635492
transform -1 0 4232 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3588 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _84_
timestamp 1624635492
transform 1 0 3496 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__84__A
timestamp 1624635492
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output69
timestamp 1624635492
transform -1 0 4600 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 4600 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output72
timestamp 1624635492
transform -1 0 4968 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1624635492
transform 1 0 4600 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 5060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output74
timestamp 1624635492
transform -1 0 5704 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output73
timestamp 1624635492
transform -1 0 5336 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5704 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_58
timestamp 1624635492
transform 1 0 6440 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1624635492
transform -1 0 6164 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output63
timestamp 1624635492
transform -1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_2  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 7452 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1624635492
transform -1 0 6808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1624635492
transform -1 0 6440 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_43 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5060 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output117
timestamp 1624635492
transform -1 0 8004 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output116
timestamp 1624635492
transform -1 0 7636 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output115
timestamp 1624635492
transform -1 0 7268 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_2  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1624635492
transform 1 0 7452 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_1_79
timestamp 1624635492
transform 1 0 8372 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80
timestamp 1624635492
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75
timestamp 1624635492
transform 1 0 8004 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output119
timestamp 1624635492
transform -1 0 9016 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output118
timestamp 1624635492
transform -1 0 8464 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 8464 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1624635492
transform 1 0 8096 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1624635492
transform 1 0 9292 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1624635492
transform -1 0 10304 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 10396 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1624635492
transform 1 0 10396 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 10856 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output121
timestamp 1624635492
transform -1 0 10028 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86
timestamp 1624635492
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_92
timestamp 1624635492
transform 1 0 9568 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1624635492
transform 1 0 11868 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 12512 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1624635492
transform 1 0 11684 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1624635492
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output120
timestamp 1624635492
transform -1 0 11592 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output122
timestamp 1624635492
transform -1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output123
timestamp 1624635492
transform -1 0 11592 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1624635492
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1624635492
transform 1 0 12788 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1624635492
transform 1 0 13064 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 14260 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1624635492
transform 1 0 13064 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1624635492
transform -1 0 14444 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1624635492
transform -1 0 15364 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1624635492
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1624635492
transform 1 0 15180 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1624635492
transform 1 0 15548 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output124
timestamp 1624635492
transform -1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output126
timestamp 1624635492
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1624635492
transform -1 0 15548 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1624635492
transform 1 0 16284 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_151
timestamp 1624635492
transform 1 0 14996 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output129
timestamp 1624635492
transform 1 0 16468 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output125
timestamp 1624635492
transform -1 0 17112 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1624635492
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1624635492
transform -1 0 17112 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output127
timestamp 1624635492
transform -1 0 17480 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1624635492
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1624635492
transform -1 0 17480 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output111
timestamp 1624635492
transform 1 0 17480 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output107
timestamp 1624635492
transform 1 0 17480 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output109
timestamp 1624635492
transform 1 0 17848 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output108
timestamp 1624635492
transform 1 0 18216 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output106
timestamp 1624635492
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output95
timestamp 1624635492
transform 1 0 18216 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1624635492
transform 1 0 2760 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1624635492
transform 1 0 2484 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output87
timestamp 1624635492
transform -1 0 1748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output89
timestamp 1624635492
transform -1 0 2116 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output91
timestamp 1624635492
transform -1 0 2484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 3312 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  output133
timestamp 1624635492
transform -1 0 3588 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__86__A
timestamp 1624635492
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__A
timestamp 1624635492
transform -1 0 4048 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1624635492
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5152 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6624 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1624635492
transform 1 0 8096 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1624635492
transform 1 0 8464 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_79
timestamp 1624635492
transform 1 0 8372 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_83
timestamp 1624635492
transform 1 0 8740 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1624635492
transform 1 0 9844 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1624635492
transform 1 0 10304 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_87 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 9108 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_98
timestamp 1624635492
transform 1 0 10120 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1624635492
transform -1 0 11132 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1624635492
transform 1 0 11132 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1624635492
transform -1 0 13156 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1624635492
transform 1 0 11408 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1624635492
transform -1 0 11960 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1624635492
transform 1 0 13156 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1624635492
transform 1 0 14444 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1624635492
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1624635492
transform 1 0 13432 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1624635492
transform 1 0 13708 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1624635492
transform 1 0 13984 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_144
timestamp 1624635492
transform 1 0 14352 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1624635492
transform -1 0 16468 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1624635492
transform -1 0 15824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1624635492
transform -1 0 16192 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1624635492
transform -1 0 15548 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1624635492
transform -1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1624635492
transform -1 0 14996 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_160
timestamp 1624635492
transform 1 0 15824 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1624635492
transform -1 0 16744 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output110
timestamp 1624635492
transform 1 0 18216 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output112
timestamp 1624635492
transform 1 0 17848 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output128
timestamp 1624635492
transform 1 0 17480 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output130
timestamp 1624635492
transform 1 0 17112 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output132
timestamp 1624635492
transform 1 0 16744 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _21_
timestamp 1624635492
transform 1 0 2484 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _82_
timestamp 1624635492
transform 1 0 2760 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output90
timestamp 1624635492
transform -1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output92
timestamp 1624635492
transform -1 0 2116 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output93
timestamp 1624635492
transform -1 0 2484 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 3864 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1624635492
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__A
timestamp 1624635492
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A
timestamp 1624635492
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_27
timestamp 1624635492
transform 1 0 3588 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1624635492
transform 1 0 6624 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_48
timestamp 1624635492
transform 1 0 5520 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5980 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_58
timestamp 1624635492
transform 1 0 6440 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 7360 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_67
timestamp 1624635492
transform 1 0 7268 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1624635492
transform -1 0 9752 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1624635492
transform 1 0 8832 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 11592 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_94
timestamp 1624635492
transform 1 0 9752 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1624635492
transform 1 0 12236 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1624635492
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1624635492
transform -1 0 11868 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1624635492
transform -1 0 12052 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_119
timestamp 1624635492
transform 1 0 12052 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_2  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1624635492
transform 1 0 14076 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1624635492
transform 1 0 13064 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1624635492
transform -1 0 14076 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1624635492
transform -1 0 13524 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1624635492
transform -1 0 13708 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_137
timestamp 1624635492
transform 1 0 13708 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_2  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1624635492
transform 1 0 14904 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1624635492
transform 1 0 15732 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1624635492
transform -1 0 17480 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1624635492
transform -1 0 17204 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1624635492
transform -1 0 16836 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1624635492
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output113
timestamp 1624635492
transform 1 0 18216 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output114
timestamp 1624635492
transform 1 0 17848 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output131
timestamp 1624635492
transform 1 0 17480 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1624635492
transform 1 0 16468 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1624635492
transform 1 0 2300 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 2300 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output76
timestamp 1624635492
transform -1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_W_FTB01_A
timestamp 1624635492
transform -1 0 2760 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__24__A
timestamp 1624635492
transform -1 0 2944 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__22__A
timestamp 1624635492
transform -1 0 3128 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 4140 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 3956 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3128 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_28
timestamp 1624635492
transform 1 0 3680 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1624635492
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1624635492
transform 1 0 4968 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1624635492
transform 1 0 5796 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_64
timestamp 1624635492
transform 1 0 6992 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_76
timestamp 1624635492
transform 1 0 8096 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 11776 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1624635492
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_87
timestamp 1624635492
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_99
timestamp 1624635492
transform 1 0 10212 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_2  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1624635492
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_116
timestamp 1624635492
transform 1 0 11776 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1624635492
transform 1 0 13064 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1624635492
transform 1 0 13984 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1624635492
transform 1 0 14352 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1624635492
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1624635492
transform 1 0 13892 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1624635492
transform -1 0 16652 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1624635492
transform -1 0 16376 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1624635492
transform -1 0 15364 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1624635492
transform 1 0 15364 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1624635492
transform 1 0 15640 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1624635492
transform -1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1624635492
transform -1 0 17848 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_2_
timestamp 1624635492
transform 1 0 16652 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output96
timestamp 1624635492
transform 1 0 18216 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output97
timestamp 1624635492
transform 1 0 17848 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_178
timestamp 1624635492
transform 1 0 17480 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1624635492
transform 1 0 2116 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp 1624635492
transform 1 0 2392 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1624635492
transform 1 0 2852 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output77
timestamp 1624635492
transform -1 0 1748 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output94
timestamp 1624635492
transform -1 0 2116 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__23__A
timestamp 1624635492
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 6348 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 3680 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_37
timestamp 1624635492
transform 1 0 4508 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 7912 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 8004 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_74
timestamp 1624635492
transform 1 0 7912 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9476 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1624635492
transform 1 0 12604 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1624635492
transform 1 0 10948 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1624635492
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 1624635492
transform 1 0 11500 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_115
timestamp 1624635492
transform 1 0 11684 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1624635492
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1624635492
transform -1 0 14260 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1624635492
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1624635492
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_128
timestamp 1624635492
transform 1 0 12880 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_136
timestamp 1624635492
transform 1 0 13616 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_143
timestamp 1624635492
transform 1 0 14260 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1624635492
transform 1 0 16008 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1624635492
transform -1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1624635492
transform -1 0 15824 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1624635492
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1624635492
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1624635492
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1624635492
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1624635492
transform -1 0 18124 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1624635492
transform 1 0 16928 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1624635492
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output98
timestamp 1624635492
transform 1 0 18216 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_181
timestamp 1624635492
transform 1 0 17756 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_185
timestamp 1624635492
transform 1 0 18124 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output79
timestamp 1624635492
transform -1 0 1748 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output78
timestamp 1624635492
transform -1 0 1748 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2024 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _26_
timestamp 1624635492
transform 1 0 1748 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1624635492
transform 1 0 1748 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_17
timestamp 1624635492
transform 1 0 2668 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__26__A
timestamp 1624635492
transform -1 0 2668 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__25__A
timestamp 1624635492
transform -1 0 2484 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1624635492
transform 1 0 2944 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 3496 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 4968 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1624635492
transform 1 0 3864 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1624635492
transform 1 0 4692 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_42
timestamp 1624635492
transform 1 0 4968 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_48
timestamp 1624635492
transform 1 0 5520 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1624635492
transform 1 0 5428 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_56
timestamp 1624635492
transform 1 0 6256 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1624635492
transform 1 0 6440 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_52
timestamp 1624635492
transform 1 0 5888 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 6256 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1624635492
transform 1 0 6440 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_2  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1624635492
transform -1 0 7452 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1624635492
transform 1 0 8004 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_69
timestamp 1624635492
transform 1 0 7452 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_81
timestamp 1624635492
transform 1 0 8556 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_69
timestamp 1624635492
transform 1 0 7452 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 10672 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__or2b_2  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1624635492
transform 1 0 9108 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 10948 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1624635492
transform 1 0 8924 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_94
timestamp 1624635492
transform 1 0 9752 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_86
timestamp 1624635492
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 11684 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1624635492
transform 1 0 11500 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624635492
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 12604 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_106
timestamp 1624635492
transform 1 0 10856 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_112
timestamp 1624635492
transform 1 0 11408 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_125
timestamp 1624635492
transform 1 0 12604 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_107
timestamp 1624635492
transform 1 0 10948 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 1624635492
transform 1 0 11500 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 13156 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14352 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624635492
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_131
timestamp 1624635492
transform 1 0 13156 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_134
timestamp 1624635492
transform 1 0 13432 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_140
timestamp 1624635492
transform 1 0 13984 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1624635492
transform 1 0 15824 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1624635492
transform 1 0 15548 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1624635492
transform 1 0 14720 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_147
timestamp 1624635492
transform 1 0 14628 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_166
timestamp 1624635492
transform 1 0 16376 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1624635492
transform 1 0 16468 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1624635492
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1624635492
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1624635492
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624635492
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_1_
timestamp 1624635492
transform 1 0 16652 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1624635492
transform -1 0 17572 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_185
timestamp 1624635492
transform 1 0 18124 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_185
timestamp 1624635492
transform 1 0 18124 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_178
timestamp 1624635492
transform 1 0 17480 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output100
timestamp 1624635492
transform 1 0 18216 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output99
timestamp 1624635492
transform 1 0 18216 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1624635492
transform -1 0 17848 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1624635492
transform -1 0 18124 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1624635492
transform -1 0 17848 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1624635492
transform -1 0 18124 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 1624635492
transform 1 0 2116 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _28_
timestamp 1624635492
transform 1 0 2392 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _85_
timestamp 1624635492
transform 1 0 2668 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output80
timestamp 1624635492
transform -1 0 1748 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output81
timestamp 1624635492
transform -1 0 2116 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__A
timestamp 1624635492
transform 1 0 2944 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4324 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__28__A
timestamp 1624635492
transform -1 0 3312 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__A
timestamp 1624635492
transform 1 0 3312 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__85__A
timestamp 1624635492
transform -1 0 3680 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_28
timestamp 1624635492
transform 1 0 3680 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_30
timestamp 1624635492
transform 1 0 3864 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_34
timestamp 1624635492
transform 1 0 4232 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _09_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 6440 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_51
timestamp 1624635492
transform 1 0 5796 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_58
timestamp 1624635492
transform 1 0 6440 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1624635492
transform 1 0 8096 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1624635492
transform 1 0 7268 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_64
timestamp 1624635492
transform 1 0 6992 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _13_
timestamp 1624635492
transform 1 0 9108 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 1624635492
transform 1 0 8924 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_92
timestamp 1624635492
transform 1 0 9568 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_104
timestamp 1624635492
transform 1 0 10672 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1624635492
transform 1 0 12420 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1624635492
transform 1 0 11592 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1624635492
transform -1 0 11592 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 14352 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1624635492
transform 1 0 13248 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1624635492
transform -1 0 14260 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1624635492
transform 1 0 16376 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1624635492
transform 1 0 17204 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output101
timestamp 1624635492
transform 1 0 18216 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1624635492
transform -1 0 18216 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _29_
timestamp 1624635492
transform 1 0 1748 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp 1624635492
transform 1 0 2852 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1624635492
transform -1 0 2852 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output82
timestamp 1624635492
transform -1 0 1748 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _10_
timestamp 1624635492
transform 1 0 3496 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _83_
timestamp 1624635492
transform 1 0 3128 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1624635492
transform 1 0 4232 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1624635492
transform -1 0 3956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__30__A
timestamp 1624635492
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_25
timestamp 1624635492
transform 1 0 3404 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_33
timestamp 1624635492
transform 1 0 4140 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_2_
timestamp 1624635492
transform 1 0 6440 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 5704 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 5244 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_47
timestamp 1624635492
transform 1 0 5428 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_50
timestamp 1624635492
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 8648 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1624635492
transform 1 0 7728 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 7544 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_67
timestamp 1624635492
transform 1 0 7268 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_81
timestamp 1624635492
transform 1 0 8556 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 11592 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1624635492
transform 1 0 12236 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624635492
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 11960 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 12052 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_118
timestamp 1624635492
transform 1 0 11960 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _14_
timestamp 1624635492
transform 1 0 13892 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 14260 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1624635492
transform 1 0 13064 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_142
timestamp 1624635492
transform 1 0 14168 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1624635492
transform 1 0 15824 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_159
timestamp 1624635492
transform 1 0 15732 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _15_
timestamp 1624635492
transform -1 0 17204 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1624635492
transform -1 0 17848 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1624635492
transform -1 0 17572 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624635492
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output102
timestamp 1624635492
transform 1 0 18216 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output103
timestamp 1624635492
transform 1 0 17848 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1624635492
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_175
timestamp 1624635492
transform 1 0 17204 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1624635492
transform 1 0 2944 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1624635492
transform 1 0 2116 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output83
timestamp 1624635492
transform -1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output84
timestamp 1624635492
transform -1 0 2116 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1624635492
transform 1 0 4784 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1624635492
transform 1 0 3864 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_39
timestamp 1624635492
transform 1 0 4692 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 5704 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_1_
timestamp 1624635492
transform 1 0 6532 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_49
timestamp 1624635492
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1624635492
transform 1 0 8188 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1624635492
transform 1 0 7360 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 9108 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 12420 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_10_123
timestamp 1624635492
transform 1 0 12420 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_2_
timestamp 1624635492
transform -1 0 13892 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624635492
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 13892 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1624635492
transform 1 0 14076 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_144
timestamp 1624635492
transform 1 0 14352 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 14904 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 14720 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1624635492
transform 1 0 17940 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1624635492
transform 1 0 17112 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output104
timestamp 1624635492
transform 1 0 18216 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1624635492
transform 1 0 16928 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1624635492
transform 1 0 16744 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 16560 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 2944 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output85
timestamp 1624635492
transform -1 0 3312 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1624635492
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 5060 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_24
timestamp 1624635492
transform 1 0 3312 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 7912 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 6072 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_43
timestamp 1624635492
transform 1 0 5060 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_53
timestamp 1624635492
transform 1 0 5980 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1624635492
transform 1 0 8556 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_74
timestamp 1624635492
transform 1 0 7912 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_77
timestamp 1624635492
transform 1 0 8188 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 10120 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_90
timestamp 1624635492
transform 1 0 9384 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_94
timestamp 1624635492
transform 1 0 9752 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_97
timestamp 1624635492
transform 1 0 10028 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 11684 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624635492
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1624635492
transform 1 0 13156 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_142
timestamp 1624635492
transform 1 0 14168 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14628 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 16284 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_146
timestamp 1624635492
transform 1 0 14536 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1624635492
transform -1 0 18124 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1624635492
transform 1 0 17020 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624635492
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output105
timestamp 1624635492
transform 1 0 18216 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1624635492
transform 1 0 16652 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1624635492
transform -1 0 16652 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_172
timestamp 1624635492
transform 1 0 16928 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_185
timestamp 1624635492
transform 1 0 18124 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 1840 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1624635492
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 3496 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 3864 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_28
timestamp 1624635492
transform 1 0 3680 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1624635492
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1624635492
transform 1 0 5796 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_44
timestamp 1624635492
transform 1 0 5152 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_48
timestamp 1624635492
transform 1 0 5520 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_62
timestamp 1624635492
transform 1 0 6808 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 7268 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_66
timestamp 1624635492
transform 1 0 7176 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1624635492
transform 1 0 8740 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9200 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1624635492
transform 1 0 10028 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_87
timestamp 1624635492
transform 1 0 9108 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1624635492
transform 1 0 11960 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_110
timestamp 1624635492
transform 1 0 11224 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_1_
timestamp 1624635492
transform 1 0 13156 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624635492
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 13064 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_130
timestamp 1624635492
transform 1 0 13064 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_142
timestamp 1624635492
transform 1 0 14168 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_144
timestamp 1624635492
transform 1 0 14352 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1624635492
transform 1 0 16192 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1624635492
transform 1 0 15088 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform -1 0 16192 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 14904 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_161
timestamp 1624635492
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1624635492
transform -1 0 18124 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1624635492
transform 1 0 17020 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1624635492
transform -1 0 18584 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_185
timestamp 1624635492
transform 1 0 18124 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform -1 0 1564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1624635492
transform 1 0 1748 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1624635492
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1624635492
transform -1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 2852 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1624635492
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1624635492
transform 1 0 2852 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1624635492
transform -1 0 2668 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _31_
timestamp 1624635492
transform 1 0 2116 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1624635492
transform 1 0 3864 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__A
timestamp 1624635492
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_1_
timestamp 1624635492
transform 1 0 3680 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1624635492
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 4508 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1624635492
transform 1 0 4416 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1624635492
transform 1 0 6440 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1624635492
transform 1 0 5428 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1624635492
transform 1 0 6072 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1624635492
transform 1 0 5244 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_42
timestamp 1624635492
transform 1 0 4968 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_46
timestamp 1624635492
transform 1 0 5336 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_56
timestamp 1624635492
transform 1 0 6256 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _12_
timestamp 1624635492
transform 1 0 6900 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 7544 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 7452 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_71
timestamp 1624635492
transform 1 0 7636 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_83
timestamp 1624635492
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_66
timestamp 1624635492
transform 1 0 7176 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_69
timestamp 1624635492
transform 1 0 7452 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1624635492
transform 1 0 9108 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1624635492
transform 1 0 10396 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1624635492
transform -1 0 10396 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1624635492
transform 1 0 9936 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_87
timestamp 1624635492
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1624635492
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_111
timestamp 1624635492
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_105
timestamp 1624635492
transform 1 0 10764 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624635492
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1624635492
transform 1 0 11224 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1624635492
transform -1 0 11132 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1624635492
transform 1 0 11684 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 12052 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 12052 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 12420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1624635492
transform 1 0 12420 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1624635492
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 13616 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_144
timestamp 1624635492
transform 1 0 14352 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_142
timestamp 1624635492
transform 1 0 14168 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_138
timestamp 1624635492
transform 1 0 13800 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_136
timestamp 1624635492
transform 1 0 13616 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 13616 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624635492
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 15456 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 15180 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1624635492
transform 1 0 15916 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform -1 0 15916 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_156
timestamp 1624635492
transform 1 0 15456 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1624635492
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1624635492
transform 1 0 16928 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1624635492
transform -1 0 17664 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1624635492
transform 1 0 17664 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624635492
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1624635492
transform -1 0 18584 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1624635492
transform -1 0 18216 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform -1 0 16836 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_170
timestamp 1624635492
transform 1 0 16744 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_181
timestamp 1624635492
transform 1 0 17756 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_189
timestamp 1624635492
transform 1 0 18492 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 4048 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1624635492
transform -1 0 2576 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1624635492
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_34
timestamp 1624635492
transform 1 0 4232 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1624635492
transform 1 0 6440 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1624635492
transform 1 0 5060 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 5888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_42
timestamp 1624635492
transform 1 0 4968 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_55
timestamp 1624635492
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 7360 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_67
timestamp 1624635492
transform 1 0 7268 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 10304 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_102
timestamp 1624635492
transform 1 0 10488 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1624635492
transform 1 0 12604 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1624635492
transform 1 0 11776 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1624635492
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624635492
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_115
timestamp 1624635492
transform 1 0 11684 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 14996 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_134
timestamp 1624635492
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_151
timestamp 1624635492
transform 1 0 14996 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1624635492
transform 1 0 16100 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1624635492
transform 1 0 16928 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624635492
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1624635492
transform -1 0 18584 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1624635492
transform -1 0 18216 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 16836 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_181
timestamp 1624635492
transform 1 0 17756 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_2_
timestamp 1624635492
transform 1 0 2668 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1624635492
transform 1 0 1840 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1624635492
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1624635492
transform 1 0 1748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform -1 0 3680 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 4784 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 3864 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_28
timestamp 1624635492
transform 1 0 3680 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_34
timestamp 1624635492
transform 1 0 4232 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 8280 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1624635492
transform 1 0 5796 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1624635492
transform -1 0 5796 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_78
timestamp 1624635492
transform 1 0 8280 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 11868 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624635492
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_87
timestamp 1624635492
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_99
timestamp 1624635492
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 13892 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 11868 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_119
timestamp 1624635492
transform 1 0 12052 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624635492
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_139
timestamp 1624635492
transform 1 0 13892 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_144
timestamp 1624635492
transform 1 0 14352 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_156
timestamp 1624635492
transform 1 0 15456 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1624635492
transform -1 0 17664 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1624635492
transform -1 0 18124 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1624635492
transform -1 0 18584 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 17848 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform -1 0 17388 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1624635492
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 16836 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_168
timestamp 1624635492
transform 1 0 16560 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_185
timestamp 1624635492
transform 1 0 18124 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 2760 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1624635492
transform 1 0 1840 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1624635492
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1624635492
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_17
timestamp 1624635492
transform 1 0 2668 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 4232 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 6440 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624635492
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1624635492
transform 1 0 5888 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_56
timestamp 1624635492
transform 1 0 6256 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1624635492
transform -1 0 9200 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_88
timestamp 1624635492
transform 1 0 9200 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_100
timestamp 1624635492
transform 1 0 10304 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624635492
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_112
timestamp 1624635492
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_115
timestamp 1624635492
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_127
timestamp 1624635492
transform 1 0 12788 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_139
timestamp 1624635492
transform 1 0 13892 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_151
timestamp 1624635492
transform 1 0 14996 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_163
timestamp 1624635492
transform 1 0 16100 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1624635492
transform -1 0 18124 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624635492
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1624635492
transform -1 0 18584 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 17848 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_172
timestamp 1624635492
transform 1 0 16928 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_185
timestamp 1624635492
transform 1 0 18124 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1624635492
transform 1 0 2208 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1624635492
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1624635492
transform 1 0 1748 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_11
timestamp 1624635492
transform 1 0 2116 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _11_
timestamp 1624635492
transform 1 0 3036 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4508 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624635492
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 3496 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 3680 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 3864 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_28
timestamp 1624635492
transform 1 0 3680 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_34
timestamp 1624635492
transform 1 0 4232 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1624635492
transform 1 0 5980 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1624635492
transform 1 0 7084 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_77
timestamp 1624635492
transform 1 0 8188 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624635492
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1624635492
transform 1 0 8924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_87
timestamp 1624635492
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_99
timestamp 1624635492
transform 1 0 10212 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_111
timestamp 1624635492
transform 1 0 11316 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_123
timestamp 1624635492
transform 1 0 12420 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624635492
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_135
timestamp 1624635492
transform 1 0 13524 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_144
timestamp 1624635492
transform 1 0 14352 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_156
timestamp 1624635492
transform 1 0 15456 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1624635492
transform -1 0 18584 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1624635492
transform -1 0 18216 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1624635492
transform -1 0 17848 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624635492
transform -1 0 17664 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_168
timestamp 1624635492
transform 1 0 16560 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_176
timestamp 1624635492
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1624635492
transform 1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1624635492
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1624635492
transform 1 0 1748 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1624635492
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1624635492
transform 1 0 2668 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1624635492
transform -1 0 2668 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1624635492
transform 1 0 2116 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _77_
timestamp 1624635492
transform -1 0 2392 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 3128 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 3128 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform -1 0 3312 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 3312 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 3496 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 3680 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 3680 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624635492
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_28
timestamp 1624635492
transform 1 0 3680 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1624635492
transform 1 0 3864 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1624635492
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1624635492
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_36
timestamp 1624635492
transform 1 0 4416 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_30
timestamp 1624635492
transform 1 0 3864 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624635492
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_42
timestamp 1624635492
transform 1 0 4968 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_54
timestamp 1624635492
transform 1 0 6072 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_58
timestamp 1624635492
transform 1 0 6440 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_48
timestamp 1624635492
transform 1 0 5520 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_60
timestamp 1624635492
transform 1 0 6624 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_70
timestamp 1624635492
transform 1 0 7544 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_82
timestamp 1624635492
transform 1 0 8648 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_72
timestamp 1624635492
transform 1 0 7728 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624635492
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_94
timestamp 1624635492
transform 1 0 9752 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1624635492
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_87
timestamp 1624635492
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_99
timestamp 1624635492
transform 1 0 10212 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624635492
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_106
timestamp 1624635492
transform 1 0 10856 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_115
timestamp 1624635492
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_111
timestamp 1624635492
transform 1 0 11316 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1624635492
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_127
timestamp 1624635492
transform 1 0 12788 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_139
timestamp 1624635492
transform 1 0 13892 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_135
timestamp 1624635492
transform 1 0 13524 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1624635492
transform 1 0 14352 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_151
timestamp 1624635492
transform 1 0 14996 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_163
timestamp 1624635492
transform 1 0 16100 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_156
timestamp 1624635492
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_168
timestamp 1624635492
transform 1 0 16560 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output150_A
timestamp 1624635492
transform 1 0 16744 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624635492
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_172
timestamp 1624635492
transform 1 0 16928 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output146_A
timestamp 1624635492
transform 1 0 16928 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1624635492
transform -1 0 17480 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624635492
transform -1 0 17296 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 17480 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform -1 0 17664 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 17664 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 17848 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 17848 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output150
timestamp 1624635492
transform 1 0 17848 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1624635492
transform -1 0 18216 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1624635492
transform -1 0 18584 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1624635492
transform -1 0 18584 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1624635492
transform -1 0 2024 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1624635492
transform 1 0 2576 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output145
timestamp 1624635492
transform -1 0 1748 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output149
timestamp 1624635492
transform -1 0 2576 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output151
timestamp 1624635492
transform -1 0 3220 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform -1 0 2208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _78_
timestamp 1624635492
transform 1 0 3220 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _79_
timestamp 1624635492
transform 1 0 3496 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1624635492
transform 1 0 3772 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform -1 0 4232 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1624635492
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1624635492
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_40
timestamp 1624635492
transform 1 0 4784 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _80_
timestamp 1624635492
transform 1 0 5980 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _81_
timestamp 1624635492
transform -1 0 6716 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624635492
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_52
timestamp 1624635492
transform 1 0 5888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_56
timestamp 1624635492
transform 1 0 6256 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_61
timestamp 1624635492
transform 1 0 6716 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_73
timestamp 1624635492
transform 1 0 7820 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_85
timestamp 1624635492
transform 1 0 8924 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_97
timestamp 1624635492
transform 1 0 10028 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624635492
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_109
timestamp 1624635492
transform 1 0 11132 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1624635492
transform 1 0 11500 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_115
timestamp 1624635492
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _71_
timestamp 1624635492
transform -1 0 13708 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _72_
timestamp 1624635492
transform -1 0 14628 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1624635492
transform -1 0 13892 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output142_A
timestamp 1624635492
transform -1 0 14076 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output144_A
timestamp 1624635492
transform 1 0 13156 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_127
timestamp 1624635492
transform 1 0 12788 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_133
timestamp 1624635492
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_141
timestamp 1624635492
transform 1 0 14076 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _73_
timestamp 1624635492
transform -1 0 15364 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _74_
timestamp 1624635492
transform -1 0 15824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output148_A
timestamp 1624635492
transform -1 0 16468 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_147
timestamp 1624635492
transform 1 0 14628 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_151
timestamp 1624635492
transform 1 0 14996 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_155
timestamp 1624635492
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_160
timestamp 1624635492
transform 1 0 15824 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_164
timestamp 1624635492
transform 1 0 16192 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624635492
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1624635492
transform -1 0 18584 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1624635492
transform -1 0 18216 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output146
timestamp 1624635492
transform 1 0 17480 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output148
timestamp 1624635492
transform 1 0 17112 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 17112 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 16836 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 16652 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1624635492
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1624635492
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1624635492
transform 1 0 2116 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1624635492
transform 1 0 2484 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1624635492
transform -1 0 3220 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624635492
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output135
timestamp 1624635492
transform -1 0 4232 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output137
timestamp 1624635492
transform -1 0 4600 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output139
timestamp 1624635492
transform -1 0 5152 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output143
timestamp 1624635492
transform -1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform -1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624635492
transform -1 0 4784 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624635492
transform 1 0 6440 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1624635492
transform 1 0 6164 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output64
timestamp 1624635492
transform -1 0 7084 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output141
timestamp 1624635492
transform -1 0 5796 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output147
timestamp 1624635492
transform -1 0 6164 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 6716 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_44
timestamp 1624635492
transform 1 0 5152 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1624635492
transform -1 0 7728 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1624635492
transform -1 0 8924 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 7912 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_65
timestamp 1624635492
transform 1 0 7084 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_74
timestamp 1624635492
transform 1 0 7912 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1624635492
transform -1 0 9108 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624635492
transform 1 0 9108 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_88
timestamp 1624635492
transform 1 0 9200 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1624635492
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_94
timestamp 1624635492
transform 1 0 9752 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1624635492
transform -1 0 9752 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1624635492
transform 1 0 9936 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_101
timestamp 1624635492
transform 1 0 10396 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1624635492
transform -1 0 10396 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1624635492
transform 1 0 10580 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_108
timestamp 1624635492
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1624635492
transform -1 0 11040 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1624635492
transform 1 0 11224 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_115
timestamp 1624635492
transform 1 0 11684 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1624635492
transform -1 0 11684 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1624635492
transform -1 0 12144 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624635492
transform 1 0 11776 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_122
timestamp 1624635492
transform 1 0 12328 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1624635492
transform -1 0 12328 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1624635492
transform 1 0 12512 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624635492
transform 1 0 14444 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1624635492
transform 1 0 13064 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output140
timestamp 1624635492
transform 1 0 14076 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output142
timestamp 1624635492
transform 1 0 13708 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output144
timestamp 1624635492
transform 1 0 13340 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1624635492
transform -1 0 12972 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_129
timestamp 1624635492
transform 1 0 12972 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1624635492
transform -1 0 16744 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1624635492
transform 1 0 15456 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output134
timestamp 1624635492
transform -1 0 14904 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output136
timestamp 1624635492
transform -1 0 15456 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output138
timestamp 1624635492
transform -1 0 16100 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 16376 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1624635492
transform -1 0 15088 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_163
timestamp 1624635492
transform 1 0 16100 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624635492
transform 1 0 17112 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1624635492
transform -1 0 18584 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1624635492
transform -1 0 18216 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1624635492
transform -1 0 17848 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1624635492
transform -1 0 17112 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1624635492
transform -1 0 17480 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
<< labels >>
rlabel metal2 s 7378 16400 7434 17200 6 IO_ISOL_N
port 0 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 SC_IN_BOT
port 1 nsew signal input
rlabel metal2 s 6090 16400 6146 17200 6 SC_IN_TOP
port 2 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 SC_OUT_BOT
port 3 nsew signal tristate
rlabel metal2 s 6734 16400 6790 17200 6 SC_OUT_TOP
port 4 nsew signal tristate
rlabel metal2 s 202 0 258 800 6 bottom_grid_pin_0_
port 5 nsew signal tristate
rlabel metal2 s 2686 0 2742 800 6 bottom_grid_pin_10_
port 6 nsew signal tristate
rlabel metal2 s 3146 0 3202 800 6 bottom_grid_pin_12_
port 7 nsew signal tristate
rlabel metal2 s 3606 0 3662 800 6 bottom_grid_pin_14_
port 8 nsew signal tristate
rlabel metal2 s 4158 0 4214 800 6 bottom_grid_pin_16_
port 9 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 bottom_grid_pin_2_
port 10 nsew signal tristate
rlabel metal2 s 1122 0 1178 800 6 bottom_grid_pin_4_
port 11 nsew signal tristate
rlabel metal2 s 1674 0 1730 800 6 bottom_grid_pin_6_
port 12 nsew signal tristate
rlabel metal2 s 2134 0 2190 800 6 bottom_grid_pin_8_
port 13 nsew signal tristate
rlabel metal2 s 4618 0 4674 800 6 ccff_head
port 14 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 ccff_tail
port 15 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 chanx_left_in[0]
port 16 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 chanx_left_in[10]
port 17 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 chanx_left_in[11]
port 18 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 chanx_left_in[12]
port 19 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 chanx_left_in[13]
port 20 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 chanx_left_in[14]
port 21 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 chanx_left_in[15]
port 22 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 chanx_left_in[16]
port 23 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 chanx_left_in[17]
port 24 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 chanx_left_in[18]
port 25 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 chanx_left_in[19]
port 26 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 chanx_left_in[1]
port 27 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[2]
port 28 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 chanx_left_in[3]
port 29 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 chanx_left_in[4]
port 30 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[5]
port 31 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[6]
port 32 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[7]
port 33 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[8]
port 34 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[9]
port 35 nsew signal input
rlabel metal3 s 0 552 800 672 6 chanx_left_out[0]
port 36 nsew signal tristate
rlabel metal3 s 0 4632 800 4752 6 chanx_left_out[10]
port 37 nsew signal tristate
rlabel metal3 s 0 5040 800 5160 6 chanx_left_out[11]
port 38 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 chanx_left_out[12]
port 39 nsew signal tristate
rlabel metal3 s 0 5992 800 6112 6 chanx_left_out[13]
port 40 nsew signal tristate
rlabel metal3 s 0 6400 800 6520 6 chanx_left_out[14]
port 41 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 chanx_left_out[15]
port 42 nsew signal tristate
rlabel metal3 s 0 7216 800 7336 6 chanx_left_out[16]
port 43 nsew signal tristate
rlabel metal3 s 0 7624 800 7744 6 chanx_left_out[17]
port 44 nsew signal tristate
rlabel metal3 s 0 8032 800 8152 6 chanx_left_out[18]
port 45 nsew signal tristate
rlabel metal3 s 0 8440 800 8560 6 chanx_left_out[19]
port 46 nsew signal tristate
rlabel metal3 s 0 960 800 1080 6 chanx_left_out[1]
port 47 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 chanx_left_out[2]
port 48 nsew signal tristate
rlabel metal3 s 0 1776 800 1896 6 chanx_left_out[3]
port 49 nsew signal tristate
rlabel metal3 s 0 2184 800 2304 6 chanx_left_out[4]
port 50 nsew signal tristate
rlabel metal3 s 0 2592 800 2712 6 chanx_left_out[5]
port 51 nsew signal tristate
rlabel metal3 s 0 3000 800 3120 6 chanx_left_out[6]
port 52 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 chanx_left_out[7]
port 53 nsew signal tristate
rlabel metal3 s 0 3816 800 3936 6 chanx_left_out[8]
port 54 nsew signal tristate
rlabel metal3 s 0 4224 800 4344 6 chanx_left_out[9]
port 55 nsew signal tristate
rlabel metal3 s 19200 8712 20000 8832 6 chanx_right_in[0]
port 56 nsew signal input
rlabel metal3 s 19200 12928 20000 13048 6 chanx_right_in[10]
port 57 nsew signal input
rlabel metal3 s 19200 13336 20000 13456 6 chanx_right_in[11]
port 58 nsew signal input
rlabel metal3 s 19200 13744 20000 13864 6 chanx_right_in[12]
port 59 nsew signal input
rlabel metal3 s 19200 14152 20000 14272 6 chanx_right_in[13]
port 60 nsew signal input
rlabel metal3 s 19200 14696 20000 14816 6 chanx_right_in[14]
port 61 nsew signal input
rlabel metal3 s 19200 15104 20000 15224 6 chanx_right_in[15]
port 62 nsew signal input
rlabel metal3 s 19200 15512 20000 15632 6 chanx_right_in[16]
port 63 nsew signal input
rlabel metal3 s 19200 15920 20000 16040 6 chanx_right_in[17]
port 64 nsew signal input
rlabel metal3 s 19200 16328 20000 16448 6 chanx_right_in[18]
port 65 nsew signal input
rlabel metal3 s 19200 16736 20000 16856 6 chanx_right_in[19]
port 66 nsew signal input
rlabel metal3 s 19200 9120 20000 9240 6 chanx_right_in[1]
port 67 nsew signal input
rlabel metal3 s 19200 9528 20000 9648 6 chanx_right_in[2]
port 68 nsew signal input
rlabel metal3 s 19200 9936 20000 10056 6 chanx_right_in[3]
port 69 nsew signal input
rlabel metal3 s 19200 10344 20000 10464 6 chanx_right_in[4]
port 70 nsew signal input
rlabel metal3 s 19200 10752 20000 10872 6 chanx_right_in[5]
port 71 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 chanx_right_in[6]
port 72 nsew signal input
rlabel metal3 s 19200 11704 20000 11824 6 chanx_right_in[7]
port 73 nsew signal input
rlabel metal3 s 19200 12112 20000 12232 6 chanx_right_in[8]
port 74 nsew signal input
rlabel metal3 s 19200 12520 20000 12640 6 chanx_right_in[9]
port 75 nsew signal input
rlabel metal3 s 19200 144 20000 264 6 chanx_right_out[0]
port 76 nsew signal tristate
rlabel metal3 s 19200 4360 20000 4480 6 chanx_right_out[10]
port 77 nsew signal tristate
rlabel metal3 s 19200 4768 20000 4888 6 chanx_right_out[11]
port 78 nsew signal tristate
rlabel metal3 s 19200 5176 20000 5296 6 chanx_right_out[12]
port 79 nsew signal tristate
rlabel metal3 s 19200 5584 20000 5704 6 chanx_right_out[13]
port 80 nsew signal tristate
rlabel metal3 s 19200 6128 20000 6248 6 chanx_right_out[14]
port 81 nsew signal tristate
rlabel metal3 s 19200 6536 20000 6656 6 chanx_right_out[15]
port 82 nsew signal tristate
rlabel metal3 s 19200 6944 20000 7064 6 chanx_right_out[16]
port 83 nsew signal tristate
rlabel metal3 s 19200 7352 20000 7472 6 chanx_right_out[17]
port 84 nsew signal tristate
rlabel metal3 s 19200 7760 20000 7880 6 chanx_right_out[18]
port 85 nsew signal tristate
rlabel metal3 s 19200 8168 20000 8288 6 chanx_right_out[19]
port 86 nsew signal tristate
rlabel metal3 s 19200 552 20000 672 6 chanx_right_out[1]
port 87 nsew signal tristate
rlabel metal3 s 19200 960 20000 1080 6 chanx_right_out[2]
port 88 nsew signal tristate
rlabel metal3 s 19200 1368 20000 1488 6 chanx_right_out[3]
port 89 nsew signal tristate
rlabel metal3 s 19200 1776 20000 1896 6 chanx_right_out[4]
port 90 nsew signal tristate
rlabel metal3 s 19200 2184 20000 2304 6 chanx_right_out[5]
port 91 nsew signal tristate
rlabel metal3 s 19200 2592 20000 2712 6 chanx_right_out[6]
port 92 nsew signal tristate
rlabel metal3 s 19200 3136 20000 3256 6 chanx_right_out[7]
port 93 nsew signal tristate
rlabel metal3 s 19200 3544 20000 3664 6 chanx_right_out[8]
port 94 nsew signal tristate
rlabel metal3 s 19200 3952 20000 4072 6 chanx_right_out[9]
port 95 nsew signal tristate
rlabel metal2 s 6642 0 6698 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
port 96 nsew signal tristate
rlabel metal2 s 7102 0 7158 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
port 97 nsew signal tristate
rlabel metal2 s 7654 0 7710 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
port 98 nsew signal tristate
rlabel metal2 s 8114 0 8170 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
port 99 nsew signal tristate
rlabel metal2 s 8666 0 8722 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
port 100 nsew signal tristate
rlabel metal2 s 9126 0 9182 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
port 101 nsew signal tristate
rlabel metal2 s 9678 0 9734 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
port 102 nsew signal tristate
rlabel metal2 s 10138 0 10194 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
port 103 nsew signal tristate
rlabel metal2 s 10598 0 10654 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
port 104 nsew signal tristate
rlabel metal2 s 11150 0 11206 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
port 105 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
port 106 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
port 107 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
port 108 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
port 109 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
port 110 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
port 111 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
port 112 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
port 113 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
port 114 nsew signal tristate
rlabel metal2 s 16118 0 16174 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
port 115 nsew signal tristate
rlabel metal2 s 16670 0 16726 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
port 116 nsew signal tristate
rlabel metal2 s 17130 0 17186 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
port 117 nsew signal tristate
rlabel metal2 s 17590 0 17646 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
port 118 nsew signal tristate
rlabel metal2 s 18142 0 18198 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
port 119 nsew signal tristate
rlabel metal2 s 18602 0 18658 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
port 120 nsew signal tristate
rlabel metal2 s 19154 0 19210 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
port 121 nsew signal tristate
rlabel metal2 s 19614 0 19670 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
port 122 nsew signal tristate
rlabel metal2 s 8022 16400 8078 17200 6 prog_clk_0_N_in
port 123 nsew signal input
rlabel metal3 s 0 144 800 264 6 prog_clk_0_W_out
port 124 nsew signal tristate
rlabel metal2 s 8666 16400 8722 17200 6 top_width_0_height_0__pin_0_
port 125 nsew signal input
rlabel metal2 s 11886 16400 11942 17200 6 top_width_0_height_0__pin_10_
port 126 nsew signal input
rlabel metal2 s 14462 16400 14518 17200 6 top_width_0_height_0__pin_11_lower
port 127 nsew signal tristate
rlabel metal2 s 3514 16400 3570 17200 6 top_width_0_height_0__pin_11_upper
port 128 nsew signal tristate
rlabel metal2 s 12530 16400 12586 17200 6 top_width_0_height_0__pin_12_
port 129 nsew signal input
rlabel metal2 s 15106 16400 15162 17200 6 top_width_0_height_0__pin_13_lower
port 130 nsew signal tristate
rlabel metal2 s 4158 16400 4214 17200 6 top_width_0_height_0__pin_13_upper
port 131 nsew signal tristate
rlabel metal2 s 13174 16400 13230 17200 6 top_width_0_height_0__pin_14_
port 132 nsew signal input
rlabel metal2 s 15750 16400 15806 17200 6 top_width_0_height_0__pin_15_lower
port 133 nsew signal tristate
rlabel metal2 s 4802 16400 4858 17200 6 top_width_0_height_0__pin_15_upper
port 134 nsew signal tristate
rlabel metal2 s 13818 16400 13874 17200 6 top_width_0_height_0__pin_16_
port 135 nsew signal input
rlabel metal2 s 16394 16400 16450 17200 6 top_width_0_height_0__pin_17_lower
port 136 nsew signal tristate
rlabel metal2 s 5446 16400 5502 17200 6 top_width_0_height_0__pin_17_upper
port 137 nsew signal tristate
rlabel metal2 s 17038 16400 17094 17200 6 top_width_0_height_0__pin_1_lower
port 138 nsew signal tristate
rlabel metal2 s 294 16400 350 17200 6 top_width_0_height_0__pin_1_upper
port 139 nsew signal tristate
rlabel metal2 s 9310 16400 9366 17200 6 top_width_0_height_0__pin_2_
port 140 nsew signal input
rlabel metal2 s 17682 16400 17738 17200 6 top_width_0_height_0__pin_3_lower
port 141 nsew signal tristate
rlabel metal2 s 938 16400 994 17200 6 top_width_0_height_0__pin_3_upper
port 142 nsew signal tristate
rlabel metal2 s 9954 16400 10010 17200 6 top_width_0_height_0__pin_4_
port 143 nsew signal input
rlabel metal2 s 18326 16400 18382 17200 6 top_width_0_height_0__pin_5_lower
port 144 nsew signal tristate
rlabel metal2 s 1582 16400 1638 17200 6 top_width_0_height_0__pin_5_upper
port 145 nsew signal tristate
rlabel metal2 s 10598 16400 10654 17200 6 top_width_0_height_0__pin_6_
port 146 nsew signal input
rlabel metal2 s 18970 16400 19026 17200 6 top_width_0_height_0__pin_7_lower
port 147 nsew signal tristate
rlabel metal2 s 2226 16400 2282 17200 6 top_width_0_height_0__pin_7_upper
port 148 nsew signal tristate
rlabel metal2 s 11242 16400 11298 17200 6 top_width_0_height_0__pin_8_
port 149 nsew signal input
rlabel metal2 s 19614 16400 19670 17200 6 top_width_0_height_0__pin_9_lower
port 150 nsew signal tristate
rlabel metal2 s 2870 16400 2926 17200 6 top_width_0_height_0__pin_9_upper
port 151 nsew signal tristate
rlabel metal4 s 15771 2128 16091 14736 6 VPWR
port 152 nsew power bidirectional
rlabel metal4 s 9840 2128 10160 14736 6 VPWR
port 153 nsew power bidirectional
rlabel metal4 s 3909 2128 4229 14736 6 VPWR
port 154 nsew power bidirectional
rlabel metal4 s 12805 2128 13125 14736 6 VGND
port 155 nsew ground bidirectional
rlabel metal4 s 6875 2128 7195 14736 6 VGND
port 156 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 17200
<< end >>
