magic
tech sky130A
magscale 1 2
timestamp 1656241038
<< viali >>
rect 1593 17289 1627 17323
rect 1961 17289 1995 17323
rect 2329 17289 2363 17323
rect 2697 17289 2731 17323
rect 3065 17289 3099 17323
rect 3433 17289 3467 17323
rect 4169 17289 4203 17323
rect 4537 17289 4571 17323
rect 4905 17289 4939 17323
rect 5273 17289 5307 17323
rect 5641 17289 5675 17323
rect 6009 17289 6043 17323
rect 6561 17289 6595 17323
rect 6929 17289 6963 17323
rect 7297 17289 7331 17323
rect 7665 17289 7699 17323
rect 8033 17289 8067 17323
rect 8401 17289 8435 17323
rect 9045 17289 9079 17323
rect 13461 17289 13495 17323
rect 14381 17289 14415 17323
rect 15577 17289 15611 17323
rect 8769 17221 8803 17255
rect 11253 17221 11287 17255
rect 13737 17221 13771 17255
rect 15209 17221 15243 17255
rect 1777 17153 1811 17187
rect 2145 17153 2179 17187
rect 2513 17153 2547 17187
rect 2881 17153 2915 17187
rect 3249 17153 3283 17187
rect 3617 17153 3651 17187
rect 4353 17153 4387 17187
rect 4721 17153 4755 17187
rect 5089 17153 5123 17187
rect 5457 17153 5491 17187
rect 5825 17153 5859 17187
rect 6193 17153 6227 17187
rect 6745 17153 6779 17187
rect 7113 17153 7147 17187
rect 7481 17153 7515 17187
rect 7849 17153 7883 17187
rect 8217 17153 8251 17187
rect 8585 17153 8619 17187
rect 9229 17153 9263 17187
rect 9597 17153 9631 17187
rect 9965 17153 9999 17187
rect 10333 17153 10367 17187
rect 10701 17153 10735 17187
rect 11069 17153 11103 17187
rect 11713 17153 11747 17187
rect 11989 17153 12023 17187
rect 12265 17153 12299 17187
rect 12541 17153 12575 17187
rect 12909 17153 12943 17187
rect 13277 17153 13311 17187
rect 13645 17153 13679 17187
rect 14289 17153 14323 17187
rect 14565 17153 14599 17187
rect 14841 17153 14875 17187
rect 15117 17153 15151 17187
rect 15393 17153 15427 17187
rect 9781 17017 9815 17051
rect 10885 17017 10919 17051
rect 11529 17017 11563 17051
rect 12081 17017 12115 17051
rect 13093 17017 13127 17051
rect 14933 17017 14967 17051
rect 9413 16949 9447 16983
rect 10149 16949 10183 16983
rect 10517 16949 10551 16983
rect 11805 16949 11839 16983
rect 12357 16949 12391 16983
rect 12725 16949 12759 16983
rect 14105 16949 14139 16983
rect 14657 16949 14691 16983
rect 9689 16745 9723 16779
rect 10057 16745 10091 16779
rect 10793 16745 10827 16779
rect 11345 16745 11379 16779
rect 11621 16745 11655 16779
rect 11897 16745 11931 16779
rect 12173 16745 12207 16779
rect 12633 16745 12667 16779
rect 13369 16745 13403 16779
rect 14105 16745 14139 16779
rect 14381 16745 14415 16779
rect 14841 16745 14875 16779
rect 14657 16677 14691 16711
rect 9321 16609 9355 16643
rect 15577 16609 15611 16643
rect 1409 16541 1443 16575
rect 1685 16541 1719 16575
rect 1961 16541 1995 16575
rect 4169 16541 4203 16575
rect 9229 16541 9263 16575
rect 15209 16541 15243 16575
rect 15485 16541 15519 16575
rect 1593 16405 1627 16439
rect 1869 16405 1903 16439
rect 3985 16405 4019 16439
rect 9045 16405 9079 16439
rect 15025 16405 15059 16439
rect 15301 16405 15335 16439
rect 1409 16201 1443 16235
rect 15393 16065 15427 16099
rect 15669 16065 15703 16099
rect 15485 15861 15519 15895
rect 5089 13889 5123 13923
rect 4629 13821 4663 13855
rect 4997 13685 5031 13719
rect 4077 12937 4111 12971
rect 5825 12937 5859 12971
rect 14473 12937 14507 12971
rect 4598 12869 4632 12903
rect 4261 12801 4295 12835
rect 6009 12801 6043 12835
rect 14289 12801 14323 12835
rect 15393 12801 15427 12835
rect 4353 12733 4387 12767
rect 5733 12665 5767 12699
rect 14105 12597 14139 12631
rect 15577 12597 15611 12631
rect 5089 12393 5123 12427
rect 7389 12393 7423 12427
rect 9321 12393 9355 12427
rect 5273 12189 5307 12223
rect 7573 12189 7607 12223
rect 9505 12189 9539 12223
rect 7205 11849 7239 11883
rect 7849 11849 7883 11883
rect 1409 11713 1443 11747
rect 1685 11713 1719 11747
rect 7389 11713 7423 11747
rect 7757 11713 7791 11747
rect 8033 11713 8067 11747
rect 8217 11645 8251 11679
rect 7573 11577 7607 11611
rect 1593 11509 1627 11543
rect 8769 11509 8803 11543
rect 8953 11305 8987 11339
rect 8217 11237 8251 11271
rect 6837 11169 6871 11203
rect 9505 11169 9539 11203
rect 8493 11101 8527 11135
rect 8769 11101 8803 11135
rect 9321 11101 9355 11135
rect 7082 11033 7116 11067
rect 9413 11033 9447 11067
rect 8309 10965 8343 10999
rect 5733 10761 5767 10795
rect 6009 10761 6043 10795
rect 7757 10761 7791 10795
rect 9229 10761 9263 10795
rect 9597 10761 9631 10795
rect 8870 10693 8904 10727
rect 3500 10625 3534 10659
rect 5917 10625 5951 10659
rect 6193 10625 6227 10659
rect 6561 10625 6595 10659
rect 6837 10625 6871 10659
rect 7297 10625 7331 10659
rect 9413 10625 9447 10659
rect 9781 10625 9815 10659
rect 10057 10625 10091 10659
rect 7021 10557 7055 10591
rect 7205 10557 7239 10591
rect 9137 10557 9171 10591
rect 6377 10489 6411 10523
rect 3571 10421 3605 10455
rect 6653 10421 6687 10455
rect 7665 10421 7699 10455
rect 9873 10421 9907 10455
rect 11253 10217 11287 10251
rect 12081 10217 12115 10251
rect 12633 10217 12667 10251
rect 13185 10217 13219 10251
rect 5089 10149 5123 10183
rect 10701 10149 10735 10183
rect 12357 10149 12391 10183
rect 5733 10081 5767 10115
rect 6101 10081 6135 10115
rect 8125 10081 8159 10115
rect 8309 10081 8343 10115
rect 9597 10081 9631 10115
rect 10333 10081 10367 10115
rect 10425 10081 10459 10115
rect 4997 10013 5031 10047
rect 5917 10013 5951 10047
rect 7757 10013 7791 10047
rect 10885 10013 10919 10047
rect 11161 10013 11195 10047
rect 11437 10013 11471 10047
rect 11713 10013 11747 10047
rect 11989 10013 12023 10047
rect 12265 10013 12299 10047
rect 12541 10013 12575 10047
rect 12817 10013 12851 10047
rect 13093 10013 13127 10047
rect 13369 10013 13403 10047
rect 5457 9945 5491 9979
rect 9505 9945 9539 9979
rect 4813 9877 4847 9911
rect 5549 9877 5583 9911
rect 8401 9877 8435 9911
rect 8769 9877 8803 9911
rect 9045 9877 9079 9911
rect 9413 9877 9447 9911
rect 9873 9877 9907 9911
rect 10241 9877 10275 9911
rect 10977 9877 11011 9911
rect 11529 9877 11563 9911
rect 11805 9877 11839 9911
rect 12909 9877 12943 9911
rect 6377 9673 6411 9707
rect 8585 9673 8619 9707
rect 10793 9673 10827 9707
rect 1409 9605 1443 9639
rect 3065 9605 3099 9639
rect 6837 9605 6871 9639
rect 5365 9537 5399 9571
rect 5917 9537 5951 9571
rect 6193 9537 6227 9571
rect 6745 9537 6779 9571
rect 7461 9537 7495 9571
rect 9045 9537 9079 9571
rect 9781 9537 9815 9571
rect 10241 9537 10275 9571
rect 10977 9537 11011 9571
rect 3249 9469 3283 9503
rect 6929 9469 6963 9503
rect 7205 9469 7239 9503
rect 8769 9469 8803 9503
rect 8953 9469 8987 9503
rect 5181 9401 5215 9435
rect 9413 9401 9447 9435
rect 10057 9401 10091 9435
rect 5733 9333 5767 9367
rect 6009 9333 6043 9367
rect 9597 9333 9631 9367
rect 6929 9129 6963 9163
rect 8401 9061 8435 9095
rect 8309 8925 8343 8959
rect 8585 8925 8619 8959
rect 9137 8925 9171 8959
rect 8064 8857 8098 8891
rect 8953 8789 8987 8823
rect 7113 8585 7147 8619
rect 7481 8585 7515 8619
rect 8033 8585 8067 8619
rect 8493 8585 8527 8619
rect 11713 8517 11747 8551
rect 1685 8449 1719 8483
rect 8401 8449 8435 8483
rect 12541 8449 12575 8483
rect 7573 8381 7607 8415
rect 7665 8381 7699 8415
rect 8677 8381 8711 8415
rect 1501 8313 1535 8347
rect 12725 8313 12759 8347
rect 5641 7497 5675 7531
rect 3249 7361 3283 7395
rect 4721 7361 4755 7395
rect 5273 7361 5307 7395
rect 5825 7361 5859 7395
rect 7573 7361 7607 7395
rect 9413 7361 9447 7395
rect 7389 7225 7423 7259
rect 3065 7157 3099 7191
rect 4537 7157 4571 7191
rect 5089 7157 5123 7191
rect 9229 7157 9263 7191
rect 1685 5185 1719 5219
rect 1501 5049 1535 5083
rect 2053 3145 2087 3179
rect 15485 3145 15519 3179
rect 1777 3009 1811 3043
rect 1869 3009 1903 3043
rect 2145 3009 2179 3043
rect 4353 3009 4387 3043
rect 15393 3009 15427 3043
rect 15669 3009 15703 3043
rect 1593 2805 1627 2839
rect 4169 2805 4203 2839
rect 8861 2805 8895 2839
rect 9137 2805 9171 2839
rect 9505 2805 9539 2839
rect 9873 2805 9907 2839
rect 10241 2805 10275 2839
rect 10609 2805 10643 2839
rect 10977 2805 11011 2839
rect 11529 2805 11563 2839
rect 11805 2805 11839 2839
rect 12081 2805 12115 2839
rect 12449 2805 12483 2839
rect 12817 2805 12851 2839
rect 13185 2805 13219 2839
rect 13553 2805 13587 2839
rect 13921 2805 13955 2839
rect 14289 2805 14323 2839
rect 14657 2805 14691 2839
rect 15025 2805 15059 2839
rect 15209 2805 15243 2839
rect 8953 2601 8987 2635
rect 9597 2601 9631 2635
rect 9965 2601 9999 2635
rect 10333 2601 10367 2635
rect 11805 2601 11839 2635
rect 12541 2601 12575 2635
rect 12909 2601 12943 2635
rect 15485 2601 15519 2635
rect 13645 2533 13679 2567
rect 14381 2533 14415 2567
rect 1777 2397 1811 2431
rect 2145 2397 2179 2431
rect 2513 2397 2547 2431
rect 2881 2397 2915 2431
rect 3249 2397 3283 2431
rect 3617 2397 3651 2431
rect 4353 2397 4387 2431
rect 4721 2397 4755 2431
rect 5089 2397 5123 2431
rect 5457 2397 5491 2431
rect 5825 2397 5859 2431
rect 6193 2397 6227 2431
rect 6929 2397 6963 2431
rect 7297 2397 7331 2431
rect 7665 2397 7699 2431
rect 8033 2397 8067 2431
rect 8401 2397 8435 2431
rect 8769 2397 8803 2431
rect 9137 2397 9171 2431
rect 9413 2397 9447 2431
rect 9781 2397 9815 2431
rect 10149 2397 10183 2431
rect 10517 2397 10551 2431
rect 10885 2397 10919 2431
rect 11253 2397 11287 2431
rect 11713 2397 11747 2431
rect 11989 2397 12023 2431
rect 12357 2397 12391 2431
rect 12725 2397 12759 2431
rect 13093 2397 13127 2431
rect 13461 2397 13495 2431
rect 13829 2397 13863 2431
rect 14289 2397 14323 2431
rect 14565 2397 14599 2431
rect 14933 2397 14967 2431
rect 15301 2397 15335 2431
rect 15669 2397 15703 2431
rect 1593 2261 1627 2295
rect 1961 2261 1995 2295
rect 2329 2261 2363 2295
rect 2697 2261 2731 2295
rect 3065 2261 3099 2295
rect 3433 2261 3467 2295
rect 4169 2261 4203 2295
rect 4537 2261 4571 2295
rect 4905 2261 4939 2295
rect 5273 2261 5307 2295
rect 5641 2261 5675 2295
rect 6009 2261 6043 2295
rect 6745 2261 6779 2295
rect 7113 2261 7147 2295
rect 7481 2261 7515 2295
rect 7849 2261 7883 2295
rect 8217 2261 8251 2295
rect 8585 2261 8619 2295
rect 9229 2261 9263 2295
rect 10701 2261 10735 2295
rect 11069 2261 11103 2295
rect 11529 2261 11563 2295
rect 12173 2261 12207 2295
rect 13277 2261 13311 2295
rect 14105 2261 14139 2295
rect 14749 2261 14783 2295
rect 15117 2261 15151 2295
<< metal1 >>
rect 9214 17688 9220 17740
rect 9272 17728 9278 17740
rect 13170 17728 13176 17740
rect 9272 17700 13176 17728
rect 9272 17688 9278 17700
rect 13170 17688 13176 17700
rect 13228 17688 13234 17740
rect 9122 17620 9128 17672
rect 9180 17660 9186 17672
rect 12526 17660 12532 17672
rect 9180 17632 12532 17660
rect 9180 17620 9186 17632
rect 12526 17620 12532 17632
rect 12584 17620 12590 17672
rect 9490 17552 9496 17604
rect 9548 17592 9554 17604
rect 12710 17592 12716 17604
rect 9548 17564 12716 17592
rect 9548 17552 9554 17564
rect 12710 17552 12716 17564
rect 12768 17552 12774 17604
rect 11330 17484 11336 17536
rect 11388 17524 11394 17536
rect 14366 17524 14372 17536
rect 11388 17496 14372 17524
rect 11388 17484 11394 17496
rect 14366 17484 14372 17496
rect 14424 17484 14430 17536
rect 1104 17434 16008 17456
rect 1104 17382 4698 17434
rect 4750 17382 4762 17434
rect 4814 17382 4826 17434
rect 4878 17382 4890 17434
rect 4942 17382 4954 17434
rect 5006 17382 8446 17434
rect 8498 17382 8510 17434
rect 8562 17382 8574 17434
rect 8626 17382 8638 17434
rect 8690 17382 8702 17434
rect 8754 17382 12194 17434
rect 12246 17382 12258 17434
rect 12310 17382 12322 17434
rect 12374 17382 12386 17434
rect 12438 17382 12450 17434
rect 12502 17382 16008 17434
rect 1104 17360 16008 17382
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 1946 17320 1952 17332
rect 1907 17292 1952 17320
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 2314 17320 2320 17332
rect 2275 17292 2320 17320
rect 2314 17280 2320 17292
rect 2372 17280 2378 17332
rect 2682 17320 2688 17332
rect 2643 17292 2688 17320
rect 2682 17280 2688 17292
rect 2740 17280 2746 17332
rect 3050 17320 3056 17332
rect 3011 17292 3056 17320
rect 3050 17280 3056 17292
rect 3108 17280 3114 17332
rect 3418 17320 3424 17332
rect 3379 17292 3424 17320
rect 3418 17280 3424 17292
rect 3476 17280 3482 17332
rect 4154 17320 4160 17332
rect 4115 17292 4160 17320
rect 4154 17280 4160 17292
rect 4212 17280 4218 17332
rect 4522 17320 4528 17332
rect 4483 17292 4528 17320
rect 4522 17280 4528 17292
rect 4580 17280 4586 17332
rect 4893 17323 4951 17329
rect 4893 17289 4905 17323
rect 4939 17320 4951 17323
rect 5074 17320 5080 17332
rect 4939 17292 5080 17320
rect 4939 17289 4951 17292
rect 4893 17283 4951 17289
rect 5074 17280 5080 17292
rect 5132 17280 5138 17332
rect 5258 17320 5264 17332
rect 5219 17292 5264 17320
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 5626 17320 5632 17332
rect 5587 17292 5632 17320
rect 5626 17280 5632 17292
rect 5684 17280 5690 17332
rect 5994 17320 6000 17332
rect 5955 17292 6000 17320
rect 5994 17280 6000 17292
rect 6052 17280 6058 17332
rect 6362 17280 6368 17332
rect 6420 17320 6426 17332
rect 6549 17323 6607 17329
rect 6549 17320 6561 17323
rect 6420 17292 6561 17320
rect 6420 17280 6426 17292
rect 6549 17289 6561 17292
rect 6595 17289 6607 17323
rect 6549 17283 6607 17289
rect 6914 17280 6920 17332
rect 6972 17320 6978 17332
rect 6972 17292 7017 17320
rect 6972 17280 6978 17292
rect 7098 17280 7104 17332
rect 7156 17320 7162 17332
rect 7285 17323 7343 17329
rect 7285 17320 7297 17323
rect 7156 17292 7297 17320
rect 7156 17280 7162 17292
rect 7285 17289 7297 17292
rect 7331 17289 7343 17323
rect 7285 17283 7343 17289
rect 7466 17280 7472 17332
rect 7524 17320 7530 17332
rect 7653 17323 7711 17329
rect 7653 17320 7665 17323
rect 7524 17292 7665 17320
rect 7524 17280 7530 17292
rect 7653 17289 7665 17292
rect 7699 17289 7711 17323
rect 7653 17283 7711 17289
rect 7834 17280 7840 17332
rect 7892 17320 7898 17332
rect 8021 17323 8079 17329
rect 8021 17320 8033 17323
rect 7892 17292 8033 17320
rect 7892 17280 7898 17292
rect 8021 17289 8033 17292
rect 8067 17289 8079 17323
rect 8021 17283 8079 17289
rect 8294 17280 8300 17332
rect 8352 17320 8358 17332
rect 8389 17323 8447 17329
rect 8389 17320 8401 17323
rect 8352 17292 8401 17320
rect 8352 17280 8358 17292
rect 8389 17289 8401 17292
rect 8435 17289 8447 17323
rect 8389 17283 8447 17289
rect 8846 17280 8852 17332
rect 8904 17320 8910 17332
rect 9033 17323 9091 17329
rect 9033 17320 9045 17323
rect 8904 17292 9045 17320
rect 8904 17280 8910 17292
rect 9033 17289 9045 17292
rect 9079 17289 9091 17323
rect 9033 17283 9091 17289
rect 9582 17280 9588 17332
rect 9640 17320 9646 17332
rect 13446 17320 13452 17332
rect 9640 17292 12388 17320
rect 13407 17292 13452 17320
rect 9640 17280 9646 17292
rect 4614 17252 4620 17264
rect 2884 17224 4620 17252
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17153 1823 17187
rect 2130 17184 2136 17196
rect 2091 17156 2136 17184
rect 1765 17147 1823 17153
rect 1780 17116 1808 17147
rect 2130 17144 2136 17156
rect 2188 17144 2194 17196
rect 2498 17184 2504 17196
rect 2459 17156 2504 17184
rect 2498 17144 2504 17156
rect 2556 17144 2562 17196
rect 2884 17193 2912 17224
rect 4614 17212 4620 17224
rect 4672 17212 4678 17264
rect 8757 17255 8815 17261
rect 4724 17224 5764 17252
rect 2869 17187 2927 17193
rect 2869 17153 2881 17187
rect 2915 17153 2927 17187
rect 2869 17147 2927 17153
rect 3237 17187 3295 17193
rect 3237 17153 3249 17187
rect 3283 17153 3295 17187
rect 3602 17184 3608 17196
rect 3563 17156 3608 17184
rect 3237 17147 3295 17153
rect 3142 17116 3148 17128
rect 1780 17088 3148 17116
rect 3142 17076 3148 17088
rect 3200 17076 3206 17128
rect 3252 17116 3280 17147
rect 3602 17144 3608 17156
rect 3660 17144 3666 17196
rect 4338 17184 4344 17196
rect 4299 17156 4344 17184
rect 4338 17144 4344 17156
rect 4396 17144 4402 17196
rect 4724 17193 4752 17224
rect 4709 17187 4767 17193
rect 4709 17153 4721 17187
rect 4755 17153 4767 17187
rect 4709 17147 4767 17153
rect 5077 17187 5135 17193
rect 5077 17153 5089 17187
rect 5123 17153 5135 17187
rect 5442 17184 5448 17196
rect 5403 17156 5448 17184
rect 5077 17147 5135 17153
rect 3252 17088 4292 17116
rect 4264 17048 4292 17088
rect 4430 17076 4436 17128
rect 4488 17116 4494 17128
rect 5092 17116 5120 17147
rect 5442 17144 5448 17156
rect 5500 17144 5506 17196
rect 4488 17088 5120 17116
rect 5736 17116 5764 17224
rect 5828 17224 8708 17252
rect 5828 17193 5856 17224
rect 5813 17187 5871 17193
rect 5813 17153 5825 17187
rect 5859 17153 5871 17187
rect 6178 17184 6184 17196
rect 6139 17156 6184 17184
rect 5813 17147 5871 17153
rect 6178 17144 6184 17156
rect 6236 17144 6242 17196
rect 6270 17144 6276 17196
rect 6328 17184 6334 17196
rect 6733 17187 6791 17193
rect 6733 17184 6745 17187
rect 6328 17156 6745 17184
rect 6328 17144 6334 17156
rect 6733 17153 6745 17156
rect 6779 17153 6791 17187
rect 6733 17147 6791 17153
rect 7101 17187 7159 17193
rect 7101 17153 7113 17187
rect 7147 17153 7159 17187
rect 7466 17184 7472 17196
rect 7427 17156 7472 17184
rect 7101 17147 7159 17153
rect 6454 17116 6460 17128
rect 5736 17088 6460 17116
rect 4488 17076 4494 17088
rect 6454 17076 6460 17088
rect 6512 17076 6518 17128
rect 5718 17048 5724 17060
rect 4264 17020 5724 17048
rect 5718 17008 5724 17020
rect 5776 17008 5782 17060
rect 7116 17048 7144 17147
rect 7466 17144 7472 17156
rect 7524 17144 7530 17196
rect 7837 17187 7895 17193
rect 7837 17153 7849 17187
rect 7883 17153 7895 17187
rect 8202 17184 8208 17196
rect 8163 17156 8208 17184
rect 7837 17147 7895 17153
rect 7852 17116 7880 17147
rect 8202 17144 8208 17156
rect 8260 17144 8266 17196
rect 8573 17187 8631 17193
rect 8573 17153 8585 17187
rect 8619 17153 8631 17187
rect 8680 17184 8708 17224
rect 8757 17221 8769 17255
rect 8803 17252 8815 17255
rect 11241 17255 11299 17261
rect 11241 17252 11253 17255
rect 8803 17224 9352 17252
rect 8803 17221 8815 17224
rect 8757 17215 8815 17221
rect 9324 17196 9352 17224
rect 10704 17224 11253 17252
rect 8846 17184 8852 17196
rect 8680 17156 8852 17184
rect 8573 17147 8631 17153
rect 8294 17116 8300 17128
rect 7852 17088 8300 17116
rect 8294 17076 8300 17088
rect 8352 17076 8358 17128
rect 8588 17116 8616 17147
rect 8846 17144 8852 17156
rect 8904 17144 8910 17196
rect 9214 17184 9220 17196
rect 9175 17156 9220 17184
rect 9214 17144 9220 17156
rect 9272 17144 9278 17196
rect 9306 17144 9312 17196
rect 9364 17184 9370 17196
rect 9585 17187 9643 17193
rect 9585 17184 9597 17187
rect 9364 17156 9597 17184
rect 9364 17144 9370 17156
rect 9585 17153 9597 17156
rect 9631 17153 9643 17187
rect 9585 17147 9643 17153
rect 9674 17144 9680 17196
rect 9732 17184 9738 17196
rect 9953 17187 10011 17193
rect 9953 17184 9965 17187
rect 9732 17156 9965 17184
rect 9732 17144 9738 17156
rect 9953 17153 9965 17156
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 10042 17144 10048 17196
rect 10100 17184 10106 17196
rect 10321 17187 10379 17193
rect 10321 17184 10333 17187
rect 10100 17156 10333 17184
rect 10100 17144 10106 17156
rect 10321 17153 10333 17156
rect 10367 17153 10379 17187
rect 10321 17147 10379 17153
rect 10410 17144 10416 17196
rect 10468 17184 10474 17196
rect 10704 17193 10732 17224
rect 11241 17221 11253 17224
rect 11287 17221 11299 17255
rect 11241 17215 11299 17221
rect 11514 17212 11520 17264
rect 11572 17252 11578 17264
rect 11572 17224 12020 17252
rect 11572 17212 11578 17224
rect 10689 17187 10747 17193
rect 10689 17184 10701 17187
rect 10468 17156 10701 17184
rect 10468 17144 10474 17156
rect 10689 17153 10701 17156
rect 10735 17153 10747 17187
rect 10689 17147 10747 17153
rect 10778 17144 10784 17196
rect 10836 17184 10842 17196
rect 11057 17187 11115 17193
rect 11057 17184 11069 17187
rect 10836 17156 11069 17184
rect 10836 17144 10842 17156
rect 11057 17153 11069 17156
rect 11103 17153 11115 17187
rect 11057 17147 11115 17153
rect 11146 17144 11152 17196
rect 11204 17184 11210 17196
rect 11992 17193 12020 17224
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 11204 17156 11713 17184
rect 11204 17144 11210 17156
rect 11701 17153 11713 17156
rect 11747 17153 11759 17187
rect 11701 17147 11759 17153
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17153 12035 17187
rect 11977 17147 12035 17153
rect 12253 17187 12311 17193
rect 12253 17153 12265 17187
rect 12299 17153 12311 17187
rect 12253 17147 12311 17153
rect 9122 17116 9128 17128
rect 8588 17088 9128 17116
rect 9122 17076 9128 17088
rect 9180 17076 9186 17128
rect 11422 17116 11428 17128
rect 9232 17088 11428 17116
rect 9232 17048 9260 17088
rect 11422 17076 11428 17088
rect 11480 17076 11486 17128
rect 11882 17076 11888 17128
rect 11940 17116 11946 17128
rect 12268 17116 12296 17147
rect 11940 17088 12296 17116
rect 12360 17116 12388 17292
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 14366 17320 14372 17332
rect 14327 17292 14372 17320
rect 14366 17280 14372 17292
rect 14424 17280 14430 17332
rect 15562 17320 15568 17332
rect 15523 17292 15568 17320
rect 15562 17280 15568 17292
rect 15620 17280 15626 17332
rect 13725 17255 13783 17261
rect 13725 17252 13737 17255
rect 13280 17224 13737 17252
rect 12434 17144 12440 17196
rect 12492 17184 12498 17196
rect 12529 17187 12587 17193
rect 12529 17184 12541 17187
rect 12492 17156 12541 17184
rect 12492 17144 12498 17156
rect 12529 17153 12541 17156
rect 12575 17153 12587 17187
rect 12529 17147 12587 17153
rect 12618 17144 12624 17196
rect 12676 17184 12682 17196
rect 12897 17187 12955 17193
rect 12897 17184 12909 17187
rect 12676 17156 12909 17184
rect 12676 17144 12682 17156
rect 12897 17153 12909 17156
rect 12943 17153 12955 17187
rect 12897 17147 12955 17153
rect 12986 17144 12992 17196
rect 13044 17184 13050 17196
rect 13280 17193 13308 17224
rect 13725 17221 13737 17224
rect 13771 17221 13783 17255
rect 13725 17215 13783 17221
rect 14090 17212 14096 17264
rect 14148 17252 14154 17264
rect 14458 17252 14464 17264
rect 14148 17224 14464 17252
rect 14148 17212 14154 17224
rect 14458 17212 14464 17224
rect 14516 17252 14522 17264
rect 15197 17255 15255 17261
rect 15197 17252 15209 17255
rect 14516 17224 14596 17252
rect 14516 17212 14522 17224
rect 13265 17187 13323 17193
rect 13265 17184 13277 17187
rect 13044 17156 13277 17184
rect 13044 17144 13050 17156
rect 13265 17153 13277 17156
rect 13311 17153 13323 17187
rect 13265 17147 13323 17153
rect 13354 17144 13360 17196
rect 13412 17184 13418 17196
rect 13633 17187 13691 17193
rect 13633 17184 13645 17187
rect 13412 17156 13645 17184
rect 13412 17144 13418 17156
rect 13633 17153 13645 17156
rect 13679 17153 13691 17187
rect 13633 17147 13691 17153
rect 13814 17144 13820 17196
rect 13872 17184 13878 17196
rect 14568 17193 14596 17224
rect 14844 17224 15209 17252
rect 14277 17187 14335 17193
rect 14277 17184 14289 17187
rect 13872 17156 14289 17184
rect 13872 17144 13878 17156
rect 14277 17153 14289 17156
rect 14323 17153 14335 17187
rect 14277 17147 14335 17153
rect 14553 17187 14611 17193
rect 14553 17153 14565 17187
rect 14599 17153 14611 17187
rect 14553 17147 14611 17153
rect 14642 17144 14648 17196
rect 14700 17184 14706 17196
rect 14844 17193 14872 17224
rect 15197 17221 15209 17224
rect 15243 17221 15255 17255
rect 15197 17215 15255 17221
rect 14829 17187 14887 17193
rect 14829 17184 14841 17187
rect 14700 17156 14841 17184
rect 14700 17144 14706 17156
rect 14829 17153 14841 17156
rect 14875 17153 14887 17187
rect 14829 17147 14887 17153
rect 14918 17144 14924 17196
rect 14976 17184 14982 17196
rect 15105 17187 15163 17193
rect 15105 17184 15117 17187
rect 14976 17156 15117 17184
rect 14976 17144 14982 17156
rect 15105 17153 15117 17156
rect 15151 17153 15163 17187
rect 15105 17147 15163 17153
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17153 15439 17187
rect 15381 17147 15439 17153
rect 12360 17088 13216 17116
rect 11940 17076 11946 17088
rect 7116 17020 9260 17048
rect 9306 17008 9312 17060
rect 9364 17048 9370 17060
rect 9769 17051 9827 17057
rect 9769 17048 9781 17051
rect 9364 17020 9781 17048
rect 9364 17008 9370 17020
rect 9769 17017 9781 17020
rect 9815 17017 9827 17051
rect 9769 17011 9827 17017
rect 9950 17008 9956 17060
rect 10008 17048 10014 17060
rect 10873 17051 10931 17057
rect 10873 17048 10885 17051
rect 10008 17020 10885 17048
rect 10008 17008 10014 17020
rect 10873 17017 10885 17020
rect 10919 17017 10931 17051
rect 10873 17011 10931 17017
rect 11054 17008 11060 17060
rect 11112 17048 11118 17060
rect 11517 17051 11575 17057
rect 11517 17048 11529 17051
rect 11112 17020 11529 17048
rect 11112 17008 11118 17020
rect 11517 17017 11529 17020
rect 11563 17017 11575 17051
rect 12069 17051 12127 17057
rect 12069 17048 12081 17051
rect 11517 17011 11575 17017
rect 11624 17020 12081 17048
rect 4338 16940 4344 16992
rect 4396 16980 4402 16992
rect 6362 16980 6368 16992
rect 4396 16952 6368 16980
rect 4396 16940 4402 16952
rect 6362 16940 6368 16952
rect 6420 16940 6426 16992
rect 9398 16980 9404 16992
rect 9359 16952 9404 16980
rect 9398 16940 9404 16952
rect 9456 16940 9462 16992
rect 10134 16980 10140 16992
rect 10095 16952 10140 16980
rect 10134 16940 10140 16952
rect 10192 16940 10198 16992
rect 10505 16983 10563 16989
rect 10505 16949 10517 16983
rect 10551 16980 10563 16983
rect 10686 16980 10692 16992
rect 10551 16952 10692 16980
rect 10551 16949 10563 16952
rect 10505 16943 10563 16949
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 10962 16940 10968 16992
rect 11020 16980 11026 16992
rect 11624 16980 11652 17020
rect 12069 17017 12081 17020
rect 12115 17017 12127 17051
rect 12069 17011 12127 17017
rect 12250 17008 12256 17060
rect 12308 17048 12314 17060
rect 13081 17051 13139 17057
rect 13081 17048 13093 17051
rect 12308 17020 13093 17048
rect 12308 17008 12314 17020
rect 13081 17017 13093 17020
rect 13127 17017 13139 17051
rect 13188 17048 13216 17088
rect 14734 17076 14740 17128
rect 14792 17116 14798 17128
rect 15396 17116 15424 17147
rect 14792 17088 15424 17116
rect 14792 17076 14798 17088
rect 14921 17051 14979 17057
rect 14921 17048 14933 17051
rect 13188 17020 14933 17048
rect 13081 17011 13139 17017
rect 14921 17017 14933 17020
rect 14967 17017 14979 17051
rect 14921 17011 14979 17017
rect 11790 16980 11796 16992
rect 11020 16952 11652 16980
rect 11751 16952 11796 16980
rect 11020 16940 11026 16952
rect 11790 16940 11796 16952
rect 11848 16940 11854 16992
rect 11974 16940 11980 16992
rect 12032 16980 12038 16992
rect 12345 16983 12403 16989
rect 12345 16980 12357 16983
rect 12032 16952 12357 16980
rect 12032 16940 12038 16952
rect 12345 16949 12357 16952
rect 12391 16949 12403 16983
rect 12710 16980 12716 16992
rect 12671 16952 12716 16980
rect 12345 16943 12403 16949
rect 12710 16940 12716 16952
rect 12768 16940 12774 16992
rect 12802 16940 12808 16992
rect 12860 16980 12866 16992
rect 14093 16983 14151 16989
rect 14093 16980 14105 16983
rect 12860 16952 14105 16980
rect 12860 16940 12866 16952
rect 14093 16949 14105 16952
rect 14139 16949 14151 16983
rect 14642 16980 14648 16992
rect 14603 16952 14648 16980
rect 14093 16943 14151 16949
rect 14642 16940 14648 16952
rect 14700 16940 14706 16992
rect 1104 16890 16008 16912
rect 1104 16838 2824 16890
rect 2876 16838 2888 16890
rect 2940 16838 2952 16890
rect 3004 16838 3016 16890
rect 3068 16838 3080 16890
rect 3132 16838 6572 16890
rect 6624 16838 6636 16890
rect 6688 16838 6700 16890
rect 6752 16838 6764 16890
rect 6816 16838 6828 16890
rect 6880 16838 10320 16890
rect 10372 16838 10384 16890
rect 10436 16838 10448 16890
rect 10500 16838 10512 16890
rect 10564 16838 10576 16890
rect 10628 16838 14068 16890
rect 14120 16838 14132 16890
rect 14184 16838 14196 16890
rect 14248 16838 14260 16890
rect 14312 16838 14324 16890
rect 14376 16838 16008 16890
rect 1104 16816 16008 16838
rect 5258 16736 5264 16788
rect 5316 16776 5322 16788
rect 9398 16776 9404 16788
rect 5316 16748 9404 16776
rect 5316 16736 5322 16748
rect 9398 16736 9404 16748
rect 9456 16736 9462 16788
rect 9674 16776 9680 16788
rect 9635 16748 9680 16776
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 10042 16776 10048 16788
rect 10003 16748 10048 16776
rect 10042 16736 10048 16748
rect 10100 16736 10106 16788
rect 10778 16776 10784 16788
rect 10739 16748 10784 16776
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 11146 16736 11152 16788
rect 11204 16776 11210 16788
rect 11333 16779 11391 16785
rect 11333 16776 11345 16779
rect 11204 16748 11345 16776
rect 11204 16736 11210 16748
rect 11333 16745 11345 16748
rect 11379 16745 11391 16779
rect 11333 16739 11391 16745
rect 11514 16736 11520 16788
rect 11572 16776 11578 16788
rect 11609 16779 11667 16785
rect 11609 16776 11621 16779
rect 11572 16748 11621 16776
rect 11572 16736 11578 16748
rect 11609 16745 11621 16748
rect 11655 16745 11667 16779
rect 11882 16776 11888 16788
rect 11843 16748 11888 16776
rect 11609 16739 11667 16745
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 12066 16736 12072 16788
rect 12124 16776 12130 16788
rect 12161 16779 12219 16785
rect 12161 16776 12173 16779
rect 12124 16748 12173 16776
rect 12124 16736 12130 16748
rect 12161 16745 12173 16748
rect 12207 16776 12219 16779
rect 12434 16776 12440 16788
rect 12207 16748 12440 16776
rect 12207 16745 12219 16748
rect 12161 16739 12219 16745
rect 12434 16736 12440 16748
rect 12492 16736 12498 16788
rect 12618 16776 12624 16788
rect 12579 16748 12624 16776
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 13354 16776 13360 16788
rect 13315 16748 13360 16776
rect 13354 16736 13360 16748
rect 13412 16736 13418 16788
rect 13814 16736 13820 16788
rect 13872 16776 13878 16788
rect 14093 16779 14151 16785
rect 14093 16776 14105 16779
rect 13872 16748 14105 16776
rect 13872 16736 13878 16748
rect 14093 16745 14105 16748
rect 14139 16745 14151 16779
rect 14093 16739 14151 16745
rect 14369 16779 14427 16785
rect 14369 16745 14381 16779
rect 14415 16776 14427 16779
rect 14458 16776 14464 16788
rect 14415 16748 14464 16776
rect 14415 16745 14427 16748
rect 14369 16739 14427 16745
rect 14458 16736 14464 16748
rect 14516 16736 14522 16788
rect 14826 16776 14832 16788
rect 14787 16748 14832 16776
rect 14826 16736 14832 16748
rect 14884 16736 14890 16788
rect 4614 16668 4620 16720
rect 4672 16708 4678 16720
rect 5534 16708 5540 16720
rect 4672 16680 5540 16708
rect 4672 16668 4678 16680
rect 5534 16668 5540 16680
rect 5592 16668 5598 16720
rect 11238 16668 11244 16720
rect 11296 16708 11302 16720
rect 12250 16708 12256 16720
rect 11296 16680 12256 16708
rect 11296 16668 11302 16680
rect 12250 16668 12256 16680
rect 12308 16668 12314 16720
rect 12342 16668 12348 16720
rect 12400 16708 12406 16720
rect 13446 16708 13452 16720
rect 12400 16680 13452 16708
rect 12400 16668 12406 16680
rect 13446 16668 13452 16680
rect 13504 16668 13510 16720
rect 14645 16711 14703 16717
rect 14645 16677 14657 16711
rect 14691 16708 14703 16711
rect 14691 16680 15240 16708
rect 14691 16677 14703 16680
rect 14645 16671 14703 16677
rect 8938 16600 8944 16652
rect 8996 16640 9002 16652
rect 9309 16643 9367 16649
rect 9309 16640 9321 16643
rect 8996 16612 9321 16640
rect 8996 16600 9002 16612
rect 1302 16532 1308 16584
rect 1360 16572 1366 16584
rect 1397 16575 1455 16581
rect 1397 16572 1409 16575
rect 1360 16544 1409 16572
rect 1360 16532 1366 16544
rect 1397 16541 1409 16544
rect 1443 16541 1455 16575
rect 1670 16572 1676 16584
rect 1583 16544 1676 16572
rect 1397 16535 1455 16541
rect 1670 16532 1676 16544
rect 1728 16572 1734 16584
rect 1949 16575 2007 16581
rect 1949 16572 1961 16575
rect 1728 16544 1961 16572
rect 1728 16532 1734 16544
rect 1949 16541 1961 16544
rect 1995 16541 2007 16575
rect 4062 16572 4068 16584
rect 1949 16535 2007 16541
rect 3252 16544 4068 16572
rect 1578 16436 1584 16448
rect 1539 16408 1584 16436
rect 1578 16396 1584 16408
rect 1636 16396 1642 16448
rect 1857 16439 1915 16445
rect 1857 16405 1869 16439
rect 1903 16436 1915 16439
rect 3252 16436 3280 16544
rect 4062 16532 4068 16544
rect 4120 16532 4126 16584
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16572 4215 16575
rect 7190 16572 7196 16584
rect 4203 16544 7196 16572
rect 4203 16541 4215 16544
rect 4157 16535 4215 16541
rect 7190 16532 7196 16544
rect 7248 16532 7254 16584
rect 9232 16581 9260 16612
rect 9309 16609 9321 16612
rect 9355 16609 9367 16643
rect 9309 16603 9367 16609
rect 9398 16600 9404 16652
rect 9456 16640 9462 16652
rect 9582 16640 9588 16652
rect 9456 16612 9588 16640
rect 9456 16600 9462 16612
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 10778 16600 10784 16652
rect 10836 16640 10842 16652
rect 11974 16640 11980 16652
rect 10836 16612 11980 16640
rect 10836 16600 10842 16612
rect 11974 16600 11980 16612
rect 12032 16600 12038 16652
rect 15212 16581 15240 16680
rect 15286 16600 15292 16652
rect 15344 16640 15350 16652
rect 15565 16643 15623 16649
rect 15565 16640 15577 16643
rect 15344 16612 15577 16640
rect 15344 16600 15350 16612
rect 9217 16575 9275 16581
rect 9217 16541 9229 16575
rect 9263 16574 9275 16575
rect 15197 16575 15255 16581
rect 9263 16546 9297 16574
rect 15197 16572 15209 16575
rect 9263 16541 9275 16546
rect 15107 16544 15209 16572
rect 9217 16535 9275 16541
rect 15197 16541 15209 16544
rect 15243 16572 15255 16575
rect 15378 16572 15384 16584
rect 15243 16544 15384 16572
rect 15243 16541 15255 16544
rect 15197 16535 15255 16541
rect 15378 16532 15384 16544
rect 15436 16532 15442 16584
rect 15488 16581 15516 16612
rect 15565 16609 15577 16612
rect 15611 16609 15623 16643
rect 15565 16603 15623 16609
rect 15473 16575 15531 16581
rect 15473 16541 15485 16575
rect 15519 16574 15531 16575
rect 15519 16546 15553 16574
rect 15519 16541 15531 16546
rect 15473 16535 15531 16541
rect 1903 16408 3280 16436
rect 1903 16405 1915 16408
rect 1857 16399 1915 16405
rect 3786 16396 3792 16448
rect 3844 16436 3850 16448
rect 3973 16439 4031 16445
rect 3973 16436 3985 16439
rect 3844 16408 3985 16436
rect 3844 16396 3850 16408
rect 3973 16405 3985 16408
rect 4019 16405 4031 16439
rect 3973 16399 4031 16405
rect 7282 16396 7288 16448
rect 7340 16436 7346 16448
rect 9033 16439 9091 16445
rect 9033 16436 9045 16439
rect 7340 16408 9045 16436
rect 7340 16396 7346 16408
rect 9033 16405 9045 16408
rect 9079 16405 9091 16439
rect 15010 16436 15016 16448
rect 14971 16408 15016 16436
rect 9033 16399 9091 16405
rect 15010 16396 15016 16408
rect 15068 16396 15074 16448
rect 15102 16396 15108 16448
rect 15160 16436 15166 16448
rect 15289 16439 15347 16445
rect 15289 16436 15301 16439
rect 15160 16408 15301 16436
rect 15160 16396 15166 16408
rect 15289 16405 15301 16408
rect 15335 16405 15347 16439
rect 15289 16399 15347 16405
rect 1104 16346 16008 16368
rect 1104 16294 4698 16346
rect 4750 16294 4762 16346
rect 4814 16294 4826 16346
rect 4878 16294 4890 16346
rect 4942 16294 4954 16346
rect 5006 16294 8446 16346
rect 8498 16294 8510 16346
rect 8562 16294 8574 16346
rect 8626 16294 8638 16346
rect 8690 16294 8702 16346
rect 8754 16294 12194 16346
rect 12246 16294 12258 16346
rect 12310 16294 12322 16346
rect 12374 16294 12386 16346
rect 12438 16294 12450 16346
rect 12502 16294 16008 16346
rect 1104 16272 16008 16294
rect 1302 16192 1308 16244
rect 1360 16232 1366 16244
rect 1397 16235 1455 16241
rect 1397 16232 1409 16235
rect 1360 16204 1409 16232
rect 1360 16192 1366 16204
rect 1397 16201 1409 16204
rect 1443 16201 1455 16235
rect 1397 16195 1455 16201
rect 1578 16192 1584 16244
rect 1636 16232 1642 16244
rect 5074 16232 5080 16244
rect 1636 16204 5080 16232
rect 1636 16192 1642 16204
rect 5074 16192 5080 16204
rect 5132 16192 5138 16244
rect 15381 16099 15439 16105
rect 15381 16065 15393 16099
rect 15427 16096 15439 16099
rect 15657 16099 15715 16105
rect 15657 16096 15669 16099
rect 15427 16068 15669 16096
rect 15427 16065 15439 16068
rect 15381 16059 15439 16065
rect 15657 16065 15669 16068
rect 15703 16096 15715 16099
rect 15930 16096 15936 16108
rect 15703 16068 15936 16096
rect 15703 16065 15715 16068
rect 15657 16059 15715 16065
rect 15930 16056 15936 16068
rect 15988 16056 15994 16108
rect 15470 15892 15476 15904
rect 15431 15864 15476 15892
rect 15470 15852 15476 15864
rect 15528 15852 15534 15904
rect 1104 15802 16008 15824
rect 1104 15750 2824 15802
rect 2876 15750 2888 15802
rect 2940 15750 2952 15802
rect 3004 15750 3016 15802
rect 3068 15750 3080 15802
rect 3132 15750 6572 15802
rect 6624 15750 6636 15802
rect 6688 15750 6700 15802
rect 6752 15750 6764 15802
rect 6816 15750 6828 15802
rect 6880 15750 10320 15802
rect 10372 15750 10384 15802
rect 10436 15750 10448 15802
rect 10500 15750 10512 15802
rect 10564 15750 10576 15802
rect 10628 15750 14068 15802
rect 14120 15750 14132 15802
rect 14184 15750 14196 15802
rect 14248 15750 14260 15802
rect 14312 15750 14324 15802
rect 14376 15750 16008 15802
rect 1104 15728 16008 15750
rect 1104 15258 16008 15280
rect 1104 15206 4698 15258
rect 4750 15206 4762 15258
rect 4814 15206 4826 15258
rect 4878 15206 4890 15258
rect 4942 15206 4954 15258
rect 5006 15206 8446 15258
rect 8498 15206 8510 15258
rect 8562 15206 8574 15258
rect 8626 15206 8638 15258
rect 8690 15206 8702 15258
rect 8754 15206 12194 15258
rect 12246 15206 12258 15258
rect 12310 15206 12322 15258
rect 12374 15206 12386 15258
rect 12438 15206 12450 15258
rect 12502 15206 16008 15258
rect 1104 15184 16008 15206
rect 1104 14714 16008 14736
rect 1104 14662 2824 14714
rect 2876 14662 2888 14714
rect 2940 14662 2952 14714
rect 3004 14662 3016 14714
rect 3068 14662 3080 14714
rect 3132 14662 6572 14714
rect 6624 14662 6636 14714
rect 6688 14662 6700 14714
rect 6752 14662 6764 14714
rect 6816 14662 6828 14714
rect 6880 14662 10320 14714
rect 10372 14662 10384 14714
rect 10436 14662 10448 14714
rect 10500 14662 10512 14714
rect 10564 14662 10576 14714
rect 10628 14662 14068 14714
rect 14120 14662 14132 14714
rect 14184 14662 14196 14714
rect 14248 14662 14260 14714
rect 14312 14662 14324 14714
rect 14376 14662 16008 14714
rect 1104 14640 16008 14662
rect 1104 14170 16008 14192
rect 1104 14118 4698 14170
rect 4750 14118 4762 14170
rect 4814 14118 4826 14170
rect 4878 14118 4890 14170
rect 4942 14118 4954 14170
rect 5006 14118 8446 14170
rect 8498 14118 8510 14170
rect 8562 14118 8574 14170
rect 8626 14118 8638 14170
rect 8690 14118 8702 14170
rect 8754 14118 12194 14170
rect 12246 14118 12258 14170
rect 12310 14118 12322 14170
rect 12374 14118 12386 14170
rect 12438 14118 12450 14170
rect 12502 14118 16008 14170
rect 1104 14096 16008 14118
rect 5074 13920 5080 13932
rect 5035 13892 5080 13920
rect 5074 13880 5080 13892
rect 5132 13880 5138 13932
rect 3510 13812 3516 13864
rect 3568 13852 3574 13864
rect 4617 13855 4675 13861
rect 4617 13852 4629 13855
rect 3568 13824 4629 13852
rect 3568 13812 3574 13824
rect 4617 13821 4629 13824
rect 4663 13821 4675 13855
rect 4617 13815 4675 13821
rect 4985 13719 5043 13725
rect 4985 13685 4997 13719
rect 5031 13716 5043 13719
rect 7650 13716 7656 13728
rect 5031 13688 7656 13716
rect 5031 13685 5043 13688
rect 4985 13679 5043 13685
rect 7650 13676 7656 13688
rect 7708 13676 7714 13728
rect 1104 13626 16008 13648
rect 1104 13574 2824 13626
rect 2876 13574 2888 13626
rect 2940 13574 2952 13626
rect 3004 13574 3016 13626
rect 3068 13574 3080 13626
rect 3132 13574 6572 13626
rect 6624 13574 6636 13626
rect 6688 13574 6700 13626
rect 6752 13574 6764 13626
rect 6816 13574 6828 13626
rect 6880 13574 10320 13626
rect 10372 13574 10384 13626
rect 10436 13574 10448 13626
rect 10500 13574 10512 13626
rect 10564 13574 10576 13626
rect 10628 13574 14068 13626
rect 14120 13574 14132 13626
rect 14184 13574 14196 13626
rect 14248 13574 14260 13626
rect 14312 13574 14324 13626
rect 14376 13574 16008 13626
rect 1104 13552 16008 13574
rect 1104 13082 16008 13104
rect 1104 13030 4698 13082
rect 4750 13030 4762 13082
rect 4814 13030 4826 13082
rect 4878 13030 4890 13082
rect 4942 13030 4954 13082
rect 5006 13030 8446 13082
rect 8498 13030 8510 13082
rect 8562 13030 8574 13082
rect 8626 13030 8638 13082
rect 8690 13030 8702 13082
rect 8754 13030 12194 13082
rect 12246 13030 12258 13082
rect 12310 13030 12322 13082
rect 12374 13030 12386 13082
rect 12438 13030 12450 13082
rect 12502 13030 16008 13082
rect 1104 13008 16008 13030
rect 3142 12928 3148 12980
rect 3200 12968 3206 12980
rect 4065 12971 4123 12977
rect 4065 12968 4077 12971
rect 3200 12940 4077 12968
rect 3200 12928 3206 12940
rect 4065 12937 4077 12940
rect 4111 12937 4123 12971
rect 4065 12931 4123 12937
rect 5718 12928 5724 12980
rect 5776 12968 5782 12980
rect 5813 12971 5871 12977
rect 5813 12968 5825 12971
rect 5776 12940 5825 12968
rect 5776 12928 5782 12940
rect 5813 12937 5825 12940
rect 5859 12937 5871 12971
rect 5813 12931 5871 12937
rect 14461 12971 14519 12977
rect 14461 12937 14473 12971
rect 14507 12968 14519 12971
rect 14734 12968 14740 12980
rect 14507 12940 14740 12968
rect 14507 12937 14519 12940
rect 14461 12931 14519 12937
rect 14734 12928 14740 12940
rect 14792 12928 14798 12980
rect 4154 12860 4160 12912
rect 4212 12900 4218 12912
rect 4586 12903 4644 12909
rect 4586 12900 4598 12903
rect 4212 12872 4598 12900
rect 4212 12860 4218 12872
rect 4586 12869 4598 12872
rect 4632 12869 4644 12903
rect 4586 12863 4644 12869
rect 7650 12860 7656 12912
rect 7708 12900 7714 12912
rect 7708 12872 15424 12900
rect 7708 12860 7714 12872
rect 4249 12835 4307 12841
rect 4249 12801 4261 12835
rect 4295 12832 4307 12835
rect 5997 12835 6055 12841
rect 4295 12804 5580 12832
rect 4295 12801 4307 12804
rect 4249 12795 4307 12801
rect 4338 12764 4344 12776
rect 4299 12736 4344 12764
rect 4338 12724 4344 12736
rect 4396 12724 4402 12776
rect 5552 12764 5580 12804
rect 5997 12801 6009 12835
rect 6043 12832 6055 12835
rect 8386 12832 8392 12844
rect 6043 12804 8392 12832
rect 6043 12801 6055 12804
rect 5997 12795 6055 12801
rect 8386 12792 8392 12804
rect 8444 12792 8450 12844
rect 15396 12841 15424 12872
rect 14277 12835 14335 12841
rect 14277 12832 14289 12835
rect 14108 12804 14289 12832
rect 7098 12764 7104 12776
rect 5552 12736 7104 12764
rect 7098 12724 7104 12736
rect 7156 12724 7162 12776
rect 5721 12699 5779 12705
rect 5721 12665 5733 12699
rect 5767 12696 5779 12699
rect 7006 12696 7012 12708
rect 5767 12668 7012 12696
rect 5767 12665 5779 12668
rect 5721 12659 5779 12665
rect 7006 12656 7012 12668
rect 7064 12656 7070 12708
rect 13906 12588 13912 12640
rect 13964 12628 13970 12640
rect 14108 12637 14136 12804
rect 14277 12801 14289 12804
rect 14323 12801 14335 12835
rect 14277 12795 14335 12801
rect 15381 12835 15439 12841
rect 15381 12801 15393 12835
rect 15427 12801 15439 12835
rect 15381 12795 15439 12801
rect 14093 12631 14151 12637
rect 14093 12628 14105 12631
rect 13964 12600 14105 12628
rect 13964 12588 13970 12600
rect 14093 12597 14105 12600
rect 14139 12597 14151 12631
rect 15562 12628 15568 12640
rect 15523 12600 15568 12628
rect 14093 12591 14151 12597
rect 15562 12588 15568 12600
rect 15620 12588 15626 12640
rect 1104 12538 16008 12560
rect 1104 12486 2824 12538
rect 2876 12486 2888 12538
rect 2940 12486 2952 12538
rect 3004 12486 3016 12538
rect 3068 12486 3080 12538
rect 3132 12486 6572 12538
rect 6624 12486 6636 12538
rect 6688 12486 6700 12538
rect 6752 12486 6764 12538
rect 6816 12486 6828 12538
rect 6880 12486 10320 12538
rect 10372 12486 10384 12538
rect 10436 12486 10448 12538
rect 10500 12486 10512 12538
rect 10564 12486 10576 12538
rect 10628 12486 14068 12538
rect 14120 12486 14132 12538
rect 14184 12486 14196 12538
rect 14248 12486 14260 12538
rect 14312 12486 14324 12538
rect 14376 12486 16008 12538
rect 1104 12464 16008 12486
rect 2498 12384 2504 12436
rect 2556 12424 2562 12436
rect 5077 12427 5135 12433
rect 5077 12424 5089 12427
rect 2556 12396 5089 12424
rect 2556 12384 2562 12396
rect 5077 12393 5089 12396
rect 5123 12393 5135 12427
rect 5077 12387 5135 12393
rect 5442 12384 5448 12436
rect 5500 12424 5506 12436
rect 7377 12427 7435 12433
rect 7377 12424 7389 12427
rect 5500 12396 7389 12424
rect 5500 12384 5506 12396
rect 7377 12393 7389 12396
rect 7423 12393 7435 12427
rect 7377 12387 7435 12393
rect 8294 12384 8300 12436
rect 8352 12424 8358 12436
rect 9309 12427 9367 12433
rect 9309 12424 9321 12427
rect 8352 12396 9321 12424
rect 8352 12384 8358 12396
rect 9309 12393 9321 12396
rect 9355 12393 9367 12427
rect 9309 12387 9367 12393
rect 5261 12223 5319 12229
rect 5261 12189 5273 12223
rect 5307 12189 5319 12223
rect 5261 12183 5319 12189
rect 7561 12223 7619 12229
rect 7561 12189 7573 12223
rect 7607 12220 7619 12223
rect 7607 12192 9260 12220
rect 7607 12189 7619 12192
rect 7561 12183 7619 12189
rect 5276 12152 5304 12183
rect 8110 12152 8116 12164
rect 5276 12124 8116 12152
rect 8110 12112 8116 12124
rect 8168 12112 8174 12164
rect 9232 12152 9260 12192
rect 9306 12180 9312 12232
rect 9364 12220 9370 12232
rect 9493 12223 9551 12229
rect 9493 12220 9505 12223
rect 9364 12192 9505 12220
rect 9364 12180 9370 12192
rect 9493 12189 9505 12192
rect 9539 12189 9551 12223
rect 9493 12183 9551 12189
rect 9766 12152 9772 12164
rect 9232 12124 9772 12152
rect 9766 12112 9772 12124
rect 9824 12112 9830 12164
rect 1104 11994 16008 12016
rect 1104 11942 4698 11994
rect 4750 11942 4762 11994
rect 4814 11942 4826 11994
rect 4878 11942 4890 11994
rect 4942 11942 4954 11994
rect 5006 11942 8446 11994
rect 8498 11942 8510 11994
rect 8562 11942 8574 11994
rect 8626 11942 8638 11994
rect 8690 11942 8702 11994
rect 8754 11942 12194 11994
rect 12246 11942 12258 11994
rect 12310 11942 12322 11994
rect 12374 11942 12386 11994
rect 12438 11942 12450 11994
rect 12502 11942 16008 11994
rect 1104 11920 16008 11942
rect 7190 11880 7196 11892
rect 7151 11852 7196 11880
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 7837 11883 7895 11889
rect 7837 11849 7849 11883
rect 7883 11849 7895 11883
rect 7837 11843 7895 11849
rect 6454 11772 6460 11824
rect 6512 11812 6518 11824
rect 7852 11812 7880 11843
rect 6512 11784 7880 11812
rect 6512 11772 6518 11784
rect 1394 11744 1400 11756
rect 1355 11716 1400 11744
rect 1394 11704 1400 11716
rect 1452 11744 1458 11756
rect 1673 11747 1731 11753
rect 1673 11744 1685 11747
rect 1452 11716 1685 11744
rect 1452 11704 1458 11716
rect 1673 11713 1685 11716
rect 1719 11713 1731 11747
rect 7374 11744 7380 11756
rect 7335 11716 7380 11744
rect 1673 11707 1731 11713
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 7742 11744 7748 11756
rect 7703 11716 7748 11744
rect 7742 11704 7748 11716
rect 7800 11704 7806 11756
rect 8018 11744 8024 11756
rect 7979 11716 8024 11744
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 5718 11636 5724 11688
rect 5776 11676 5782 11688
rect 8202 11676 8208 11688
rect 5776 11648 8208 11676
rect 5776 11636 5782 11648
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 6362 11568 6368 11620
rect 6420 11608 6426 11620
rect 7561 11611 7619 11617
rect 7561 11608 7573 11611
rect 6420 11580 7573 11608
rect 6420 11568 6426 11580
rect 7561 11577 7573 11580
rect 7607 11577 7619 11611
rect 7561 11571 7619 11577
rect 1581 11543 1639 11549
rect 1581 11509 1593 11543
rect 1627 11540 1639 11543
rect 5902 11540 5908 11552
rect 1627 11512 5908 11540
rect 1627 11509 1639 11512
rect 1581 11503 1639 11509
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 8757 11543 8815 11549
rect 8757 11509 8769 11543
rect 8803 11540 8815 11543
rect 8846 11540 8852 11552
rect 8803 11512 8852 11540
rect 8803 11509 8815 11512
rect 8757 11503 8815 11509
rect 8846 11500 8852 11512
rect 8904 11500 8910 11552
rect 1104 11450 16008 11472
rect 1104 11398 2824 11450
rect 2876 11398 2888 11450
rect 2940 11398 2952 11450
rect 3004 11398 3016 11450
rect 3068 11398 3080 11450
rect 3132 11398 6572 11450
rect 6624 11398 6636 11450
rect 6688 11398 6700 11450
rect 6752 11398 6764 11450
rect 6816 11398 6828 11450
rect 6880 11398 10320 11450
rect 10372 11398 10384 11450
rect 10436 11398 10448 11450
rect 10500 11398 10512 11450
rect 10564 11398 10576 11450
rect 10628 11398 14068 11450
rect 14120 11398 14132 11450
rect 14184 11398 14196 11450
rect 14248 11398 14260 11450
rect 14312 11398 14324 11450
rect 14376 11398 16008 11450
rect 1104 11376 16008 11398
rect 7006 11296 7012 11348
rect 7064 11336 7070 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 7064 11308 8953 11336
rect 7064 11296 7070 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 8941 11299 8999 11305
rect 8202 11268 8208 11280
rect 8163 11240 8208 11268
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 10870 11268 10876 11280
rect 8496 11240 10876 11268
rect 4338 11160 4344 11212
rect 4396 11200 4402 11212
rect 6825 11203 6883 11209
rect 6825 11200 6837 11203
rect 4396 11172 6837 11200
rect 4396 11160 4402 11172
rect 6825 11169 6837 11172
rect 6871 11169 6883 11203
rect 6825 11163 6883 11169
rect 6840 11132 6868 11163
rect 8496 11141 8524 11240
rect 10870 11228 10876 11240
rect 10928 11228 10934 11280
rect 9490 11200 9496 11212
rect 9451 11172 9496 11200
rect 9490 11160 9496 11172
rect 9548 11160 9554 11212
rect 8481 11135 8539 11141
rect 6840 11104 8294 11132
rect 4338 11024 4344 11076
rect 4396 11064 4402 11076
rect 4396 11036 6868 11064
rect 4396 11024 4402 11036
rect 6840 10996 6868 11036
rect 6914 11024 6920 11076
rect 6972 11064 6978 11076
rect 7070 11067 7128 11073
rect 7070 11064 7082 11067
rect 6972 11036 7082 11064
rect 6972 11024 6978 11036
rect 7070 11033 7082 11036
rect 7116 11033 7128 11067
rect 8266 11064 8294 11104
rect 8481 11101 8493 11135
rect 8527 11101 8539 11135
rect 8481 11095 8539 11101
rect 8757 11135 8815 11141
rect 8757 11101 8769 11135
rect 8803 11132 8815 11135
rect 9309 11135 9367 11141
rect 9309 11132 9321 11135
rect 8803 11104 9321 11132
rect 8803 11101 8815 11104
rect 8757 11095 8815 11101
rect 9309 11101 9321 11104
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 9122 11064 9128 11076
rect 7070 11027 7128 11033
rect 7208 11036 8156 11064
rect 8266 11036 9128 11064
rect 7208 10996 7236 11036
rect 6840 10968 7236 10996
rect 8128 10996 8156 11036
rect 9122 11024 9128 11036
rect 9180 11024 9186 11076
rect 9398 11064 9404 11076
rect 9359 11036 9404 11064
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 8297 10999 8355 11005
rect 8297 10996 8309 10999
rect 8128 10968 8309 10996
rect 8297 10965 8309 10968
rect 8343 10965 8355 10999
rect 8297 10959 8355 10965
rect 9214 10956 9220 11008
rect 9272 10996 9278 11008
rect 9582 10996 9588 11008
rect 9272 10968 9588 10996
rect 9272 10956 9278 10968
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 1104 10906 16008 10928
rect 1104 10854 4698 10906
rect 4750 10854 4762 10906
rect 4814 10854 4826 10906
rect 4878 10854 4890 10906
rect 4942 10854 4954 10906
rect 5006 10854 8446 10906
rect 8498 10854 8510 10906
rect 8562 10854 8574 10906
rect 8626 10854 8638 10906
rect 8690 10854 8702 10906
rect 8754 10854 12194 10906
rect 12246 10854 12258 10906
rect 12310 10854 12322 10906
rect 12374 10854 12386 10906
rect 12438 10854 12450 10906
rect 12502 10854 16008 10906
rect 1104 10832 16008 10854
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 5721 10795 5779 10801
rect 5721 10792 5733 10795
rect 5592 10764 5733 10792
rect 5592 10752 5598 10764
rect 5721 10761 5733 10764
rect 5767 10761 5779 10795
rect 5721 10755 5779 10761
rect 5997 10795 6055 10801
rect 5997 10761 6009 10795
rect 6043 10761 6055 10795
rect 5997 10755 6055 10761
rect 3602 10684 3608 10736
rect 3660 10724 3666 10736
rect 6012 10724 6040 10755
rect 7650 10752 7656 10804
rect 7708 10792 7714 10804
rect 7745 10795 7803 10801
rect 7745 10792 7757 10795
rect 7708 10764 7757 10792
rect 7708 10752 7714 10764
rect 7745 10761 7757 10764
rect 7791 10761 7803 10795
rect 7745 10755 7803 10761
rect 8938 10752 8944 10804
rect 8996 10792 9002 10804
rect 9217 10795 9275 10801
rect 9217 10792 9229 10795
rect 8996 10764 9229 10792
rect 8996 10752 9002 10764
rect 9217 10761 9229 10764
rect 9263 10761 9275 10795
rect 9217 10755 9275 10761
rect 9585 10795 9643 10801
rect 9585 10761 9597 10795
rect 9631 10761 9643 10795
rect 9585 10755 9643 10761
rect 3660 10696 6040 10724
rect 6104 10696 7604 10724
rect 3660 10684 3666 10696
rect 3510 10665 3516 10668
rect 3488 10659 3516 10665
rect 3488 10625 3500 10659
rect 3488 10619 3516 10625
rect 3510 10616 3516 10619
rect 3568 10616 3574 10668
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 5905 10659 5963 10665
rect 5905 10656 5917 10659
rect 5592 10628 5917 10656
rect 5592 10616 5598 10628
rect 5905 10625 5917 10628
rect 5951 10625 5963 10659
rect 5905 10619 5963 10625
rect 5994 10616 6000 10668
rect 6052 10656 6058 10668
rect 6104 10656 6132 10696
rect 6052 10628 6132 10656
rect 6181 10659 6239 10665
rect 6052 10616 6058 10628
rect 6181 10625 6193 10659
rect 6227 10625 6239 10659
rect 6181 10619 6239 10625
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10625 6607 10659
rect 6822 10656 6828 10668
rect 6783 10628 6828 10656
rect 6549 10619 6607 10625
rect 5626 10548 5632 10600
rect 5684 10588 5690 10600
rect 6196 10588 6224 10619
rect 5684 10560 6224 10588
rect 5684 10548 5690 10560
rect 5074 10480 5080 10532
rect 5132 10520 5138 10532
rect 6365 10523 6423 10529
rect 6365 10520 6377 10523
rect 5132 10492 6377 10520
rect 5132 10480 5138 10492
rect 6365 10489 6377 10492
rect 6411 10489 6423 10523
rect 6564 10520 6592 10619
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 7098 10656 7104 10668
rect 7024 10628 7104 10656
rect 7024 10597 7052 10628
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 7282 10616 7288 10668
rect 7340 10656 7346 10668
rect 7466 10656 7472 10668
rect 7340 10628 7472 10656
rect 7340 10616 7346 10628
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 7576 10656 7604 10696
rect 8846 10684 8852 10736
rect 8904 10733 8910 10736
rect 8904 10724 8916 10733
rect 9600 10724 9628 10755
rect 12066 10724 12072 10736
rect 8904 10696 8949 10724
rect 9048 10696 9628 10724
rect 9784 10696 12072 10724
rect 8904 10687 8916 10696
rect 8904 10684 8910 10687
rect 9048 10656 9076 10696
rect 7576 10628 9076 10656
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10656 9459 10659
rect 9582 10656 9588 10668
rect 9447 10628 9588 10656
rect 9447 10625 9459 10628
rect 9401 10619 9459 10625
rect 9582 10616 9588 10628
rect 9640 10616 9646 10668
rect 9784 10665 9812 10696
rect 12066 10684 12072 10696
rect 12124 10684 12130 10736
rect 9769 10659 9827 10665
rect 9769 10625 9781 10659
rect 9815 10625 9827 10659
rect 9769 10619 9827 10625
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10656 10103 10659
rect 11238 10656 11244 10668
rect 10091 10628 11244 10656
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10557 7067 10591
rect 7190 10588 7196 10600
rect 7151 10560 7196 10588
rect 7009 10551 7067 10557
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 9122 10548 9128 10600
rect 9180 10588 9186 10600
rect 11146 10588 11152 10600
rect 9180 10560 11152 10588
rect 9180 10548 9186 10560
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 11054 10520 11060 10532
rect 6564 10492 8248 10520
rect 6365 10483 6423 10489
rect 3559 10455 3617 10461
rect 3559 10421 3571 10455
rect 3605 10452 3617 10455
rect 5810 10452 5816 10464
rect 3605 10424 5816 10452
rect 3605 10421 3617 10424
rect 3559 10415 3617 10421
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 6454 10412 6460 10464
rect 6512 10452 6518 10464
rect 6641 10455 6699 10461
rect 6641 10452 6653 10455
rect 6512 10424 6653 10452
rect 6512 10412 6518 10424
rect 6641 10421 6653 10424
rect 6687 10421 6699 10455
rect 7650 10452 7656 10464
rect 7611 10424 7656 10452
rect 6641 10415 6699 10421
rect 7650 10412 7656 10424
rect 7708 10412 7714 10464
rect 8220 10452 8248 10492
rect 9784 10492 11060 10520
rect 9784 10452 9812 10492
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 8220 10424 9812 10452
rect 9861 10455 9919 10461
rect 9861 10421 9873 10455
rect 9907 10452 9919 10455
rect 9950 10452 9956 10464
rect 9907 10424 9956 10452
rect 9907 10421 9919 10424
rect 9861 10415 9919 10421
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 11698 10412 11704 10464
rect 11756 10452 11762 10464
rect 14642 10452 14648 10464
rect 11756 10424 14648 10452
rect 11756 10412 11762 10424
rect 14642 10412 14648 10424
rect 14700 10412 14706 10464
rect 1104 10362 16008 10384
rect 1104 10310 2824 10362
rect 2876 10310 2888 10362
rect 2940 10310 2952 10362
rect 3004 10310 3016 10362
rect 3068 10310 3080 10362
rect 3132 10310 6572 10362
rect 6624 10310 6636 10362
rect 6688 10310 6700 10362
rect 6752 10310 6764 10362
rect 6816 10310 6828 10362
rect 6880 10310 10320 10362
rect 10372 10310 10384 10362
rect 10436 10310 10448 10362
rect 10500 10310 10512 10362
rect 10564 10310 10576 10362
rect 10628 10310 14068 10362
rect 14120 10310 14132 10362
rect 14184 10310 14196 10362
rect 14248 10310 14260 10362
rect 14312 10310 14324 10362
rect 14376 10310 16008 10362
rect 1104 10288 16008 10310
rect 8110 10208 8116 10260
rect 8168 10248 8174 10260
rect 11241 10251 11299 10257
rect 8168 10220 10824 10248
rect 8168 10208 8174 10220
rect 3234 10140 3240 10192
rect 3292 10180 3298 10192
rect 5077 10183 5135 10189
rect 5077 10180 5089 10183
rect 3292 10152 5089 10180
rect 3292 10140 3298 10152
rect 5077 10149 5089 10152
rect 5123 10149 5135 10183
rect 5077 10143 5135 10149
rect 5534 10140 5540 10192
rect 5592 10180 5598 10192
rect 6362 10180 6368 10192
rect 5592 10152 6368 10180
rect 5592 10140 5598 10152
rect 6362 10140 6368 10152
rect 6420 10140 6426 10192
rect 7650 10140 7656 10192
rect 7708 10180 7714 10192
rect 7708 10152 9812 10180
rect 7708 10140 7714 10152
rect 5718 10112 5724 10124
rect 5679 10084 5724 10112
rect 5718 10072 5724 10084
rect 5776 10072 5782 10124
rect 5810 10072 5816 10124
rect 5868 10112 5874 10124
rect 6089 10115 6147 10121
rect 6089 10112 6101 10115
rect 5868 10084 6101 10112
rect 5868 10072 5874 10084
rect 6089 10081 6101 10084
rect 6135 10081 6147 10115
rect 6089 10075 6147 10081
rect 7098 10072 7104 10124
rect 7156 10112 7162 10124
rect 8113 10115 8171 10121
rect 8113 10112 8125 10115
rect 7156 10084 8125 10112
rect 7156 10072 7162 10084
rect 8113 10081 8125 10084
rect 8159 10081 8171 10115
rect 8294 10112 8300 10124
rect 8255 10084 8300 10112
rect 8113 10075 8171 10081
rect 8294 10072 8300 10084
rect 8352 10072 8358 10124
rect 8386 10072 8392 10124
rect 8444 10112 8450 10124
rect 8444 10084 9444 10112
rect 8444 10072 8450 10084
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10044 5043 10047
rect 5258 10044 5264 10056
rect 5031 10016 5264 10044
rect 5031 10013 5043 10016
rect 4985 10007 5043 10013
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 5902 10044 5908 10056
rect 5863 10016 5908 10044
rect 5902 10004 5908 10016
rect 5960 10004 5966 10056
rect 7742 10044 7748 10056
rect 7703 10016 7748 10044
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 9416 10044 9444 10084
rect 9490 10072 9496 10124
rect 9548 10112 9554 10124
rect 9585 10115 9643 10121
rect 9585 10112 9597 10115
rect 9548 10084 9597 10112
rect 9548 10072 9554 10084
rect 9585 10081 9597 10084
rect 9631 10112 9643 10115
rect 9784 10112 9812 10152
rect 10042 10140 10048 10192
rect 10100 10180 10106 10192
rect 10689 10183 10747 10189
rect 10689 10180 10701 10183
rect 10100 10152 10701 10180
rect 10100 10140 10106 10152
rect 10689 10149 10701 10152
rect 10735 10149 10747 10183
rect 10796 10180 10824 10220
rect 11241 10217 11253 10251
rect 11287 10248 11299 10251
rect 11422 10248 11428 10260
rect 11287 10220 11428 10248
rect 11287 10217 11299 10220
rect 11241 10211 11299 10217
rect 11422 10208 11428 10220
rect 11480 10208 11486 10260
rect 12069 10251 12127 10257
rect 12069 10248 12081 10251
rect 11532 10220 12081 10248
rect 11532 10180 11560 10220
rect 12069 10217 12081 10220
rect 12115 10217 12127 10251
rect 12069 10211 12127 10217
rect 12526 10208 12532 10260
rect 12584 10248 12590 10260
rect 12621 10251 12679 10257
rect 12621 10248 12633 10251
rect 12584 10220 12633 10248
rect 12584 10208 12590 10220
rect 12621 10217 12633 10220
rect 12667 10217 12679 10251
rect 13170 10248 13176 10260
rect 13131 10220 13176 10248
rect 12621 10211 12679 10217
rect 13170 10208 13176 10220
rect 13228 10208 13234 10260
rect 10796 10152 11560 10180
rect 10689 10143 10747 10149
rect 11606 10140 11612 10192
rect 11664 10180 11670 10192
rect 12345 10183 12403 10189
rect 12345 10180 12357 10183
rect 11664 10152 12357 10180
rect 11664 10140 11670 10152
rect 12345 10149 12357 10152
rect 12391 10149 12403 10183
rect 15010 10180 15016 10192
rect 12345 10143 12403 10149
rect 12544 10152 15016 10180
rect 10321 10115 10379 10121
rect 10321 10112 10333 10115
rect 9631 10084 9720 10112
rect 9784 10084 10333 10112
rect 9631 10081 9643 10084
rect 9585 10075 9643 10081
rect 9692 10044 9720 10084
rect 10321 10081 10333 10084
rect 10367 10081 10379 10115
rect 10321 10075 10379 10081
rect 10413 10115 10471 10121
rect 10413 10081 10425 10115
rect 10459 10081 10471 10115
rect 10413 10075 10471 10081
rect 10428 10044 10456 10075
rect 11238 10072 11244 10124
rect 11296 10112 11302 10124
rect 11296 10084 12296 10112
rect 11296 10072 11302 10084
rect 9416 10016 9628 10044
rect 9692 10016 10456 10044
rect 10873 10047 10931 10053
rect 5445 9979 5503 9985
rect 5445 9945 5457 9979
rect 5491 9976 5503 9979
rect 5810 9976 5816 9988
rect 5491 9948 5816 9976
rect 5491 9945 5503 9948
rect 5445 9939 5503 9945
rect 5810 9936 5816 9948
rect 5868 9936 5874 9988
rect 7558 9936 7564 9988
rect 7616 9976 7622 9988
rect 9214 9976 9220 9988
rect 7616 9948 9220 9976
rect 7616 9936 7622 9948
rect 9214 9936 9220 9948
rect 9272 9976 9278 9988
rect 9493 9979 9551 9985
rect 9493 9976 9505 9979
rect 9272 9948 9505 9976
rect 9272 9936 9278 9948
rect 9493 9945 9505 9948
rect 9539 9945 9551 9979
rect 9600 9976 9628 10016
rect 10873 10013 10885 10047
rect 10919 10044 10931 10047
rect 10962 10044 10968 10056
rect 10919 10016 10968 10044
rect 10919 10013 10931 10016
rect 10873 10007 10931 10013
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 11149 10047 11207 10053
rect 11149 10013 11161 10047
rect 11195 10044 11207 10047
rect 11330 10044 11336 10056
rect 11195 10016 11336 10044
rect 11195 10013 11207 10016
rect 11149 10007 11207 10013
rect 11330 10004 11336 10016
rect 11388 10004 11394 10056
rect 11425 10047 11483 10053
rect 11425 10013 11437 10047
rect 11471 10044 11483 10047
rect 11514 10044 11520 10056
rect 11471 10016 11520 10044
rect 11471 10013 11483 10016
rect 11425 10007 11483 10013
rect 11514 10004 11520 10016
rect 11572 10004 11578 10056
rect 11698 10044 11704 10056
rect 11659 10016 11704 10044
rect 11698 10004 11704 10016
rect 11756 10004 11762 10056
rect 12268 10053 12296 10084
rect 12544 10053 12572 10152
rect 15010 10140 15016 10152
rect 15068 10140 15074 10192
rect 15470 10112 15476 10124
rect 13096 10084 15476 10112
rect 11977 10047 12035 10053
rect 11977 10013 11989 10047
rect 12023 10013 12035 10047
rect 11977 10007 12035 10013
rect 12253 10047 12311 10053
rect 12253 10013 12265 10047
rect 12299 10013 12311 10047
rect 12253 10007 12311 10013
rect 12529 10047 12587 10053
rect 12529 10013 12541 10047
rect 12575 10013 12587 10047
rect 12529 10007 12587 10013
rect 12805 10047 12863 10053
rect 12805 10013 12817 10047
rect 12851 10044 12863 10047
rect 12986 10044 12992 10056
rect 12851 10016 12992 10044
rect 12851 10013 12863 10016
rect 12805 10007 12863 10013
rect 10318 9976 10324 9988
rect 9600 9948 10324 9976
rect 9493 9939 9551 9945
rect 10318 9936 10324 9948
rect 10376 9936 10382 9988
rect 11992 9976 12020 10007
rect 12986 10004 12992 10016
rect 13044 10004 13050 10056
rect 13096 10053 13124 10084
rect 15470 10072 15476 10084
rect 15528 10072 15534 10124
rect 13081 10047 13139 10053
rect 13081 10013 13093 10047
rect 13127 10013 13139 10047
rect 13354 10044 13360 10056
rect 13315 10016 13360 10044
rect 13081 10007 13139 10013
rect 13354 10004 13360 10016
rect 13412 10004 13418 10056
rect 15102 9976 15108 9988
rect 11992 9948 15108 9976
rect 15102 9936 15108 9948
rect 15160 9936 15166 9988
rect 3694 9868 3700 9920
rect 3752 9908 3758 9920
rect 4801 9911 4859 9917
rect 4801 9908 4813 9911
rect 3752 9880 4813 9908
rect 3752 9868 3758 9880
rect 4801 9877 4813 9880
rect 4847 9877 4859 9911
rect 5534 9908 5540 9920
rect 5495 9880 5540 9908
rect 4801 9871 4859 9877
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 7282 9868 7288 9920
rect 7340 9908 7346 9920
rect 8386 9908 8392 9920
rect 7340 9880 8392 9908
rect 7340 9868 7346 9880
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 8720 9880 8769 9908
rect 8720 9868 8726 9880
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 8757 9871 8815 9877
rect 8938 9868 8944 9920
rect 8996 9908 9002 9920
rect 9033 9911 9091 9917
rect 9033 9908 9045 9911
rect 8996 9880 9045 9908
rect 8996 9868 9002 9880
rect 9033 9877 9045 9880
rect 9079 9877 9091 9911
rect 9033 9871 9091 9877
rect 9306 9868 9312 9920
rect 9364 9908 9370 9920
rect 9401 9911 9459 9917
rect 9401 9908 9413 9911
rect 9364 9880 9413 9908
rect 9364 9868 9370 9880
rect 9401 9877 9413 9880
rect 9447 9877 9459 9911
rect 9858 9908 9864 9920
rect 9819 9880 9864 9908
rect 9401 9871 9459 9877
rect 9858 9868 9864 9880
rect 9916 9868 9922 9920
rect 10226 9908 10232 9920
rect 10187 9880 10232 9908
rect 10226 9868 10232 9880
rect 10284 9868 10290 9920
rect 10870 9868 10876 9920
rect 10928 9908 10934 9920
rect 10965 9911 11023 9917
rect 10965 9908 10977 9911
rect 10928 9880 10977 9908
rect 10928 9868 10934 9880
rect 10965 9877 10977 9880
rect 11011 9877 11023 9911
rect 10965 9871 11023 9877
rect 11422 9868 11428 9920
rect 11480 9908 11486 9920
rect 11517 9911 11575 9917
rect 11517 9908 11529 9911
rect 11480 9880 11529 9908
rect 11480 9868 11486 9880
rect 11517 9877 11529 9880
rect 11563 9877 11575 9911
rect 11517 9871 11575 9877
rect 11698 9868 11704 9920
rect 11756 9908 11762 9920
rect 11793 9911 11851 9917
rect 11793 9908 11805 9911
rect 11756 9880 11805 9908
rect 11756 9868 11762 9880
rect 11793 9877 11805 9880
rect 11839 9877 11851 9911
rect 11793 9871 11851 9877
rect 12897 9911 12955 9917
rect 12897 9877 12909 9911
rect 12943 9908 12955 9911
rect 13078 9908 13084 9920
rect 12943 9880 13084 9908
rect 12943 9877 12955 9880
rect 12897 9871 12955 9877
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 1104 9818 16008 9840
rect 1104 9766 4698 9818
rect 4750 9766 4762 9818
rect 4814 9766 4826 9818
rect 4878 9766 4890 9818
rect 4942 9766 4954 9818
rect 5006 9766 8446 9818
rect 8498 9766 8510 9818
rect 8562 9766 8574 9818
rect 8626 9766 8638 9818
rect 8690 9766 8702 9818
rect 8754 9766 12194 9818
rect 12246 9766 12258 9818
rect 12310 9766 12322 9818
rect 12374 9766 12386 9818
rect 12438 9766 12450 9818
rect 12502 9766 16008 9818
rect 1104 9744 16008 9766
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 6365 9707 6423 9713
rect 6365 9704 6377 9707
rect 5868 9676 6377 9704
rect 5868 9664 5874 9676
rect 6365 9673 6377 9676
rect 6411 9673 6423 9707
rect 6365 9667 6423 9673
rect 8573 9707 8631 9713
rect 8573 9673 8585 9707
rect 8619 9704 8631 9707
rect 8662 9704 8668 9716
rect 8619 9676 8668 9704
rect 8619 9673 8631 9676
rect 8573 9667 8631 9673
rect 8662 9664 8668 9676
rect 8720 9704 8726 9716
rect 9490 9704 9496 9716
rect 8720 9676 9496 9704
rect 8720 9664 8726 9676
rect 9490 9664 9496 9676
rect 9548 9664 9554 9716
rect 10781 9707 10839 9713
rect 10781 9673 10793 9707
rect 10827 9673 10839 9707
rect 10781 9667 10839 9673
rect 1397 9639 1455 9645
rect 1397 9605 1409 9639
rect 1443 9636 1455 9639
rect 1486 9636 1492 9648
rect 1443 9608 1492 9636
rect 1443 9605 1455 9608
rect 1397 9599 1455 9605
rect 1486 9596 1492 9608
rect 1544 9596 1550 9648
rect 3053 9639 3111 9645
rect 3053 9605 3065 9639
rect 3099 9636 3111 9639
rect 3510 9636 3516 9648
rect 3099 9608 3516 9636
rect 3099 9605 3111 9608
rect 3053 9599 3111 9605
rect 3510 9596 3516 9608
rect 3568 9596 3574 9648
rect 6825 9639 6883 9645
rect 6825 9605 6837 9639
rect 6871 9636 6883 9639
rect 8938 9636 8944 9648
rect 6871 9608 8944 9636
rect 6871 9605 6883 9608
rect 6825 9599 6883 9605
rect 8938 9596 8944 9608
rect 8996 9596 9002 9648
rect 10796 9636 10824 9667
rect 11514 9664 11520 9716
rect 11572 9704 11578 9716
rect 13722 9704 13728 9716
rect 11572 9676 13728 9704
rect 11572 9664 11578 9676
rect 13722 9664 13728 9676
rect 13780 9664 13786 9716
rect 9324 9608 10824 9636
rect 5350 9568 5356 9580
rect 5311 9540 5356 9568
rect 5350 9528 5356 9540
rect 5408 9528 5414 9580
rect 5905 9571 5963 9577
rect 5905 9537 5917 9571
rect 5951 9568 5963 9571
rect 6086 9568 6092 9580
rect 5951 9540 6092 9568
rect 5951 9537 5963 9540
rect 5905 9531 5963 9537
rect 6086 9528 6092 9540
rect 6144 9528 6150 9580
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9537 6239 9571
rect 6181 9531 6239 9537
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9568 6791 9571
rect 7006 9568 7012 9580
rect 6779 9540 7012 9568
rect 6779 9537 6791 9540
rect 6733 9531 6791 9537
rect 3237 9503 3295 9509
rect 3237 9469 3249 9503
rect 3283 9500 3295 9503
rect 3418 9500 3424 9512
rect 3283 9472 3424 9500
rect 3283 9469 3295 9472
rect 3237 9463 3295 9469
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 2130 9392 2136 9444
rect 2188 9432 2194 9444
rect 5169 9435 5227 9441
rect 5169 9432 5181 9435
rect 2188 9404 5181 9432
rect 2188 9392 2194 9404
rect 5169 9401 5181 9404
rect 5215 9401 5227 9435
rect 6196 9432 6224 9531
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 7098 9528 7104 9580
rect 7156 9568 7162 9580
rect 7449 9571 7507 9577
rect 7449 9568 7461 9571
rect 7156 9540 7461 9568
rect 7156 9528 7162 9540
rect 7449 9537 7461 9540
rect 7495 9568 7507 9571
rect 8680 9568 8800 9572
rect 7495 9544 8800 9568
rect 7495 9540 8708 9544
rect 7495 9537 7507 9540
rect 7449 9531 7507 9537
rect 6914 9500 6920 9512
rect 6875 9472 6920 9500
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 7193 9503 7251 9509
rect 7193 9469 7205 9503
rect 7239 9469 7251 9503
rect 7193 9463 7251 9469
rect 7098 9432 7104 9444
rect 6196 9404 7104 9432
rect 5169 9395 5227 9401
rect 7098 9392 7104 9404
rect 7156 9392 7162 9444
rect 5718 9364 5724 9376
rect 5679 9336 5724 9364
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 5994 9364 6000 9376
rect 5955 9336 6000 9364
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 7208 9364 7236 9463
rect 8294 9460 8300 9512
rect 8352 9500 8358 9512
rect 8570 9500 8576 9512
rect 8352 9472 8576 9500
rect 8352 9460 8358 9472
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 8772 9509 8800 9544
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9568 9091 9571
rect 9214 9568 9220 9580
rect 9079 9540 9220 9568
rect 9079 9537 9091 9540
rect 9033 9531 9091 9537
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 8757 9503 8815 9509
rect 8757 9469 8769 9503
rect 8803 9469 8815 9503
rect 8757 9463 8815 9469
rect 8938 9460 8944 9512
rect 8996 9500 9002 9512
rect 8996 9472 9041 9500
rect 8996 9460 9002 9472
rect 8202 9392 8208 9444
rect 8260 9432 8266 9444
rect 9324 9432 9352 9608
rect 9582 9568 9588 9580
rect 9416 9540 9588 9568
rect 9416 9441 9444 9540
rect 9582 9528 9588 9540
rect 9640 9528 9646 9580
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 10229 9571 10287 9577
rect 10229 9537 10241 9571
rect 10275 9568 10287 9571
rect 10965 9571 11023 9577
rect 10275 9540 10916 9568
rect 10275 9537 10287 9540
rect 10229 9531 10287 9537
rect 9784 9500 9812 9531
rect 10778 9500 10784 9512
rect 9784 9472 10784 9500
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 10888 9500 10916 9540
rect 10965 9537 10977 9571
rect 11011 9568 11023 9571
rect 11882 9568 11888 9580
rect 11011 9540 11888 9568
rect 11011 9537 11023 9540
rect 10965 9531 11023 9537
rect 11882 9528 11888 9540
rect 11940 9528 11946 9580
rect 11974 9500 11980 9512
rect 10888 9472 11980 9500
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 8260 9404 8800 9432
rect 8260 9392 8266 9404
rect 8294 9364 8300 9376
rect 7208 9336 8300 9364
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 8772 9364 8800 9404
rect 8956 9404 9352 9432
rect 9401 9435 9459 9441
rect 8956 9364 8984 9404
rect 9401 9401 9413 9435
rect 9447 9401 9459 9435
rect 9401 9395 9459 9401
rect 10045 9435 10103 9441
rect 10045 9401 10057 9435
rect 10091 9432 10103 9435
rect 10226 9432 10232 9444
rect 10091 9404 10232 9432
rect 10091 9401 10103 9404
rect 10045 9395 10103 9401
rect 10226 9392 10232 9404
rect 10284 9392 10290 9444
rect 8772 9336 8984 9364
rect 9030 9324 9036 9376
rect 9088 9364 9094 9376
rect 9214 9364 9220 9376
rect 9088 9336 9220 9364
rect 9088 9324 9094 9336
rect 9214 9324 9220 9336
rect 9272 9324 9278 9376
rect 9582 9364 9588 9376
rect 9543 9336 9588 9364
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 1104 9274 16008 9296
rect 1104 9222 2824 9274
rect 2876 9222 2888 9274
rect 2940 9222 2952 9274
rect 3004 9222 3016 9274
rect 3068 9222 3080 9274
rect 3132 9222 6572 9274
rect 6624 9222 6636 9274
rect 6688 9222 6700 9274
rect 6752 9222 6764 9274
rect 6816 9222 6828 9274
rect 6880 9222 10320 9274
rect 10372 9222 10384 9274
rect 10436 9222 10448 9274
rect 10500 9222 10512 9274
rect 10564 9222 10576 9274
rect 10628 9222 14068 9274
rect 14120 9222 14132 9274
rect 14184 9222 14196 9274
rect 14248 9222 14260 9274
rect 14312 9222 14324 9274
rect 14376 9222 16008 9274
rect 1104 9200 16008 9222
rect 6914 9160 6920 9172
rect 6875 9132 6920 9160
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 9674 9160 9680 9172
rect 7156 9132 9680 9160
rect 7156 9120 7162 9132
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 8386 9092 8392 9104
rect 8347 9064 8392 9092
rect 8386 9052 8392 9064
rect 8444 9052 8450 9104
rect 8570 9052 8576 9104
rect 8628 9092 8634 9104
rect 8938 9092 8944 9104
rect 8628 9064 8944 9092
rect 8628 9052 8634 9064
rect 8938 9052 8944 9064
rect 8996 9052 9002 9104
rect 10134 9024 10140 9036
rect 8220 8996 10140 9024
rect 6086 8916 6092 8968
rect 6144 8956 6150 8968
rect 8220 8956 8248 8996
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 6144 8928 8248 8956
rect 6144 8916 6150 8928
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 8573 8959 8631 8965
rect 8352 8928 8397 8956
rect 8352 8916 8358 8928
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 9030 8956 9036 8968
rect 8619 8928 9036 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8956 9183 8959
rect 10686 8956 10692 8968
rect 9171 8928 10692 8956
rect 9171 8925 9183 8928
rect 9125 8919 9183 8925
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 8052 8891 8110 8897
rect 8052 8857 8064 8891
rect 8098 8888 8110 8891
rect 8478 8888 8484 8900
rect 8098 8860 8484 8888
rect 8098 8857 8110 8860
rect 8052 8851 8110 8857
rect 8478 8848 8484 8860
rect 8536 8848 8542 8900
rect 9582 8888 9588 8900
rect 8772 8860 9588 8888
rect 6178 8780 6184 8832
rect 6236 8820 6242 8832
rect 8772 8820 8800 8860
rect 9582 8848 9588 8860
rect 9640 8848 9646 8900
rect 9766 8848 9772 8900
rect 9824 8888 9830 8900
rect 12618 8888 12624 8900
rect 9824 8860 12624 8888
rect 9824 8848 9830 8860
rect 12618 8848 12624 8860
rect 12676 8848 12682 8900
rect 8938 8820 8944 8832
rect 6236 8792 8800 8820
rect 8899 8792 8944 8820
rect 6236 8780 6242 8792
rect 8938 8780 8944 8792
rect 8996 8780 9002 8832
rect 1104 8730 16008 8752
rect 1104 8678 4698 8730
rect 4750 8678 4762 8730
rect 4814 8678 4826 8730
rect 4878 8678 4890 8730
rect 4942 8678 4954 8730
rect 5006 8678 8446 8730
rect 8498 8678 8510 8730
rect 8562 8678 8574 8730
rect 8626 8678 8638 8730
rect 8690 8678 8702 8730
rect 8754 8678 12194 8730
rect 12246 8678 12258 8730
rect 12310 8678 12322 8730
rect 12374 8678 12386 8730
rect 12438 8678 12450 8730
rect 12502 8678 16008 8730
rect 1104 8656 16008 8678
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 7101 8619 7159 8625
rect 7101 8616 7113 8619
rect 5592 8588 7113 8616
rect 5592 8576 5598 8588
rect 7101 8585 7113 8588
rect 7147 8585 7159 8619
rect 7101 8579 7159 8585
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 7515 8588 8033 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 8021 8585 8033 8588
rect 8067 8585 8079 8619
rect 8021 8579 8079 8585
rect 8481 8619 8539 8625
rect 8481 8585 8493 8619
rect 8527 8616 8539 8619
rect 8846 8616 8852 8628
rect 8527 8588 8852 8616
rect 8527 8585 8539 8588
rect 8481 8579 8539 8585
rect 8846 8576 8852 8588
rect 8904 8576 8910 8628
rect 8294 8508 8300 8560
rect 8352 8548 8358 8560
rect 11146 8548 11152 8560
rect 8352 8520 11152 8548
rect 8352 8508 8358 8520
rect 11146 8508 11152 8520
rect 11204 8548 11210 8560
rect 11701 8551 11759 8557
rect 11701 8548 11713 8551
rect 11204 8520 11713 8548
rect 11204 8508 11210 8520
rect 11701 8517 11713 8520
rect 11747 8517 11759 8551
rect 11701 8511 11759 8517
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 3510 8480 3516 8492
rect 1719 8452 3516 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 6914 8440 6920 8492
rect 6972 8480 6978 8492
rect 8386 8480 8392 8492
rect 6972 8452 7696 8480
rect 8347 8452 8392 8480
rect 6972 8440 6978 8452
rect 7668 8421 7696 8452
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 9858 8480 9864 8492
rect 8496 8452 9864 8480
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8381 7619 8415
rect 7561 8375 7619 8381
rect 7653 8415 7711 8421
rect 7653 8381 7665 8415
rect 7699 8381 7711 8415
rect 8496 8412 8524 8452
rect 9858 8440 9864 8452
rect 9916 8440 9922 8492
rect 12529 8483 12587 8489
rect 12529 8449 12541 8483
rect 12575 8480 12587 8483
rect 12575 8452 12756 8480
rect 12575 8449 12587 8452
rect 12529 8443 12587 8449
rect 7653 8375 7711 8381
rect 7760 8384 8524 8412
rect 8665 8415 8723 8421
rect 1486 8344 1492 8356
rect 1447 8316 1492 8344
rect 1486 8304 1492 8316
rect 1544 8304 1550 8356
rect 7576 8344 7604 8375
rect 7760 8344 7788 8384
rect 8665 8381 8677 8415
rect 8711 8412 8723 8415
rect 9490 8412 9496 8424
rect 8711 8384 9496 8412
rect 8711 8381 8723 8384
rect 8665 8375 8723 8381
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 12728 8356 12756 8452
rect 7576 8316 7788 8344
rect 8294 8304 8300 8356
rect 8352 8344 8358 8356
rect 8938 8344 8944 8356
rect 8352 8316 8944 8344
rect 8352 8304 8358 8316
rect 8938 8304 8944 8316
rect 8996 8304 9002 8356
rect 9766 8344 9772 8356
rect 9048 8316 9772 8344
rect 8386 8236 8392 8288
rect 8444 8276 8450 8288
rect 9048 8276 9076 8316
rect 9766 8304 9772 8316
rect 9824 8304 9830 8356
rect 12710 8344 12716 8356
rect 12671 8316 12716 8344
rect 12710 8304 12716 8316
rect 12768 8304 12774 8356
rect 8444 8248 9076 8276
rect 8444 8236 8450 8248
rect 1104 8186 16008 8208
rect 1104 8134 2824 8186
rect 2876 8134 2888 8186
rect 2940 8134 2952 8186
rect 3004 8134 3016 8186
rect 3068 8134 3080 8186
rect 3132 8134 6572 8186
rect 6624 8134 6636 8186
rect 6688 8134 6700 8186
rect 6752 8134 6764 8186
rect 6816 8134 6828 8186
rect 6880 8134 10320 8186
rect 10372 8134 10384 8186
rect 10436 8134 10448 8186
rect 10500 8134 10512 8186
rect 10564 8134 10576 8186
rect 10628 8134 14068 8186
rect 14120 8134 14132 8186
rect 14184 8134 14196 8186
rect 14248 8134 14260 8186
rect 14312 8134 14324 8186
rect 14376 8134 16008 8186
rect 1104 8112 16008 8134
rect 1104 7642 16008 7664
rect 1104 7590 4698 7642
rect 4750 7590 4762 7642
rect 4814 7590 4826 7642
rect 4878 7590 4890 7642
rect 4942 7590 4954 7642
rect 5006 7590 8446 7642
rect 8498 7590 8510 7642
rect 8562 7590 8574 7642
rect 8626 7590 8638 7642
rect 8690 7590 8702 7642
rect 8754 7590 12194 7642
rect 12246 7590 12258 7642
rect 12310 7590 12322 7642
rect 12374 7590 12386 7642
rect 12438 7590 12450 7642
rect 12502 7590 16008 7642
rect 1104 7568 16008 7590
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 5629 7531 5687 7537
rect 5629 7528 5641 7531
rect 4212 7500 5641 7528
rect 4212 7488 4218 7500
rect 5629 7497 5641 7500
rect 5675 7497 5687 7531
rect 7466 7528 7472 7540
rect 5629 7491 5687 7497
rect 5736 7500 7472 7528
rect 5736 7460 5764 7500
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 4724 7432 5764 7460
rect 3234 7392 3240 7404
rect 3195 7364 3240 7392
rect 3234 7352 3240 7364
rect 3292 7352 3298 7404
rect 4724 7401 4752 7432
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7361 4767 7395
rect 4709 7355 4767 7361
rect 5261 7395 5319 7401
rect 5261 7361 5273 7395
rect 5307 7361 5319 7395
rect 5261 7355 5319 7361
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 7282 7392 7288 7404
rect 5859 7364 7288 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 5276 7324 5304 7355
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7558 7392 7564 7404
rect 7519 7364 7564 7392
rect 7558 7352 7564 7364
rect 7616 7352 7622 7404
rect 9398 7392 9404 7404
rect 9359 7364 9404 7392
rect 9398 7352 9404 7364
rect 9456 7352 9462 7404
rect 8846 7324 8852 7336
rect 5276 7296 8852 7324
rect 8846 7284 8852 7296
rect 8904 7284 8910 7336
rect 5166 7216 5172 7268
rect 5224 7256 5230 7268
rect 7377 7259 7435 7265
rect 7377 7256 7389 7259
rect 5224 7228 7389 7256
rect 5224 7216 5230 7228
rect 7377 7225 7389 7228
rect 7423 7225 7435 7259
rect 7377 7219 7435 7225
rect 3053 7191 3111 7197
rect 3053 7157 3065 7191
rect 3099 7188 3111 7191
rect 3142 7188 3148 7200
rect 3099 7160 3148 7188
rect 3099 7157 3111 7160
rect 3053 7151 3111 7157
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 3326 7148 3332 7200
rect 3384 7188 3390 7200
rect 4525 7191 4583 7197
rect 4525 7188 4537 7191
rect 3384 7160 4537 7188
rect 3384 7148 3390 7160
rect 4525 7157 4537 7160
rect 4571 7157 4583 7191
rect 4525 7151 4583 7157
rect 4614 7148 4620 7200
rect 4672 7188 4678 7200
rect 5077 7191 5135 7197
rect 5077 7188 5089 7191
rect 4672 7160 5089 7188
rect 4672 7148 4678 7160
rect 5077 7157 5089 7160
rect 5123 7157 5135 7191
rect 5077 7151 5135 7157
rect 7650 7148 7656 7200
rect 7708 7188 7714 7200
rect 9217 7191 9275 7197
rect 9217 7188 9229 7191
rect 7708 7160 9229 7188
rect 7708 7148 7714 7160
rect 9217 7157 9229 7160
rect 9263 7157 9275 7191
rect 9217 7151 9275 7157
rect 1104 7098 16008 7120
rect 1104 7046 2824 7098
rect 2876 7046 2888 7098
rect 2940 7046 2952 7098
rect 3004 7046 3016 7098
rect 3068 7046 3080 7098
rect 3132 7046 6572 7098
rect 6624 7046 6636 7098
rect 6688 7046 6700 7098
rect 6752 7046 6764 7098
rect 6816 7046 6828 7098
rect 6880 7046 10320 7098
rect 10372 7046 10384 7098
rect 10436 7046 10448 7098
rect 10500 7046 10512 7098
rect 10564 7046 10576 7098
rect 10628 7046 14068 7098
rect 14120 7046 14132 7098
rect 14184 7046 14196 7098
rect 14248 7046 14260 7098
rect 14312 7046 14324 7098
rect 14376 7046 16008 7098
rect 1104 7024 16008 7046
rect 1104 6554 16008 6576
rect 1104 6502 4698 6554
rect 4750 6502 4762 6554
rect 4814 6502 4826 6554
rect 4878 6502 4890 6554
rect 4942 6502 4954 6554
rect 5006 6502 8446 6554
rect 8498 6502 8510 6554
rect 8562 6502 8574 6554
rect 8626 6502 8638 6554
rect 8690 6502 8702 6554
rect 8754 6502 12194 6554
rect 12246 6502 12258 6554
rect 12310 6502 12322 6554
rect 12374 6502 12386 6554
rect 12438 6502 12450 6554
rect 12502 6502 16008 6554
rect 1104 6480 16008 6502
rect 1104 6010 16008 6032
rect 1104 5958 2824 6010
rect 2876 5958 2888 6010
rect 2940 5958 2952 6010
rect 3004 5958 3016 6010
rect 3068 5958 3080 6010
rect 3132 5958 6572 6010
rect 6624 5958 6636 6010
rect 6688 5958 6700 6010
rect 6752 5958 6764 6010
rect 6816 5958 6828 6010
rect 6880 5958 10320 6010
rect 10372 5958 10384 6010
rect 10436 5958 10448 6010
rect 10500 5958 10512 6010
rect 10564 5958 10576 6010
rect 10628 5958 14068 6010
rect 14120 5958 14132 6010
rect 14184 5958 14196 6010
rect 14248 5958 14260 6010
rect 14312 5958 14324 6010
rect 14376 5958 16008 6010
rect 1104 5936 16008 5958
rect 1104 5466 16008 5488
rect 1104 5414 4698 5466
rect 4750 5414 4762 5466
rect 4814 5414 4826 5466
rect 4878 5414 4890 5466
rect 4942 5414 4954 5466
rect 5006 5414 8446 5466
rect 8498 5414 8510 5466
rect 8562 5414 8574 5466
rect 8626 5414 8638 5466
rect 8690 5414 8702 5466
rect 8754 5414 12194 5466
rect 12246 5414 12258 5466
rect 12310 5414 12322 5466
rect 12374 5414 12386 5466
rect 12438 5414 12450 5466
rect 12502 5414 16008 5466
rect 1104 5392 16008 5414
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 3142 5216 3148 5228
rect 1719 5188 3148 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 1486 5080 1492 5092
rect 1447 5052 1492 5080
rect 1486 5040 1492 5052
rect 1544 5040 1550 5092
rect 1104 4922 16008 4944
rect 1104 4870 2824 4922
rect 2876 4870 2888 4922
rect 2940 4870 2952 4922
rect 3004 4870 3016 4922
rect 3068 4870 3080 4922
rect 3132 4870 6572 4922
rect 6624 4870 6636 4922
rect 6688 4870 6700 4922
rect 6752 4870 6764 4922
rect 6816 4870 6828 4922
rect 6880 4870 10320 4922
rect 10372 4870 10384 4922
rect 10436 4870 10448 4922
rect 10500 4870 10512 4922
rect 10564 4870 10576 4922
rect 10628 4870 14068 4922
rect 14120 4870 14132 4922
rect 14184 4870 14196 4922
rect 14248 4870 14260 4922
rect 14312 4870 14324 4922
rect 14376 4870 16008 4922
rect 1104 4848 16008 4870
rect 1104 4378 16008 4400
rect 1104 4326 4698 4378
rect 4750 4326 4762 4378
rect 4814 4326 4826 4378
rect 4878 4326 4890 4378
rect 4942 4326 4954 4378
rect 5006 4326 8446 4378
rect 8498 4326 8510 4378
rect 8562 4326 8574 4378
rect 8626 4326 8638 4378
rect 8690 4326 8702 4378
rect 8754 4326 12194 4378
rect 12246 4326 12258 4378
rect 12310 4326 12322 4378
rect 12374 4326 12386 4378
rect 12438 4326 12450 4378
rect 12502 4326 16008 4378
rect 1104 4304 16008 4326
rect 7742 4088 7748 4140
rect 7800 4128 7806 4140
rect 12710 4128 12716 4140
rect 7800 4100 12716 4128
rect 7800 4088 7806 4100
rect 12710 4088 12716 4100
rect 12768 4088 12774 4140
rect 9214 4020 9220 4072
rect 9272 4060 9278 4072
rect 10134 4060 10140 4072
rect 9272 4032 10140 4060
rect 9272 4020 9278 4032
rect 10134 4020 10140 4032
rect 10192 4020 10198 4072
rect 6362 3952 6368 4004
rect 6420 3992 6426 4004
rect 9766 3992 9772 4004
rect 6420 3964 9772 3992
rect 6420 3952 6426 3964
rect 9766 3952 9772 3964
rect 9824 3952 9830 4004
rect 1104 3834 16008 3856
rect 1104 3782 2824 3834
rect 2876 3782 2888 3834
rect 2940 3782 2952 3834
rect 3004 3782 3016 3834
rect 3068 3782 3080 3834
rect 3132 3782 6572 3834
rect 6624 3782 6636 3834
rect 6688 3782 6700 3834
rect 6752 3782 6764 3834
rect 6816 3782 6828 3834
rect 6880 3782 10320 3834
rect 10372 3782 10384 3834
rect 10436 3782 10448 3834
rect 10500 3782 10512 3834
rect 10564 3782 10576 3834
rect 10628 3782 14068 3834
rect 14120 3782 14132 3834
rect 14184 3782 14196 3834
rect 14248 3782 14260 3834
rect 14312 3782 14324 3834
rect 14376 3782 16008 3834
rect 1104 3760 16008 3782
rect 1104 3290 16008 3312
rect 1104 3238 4698 3290
rect 4750 3238 4762 3290
rect 4814 3238 4826 3290
rect 4878 3238 4890 3290
rect 4942 3238 4954 3290
rect 5006 3238 8446 3290
rect 8498 3238 8510 3290
rect 8562 3238 8574 3290
rect 8626 3238 8638 3290
rect 8690 3238 8702 3290
rect 8754 3238 12194 3290
rect 12246 3238 12258 3290
rect 12310 3238 12322 3290
rect 12374 3238 12386 3290
rect 12438 3238 12450 3290
rect 12502 3238 16008 3290
rect 1104 3216 16008 3238
rect 2041 3179 2099 3185
rect 2041 3145 2053 3179
rect 2087 3176 2099 3179
rect 3418 3176 3424 3188
rect 2087 3148 3424 3176
rect 2087 3145 2099 3148
rect 2041 3139 2099 3145
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 8754 3136 8760 3188
rect 8812 3176 8818 3188
rect 13078 3176 13084 3188
rect 8812 3148 13084 3176
rect 8812 3136 8818 3148
rect 13078 3136 13084 3148
rect 13136 3136 13142 3188
rect 13354 3136 13360 3188
rect 13412 3176 13418 3188
rect 15473 3179 15531 3185
rect 15473 3176 15485 3179
rect 13412 3148 15485 3176
rect 13412 3136 13418 3148
rect 15473 3145 15485 3148
rect 15519 3145 15531 3179
rect 15473 3139 15531 3145
rect 3326 3108 3332 3120
rect 1780 3080 3332 3108
rect 1780 3049 1808 3080
rect 3326 3068 3332 3080
rect 3384 3068 3390 3120
rect 1765 3043 1823 3049
rect 1765 3009 1777 3043
rect 1811 3009 1823 3043
rect 1765 3003 1823 3009
rect 1854 3000 1860 3052
rect 1912 3040 1918 3052
rect 2133 3043 2191 3049
rect 2133 3040 2145 3043
rect 1912 3012 2145 3040
rect 1912 3000 1918 3012
rect 2133 3009 2145 3012
rect 2179 3009 2191 3043
rect 2133 3003 2191 3009
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3040 4399 3043
rect 6454 3040 6460 3052
rect 4387 3012 6460 3040
rect 4387 3009 4399 3012
rect 4341 3003 4399 3009
rect 6454 3000 6460 3012
rect 6512 3000 6518 3052
rect 15381 3043 15439 3049
rect 15381 3009 15393 3043
rect 15427 3040 15439 3043
rect 15657 3043 15715 3049
rect 15657 3040 15669 3043
rect 15427 3012 15669 3040
rect 15427 3009 15439 3012
rect 15381 3003 15439 3009
rect 15657 3009 15669 3012
rect 15703 3040 15715 3043
rect 15746 3040 15752 3052
rect 15703 3012 15752 3040
rect 15703 3009 15715 3012
rect 15657 3003 15715 3009
rect 15746 3000 15752 3012
rect 15804 3000 15810 3052
rect 8662 2932 8668 2984
rect 8720 2972 8726 2984
rect 10870 2972 10876 2984
rect 8720 2944 10876 2972
rect 8720 2932 8726 2944
rect 10870 2932 10876 2944
rect 10928 2932 10934 2984
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 1452 2808 1593 2836
rect 1452 2796 1458 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 3970 2796 3976 2848
rect 4028 2836 4034 2848
rect 4157 2839 4215 2845
rect 4157 2836 4169 2839
rect 4028 2808 4169 2836
rect 4028 2796 4034 2808
rect 4157 2805 4169 2808
rect 4203 2805 4215 2839
rect 8846 2836 8852 2848
rect 8807 2808 8852 2836
rect 4157 2799 4215 2805
rect 8846 2796 8852 2808
rect 8904 2796 8910 2848
rect 9122 2836 9128 2848
rect 9083 2808 9128 2836
rect 9122 2796 9128 2808
rect 9180 2796 9186 2848
rect 9490 2836 9496 2848
rect 9451 2808 9496 2836
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 9858 2836 9864 2848
rect 9819 2808 9864 2836
rect 9858 2796 9864 2808
rect 9916 2796 9922 2848
rect 10226 2836 10232 2848
rect 10187 2808 10232 2836
rect 10226 2796 10232 2808
rect 10284 2796 10290 2848
rect 10597 2839 10655 2845
rect 10597 2805 10609 2839
rect 10643 2836 10655 2839
rect 10686 2836 10692 2848
rect 10643 2808 10692 2836
rect 10643 2805 10655 2808
rect 10597 2799 10655 2805
rect 10686 2796 10692 2808
rect 10744 2796 10750 2848
rect 10962 2836 10968 2848
rect 10923 2808 10968 2836
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 11330 2796 11336 2848
rect 11388 2836 11394 2848
rect 11517 2839 11575 2845
rect 11517 2836 11529 2839
rect 11388 2808 11529 2836
rect 11388 2796 11394 2808
rect 11517 2805 11529 2808
rect 11563 2805 11575 2839
rect 11790 2836 11796 2848
rect 11751 2808 11796 2836
rect 11517 2799 11575 2805
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 12066 2836 12072 2848
rect 12027 2808 12072 2836
rect 12066 2796 12072 2808
rect 12124 2796 12130 2848
rect 12437 2839 12495 2845
rect 12437 2805 12449 2839
rect 12483 2836 12495 2839
rect 12526 2836 12532 2848
rect 12483 2808 12532 2836
rect 12483 2805 12495 2808
rect 12437 2799 12495 2805
rect 12526 2796 12532 2808
rect 12584 2796 12590 2848
rect 12802 2836 12808 2848
rect 12763 2808 12808 2836
rect 12802 2796 12808 2808
rect 12860 2796 12866 2848
rect 13170 2836 13176 2848
rect 13131 2808 13176 2836
rect 13170 2796 13176 2808
rect 13228 2796 13234 2848
rect 13541 2839 13599 2845
rect 13541 2805 13553 2839
rect 13587 2836 13599 2839
rect 13814 2836 13820 2848
rect 13587 2808 13820 2836
rect 13587 2805 13599 2808
rect 13541 2799 13599 2805
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 14277 2839 14335 2845
rect 13964 2808 14009 2836
rect 13964 2796 13970 2808
rect 14277 2805 14289 2839
rect 14323 2836 14335 2839
rect 14458 2836 14464 2848
rect 14323 2808 14464 2836
rect 14323 2805 14335 2808
rect 14277 2799 14335 2805
rect 14458 2796 14464 2808
rect 14516 2796 14522 2848
rect 14642 2836 14648 2848
rect 14603 2808 14648 2836
rect 14642 2796 14648 2808
rect 14700 2796 14706 2848
rect 15010 2836 15016 2848
rect 14971 2808 15016 2836
rect 15010 2796 15016 2808
rect 15068 2796 15074 2848
rect 15197 2839 15255 2845
rect 15197 2805 15209 2839
rect 15243 2836 15255 2839
rect 15378 2836 15384 2848
rect 15243 2808 15384 2836
rect 15243 2805 15255 2808
rect 15197 2799 15255 2805
rect 15378 2796 15384 2808
rect 15436 2796 15442 2848
rect 1104 2746 16008 2768
rect 1104 2694 2824 2746
rect 2876 2694 2888 2746
rect 2940 2694 2952 2746
rect 3004 2694 3016 2746
rect 3068 2694 3080 2746
rect 3132 2694 6572 2746
rect 6624 2694 6636 2746
rect 6688 2694 6700 2746
rect 6752 2694 6764 2746
rect 6816 2694 6828 2746
rect 6880 2694 10320 2746
rect 10372 2694 10384 2746
rect 10436 2694 10448 2746
rect 10500 2694 10512 2746
rect 10564 2694 10576 2746
rect 10628 2694 14068 2746
rect 14120 2694 14132 2746
rect 14184 2694 14196 2746
rect 14248 2694 14260 2746
rect 14312 2694 14324 2746
rect 14376 2694 16008 2746
rect 1104 2672 16008 2694
rect 4614 2632 4620 2644
rect 2148 2604 4620 2632
rect 2148 2437 2176 2604
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 7248 2604 8953 2632
rect 7248 2592 7254 2604
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 9582 2632 9588 2644
rect 9543 2604 9588 2632
rect 8941 2595 8999 2601
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 9766 2592 9772 2644
rect 9824 2632 9830 2644
rect 9953 2635 10011 2641
rect 9953 2632 9965 2635
rect 9824 2604 9965 2632
rect 9824 2592 9830 2604
rect 9953 2601 9965 2604
rect 9999 2601 10011 2635
rect 9953 2595 10011 2601
rect 10134 2592 10140 2644
rect 10192 2632 10198 2644
rect 10321 2635 10379 2641
rect 10321 2632 10333 2635
rect 10192 2604 10333 2632
rect 10192 2592 10198 2604
rect 10321 2601 10333 2604
rect 10367 2601 10379 2635
rect 10321 2595 10379 2601
rect 11514 2592 11520 2644
rect 11572 2632 11578 2644
rect 11793 2635 11851 2641
rect 11793 2632 11805 2635
rect 11572 2604 11805 2632
rect 11572 2592 11578 2604
rect 11793 2601 11805 2604
rect 11839 2601 11851 2635
rect 11793 2595 11851 2601
rect 12529 2635 12587 2641
rect 12529 2601 12541 2635
rect 12575 2632 12587 2635
rect 12618 2632 12624 2644
rect 12575 2604 12624 2632
rect 12575 2601 12587 2604
rect 12529 2595 12587 2601
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 12894 2632 12900 2644
rect 12855 2604 12900 2632
rect 12894 2592 12900 2604
rect 12952 2592 12958 2644
rect 12986 2592 12992 2644
rect 13044 2632 13050 2644
rect 15473 2635 15531 2641
rect 15473 2632 15485 2635
rect 13044 2604 13768 2632
rect 13044 2592 13050 2604
rect 3694 2564 3700 2576
rect 2424 2536 3700 2564
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2397 2191 2431
rect 2133 2391 2191 2397
rect 1780 2360 1808 2391
rect 2424 2360 2452 2536
rect 3694 2524 3700 2536
rect 3752 2524 3758 2576
rect 8294 2564 8300 2576
rect 4724 2536 8300 2564
rect 4154 2496 4160 2508
rect 2884 2468 4160 2496
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2428 2559 2431
rect 2774 2428 2780 2440
rect 2547 2400 2780 2428
rect 2547 2397 2559 2400
rect 2501 2391 2559 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 2884 2437 2912 2468
rect 4154 2456 4160 2468
rect 4212 2456 4218 2508
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2428 3295 2431
rect 3510 2428 3516 2440
rect 3283 2400 3516 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2397 3663 2431
rect 4338 2428 4344 2440
rect 4299 2400 4344 2428
rect 3605 2391 3663 2397
rect 1780 2332 2452 2360
rect 3620 2360 3648 2391
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 4724 2437 4752 2536
rect 8294 2524 8300 2536
rect 8352 2524 8358 2576
rect 11698 2564 11704 2576
rect 8404 2536 11704 2564
rect 8404 2496 8432 2536
rect 11698 2524 11704 2536
rect 11756 2524 11762 2576
rect 11974 2524 11980 2576
rect 12032 2564 12038 2576
rect 13633 2567 13691 2573
rect 13633 2564 13645 2567
rect 12032 2536 13645 2564
rect 12032 2524 12038 2536
rect 13633 2533 13645 2536
rect 13679 2533 13691 2567
rect 13740 2564 13768 2604
rect 14200 2604 15485 2632
rect 14200 2564 14228 2604
rect 15473 2601 15485 2604
rect 15519 2601 15531 2635
rect 15473 2595 15531 2601
rect 13740 2536 14228 2564
rect 14369 2567 14427 2573
rect 13633 2527 13691 2533
rect 14369 2533 14381 2567
rect 14415 2533 14427 2567
rect 14369 2527 14427 2533
rect 11606 2496 11612 2508
rect 8312 2468 8432 2496
rect 8680 2468 11612 2496
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 5077 2431 5135 2437
rect 5077 2397 5089 2431
rect 5123 2428 5135 2431
rect 5166 2428 5172 2440
rect 5123 2400 5172 2428
rect 5123 2397 5135 2400
rect 5077 2391 5135 2397
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 5442 2428 5448 2440
rect 5403 2400 5448 2428
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 5810 2428 5816 2440
rect 5771 2400 5816 2428
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 6181 2431 6239 2437
rect 6181 2397 6193 2431
rect 6227 2428 6239 2431
rect 6454 2428 6460 2440
rect 6227 2400 6460 2428
rect 6227 2397 6239 2400
rect 6181 2391 6239 2397
rect 6454 2388 6460 2400
rect 6512 2388 6518 2440
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2428 7343 2431
rect 7466 2428 7472 2440
rect 7331 2400 7472 2428
rect 7331 2397 7343 2400
rect 7285 2391 7343 2397
rect 4982 2360 4988 2372
rect 3620 2332 4988 2360
rect 4982 2320 4988 2332
rect 5040 2320 5046 2372
rect 6932 2360 6960 2391
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 7650 2428 7656 2440
rect 7611 2400 7656 2428
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 8021 2431 8079 2437
rect 8021 2397 8033 2431
rect 8067 2428 8079 2431
rect 8312 2428 8340 2468
rect 8067 2400 8340 2428
rect 8389 2431 8447 2437
rect 8067 2397 8079 2400
rect 8021 2391 8079 2397
rect 8389 2397 8401 2431
rect 8435 2428 8447 2431
rect 8680 2428 8708 2468
rect 11606 2456 11612 2468
rect 11664 2456 11670 2508
rect 11882 2456 11888 2508
rect 11940 2496 11946 2508
rect 14384 2496 14412 2527
rect 11940 2468 14412 2496
rect 11940 2456 11946 2468
rect 8435 2400 8708 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 8754 2388 8760 2440
rect 8812 2428 8818 2440
rect 9125 2431 9183 2437
rect 8812 2400 8857 2428
rect 8812 2388 8818 2400
rect 9125 2397 9137 2431
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 8662 2360 8668 2372
rect 6932 2332 8668 2360
rect 8662 2320 8668 2332
rect 8720 2320 8726 2372
rect 8846 2320 8852 2372
rect 8904 2360 8910 2372
rect 9140 2360 9168 2391
rect 9214 2388 9220 2440
rect 9272 2428 9278 2440
rect 9401 2431 9459 2437
rect 9401 2428 9413 2431
rect 9272 2400 9413 2428
rect 9272 2388 9278 2400
rect 9401 2397 9413 2400
rect 9447 2397 9459 2431
rect 9401 2391 9459 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9732 2400 9781 2428
rect 9732 2388 9738 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 9858 2388 9864 2440
rect 9916 2428 9922 2440
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 9916 2400 10149 2428
rect 9916 2388 9922 2400
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 10137 2391 10195 2397
rect 10226 2388 10232 2440
rect 10284 2428 10290 2440
rect 10505 2431 10563 2437
rect 10505 2428 10517 2431
rect 10284 2400 10517 2428
rect 10284 2388 10290 2400
rect 10505 2397 10517 2400
rect 10551 2397 10563 2431
rect 10505 2391 10563 2397
rect 10594 2388 10600 2440
rect 10652 2428 10658 2440
rect 10873 2431 10931 2437
rect 10873 2428 10885 2431
rect 10652 2400 10885 2428
rect 10652 2388 10658 2400
rect 10873 2397 10885 2400
rect 10919 2397 10931 2431
rect 10873 2391 10931 2397
rect 11054 2388 11060 2440
rect 11112 2428 11118 2440
rect 11241 2431 11299 2437
rect 11241 2428 11253 2431
rect 11112 2400 11253 2428
rect 11112 2388 11118 2400
rect 11241 2397 11253 2400
rect 11287 2397 11299 2431
rect 11241 2391 11299 2397
rect 11330 2388 11336 2440
rect 11388 2428 11394 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11388 2400 11713 2428
rect 11388 2388 11394 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 11790 2388 11796 2440
rect 11848 2428 11854 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11848 2400 11989 2428
rect 11848 2388 11854 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 12066 2388 12072 2440
rect 12124 2428 12130 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 12124 2400 12357 2428
rect 12124 2388 12130 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 12526 2388 12532 2440
rect 12584 2428 12590 2440
rect 12713 2431 12771 2437
rect 12713 2428 12725 2431
rect 12584 2400 12725 2428
rect 12584 2388 12590 2400
rect 12713 2397 12725 2400
rect 12759 2397 12771 2431
rect 12713 2391 12771 2397
rect 12802 2388 12808 2440
rect 12860 2428 12866 2440
rect 13081 2431 13139 2437
rect 13081 2428 13093 2431
rect 12860 2400 13093 2428
rect 12860 2388 12866 2400
rect 13081 2397 13093 2400
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 13170 2388 13176 2440
rect 13228 2428 13234 2440
rect 13449 2431 13507 2437
rect 13449 2428 13461 2431
rect 13228 2400 13461 2428
rect 13228 2388 13234 2400
rect 13449 2397 13461 2400
rect 13495 2397 13507 2431
rect 13814 2428 13820 2440
rect 13775 2400 13820 2428
rect 13449 2391 13507 2397
rect 13814 2388 13820 2400
rect 13872 2388 13878 2440
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 13964 2400 14289 2428
rect 13964 2388 13970 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 14366 2388 14372 2440
rect 14424 2428 14430 2440
rect 14553 2431 14611 2437
rect 14553 2428 14565 2431
rect 14424 2400 14565 2428
rect 14424 2388 14430 2400
rect 14553 2397 14565 2400
rect 14599 2397 14611 2431
rect 14553 2391 14611 2397
rect 14642 2388 14648 2440
rect 14700 2428 14706 2440
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 14700 2400 14933 2428
rect 14700 2388 14706 2400
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 14921 2391 14979 2397
rect 15194 2388 15200 2440
rect 15252 2428 15258 2440
rect 15289 2431 15347 2437
rect 15289 2428 15301 2431
rect 15252 2400 15301 2428
rect 15252 2388 15258 2400
rect 15289 2397 15301 2400
rect 15335 2397 15347 2431
rect 15289 2391 15347 2397
rect 15378 2388 15384 2440
rect 15436 2428 15442 2440
rect 15657 2431 15715 2437
rect 15657 2428 15669 2431
rect 15436 2400 15669 2428
rect 15436 2388 15442 2400
rect 15657 2397 15669 2400
rect 15703 2397 15715 2431
rect 15657 2391 15715 2397
rect 8904 2332 9168 2360
rect 8904 2320 8910 2332
rect 10778 2320 10784 2372
rect 10836 2360 10842 2372
rect 10836 2332 13032 2360
rect 10836 2320 10842 2332
rect 1581 2295 1639 2301
rect 1581 2261 1593 2295
rect 1627 2292 1639 2295
rect 1762 2292 1768 2304
rect 1627 2264 1768 2292
rect 1627 2261 1639 2264
rect 1581 2255 1639 2261
rect 1762 2252 1768 2264
rect 1820 2252 1826 2304
rect 1949 2295 2007 2301
rect 1949 2261 1961 2295
rect 1995 2292 2007 2295
rect 2130 2292 2136 2304
rect 1995 2264 2136 2292
rect 1995 2261 2007 2264
rect 1949 2255 2007 2261
rect 2130 2252 2136 2264
rect 2188 2252 2194 2304
rect 2317 2295 2375 2301
rect 2317 2261 2329 2295
rect 2363 2292 2375 2295
rect 2498 2292 2504 2304
rect 2363 2264 2504 2292
rect 2363 2261 2375 2264
rect 2317 2255 2375 2261
rect 2498 2252 2504 2264
rect 2556 2252 2562 2304
rect 2685 2295 2743 2301
rect 2685 2261 2697 2295
rect 2731 2292 2743 2295
rect 2866 2292 2872 2304
rect 2731 2264 2872 2292
rect 2731 2261 2743 2264
rect 2685 2255 2743 2261
rect 2866 2252 2872 2264
rect 2924 2252 2930 2304
rect 3053 2295 3111 2301
rect 3053 2261 3065 2295
rect 3099 2292 3111 2295
rect 3234 2292 3240 2304
rect 3099 2264 3240 2292
rect 3099 2261 3111 2264
rect 3053 2255 3111 2261
rect 3234 2252 3240 2264
rect 3292 2252 3298 2304
rect 3421 2295 3479 2301
rect 3421 2261 3433 2295
rect 3467 2292 3479 2295
rect 3602 2292 3608 2304
rect 3467 2264 3608 2292
rect 3467 2261 3479 2264
rect 3421 2255 3479 2261
rect 3602 2252 3608 2264
rect 3660 2252 3666 2304
rect 4157 2295 4215 2301
rect 4157 2261 4169 2295
rect 4203 2292 4215 2295
rect 4338 2292 4344 2304
rect 4203 2264 4344 2292
rect 4203 2261 4215 2264
rect 4157 2255 4215 2261
rect 4338 2252 4344 2264
rect 4396 2252 4402 2304
rect 4525 2295 4583 2301
rect 4525 2261 4537 2295
rect 4571 2292 4583 2295
rect 4614 2292 4620 2304
rect 4571 2264 4620 2292
rect 4571 2261 4583 2264
rect 4525 2255 4583 2261
rect 4614 2252 4620 2264
rect 4672 2252 4678 2304
rect 4893 2295 4951 2301
rect 4893 2261 4905 2295
rect 4939 2292 4951 2295
rect 5074 2292 5080 2304
rect 4939 2264 5080 2292
rect 4939 2261 4951 2264
rect 4893 2255 4951 2261
rect 5074 2252 5080 2264
rect 5132 2252 5138 2304
rect 5261 2295 5319 2301
rect 5261 2261 5273 2295
rect 5307 2292 5319 2295
rect 5442 2292 5448 2304
rect 5307 2264 5448 2292
rect 5307 2261 5319 2264
rect 5261 2255 5319 2261
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 5629 2295 5687 2301
rect 5629 2261 5641 2295
rect 5675 2292 5687 2295
rect 5810 2292 5816 2304
rect 5675 2264 5816 2292
rect 5675 2261 5687 2264
rect 5629 2255 5687 2261
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 5997 2295 6055 2301
rect 5997 2261 6009 2295
rect 6043 2292 6055 2295
rect 6178 2292 6184 2304
rect 6043 2264 6184 2292
rect 6043 2261 6055 2264
rect 5997 2255 6055 2261
rect 6178 2252 6184 2264
rect 6236 2252 6242 2304
rect 6546 2252 6552 2304
rect 6604 2292 6610 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6604 2264 6745 2292
rect 6604 2252 6610 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 6914 2252 6920 2304
rect 6972 2292 6978 2304
rect 7101 2295 7159 2301
rect 7101 2292 7113 2295
rect 6972 2264 7113 2292
rect 6972 2252 6978 2264
rect 7101 2261 7113 2264
rect 7147 2261 7159 2295
rect 7101 2255 7159 2261
rect 7282 2252 7288 2304
rect 7340 2292 7346 2304
rect 7469 2295 7527 2301
rect 7469 2292 7481 2295
rect 7340 2264 7481 2292
rect 7340 2252 7346 2264
rect 7469 2261 7481 2264
rect 7515 2261 7527 2295
rect 7469 2255 7527 2261
rect 7650 2252 7656 2304
rect 7708 2292 7714 2304
rect 7837 2295 7895 2301
rect 7837 2292 7849 2295
rect 7708 2264 7849 2292
rect 7708 2252 7714 2264
rect 7837 2261 7849 2264
rect 7883 2261 7895 2295
rect 7837 2255 7895 2261
rect 8018 2252 8024 2304
rect 8076 2292 8082 2304
rect 8205 2295 8263 2301
rect 8205 2292 8217 2295
rect 8076 2264 8217 2292
rect 8076 2252 8082 2264
rect 8205 2261 8217 2264
rect 8251 2261 8263 2295
rect 8205 2255 8263 2261
rect 8294 2252 8300 2304
rect 8352 2292 8358 2304
rect 8573 2295 8631 2301
rect 8573 2292 8585 2295
rect 8352 2264 8585 2292
rect 8352 2252 8358 2264
rect 8573 2261 8585 2264
rect 8619 2261 8631 2295
rect 9214 2292 9220 2304
rect 9175 2264 9220 2292
rect 8573 2255 8631 2261
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 10686 2292 10692 2304
rect 10647 2264 10692 2292
rect 10686 2252 10692 2264
rect 10744 2252 10750 2304
rect 11054 2292 11060 2304
rect 11015 2264 11060 2292
rect 11054 2252 11060 2264
rect 11112 2252 11118 2304
rect 11514 2292 11520 2304
rect 11475 2264 11520 2292
rect 11514 2252 11520 2264
rect 11572 2252 11578 2304
rect 11974 2252 11980 2304
rect 12032 2292 12038 2304
rect 12161 2295 12219 2301
rect 12161 2292 12173 2295
rect 12032 2264 12173 2292
rect 12032 2252 12038 2264
rect 12161 2261 12173 2264
rect 12207 2261 12219 2295
rect 13004 2292 13032 2332
rect 13265 2295 13323 2301
rect 13265 2292 13277 2295
rect 13004 2264 13277 2292
rect 12161 2255 12219 2261
rect 13265 2261 13277 2264
rect 13311 2261 13323 2295
rect 13265 2255 13323 2261
rect 13722 2252 13728 2304
rect 13780 2292 13786 2304
rect 14093 2295 14151 2301
rect 14093 2292 14105 2295
rect 13780 2264 14105 2292
rect 13780 2252 13786 2264
rect 14093 2261 14105 2264
rect 14139 2261 14151 2295
rect 14734 2292 14740 2304
rect 14695 2264 14740 2292
rect 14093 2255 14151 2261
rect 14734 2252 14740 2264
rect 14792 2252 14798 2304
rect 15102 2292 15108 2304
rect 15063 2264 15108 2292
rect 15102 2252 15108 2264
rect 15160 2252 15166 2304
rect 1104 2202 16008 2224
rect 1104 2150 4698 2202
rect 4750 2150 4762 2202
rect 4814 2150 4826 2202
rect 4878 2150 4890 2202
rect 4942 2150 4954 2202
rect 5006 2150 8446 2202
rect 8498 2150 8510 2202
rect 8562 2150 8574 2202
rect 8626 2150 8638 2202
rect 8690 2150 8702 2202
rect 8754 2150 12194 2202
rect 12246 2150 12258 2202
rect 12310 2150 12322 2202
rect 12374 2150 12386 2202
rect 12438 2150 12450 2202
rect 12502 2150 16008 2202
rect 1104 2128 16008 2150
rect 5534 2048 5540 2100
rect 5592 2088 5598 2100
rect 10686 2088 10692 2100
rect 5592 2060 10692 2088
rect 5592 2048 5598 2060
rect 10686 2048 10692 2060
rect 10744 2048 10750 2100
rect 11146 2048 11152 2100
rect 11204 2088 11210 2100
rect 15102 2088 15108 2100
rect 11204 2060 15108 2088
rect 11204 2048 11210 2060
rect 15102 2048 15108 2060
rect 15160 2048 15166 2100
rect 3510 1980 3516 2032
rect 3568 2020 3574 2032
rect 5994 2020 6000 2032
rect 3568 1992 6000 2020
rect 3568 1980 3574 1992
rect 5994 1980 6000 1992
rect 6052 1980 6058 2032
rect 7466 1980 7472 2032
rect 7524 2020 7530 2032
rect 11422 2020 11428 2032
rect 7524 1992 11428 2020
rect 7524 1980 7530 1992
rect 11422 1980 11428 1992
rect 11480 1980 11486 2032
rect 5350 1912 5356 1964
rect 5408 1952 5414 1964
rect 9214 1952 9220 1964
rect 5408 1924 9220 1952
rect 5408 1912 5414 1924
rect 9214 1912 9220 1924
rect 9272 1912 9278 1964
rect 9306 1912 9312 1964
rect 9364 1952 9370 1964
rect 14734 1952 14740 1964
rect 9364 1924 14740 1952
rect 9364 1912 9370 1924
rect 14734 1912 14740 1924
rect 14792 1912 14798 1964
rect 2774 1844 2780 1896
rect 2832 1884 2838 1896
rect 5718 1884 5724 1896
rect 2832 1856 5724 1884
rect 2832 1844 2838 1856
rect 5718 1844 5724 1856
rect 5776 1844 5782 1896
rect 9030 1844 9036 1896
rect 9088 1884 9094 1896
rect 11974 1884 11980 1896
rect 9088 1856 11980 1884
rect 9088 1844 9094 1856
rect 11974 1844 11980 1856
rect 12032 1844 12038 1896
rect 6454 1776 6460 1828
rect 6512 1816 6518 1828
rect 6512 1788 6914 1816
rect 6512 1776 6518 1788
rect 6886 1748 6914 1788
rect 7374 1776 7380 1828
rect 7432 1816 7438 1828
rect 11054 1816 11060 1828
rect 7432 1788 11060 1816
rect 7432 1776 7438 1788
rect 11054 1776 11060 1788
rect 11112 1776 11118 1828
rect 10042 1748 10048 1760
rect 6886 1720 10048 1748
rect 10042 1708 10048 1720
rect 10100 1708 10106 1760
<< via1 >>
rect 9220 17688 9272 17740
rect 13176 17688 13228 17740
rect 9128 17620 9180 17672
rect 12532 17620 12584 17672
rect 9496 17552 9548 17604
rect 12716 17552 12768 17604
rect 11336 17484 11388 17536
rect 14372 17484 14424 17536
rect 4698 17382 4750 17434
rect 4762 17382 4814 17434
rect 4826 17382 4878 17434
rect 4890 17382 4942 17434
rect 4954 17382 5006 17434
rect 8446 17382 8498 17434
rect 8510 17382 8562 17434
rect 8574 17382 8626 17434
rect 8638 17382 8690 17434
rect 8702 17382 8754 17434
rect 12194 17382 12246 17434
rect 12258 17382 12310 17434
rect 12322 17382 12374 17434
rect 12386 17382 12438 17434
rect 12450 17382 12502 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 1952 17323 2004 17332
rect 1952 17289 1961 17323
rect 1961 17289 1995 17323
rect 1995 17289 2004 17323
rect 1952 17280 2004 17289
rect 2320 17323 2372 17332
rect 2320 17289 2329 17323
rect 2329 17289 2363 17323
rect 2363 17289 2372 17323
rect 2320 17280 2372 17289
rect 2688 17323 2740 17332
rect 2688 17289 2697 17323
rect 2697 17289 2731 17323
rect 2731 17289 2740 17323
rect 2688 17280 2740 17289
rect 3056 17323 3108 17332
rect 3056 17289 3065 17323
rect 3065 17289 3099 17323
rect 3099 17289 3108 17323
rect 3056 17280 3108 17289
rect 3424 17323 3476 17332
rect 3424 17289 3433 17323
rect 3433 17289 3467 17323
rect 3467 17289 3476 17323
rect 3424 17280 3476 17289
rect 4160 17323 4212 17332
rect 4160 17289 4169 17323
rect 4169 17289 4203 17323
rect 4203 17289 4212 17323
rect 4160 17280 4212 17289
rect 4528 17323 4580 17332
rect 4528 17289 4537 17323
rect 4537 17289 4571 17323
rect 4571 17289 4580 17323
rect 4528 17280 4580 17289
rect 5080 17280 5132 17332
rect 5264 17323 5316 17332
rect 5264 17289 5273 17323
rect 5273 17289 5307 17323
rect 5307 17289 5316 17323
rect 5264 17280 5316 17289
rect 5632 17323 5684 17332
rect 5632 17289 5641 17323
rect 5641 17289 5675 17323
rect 5675 17289 5684 17323
rect 5632 17280 5684 17289
rect 6000 17323 6052 17332
rect 6000 17289 6009 17323
rect 6009 17289 6043 17323
rect 6043 17289 6052 17323
rect 6000 17280 6052 17289
rect 6368 17280 6420 17332
rect 6920 17323 6972 17332
rect 6920 17289 6929 17323
rect 6929 17289 6963 17323
rect 6963 17289 6972 17323
rect 6920 17280 6972 17289
rect 7104 17280 7156 17332
rect 7472 17280 7524 17332
rect 7840 17280 7892 17332
rect 8300 17280 8352 17332
rect 8852 17280 8904 17332
rect 9588 17280 9640 17332
rect 13452 17323 13504 17332
rect 2136 17187 2188 17196
rect 2136 17153 2145 17187
rect 2145 17153 2179 17187
rect 2179 17153 2188 17187
rect 2136 17144 2188 17153
rect 2504 17187 2556 17196
rect 2504 17153 2513 17187
rect 2513 17153 2547 17187
rect 2547 17153 2556 17187
rect 2504 17144 2556 17153
rect 4620 17212 4672 17264
rect 3608 17187 3660 17196
rect 3148 17076 3200 17128
rect 3608 17153 3617 17187
rect 3617 17153 3651 17187
rect 3651 17153 3660 17187
rect 3608 17144 3660 17153
rect 4344 17187 4396 17196
rect 4344 17153 4353 17187
rect 4353 17153 4387 17187
rect 4387 17153 4396 17187
rect 4344 17144 4396 17153
rect 5448 17187 5500 17196
rect 4436 17076 4488 17128
rect 5448 17153 5457 17187
rect 5457 17153 5491 17187
rect 5491 17153 5500 17187
rect 5448 17144 5500 17153
rect 6184 17187 6236 17196
rect 6184 17153 6193 17187
rect 6193 17153 6227 17187
rect 6227 17153 6236 17187
rect 6184 17144 6236 17153
rect 6276 17144 6328 17196
rect 7472 17187 7524 17196
rect 6460 17076 6512 17128
rect 5724 17008 5776 17060
rect 7472 17153 7481 17187
rect 7481 17153 7515 17187
rect 7515 17153 7524 17187
rect 7472 17144 7524 17153
rect 8208 17187 8260 17196
rect 8208 17153 8217 17187
rect 8217 17153 8251 17187
rect 8251 17153 8260 17187
rect 8208 17144 8260 17153
rect 8300 17076 8352 17128
rect 8852 17144 8904 17196
rect 9220 17187 9272 17196
rect 9220 17153 9229 17187
rect 9229 17153 9263 17187
rect 9263 17153 9272 17187
rect 9220 17144 9272 17153
rect 9312 17144 9364 17196
rect 9680 17144 9732 17196
rect 10048 17144 10100 17196
rect 10416 17144 10468 17196
rect 11520 17212 11572 17264
rect 10784 17144 10836 17196
rect 11152 17144 11204 17196
rect 9128 17076 9180 17128
rect 11428 17076 11480 17128
rect 11888 17076 11940 17128
rect 13452 17289 13461 17323
rect 13461 17289 13495 17323
rect 13495 17289 13504 17323
rect 13452 17280 13504 17289
rect 14372 17323 14424 17332
rect 14372 17289 14381 17323
rect 14381 17289 14415 17323
rect 14415 17289 14424 17323
rect 14372 17280 14424 17289
rect 15568 17323 15620 17332
rect 15568 17289 15577 17323
rect 15577 17289 15611 17323
rect 15611 17289 15620 17323
rect 15568 17280 15620 17289
rect 12440 17144 12492 17196
rect 12624 17144 12676 17196
rect 12992 17144 13044 17196
rect 14096 17212 14148 17264
rect 14464 17212 14516 17264
rect 13360 17144 13412 17196
rect 13820 17144 13872 17196
rect 14648 17144 14700 17196
rect 14924 17144 14976 17196
rect 9312 17008 9364 17060
rect 9956 17008 10008 17060
rect 11060 17008 11112 17060
rect 4344 16940 4396 16992
rect 6368 16940 6420 16992
rect 9404 16983 9456 16992
rect 9404 16949 9413 16983
rect 9413 16949 9447 16983
rect 9447 16949 9456 16983
rect 9404 16940 9456 16949
rect 10140 16983 10192 16992
rect 10140 16949 10149 16983
rect 10149 16949 10183 16983
rect 10183 16949 10192 16983
rect 10140 16940 10192 16949
rect 10692 16940 10744 16992
rect 10968 16940 11020 16992
rect 12256 17008 12308 17060
rect 14740 17076 14792 17128
rect 11796 16983 11848 16992
rect 11796 16949 11805 16983
rect 11805 16949 11839 16983
rect 11839 16949 11848 16983
rect 11796 16940 11848 16949
rect 11980 16940 12032 16992
rect 12716 16983 12768 16992
rect 12716 16949 12725 16983
rect 12725 16949 12759 16983
rect 12759 16949 12768 16983
rect 12716 16940 12768 16949
rect 12808 16940 12860 16992
rect 14648 16983 14700 16992
rect 14648 16949 14657 16983
rect 14657 16949 14691 16983
rect 14691 16949 14700 16983
rect 14648 16940 14700 16949
rect 2824 16838 2876 16890
rect 2888 16838 2940 16890
rect 2952 16838 3004 16890
rect 3016 16838 3068 16890
rect 3080 16838 3132 16890
rect 6572 16838 6624 16890
rect 6636 16838 6688 16890
rect 6700 16838 6752 16890
rect 6764 16838 6816 16890
rect 6828 16838 6880 16890
rect 10320 16838 10372 16890
rect 10384 16838 10436 16890
rect 10448 16838 10500 16890
rect 10512 16838 10564 16890
rect 10576 16838 10628 16890
rect 14068 16838 14120 16890
rect 14132 16838 14184 16890
rect 14196 16838 14248 16890
rect 14260 16838 14312 16890
rect 14324 16838 14376 16890
rect 5264 16736 5316 16788
rect 9404 16736 9456 16788
rect 9680 16779 9732 16788
rect 9680 16745 9689 16779
rect 9689 16745 9723 16779
rect 9723 16745 9732 16779
rect 9680 16736 9732 16745
rect 10048 16779 10100 16788
rect 10048 16745 10057 16779
rect 10057 16745 10091 16779
rect 10091 16745 10100 16779
rect 10048 16736 10100 16745
rect 10784 16779 10836 16788
rect 10784 16745 10793 16779
rect 10793 16745 10827 16779
rect 10827 16745 10836 16779
rect 10784 16736 10836 16745
rect 11152 16736 11204 16788
rect 11520 16736 11572 16788
rect 11888 16779 11940 16788
rect 11888 16745 11897 16779
rect 11897 16745 11931 16779
rect 11931 16745 11940 16779
rect 11888 16736 11940 16745
rect 12072 16736 12124 16788
rect 12440 16736 12492 16788
rect 12624 16779 12676 16788
rect 12624 16745 12633 16779
rect 12633 16745 12667 16779
rect 12667 16745 12676 16779
rect 12624 16736 12676 16745
rect 13360 16779 13412 16788
rect 13360 16745 13369 16779
rect 13369 16745 13403 16779
rect 13403 16745 13412 16779
rect 13360 16736 13412 16745
rect 13820 16736 13872 16788
rect 14464 16736 14516 16788
rect 14832 16779 14884 16788
rect 14832 16745 14841 16779
rect 14841 16745 14875 16779
rect 14875 16745 14884 16779
rect 14832 16736 14884 16745
rect 4620 16668 4672 16720
rect 5540 16668 5592 16720
rect 11244 16668 11296 16720
rect 12256 16668 12308 16720
rect 12348 16668 12400 16720
rect 13452 16668 13504 16720
rect 8944 16600 8996 16652
rect 1308 16532 1360 16584
rect 1676 16575 1728 16584
rect 1676 16541 1685 16575
rect 1685 16541 1719 16575
rect 1719 16541 1728 16575
rect 1676 16532 1728 16541
rect 1584 16439 1636 16448
rect 1584 16405 1593 16439
rect 1593 16405 1627 16439
rect 1627 16405 1636 16439
rect 1584 16396 1636 16405
rect 4068 16532 4120 16584
rect 7196 16532 7248 16584
rect 9404 16600 9456 16652
rect 9588 16600 9640 16652
rect 10784 16600 10836 16652
rect 11980 16600 12032 16652
rect 15292 16600 15344 16652
rect 15384 16532 15436 16584
rect 3792 16396 3844 16448
rect 7288 16396 7340 16448
rect 15016 16439 15068 16448
rect 15016 16405 15025 16439
rect 15025 16405 15059 16439
rect 15059 16405 15068 16439
rect 15016 16396 15068 16405
rect 15108 16396 15160 16448
rect 4698 16294 4750 16346
rect 4762 16294 4814 16346
rect 4826 16294 4878 16346
rect 4890 16294 4942 16346
rect 4954 16294 5006 16346
rect 8446 16294 8498 16346
rect 8510 16294 8562 16346
rect 8574 16294 8626 16346
rect 8638 16294 8690 16346
rect 8702 16294 8754 16346
rect 12194 16294 12246 16346
rect 12258 16294 12310 16346
rect 12322 16294 12374 16346
rect 12386 16294 12438 16346
rect 12450 16294 12502 16346
rect 1308 16192 1360 16244
rect 1584 16192 1636 16244
rect 5080 16192 5132 16244
rect 15936 16056 15988 16108
rect 15476 15895 15528 15904
rect 15476 15861 15485 15895
rect 15485 15861 15519 15895
rect 15519 15861 15528 15895
rect 15476 15852 15528 15861
rect 2824 15750 2876 15802
rect 2888 15750 2940 15802
rect 2952 15750 3004 15802
rect 3016 15750 3068 15802
rect 3080 15750 3132 15802
rect 6572 15750 6624 15802
rect 6636 15750 6688 15802
rect 6700 15750 6752 15802
rect 6764 15750 6816 15802
rect 6828 15750 6880 15802
rect 10320 15750 10372 15802
rect 10384 15750 10436 15802
rect 10448 15750 10500 15802
rect 10512 15750 10564 15802
rect 10576 15750 10628 15802
rect 14068 15750 14120 15802
rect 14132 15750 14184 15802
rect 14196 15750 14248 15802
rect 14260 15750 14312 15802
rect 14324 15750 14376 15802
rect 4698 15206 4750 15258
rect 4762 15206 4814 15258
rect 4826 15206 4878 15258
rect 4890 15206 4942 15258
rect 4954 15206 5006 15258
rect 8446 15206 8498 15258
rect 8510 15206 8562 15258
rect 8574 15206 8626 15258
rect 8638 15206 8690 15258
rect 8702 15206 8754 15258
rect 12194 15206 12246 15258
rect 12258 15206 12310 15258
rect 12322 15206 12374 15258
rect 12386 15206 12438 15258
rect 12450 15206 12502 15258
rect 2824 14662 2876 14714
rect 2888 14662 2940 14714
rect 2952 14662 3004 14714
rect 3016 14662 3068 14714
rect 3080 14662 3132 14714
rect 6572 14662 6624 14714
rect 6636 14662 6688 14714
rect 6700 14662 6752 14714
rect 6764 14662 6816 14714
rect 6828 14662 6880 14714
rect 10320 14662 10372 14714
rect 10384 14662 10436 14714
rect 10448 14662 10500 14714
rect 10512 14662 10564 14714
rect 10576 14662 10628 14714
rect 14068 14662 14120 14714
rect 14132 14662 14184 14714
rect 14196 14662 14248 14714
rect 14260 14662 14312 14714
rect 14324 14662 14376 14714
rect 4698 14118 4750 14170
rect 4762 14118 4814 14170
rect 4826 14118 4878 14170
rect 4890 14118 4942 14170
rect 4954 14118 5006 14170
rect 8446 14118 8498 14170
rect 8510 14118 8562 14170
rect 8574 14118 8626 14170
rect 8638 14118 8690 14170
rect 8702 14118 8754 14170
rect 12194 14118 12246 14170
rect 12258 14118 12310 14170
rect 12322 14118 12374 14170
rect 12386 14118 12438 14170
rect 12450 14118 12502 14170
rect 5080 13923 5132 13932
rect 5080 13889 5089 13923
rect 5089 13889 5123 13923
rect 5123 13889 5132 13923
rect 5080 13880 5132 13889
rect 3516 13812 3568 13864
rect 7656 13676 7708 13728
rect 2824 13574 2876 13626
rect 2888 13574 2940 13626
rect 2952 13574 3004 13626
rect 3016 13574 3068 13626
rect 3080 13574 3132 13626
rect 6572 13574 6624 13626
rect 6636 13574 6688 13626
rect 6700 13574 6752 13626
rect 6764 13574 6816 13626
rect 6828 13574 6880 13626
rect 10320 13574 10372 13626
rect 10384 13574 10436 13626
rect 10448 13574 10500 13626
rect 10512 13574 10564 13626
rect 10576 13574 10628 13626
rect 14068 13574 14120 13626
rect 14132 13574 14184 13626
rect 14196 13574 14248 13626
rect 14260 13574 14312 13626
rect 14324 13574 14376 13626
rect 4698 13030 4750 13082
rect 4762 13030 4814 13082
rect 4826 13030 4878 13082
rect 4890 13030 4942 13082
rect 4954 13030 5006 13082
rect 8446 13030 8498 13082
rect 8510 13030 8562 13082
rect 8574 13030 8626 13082
rect 8638 13030 8690 13082
rect 8702 13030 8754 13082
rect 12194 13030 12246 13082
rect 12258 13030 12310 13082
rect 12322 13030 12374 13082
rect 12386 13030 12438 13082
rect 12450 13030 12502 13082
rect 3148 12928 3200 12980
rect 5724 12928 5776 12980
rect 14740 12928 14792 12980
rect 4160 12860 4212 12912
rect 7656 12860 7708 12912
rect 4344 12767 4396 12776
rect 4344 12733 4353 12767
rect 4353 12733 4387 12767
rect 4387 12733 4396 12767
rect 4344 12724 4396 12733
rect 8392 12792 8444 12844
rect 7104 12724 7156 12776
rect 7012 12656 7064 12708
rect 13912 12588 13964 12640
rect 15568 12631 15620 12640
rect 15568 12597 15577 12631
rect 15577 12597 15611 12631
rect 15611 12597 15620 12631
rect 15568 12588 15620 12597
rect 2824 12486 2876 12538
rect 2888 12486 2940 12538
rect 2952 12486 3004 12538
rect 3016 12486 3068 12538
rect 3080 12486 3132 12538
rect 6572 12486 6624 12538
rect 6636 12486 6688 12538
rect 6700 12486 6752 12538
rect 6764 12486 6816 12538
rect 6828 12486 6880 12538
rect 10320 12486 10372 12538
rect 10384 12486 10436 12538
rect 10448 12486 10500 12538
rect 10512 12486 10564 12538
rect 10576 12486 10628 12538
rect 14068 12486 14120 12538
rect 14132 12486 14184 12538
rect 14196 12486 14248 12538
rect 14260 12486 14312 12538
rect 14324 12486 14376 12538
rect 2504 12384 2556 12436
rect 5448 12384 5500 12436
rect 8300 12384 8352 12436
rect 8116 12112 8168 12164
rect 9312 12180 9364 12232
rect 9772 12112 9824 12164
rect 4698 11942 4750 11994
rect 4762 11942 4814 11994
rect 4826 11942 4878 11994
rect 4890 11942 4942 11994
rect 4954 11942 5006 11994
rect 8446 11942 8498 11994
rect 8510 11942 8562 11994
rect 8574 11942 8626 11994
rect 8638 11942 8690 11994
rect 8702 11942 8754 11994
rect 12194 11942 12246 11994
rect 12258 11942 12310 11994
rect 12322 11942 12374 11994
rect 12386 11942 12438 11994
rect 12450 11942 12502 11994
rect 7196 11883 7248 11892
rect 7196 11849 7205 11883
rect 7205 11849 7239 11883
rect 7239 11849 7248 11883
rect 7196 11840 7248 11849
rect 6460 11772 6512 11824
rect 1400 11747 1452 11756
rect 1400 11713 1409 11747
rect 1409 11713 1443 11747
rect 1443 11713 1452 11747
rect 1400 11704 1452 11713
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 7748 11747 7800 11756
rect 7748 11713 7757 11747
rect 7757 11713 7791 11747
rect 7791 11713 7800 11747
rect 7748 11704 7800 11713
rect 8024 11747 8076 11756
rect 8024 11713 8033 11747
rect 8033 11713 8067 11747
rect 8067 11713 8076 11747
rect 8024 11704 8076 11713
rect 5724 11636 5776 11688
rect 8208 11679 8260 11688
rect 8208 11645 8217 11679
rect 8217 11645 8251 11679
rect 8251 11645 8260 11679
rect 8208 11636 8260 11645
rect 6368 11568 6420 11620
rect 5908 11500 5960 11552
rect 8852 11500 8904 11552
rect 2824 11398 2876 11450
rect 2888 11398 2940 11450
rect 2952 11398 3004 11450
rect 3016 11398 3068 11450
rect 3080 11398 3132 11450
rect 6572 11398 6624 11450
rect 6636 11398 6688 11450
rect 6700 11398 6752 11450
rect 6764 11398 6816 11450
rect 6828 11398 6880 11450
rect 10320 11398 10372 11450
rect 10384 11398 10436 11450
rect 10448 11398 10500 11450
rect 10512 11398 10564 11450
rect 10576 11398 10628 11450
rect 14068 11398 14120 11450
rect 14132 11398 14184 11450
rect 14196 11398 14248 11450
rect 14260 11398 14312 11450
rect 14324 11398 14376 11450
rect 7012 11296 7064 11348
rect 8208 11271 8260 11280
rect 8208 11237 8217 11271
rect 8217 11237 8251 11271
rect 8251 11237 8260 11271
rect 8208 11228 8260 11237
rect 4344 11160 4396 11212
rect 10876 11228 10928 11280
rect 9496 11203 9548 11212
rect 9496 11169 9505 11203
rect 9505 11169 9539 11203
rect 9539 11169 9548 11203
rect 9496 11160 9548 11169
rect 4344 11024 4396 11076
rect 6920 11024 6972 11076
rect 9128 11024 9180 11076
rect 9404 11067 9456 11076
rect 9404 11033 9413 11067
rect 9413 11033 9447 11067
rect 9447 11033 9456 11067
rect 9404 11024 9456 11033
rect 9220 10956 9272 11008
rect 9588 10956 9640 11008
rect 4698 10854 4750 10906
rect 4762 10854 4814 10906
rect 4826 10854 4878 10906
rect 4890 10854 4942 10906
rect 4954 10854 5006 10906
rect 8446 10854 8498 10906
rect 8510 10854 8562 10906
rect 8574 10854 8626 10906
rect 8638 10854 8690 10906
rect 8702 10854 8754 10906
rect 12194 10854 12246 10906
rect 12258 10854 12310 10906
rect 12322 10854 12374 10906
rect 12386 10854 12438 10906
rect 12450 10854 12502 10906
rect 5540 10752 5592 10804
rect 3608 10684 3660 10736
rect 7656 10752 7708 10804
rect 8944 10752 8996 10804
rect 3516 10659 3568 10668
rect 3516 10625 3534 10659
rect 3534 10625 3568 10659
rect 3516 10616 3568 10625
rect 5540 10616 5592 10668
rect 6000 10616 6052 10668
rect 6828 10659 6880 10668
rect 5632 10548 5684 10600
rect 5080 10480 5132 10532
rect 6828 10625 6837 10659
rect 6837 10625 6871 10659
rect 6871 10625 6880 10659
rect 6828 10616 6880 10625
rect 7104 10616 7156 10668
rect 7288 10659 7340 10668
rect 7288 10625 7297 10659
rect 7297 10625 7331 10659
rect 7331 10625 7340 10659
rect 7288 10616 7340 10625
rect 7472 10616 7524 10668
rect 8852 10727 8904 10736
rect 8852 10693 8870 10727
rect 8870 10693 8904 10727
rect 8852 10684 8904 10693
rect 9588 10616 9640 10668
rect 12072 10684 12124 10736
rect 11244 10616 11296 10668
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 9128 10591 9180 10600
rect 9128 10557 9137 10591
rect 9137 10557 9171 10591
rect 9171 10557 9180 10591
rect 9128 10548 9180 10557
rect 11152 10548 11204 10600
rect 5816 10412 5868 10464
rect 6460 10412 6512 10464
rect 7656 10455 7708 10464
rect 7656 10421 7665 10455
rect 7665 10421 7699 10455
rect 7699 10421 7708 10455
rect 7656 10412 7708 10421
rect 11060 10480 11112 10532
rect 9956 10412 10008 10464
rect 11704 10412 11756 10464
rect 14648 10412 14700 10464
rect 2824 10310 2876 10362
rect 2888 10310 2940 10362
rect 2952 10310 3004 10362
rect 3016 10310 3068 10362
rect 3080 10310 3132 10362
rect 6572 10310 6624 10362
rect 6636 10310 6688 10362
rect 6700 10310 6752 10362
rect 6764 10310 6816 10362
rect 6828 10310 6880 10362
rect 10320 10310 10372 10362
rect 10384 10310 10436 10362
rect 10448 10310 10500 10362
rect 10512 10310 10564 10362
rect 10576 10310 10628 10362
rect 14068 10310 14120 10362
rect 14132 10310 14184 10362
rect 14196 10310 14248 10362
rect 14260 10310 14312 10362
rect 14324 10310 14376 10362
rect 8116 10208 8168 10260
rect 3240 10140 3292 10192
rect 5540 10140 5592 10192
rect 6368 10140 6420 10192
rect 7656 10140 7708 10192
rect 5724 10115 5776 10124
rect 5724 10081 5733 10115
rect 5733 10081 5767 10115
rect 5767 10081 5776 10115
rect 5724 10072 5776 10081
rect 5816 10072 5868 10124
rect 7104 10072 7156 10124
rect 8300 10115 8352 10124
rect 8300 10081 8309 10115
rect 8309 10081 8343 10115
rect 8343 10081 8352 10115
rect 8300 10072 8352 10081
rect 8392 10072 8444 10124
rect 5264 10004 5316 10056
rect 5908 10047 5960 10056
rect 5908 10013 5917 10047
rect 5917 10013 5951 10047
rect 5951 10013 5960 10047
rect 5908 10004 5960 10013
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 9496 10072 9548 10124
rect 10048 10140 10100 10192
rect 11428 10208 11480 10260
rect 12532 10208 12584 10260
rect 13176 10251 13228 10260
rect 13176 10217 13185 10251
rect 13185 10217 13219 10251
rect 13219 10217 13228 10251
rect 13176 10208 13228 10217
rect 11612 10140 11664 10192
rect 11244 10072 11296 10124
rect 5816 9936 5868 9988
rect 7564 9936 7616 9988
rect 9220 9936 9272 9988
rect 10968 10004 11020 10056
rect 11336 10004 11388 10056
rect 11520 10004 11572 10056
rect 11704 10047 11756 10056
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 15016 10140 15068 10192
rect 10324 9936 10376 9988
rect 12992 10004 13044 10056
rect 15476 10072 15528 10124
rect 13360 10047 13412 10056
rect 13360 10013 13369 10047
rect 13369 10013 13403 10047
rect 13403 10013 13412 10047
rect 13360 10004 13412 10013
rect 15108 9936 15160 9988
rect 3700 9868 3752 9920
rect 5540 9911 5592 9920
rect 5540 9877 5549 9911
rect 5549 9877 5583 9911
rect 5583 9877 5592 9911
rect 5540 9868 5592 9877
rect 7288 9868 7340 9920
rect 8392 9911 8444 9920
rect 8392 9877 8401 9911
rect 8401 9877 8435 9911
rect 8435 9877 8444 9911
rect 8392 9868 8444 9877
rect 8668 9868 8720 9920
rect 8944 9868 8996 9920
rect 9312 9868 9364 9920
rect 9864 9911 9916 9920
rect 9864 9877 9873 9911
rect 9873 9877 9907 9911
rect 9907 9877 9916 9911
rect 9864 9868 9916 9877
rect 10232 9911 10284 9920
rect 10232 9877 10241 9911
rect 10241 9877 10275 9911
rect 10275 9877 10284 9911
rect 10232 9868 10284 9877
rect 10876 9868 10928 9920
rect 11428 9868 11480 9920
rect 11704 9868 11756 9920
rect 13084 9868 13136 9920
rect 4698 9766 4750 9818
rect 4762 9766 4814 9818
rect 4826 9766 4878 9818
rect 4890 9766 4942 9818
rect 4954 9766 5006 9818
rect 8446 9766 8498 9818
rect 8510 9766 8562 9818
rect 8574 9766 8626 9818
rect 8638 9766 8690 9818
rect 8702 9766 8754 9818
rect 12194 9766 12246 9818
rect 12258 9766 12310 9818
rect 12322 9766 12374 9818
rect 12386 9766 12438 9818
rect 12450 9766 12502 9818
rect 5816 9664 5868 9716
rect 8668 9664 8720 9716
rect 9496 9664 9548 9716
rect 1492 9596 1544 9648
rect 3516 9596 3568 9648
rect 8944 9596 8996 9648
rect 11520 9664 11572 9716
rect 13728 9664 13780 9716
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 6092 9528 6144 9580
rect 3424 9460 3476 9512
rect 2136 9392 2188 9444
rect 7012 9528 7064 9580
rect 7104 9528 7156 9580
rect 6920 9503 6972 9512
rect 6920 9469 6929 9503
rect 6929 9469 6963 9503
rect 6963 9469 6972 9503
rect 6920 9460 6972 9469
rect 7104 9392 7156 9444
rect 5724 9367 5776 9376
rect 5724 9333 5733 9367
rect 5733 9333 5767 9367
rect 5767 9333 5776 9367
rect 5724 9324 5776 9333
rect 6000 9367 6052 9376
rect 6000 9333 6009 9367
rect 6009 9333 6043 9367
rect 6043 9333 6052 9367
rect 6000 9324 6052 9333
rect 8300 9460 8352 9512
rect 8576 9460 8628 9512
rect 9220 9528 9272 9580
rect 8944 9503 8996 9512
rect 8944 9469 8953 9503
rect 8953 9469 8987 9503
rect 8987 9469 8996 9503
rect 8944 9460 8996 9469
rect 8208 9392 8260 9444
rect 9588 9528 9640 9580
rect 10784 9460 10836 9512
rect 11888 9528 11940 9580
rect 11980 9460 12032 9512
rect 8300 9324 8352 9376
rect 10232 9392 10284 9444
rect 9036 9324 9088 9376
rect 9220 9324 9272 9376
rect 9588 9367 9640 9376
rect 9588 9333 9597 9367
rect 9597 9333 9631 9367
rect 9631 9333 9640 9367
rect 9588 9324 9640 9333
rect 2824 9222 2876 9274
rect 2888 9222 2940 9274
rect 2952 9222 3004 9274
rect 3016 9222 3068 9274
rect 3080 9222 3132 9274
rect 6572 9222 6624 9274
rect 6636 9222 6688 9274
rect 6700 9222 6752 9274
rect 6764 9222 6816 9274
rect 6828 9222 6880 9274
rect 10320 9222 10372 9274
rect 10384 9222 10436 9274
rect 10448 9222 10500 9274
rect 10512 9222 10564 9274
rect 10576 9222 10628 9274
rect 14068 9222 14120 9274
rect 14132 9222 14184 9274
rect 14196 9222 14248 9274
rect 14260 9222 14312 9274
rect 14324 9222 14376 9274
rect 6920 9163 6972 9172
rect 6920 9129 6929 9163
rect 6929 9129 6963 9163
rect 6963 9129 6972 9163
rect 6920 9120 6972 9129
rect 7104 9120 7156 9172
rect 9680 9120 9732 9172
rect 8392 9095 8444 9104
rect 8392 9061 8401 9095
rect 8401 9061 8435 9095
rect 8435 9061 8444 9095
rect 8392 9052 8444 9061
rect 8576 9052 8628 9104
rect 8944 9052 8996 9104
rect 6092 8916 6144 8968
rect 10140 8984 10192 9036
rect 8300 8959 8352 8968
rect 8300 8925 8309 8959
rect 8309 8925 8343 8959
rect 8343 8925 8352 8959
rect 8300 8916 8352 8925
rect 9036 8916 9088 8968
rect 10692 8916 10744 8968
rect 8484 8848 8536 8900
rect 6184 8780 6236 8832
rect 9588 8848 9640 8900
rect 9772 8848 9824 8900
rect 12624 8848 12676 8900
rect 8944 8823 8996 8832
rect 8944 8789 8953 8823
rect 8953 8789 8987 8823
rect 8987 8789 8996 8823
rect 8944 8780 8996 8789
rect 4698 8678 4750 8730
rect 4762 8678 4814 8730
rect 4826 8678 4878 8730
rect 4890 8678 4942 8730
rect 4954 8678 5006 8730
rect 8446 8678 8498 8730
rect 8510 8678 8562 8730
rect 8574 8678 8626 8730
rect 8638 8678 8690 8730
rect 8702 8678 8754 8730
rect 12194 8678 12246 8730
rect 12258 8678 12310 8730
rect 12322 8678 12374 8730
rect 12386 8678 12438 8730
rect 12450 8678 12502 8730
rect 5540 8576 5592 8628
rect 8852 8576 8904 8628
rect 8300 8508 8352 8560
rect 11152 8508 11204 8560
rect 3516 8440 3568 8492
rect 6920 8440 6972 8492
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 9864 8440 9916 8492
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 9496 8372 9548 8424
rect 8300 8304 8352 8356
rect 8944 8304 8996 8356
rect 8392 8236 8444 8288
rect 9772 8304 9824 8356
rect 12716 8347 12768 8356
rect 12716 8313 12725 8347
rect 12725 8313 12759 8347
rect 12759 8313 12768 8347
rect 12716 8304 12768 8313
rect 2824 8134 2876 8186
rect 2888 8134 2940 8186
rect 2952 8134 3004 8186
rect 3016 8134 3068 8186
rect 3080 8134 3132 8186
rect 6572 8134 6624 8186
rect 6636 8134 6688 8186
rect 6700 8134 6752 8186
rect 6764 8134 6816 8186
rect 6828 8134 6880 8186
rect 10320 8134 10372 8186
rect 10384 8134 10436 8186
rect 10448 8134 10500 8186
rect 10512 8134 10564 8186
rect 10576 8134 10628 8186
rect 14068 8134 14120 8186
rect 14132 8134 14184 8186
rect 14196 8134 14248 8186
rect 14260 8134 14312 8186
rect 14324 8134 14376 8186
rect 4698 7590 4750 7642
rect 4762 7590 4814 7642
rect 4826 7590 4878 7642
rect 4890 7590 4942 7642
rect 4954 7590 5006 7642
rect 8446 7590 8498 7642
rect 8510 7590 8562 7642
rect 8574 7590 8626 7642
rect 8638 7590 8690 7642
rect 8702 7590 8754 7642
rect 12194 7590 12246 7642
rect 12258 7590 12310 7642
rect 12322 7590 12374 7642
rect 12386 7590 12438 7642
rect 12450 7590 12502 7642
rect 4160 7488 4212 7540
rect 7472 7488 7524 7540
rect 3240 7395 3292 7404
rect 3240 7361 3249 7395
rect 3249 7361 3283 7395
rect 3283 7361 3292 7395
rect 3240 7352 3292 7361
rect 7288 7352 7340 7404
rect 7564 7395 7616 7404
rect 7564 7361 7573 7395
rect 7573 7361 7607 7395
rect 7607 7361 7616 7395
rect 7564 7352 7616 7361
rect 9404 7395 9456 7404
rect 9404 7361 9413 7395
rect 9413 7361 9447 7395
rect 9447 7361 9456 7395
rect 9404 7352 9456 7361
rect 8852 7284 8904 7336
rect 5172 7216 5224 7268
rect 3148 7148 3200 7200
rect 3332 7148 3384 7200
rect 4620 7148 4672 7200
rect 7656 7148 7708 7200
rect 2824 7046 2876 7098
rect 2888 7046 2940 7098
rect 2952 7046 3004 7098
rect 3016 7046 3068 7098
rect 3080 7046 3132 7098
rect 6572 7046 6624 7098
rect 6636 7046 6688 7098
rect 6700 7046 6752 7098
rect 6764 7046 6816 7098
rect 6828 7046 6880 7098
rect 10320 7046 10372 7098
rect 10384 7046 10436 7098
rect 10448 7046 10500 7098
rect 10512 7046 10564 7098
rect 10576 7046 10628 7098
rect 14068 7046 14120 7098
rect 14132 7046 14184 7098
rect 14196 7046 14248 7098
rect 14260 7046 14312 7098
rect 14324 7046 14376 7098
rect 4698 6502 4750 6554
rect 4762 6502 4814 6554
rect 4826 6502 4878 6554
rect 4890 6502 4942 6554
rect 4954 6502 5006 6554
rect 8446 6502 8498 6554
rect 8510 6502 8562 6554
rect 8574 6502 8626 6554
rect 8638 6502 8690 6554
rect 8702 6502 8754 6554
rect 12194 6502 12246 6554
rect 12258 6502 12310 6554
rect 12322 6502 12374 6554
rect 12386 6502 12438 6554
rect 12450 6502 12502 6554
rect 2824 5958 2876 6010
rect 2888 5958 2940 6010
rect 2952 5958 3004 6010
rect 3016 5958 3068 6010
rect 3080 5958 3132 6010
rect 6572 5958 6624 6010
rect 6636 5958 6688 6010
rect 6700 5958 6752 6010
rect 6764 5958 6816 6010
rect 6828 5958 6880 6010
rect 10320 5958 10372 6010
rect 10384 5958 10436 6010
rect 10448 5958 10500 6010
rect 10512 5958 10564 6010
rect 10576 5958 10628 6010
rect 14068 5958 14120 6010
rect 14132 5958 14184 6010
rect 14196 5958 14248 6010
rect 14260 5958 14312 6010
rect 14324 5958 14376 6010
rect 4698 5414 4750 5466
rect 4762 5414 4814 5466
rect 4826 5414 4878 5466
rect 4890 5414 4942 5466
rect 4954 5414 5006 5466
rect 8446 5414 8498 5466
rect 8510 5414 8562 5466
rect 8574 5414 8626 5466
rect 8638 5414 8690 5466
rect 8702 5414 8754 5466
rect 12194 5414 12246 5466
rect 12258 5414 12310 5466
rect 12322 5414 12374 5466
rect 12386 5414 12438 5466
rect 12450 5414 12502 5466
rect 3148 5176 3200 5228
rect 1492 5083 1544 5092
rect 1492 5049 1501 5083
rect 1501 5049 1535 5083
rect 1535 5049 1544 5083
rect 1492 5040 1544 5049
rect 2824 4870 2876 4922
rect 2888 4870 2940 4922
rect 2952 4870 3004 4922
rect 3016 4870 3068 4922
rect 3080 4870 3132 4922
rect 6572 4870 6624 4922
rect 6636 4870 6688 4922
rect 6700 4870 6752 4922
rect 6764 4870 6816 4922
rect 6828 4870 6880 4922
rect 10320 4870 10372 4922
rect 10384 4870 10436 4922
rect 10448 4870 10500 4922
rect 10512 4870 10564 4922
rect 10576 4870 10628 4922
rect 14068 4870 14120 4922
rect 14132 4870 14184 4922
rect 14196 4870 14248 4922
rect 14260 4870 14312 4922
rect 14324 4870 14376 4922
rect 4698 4326 4750 4378
rect 4762 4326 4814 4378
rect 4826 4326 4878 4378
rect 4890 4326 4942 4378
rect 4954 4326 5006 4378
rect 8446 4326 8498 4378
rect 8510 4326 8562 4378
rect 8574 4326 8626 4378
rect 8638 4326 8690 4378
rect 8702 4326 8754 4378
rect 12194 4326 12246 4378
rect 12258 4326 12310 4378
rect 12322 4326 12374 4378
rect 12386 4326 12438 4378
rect 12450 4326 12502 4378
rect 7748 4088 7800 4140
rect 12716 4088 12768 4140
rect 9220 4020 9272 4072
rect 10140 4020 10192 4072
rect 6368 3952 6420 4004
rect 9772 3952 9824 4004
rect 2824 3782 2876 3834
rect 2888 3782 2940 3834
rect 2952 3782 3004 3834
rect 3016 3782 3068 3834
rect 3080 3782 3132 3834
rect 6572 3782 6624 3834
rect 6636 3782 6688 3834
rect 6700 3782 6752 3834
rect 6764 3782 6816 3834
rect 6828 3782 6880 3834
rect 10320 3782 10372 3834
rect 10384 3782 10436 3834
rect 10448 3782 10500 3834
rect 10512 3782 10564 3834
rect 10576 3782 10628 3834
rect 14068 3782 14120 3834
rect 14132 3782 14184 3834
rect 14196 3782 14248 3834
rect 14260 3782 14312 3834
rect 14324 3782 14376 3834
rect 4698 3238 4750 3290
rect 4762 3238 4814 3290
rect 4826 3238 4878 3290
rect 4890 3238 4942 3290
rect 4954 3238 5006 3290
rect 8446 3238 8498 3290
rect 8510 3238 8562 3290
rect 8574 3238 8626 3290
rect 8638 3238 8690 3290
rect 8702 3238 8754 3290
rect 12194 3238 12246 3290
rect 12258 3238 12310 3290
rect 12322 3238 12374 3290
rect 12386 3238 12438 3290
rect 12450 3238 12502 3290
rect 3424 3136 3476 3188
rect 8760 3136 8812 3188
rect 13084 3136 13136 3188
rect 13360 3136 13412 3188
rect 3332 3068 3384 3120
rect 1860 3043 1912 3052
rect 1860 3009 1869 3043
rect 1869 3009 1903 3043
rect 1903 3009 1912 3043
rect 1860 3000 1912 3009
rect 6460 3000 6512 3052
rect 15752 3000 15804 3052
rect 8668 2932 8720 2984
rect 10876 2932 10928 2984
rect 1400 2796 1452 2848
rect 3976 2796 4028 2848
rect 8852 2839 8904 2848
rect 8852 2805 8861 2839
rect 8861 2805 8895 2839
rect 8895 2805 8904 2839
rect 8852 2796 8904 2805
rect 9128 2839 9180 2848
rect 9128 2805 9137 2839
rect 9137 2805 9171 2839
rect 9171 2805 9180 2839
rect 9128 2796 9180 2805
rect 9496 2839 9548 2848
rect 9496 2805 9505 2839
rect 9505 2805 9539 2839
rect 9539 2805 9548 2839
rect 9496 2796 9548 2805
rect 9864 2839 9916 2848
rect 9864 2805 9873 2839
rect 9873 2805 9907 2839
rect 9907 2805 9916 2839
rect 9864 2796 9916 2805
rect 10232 2839 10284 2848
rect 10232 2805 10241 2839
rect 10241 2805 10275 2839
rect 10275 2805 10284 2839
rect 10232 2796 10284 2805
rect 10692 2796 10744 2848
rect 10968 2839 11020 2848
rect 10968 2805 10977 2839
rect 10977 2805 11011 2839
rect 11011 2805 11020 2839
rect 10968 2796 11020 2805
rect 11336 2796 11388 2848
rect 11796 2839 11848 2848
rect 11796 2805 11805 2839
rect 11805 2805 11839 2839
rect 11839 2805 11848 2839
rect 11796 2796 11848 2805
rect 12072 2839 12124 2848
rect 12072 2805 12081 2839
rect 12081 2805 12115 2839
rect 12115 2805 12124 2839
rect 12072 2796 12124 2805
rect 12532 2796 12584 2848
rect 12808 2839 12860 2848
rect 12808 2805 12817 2839
rect 12817 2805 12851 2839
rect 12851 2805 12860 2839
rect 12808 2796 12860 2805
rect 13176 2839 13228 2848
rect 13176 2805 13185 2839
rect 13185 2805 13219 2839
rect 13219 2805 13228 2839
rect 13176 2796 13228 2805
rect 13820 2796 13872 2848
rect 13912 2839 13964 2848
rect 13912 2805 13921 2839
rect 13921 2805 13955 2839
rect 13955 2805 13964 2839
rect 13912 2796 13964 2805
rect 14464 2796 14516 2848
rect 14648 2839 14700 2848
rect 14648 2805 14657 2839
rect 14657 2805 14691 2839
rect 14691 2805 14700 2839
rect 14648 2796 14700 2805
rect 15016 2839 15068 2848
rect 15016 2805 15025 2839
rect 15025 2805 15059 2839
rect 15059 2805 15068 2839
rect 15016 2796 15068 2805
rect 15384 2796 15436 2848
rect 2824 2694 2876 2746
rect 2888 2694 2940 2746
rect 2952 2694 3004 2746
rect 3016 2694 3068 2746
rect 3080 2694 3132 2746
rect 6572 2694 6624 2746
rect 6636 2694 6688 2746
rect 6700 2694 6752 2746
rect 6764 2694 6816 2746
rect 6828 2694 6880 2746
rect 10320 2694 10372 2746
rect 10384 2694 10436 2746
rect 10448 2694 10500 2746
rect 10512 2694 10564 2746
rect 10576 2694 10628 2746
rect 14068 2694 14120 2746
rect 14132 2694 14184 2746
rect 14196 2694 14248 2746
rect 14260 2694 14312 2746
rect 14324 2694 14376 2746
rect 4620 2592 4672 2644
rect 7196 2592 7248 2644
rect 9588 2635 9640 2644
rect 9588 2601 9597 2635
rect 9597 2601 9631 2635
rect 9631 2601 9640 2635
rect 9588 2592 9640 2601
rect 9772 2592 9824 2644
rect 10140 2592 10192 2644
rect 11520 2592 11572 2644
rect 12624 2592 12676 2644
rect 12900 2635 12952 2644
rect 12900 2601 12909 2635
rect 12909 2601 12943 2635
rect 12943 2601 12952 2635
rect 12900 2592 12952 2601
rect 12992 2592 13044 2644
rect 3700 2524 3752 2576
rect 2780 2388 2832 2440
rect 4160 2456 4212 2508
rect 3516 2388 3568 2440
rect 4344 2431 4396 2440
rect 4344 2397 4353 2431
rect 4353 2397 4387 2431
rect 4387 2397 4396 2431
rect 4344 2388 4396 2397
rect 8300 2524 8352 2576
rect 11704 2524 11756 2576
rect 11980 2524 12032 2576
rect 5172 2388 5224 2440
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 6460 2388 6512 2440
rect 4988 2320 5040 2372
rect 7472 2388 7524 2440
rect 7656 2431 7708 2440
rect 7656 2397 7665 2431
rect 7665 2397 7699 2431
rect 7699 2397 7708 2431
rect 7656 2388 7708 2397
rect 11612 2456 11664 2508
rect 11888 2456 11940 2508
rect 8760 2431 8812 2440
rect 8760 2397 8769 2431
rect 8769 2397 8803 2431
rect 8803 2397 8812 2431
rect 8760 2388 8812 2397
rect 8668 2320 8720 2372
rect 8852 2320 8904 2372
rect 9220 2388 9272 2440
rect 9680 2388 9732 2440
rect 9864 2388 9916 2440
rect 10232 2388 10284 2440
rect 10600 2388 10652 2440
rect 11060 2388 11112 2440
rect 11336 2388 11388 2440
rect 11796 2388 11848 2440
rect 12072 2388 12124 2440
rect 12532 2388 12584 2440
rect 12808 2388 12860 2440
rect 13176 2388 13228 2440
rect 13820 2431 13872 2440
rect 13820 2397 13829 2431
rect 13829 2397 13863 2431
rect 13863 2397 13872 2431
rect 13820 2388 13872 2397
rect 13912 2388 13964 2440
rect 14372 2388 14424 2440
rect 14648 2388 14700 2440
rect 15200 2388 15252 2440
rect 15384 2388 15436 2440
rect 10784 2320 10836 2372
rect 1768 2252 1820 2304
rect 2136 2252 2188 2304
rect 2504 2252 2556 2304
rect 2872 2252 2924 2304
rect 3240 2252 3292 2304
rect 3608 2252 3660 2304
rect 4344 2252 4396 2304
rect 4620 2252 4672 2304
rect 5080 2252 5132 2304
rect 5448 2252 5500 2304
rect 5816 2252 5868 2304
rect 6184 2252 6236 2304
rect 6552 2252 6604 2304
rect 6920 2252 6972 2304
rect 7288 2252 7340 2304
rect 7656 2252 7708 2304
rect 8024 2252 8076 2304
rect 8300 2252 8352 2304
rect 9220 2295 9272 2304
rect 9220 2261 9229 2295
rect 9229 2261 9263 2295
rect 9263 2261 9272 2295
rect 9220 2252 9272 2261
rect 10692 2295 10744 2304
rect 10692 2261 10701 2295
rect 10701 2261 10735 2295
rect 10735 2261 10744 2295
rect 10692 2252 10744 2261
rect 11060 2295 11112 2304
rect 11060 2261 11069 2295
rect 11069 2261 11103 2295
rect 11103 2261 11112 2295
rect 11060 2252 11112 2261
rect 11520 2295 11572 2304
rect 11520 2261 11529 2295
rect 11529 2261 11563 2295
rect 11563 2261 11572 2295
rect 11520 2252 11572 2261
rect 11980 2252 12032 2304
rect 13728 2252 13780 2304
rect 14740 2295 14792 2304
rect 14740 2261 14749 2295
rect 14749 2261 14783 2295
rect 14783 2261 14792 2295
rect 14740 2252 14792 2261
rect 15108 2295 15160 2304
rect 15108 2261 15117 2295
rect 15117 2261 15151 2295
rect 15151 2261 15160 2295
rect 15108 2252 15160 2261
rect 4698 2150 4750 2202
rect 4762 2150 4814 2202
rect 4826 2150 4878 2202
rect 4890 2150 4942 2202
rect 4954 2150 5006 2202
rect 8446 2150 8498 2202
rect 8510 2150 8562 2202
rect 8574 2150 8626 2202
rect 8638 2150 8690 2202
rect 8702 2150 8754 2202
rect 12194 2150 12246 2202
rect 12258 2150 12310 2202
rect 12322 2150 12374 2202
rect 12386 2150 12438 2202
rect 12450 2150 12502 2202
rect 5540 2048 5592 2100
rect 10692 2048 10744 2100
rect 11152 2048 11204 2100
rect 15108 2048 15160 2100
rect 3516 1980 3568 2032
rect 6000 1980 6052 2032
rect 7472 1980 7524 2032
rect 11428 1980 11480 2032
rect 5356 1912 5408 1964
rect 9220 1912 9272 1964
rect 9312 1912 9364 1964
rect 14740 1912 14792 1964
rect 2780 1844 2832 1896
rect 5724 1844 5776 1896
rect 9036 1844 9088 1896
rect 11980 1844 12032 1896
rect 6460 1776 6512 1828
rect 7380 1776 7432 1828
rect 11060 1776 11112 1828
rect 10048 1708 10100 1760
<< metal2 >>
rect 1214 19200 1270 20000
rect 1582 19200 1638 20000
rect 1950 19200 2006 20000
rect 2318 19200 2374 20000
rect 2686 19200 2742 20000
rect 3054 19200 3110 20000
rect 3422 19200 3478 20000
rect 3790 19200 3846 20000
rect 4158 19200 4214 20000
rect 4526 19200 4582 20000
rect 4894 19200 4950 20000
rect 5262 19200 5318 20000
rect 5630 19200 5686 20000
rect 5998 19200 6054 20000
rect 6366 19200 6422 20000
rect 6734 19200 6790 20000
rect 7102 19200 7158 20000
rect 7470 19200 7526 20000
rect 7838 19200 7894 20000
rect 8206 19200 8262 20000
rect 8574 19200 8630 20000
rect 8680 19230 8892 19258
rect 1228 16574 1256 19200
rect 1596 17338 1624 19200
rect 1674 18184 1730 18193
rect 1674 18119 1730 18128
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1688 16590 1716 18119
rect 1964 17338 1992 19200
rect 2332 17338 2360 19200
rect 2700 17338 2728 19200
rect 3068 17338 3096 19200
rect 3436 17338 3464 19200
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 2320 17332 2372 17338
rect 2320 17274 2372 17280
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 3608 17196 3660 17202
rect 3608 17138 3660 17144
rect 1308 16584 1360 16590
rect 1228 16546 1308 16574
rect 1308 16526 1360 16532
rect 1676 16584 1728 16590
rect 1676 16526 1728 16532
rect 1320 16250 1348 16526
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1596 16250 1624 16390
rect 1308 16244 1360 16250
rect 1308 16186 1360 16192
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1490 14920 1546 14929
rect 1490 14855 1546 14864
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1412 11665 1440 11698
rect 1398 11656 1454 11665
rect 1398 11591 1454 11600
rect 1504 9654 1532 14855
rect 1492 9648 1544 9654
rect 1492 9590 1544 9596
rect 2148 9450 2176 17138
rect 2516 12442 2544 17138
rect 3148 17128 3200 17134
rect 3148 17070 3200 17076
rect 2824 16892 3132 16901
rect 2824 16890 2830 16892
rect 2886 16890 2910 16892
rect 2966 16890 2990 16892
rect 3046 16890 3070 16892
rect 3126 16890 3132 16892
rect 2886 16838 2888 16890
rect 3068 16838 3070 16890
rect 2824 16836 2830 16838
rect 2886 16836 2910 16838
rect 2966 16836 2990 16838
rect 3046 16836 3070 16838
rect 3126 16836 3132 16838
rect 2824 16827 3132 16836
rect 2824 15804 3132 15813
rect 2824 15802 2830 15804
rect 2886 15802 2910 15804
rect 2966 15802 2990 15804
rect 3046 15802 3070 15804
rect 3126 15802 3132 15804
rect 2886 15750 2888 15802
rect 3068 15750 3070 15802
rect 2824 15748 2830 15750
rect 2886 15748 2910 15750
rect 2966 15748 2990 15750
rect 3046 15748 3070 15750
rect 3126 15748 3132 15750
rect 2824 15739 3132 15748
rect 2824 14716 3132 14725
rect 2824 14714 2830 14716
rect 2886 14714 2910 14716
rect 2966 14714 2990 14716
rect 3046 14714 3070 14716
rect 3126 14714 3132 14716
rect 2886 14662 2888 14714
rect 3068 14662 3070 14714
rect 2824 14660 2830 14662
rect 2886 14660 2910 14662
rect 2966 14660 2990 14662
rect 3046 14660 3070 14662
rect 3126 14660 3132 14662
rect 2824 14651 3132 14660
rect 2824 13628 3132 13637
rect 2824 13626 2830 13628
rect 2886 13626 2910 13628
rect 2966 13626 2990 13628
rect 3046 13626 3070 13628
rect 3126 13626 3132 13628
rect 2886 13574 2888 13626
rect 3068 13574 3070 13626
rect 2824 13572 2830 13574
rect 2886 13572 2910 13574
rect 2966 13572 2990 13574
rect 3046 13572 3070 13574
rect 3126 13572 3132 13574
rect 2824 13563 3132 13572
rect 3160 12986 3188 17070
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 2824 12540 3132 12549
rect 2824 12538 2830 12540
rect 2886 12538 2910 12540
rect 2966 12538 2990 12540
rect 3046 12538 3070 12540
rect 3126 12538 3132 12540
rect 2886 12486 2888 12538
rect 3068 12486 3070 12538
rect 2824 12484 2830 12486
rect 2886 12484 2910 12486
rect 2966 12484 2990 12486
rect 3046 12484 3070 12486
rect 3126 12484 3132 12486
rect 2824 12475 3132 12484
rect 2504 12436 2556 12442
rect 2504 12378 2556 12384
rect 2824 11452 3132 11461
rect 2824 11450 2830 11452
rect 2886 11450 2910 11452
rect 2966 11450 2990 11452
rect 3046 11450 3070 11452
rect 3126 11450 3132 11452
rect 2886 11398 2888 11450
rect 3068 11398 3070 11450
rect 2824 11396 2830 11398
rect 2886 11396 2910 11398
rect 2966 11396 2990 11398
rect 3046 11396 3070 11398
rect 3126 11396 3132 11398
rect 2824 11387 3132 11396
rect 3528 10674 3556 13806
rect 3620 10742 3648 17138
rect 3804 16454 3832 19200
rect 4172 17338 4200 19200
rect 4540 17338 4568 19200
rect 4908 17626 4936 19200
rect 4908 17598 5120 17626
rect 4698 17436 5006 17445
rect 4698 17434 4704 17436
rect 4760 17434 4784 17436
rect 4840 17434 4864 17436
rect 4920 17434 4944 17436
rect 5000 17434 5006 17436
rect 4760 17382 4762 17434
rect 4942 17382 4944 17434
rect 4698 17380 4704 17382
rect 4760 17380 4784 17382
rect 4840 17380 4864 17382
rect 4920 17380 4944 17382
rect 5000 17380 5006 17382
rect 4698 17371 5006 17380
rect 5092 17338 5120 17598
rect 5276 17338 5304 19200
rect 5644 17338 5672 19200
rect 6012 17338 6040 19200
rect 6380 17338 6408 19200
rect 6748 17898 6776 19200
rect 6748 17870 6960 17898
rect 6932 17338 6960 17870
rect 7116 17338 7144 19200
rect 7484 17338 7512 19200
rect 7852 17338 7880 19200
rect 8220 17354 8248 19200
rect 8588 19122 8616 19200
rect 8680 19122 8708 19230
rect 8588 19094 8708 19122
rect 8446 17436 8754 17445
rect 8446 17434 8452 17436
rect 8508 17434 8532 17436
rect 8588 17434 8612 17436
rect 8668 17434 8692 17436
rect 8748 17434 8754 17436
rect 8508 17382 8510 17434
rect 8690 17382 8692 17434
rect 8446 17380 8452 17382
rect 8508 17380 8532 17382
rect 8588 17380 8612 17382
rect 8668 17380 8692 17382
rect 8748 17380 8754 17382
rect 8446 17371 8754 17380
rect 8220 17338 8340 17354
rect 8864 17338 8892 19230
rect 8942 19200 8998 20000
rect 9310 19200 9366 20000
rect 9678 19200 9734 20000
rect 10046 19200 10102 20000
rect 10414 19200 10470 20000
rect 10782 19200 10838 20000
rect 11150 19200 11206 20000
rect 11518 19200 11574 20000
rect 11886 19200 11942 20000
rect 12254 19200 12310 20000
rect 12622 19200 12678 20000
rect 12990 19200 13046 20000
rect 13358 19200 13414 20000
rect 13726 19200 13782 20000
rect 14094 19200 14150 20000
rect 14462 19200 14518 20000
rect 14830 19200 14886 20000
rect 15198 19200 15254 20000
rect 15566 19200 15622 20000
rect 15934 19200 15990 20000
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4528 17332 4580 17338
rect 4528 17274 4580 17280
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5632 17332 5684 17338
rect 5632 17274 5684 17280
rect 6000 17332 6052 17338
rect 6000 17274 6052 17280
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7472 17332 7524 17338
rect 7472 17274 7524 17280
rect 7840 17332 7892 17338
rect 8220 17332 8352 17338
rect 8220 17326 8300 17332
rect 7840 17274 7892 17280
rect 8300 17274 8352 17280
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4356 16998 4384 17138
rect 4436 17128 4488 17134
rect 4436 17070 4488 17076
rect 4344 16992 4396 16998
rect 4344 16934 4396 16940
rect 4068 16584 4120 16590
rect 4120 16544 4200 16572
rect 4068 16526 4120 16532
rect 3792 16448 3844 16454
rect 3792 16390 3844 16396
rect 4172 12918 4200 16544
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4356 11218 4384 12718
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 3608 10736 3660 10742
rect 3608 10678 3660 10684
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 2824 10364 3132 10373
rect 2824 10362 2830 10364
rect 2886 10362 2910 10364
rect 2966 10362 2990 10364
rect 3046 10362 3070 10364
rect 3126 10362 3132 10364
rect 2886 10310 2888 10362
rect 3068 10310 3070 10362
rect 2824 10308 2830 10310
rect 2886 10308 2910 10310
rect 2966 10308 2990 10310
rect 3046 10308 3070 10310
rect 3126 10308 3132 10310
rect 2824 10299 3132 10308
rect 3240 10192 3292 10198
rect 3240 10134 3292 10140
rect 2136 9444 2188 9450
rect 2136 9386 2188 9392
rect 2824 9276 3132 9285
rect 2824 9274 2830 9276
rect 2886 9274 2910 9276
rect 2966 9274 2990 9276
rect 3046 9274 3070 9276
rect 3126 9274 3132 9276
rect 2886 9222 2888 9274
rect 3068 9222 3070 9274
rect 2824 9220 2830 9222
rect 2886 9220 2910 9222
rect 2966 9220 2990 9222
rect 3046 9220 3070 9222
rect 3126 9220 3132 9222
rect 2824 9211 3132 9220
rect 1490 8392 1546 8401
rect 1490 8327 1492 8336
rect 1544 8327 1546 8336
rect 1492 8298 1544 8304
rect 2824 8188 3132 8197
rect 2824 8186 2830 8188
rect 2886 8186 2910 8188
rect 2966 8186 2990 8188
rect 3046 8186 3070 8188
rect 3126 8186 3132 8188
rect 2886 8134 2888 8186
rect 3068 8134 3070 8186
rect 2824 8132 2830 8134
rect 2886 8132 2910 8134
rect 2966 8132 2990 8134
rect 3046 8132 3070 8134
rect 3126 8132 3132 8134
rect 2824 8123 3132 8132
rect 3252 7410 3280 10134
rect 3528 9654 3556 10610
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3516 9648 3568 9654
rect 3516 9590 3568 9596
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 2824 7100 3132 7109
rect 2824 7098 2830 7100
rect 2886 7098 2910 7100
rect 2966 7098 2990 7100
rect 3046 7098 3070 7100
rect 3126 7098 3132 7100
rect 2886 7046 2888 7098
rect 3068 7046 3070 7098
rect 2824 7044 2830 7046
rect 2886 7044 2910 7046
rect 2966 7044 2990 7046
rect 3046 7044 3070 7046
rect 3126 7044 3132 7046
rect 2824 7035 3132 7044
rect 2824 6012 3132 6021
rect 2824 6010 2830 6012
rect 2886 6010 2910 6012
rect 2966 6010 2990 6012
rect 3046 6010 3070 6012
rect 3126 6010 3132 6012
rect 2886 5958 2888 6010
rect 3068 5958 3070 6010
rect 2824 5956 2830 5958
rect 2886 5956 2910 5958
rect 2966 5956 2990 5958
rect 3046 5956 3070 5958
rect 3126 5956 3132 5958
rect 2824 5947 3132 5956
rect 3160 5234 3188 7142
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 1490 5128 1546 5137
rect 1490 5063 1492 5072
rect 1544 5063 1546 5072
rect 1492 5034 1544 5040
rect 2824 4924 3132 4933
rect 2824 4922 2830 4924
rect 2886 4922 2910 4924
rect 2966 4922 2990 4924
rect 3046 4922 3070 4924
rect 3126 4922 3132 4924
rect 2886 4870 2888 4922
rect 3068 4870 3070 4922
rect 2824 4868 2830 4870
rect 2886 4868 2910 4870
rect 2966 4868 2990 4870
rect 3046 4868 3070 4870
rect 3126 4868 3132 4870
rect 2824 4859 3132 4868
rect 2824 3836 3132 3845
rect 2824 3834 2830 3836
rect 2886 3834 2910 3836
rect 2966 3834 2990 3836
rect 3046 3834 3070 3836
rect 3126 3834 3132 3836
rect 2886 3782 2888 3834
rect 3068 3782 3070 3834
rect 2824 3780 2830 3782
rect 2886 3780 2910 3782
rect 2966 3780 2990 3782
rect 3046 3780 3070 3782
rect 3126 3780 3132 3782
rect 2824 3771 3132 3780
rect 3344 3126 3372 7142
rect 3436 3194 3464 9454
rect 3528 8498 3556 9590
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3332 3120 3384 3126
rect 3332 3062 3384 3068
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1412 800 1440 2790
rect 1768 2304 1820 2310
rect 1768 2246 1820 2252
rect 1780 800 1808 2246
rect 1872 1873 1900 2994
rect 2824 2748 3132 2757
rect 2824 2746 2830 2748
rect 2886 2746 2910 2748
rect 2966 2746 2990 2748
rect 3046 2746 3070 2748
rect 3126 2746 3132 2748
rect 2886 2694 2888 2746
rect 3068 2694 3070 2746
rect 2824 2692 2830 2694
rect 2886 2692 2910 2694
rect 2966 2692 2990 2694
rect 3046 2692 3070 2694
rect 3126 2692 3132 2694
rect 2824 2683 3132 2692
rect 3712 2582 3740 9862
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 3700 2576 3752 2582
rect 3700 2518 3752 2524
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 1858 1864 1914 1873
rect 1858 1799 1914 1808
rect 2148 800 2176 2246
rect 2516 800 2544 2246
rect 2792 1902 2820 2382
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 2780 1896 2832 1902
rect 2780 1838 2832 1844
rect 2884 800 2912 2246
rect 3252 800 3280 2246
rect 3528 2038 3556 2382
rect 3608 2304 3660 2310
rect 3608 2246 3660 2252
rect 3516 2032 3568 2038
rect 3516 1974 3568 1980
rect 3620 800 3648 2246
rect 3988 800 4016 2790
rect 4172 2514 4200 7482
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 4356 2446 4384 11018
rect 4448 9489 4476 17070
rect 4632 16726 4660 17206
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6276 17196 6328 17202
rect 6276 17138 6328 17144
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 8852 17196 8904 17202
rect 8852 17138 8904 17144
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 4620 16720 4672 16726
rect 4620 16662 4672 16668
rect 4698 16348 5006 16357
rect 4698 16346 4704 16348
rect 4760 16346 4784 16348
rect 4840 16346 4864 16348
rect 4920 16346 4944 16348
rect 5000 16346 5006 16348
rect 4760 16294 4762 16346
rect 4942 16294 4944 16346
rect 4698 16292 4704 16294
rect 4760 16292 4784 16294
rect 4840 16292 4864 16294
rect 4920 16292 4944 16294
rect 5000 16292 5006 16294
rect 4698 16283 5006 16292
rect 5080 16244 5132 16250
rect 5080 16186 5132 16192
rect 4698 15260 5006 15269
rect 4698 15258 4704 15260
rect 4760 15258 4784 15260
rect 4840 15258 4864 15260
rect 4920 15258 4944 15260
rect 5000 15258 5006 15260
rect 4760 15206 4762 15258
rect 4942 15206 4944 15258
rect 4698 15204 4704 15206
rect 4760 15204 4784 15206
rect 4840 15204 4864 15206
rect 4920 15204 4944 15206
rect 5000 15204 5006 15206
rect 4698 15195 5006 15204
rect 4698 14172 5006 14181
rect 4698 14170 4704 14172
rect 4760 14170 4784 14172
rect 4840 14170 4864 14172
rect 4920 14170 4944 14172
rect 5000 14170 5006 14172
rect 4760 14118 4762 14170
rect 4942 14118 4944 14170
rect 4698 14116 4704 14118
rect 4760 14116 4784 14118
rect 4840 14116 4864 14118
rect 4920 14116 4944 14118
rect 5000 14116 5006 14118
rect 4698 14107 5006 14116
rect 5092 13938 5120 16186
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 4698 13084 5006 13093
rect 4698 13082 4704 13084
rect 4760 13082 4784 13084
rect 4840 13082 4864 13084
rect 4920 13082 4944 13084
rect 5000 13082 5006 13084
rect 4760 13030 4762 13082
rect 4942 13030 4944 13082
rect 4698 13028 4704 13030
rect 4760 13028 4784 13030
rect 4840 13028 4864 13030
rect 4920 13028 4944 13030
rect 5000 13028 5006 13030
rect 4698 13019 5006 13028
rect 4698 11996 5006 12005
rect 4698 11994 4704 11996
rect 4760 11994 4784 11996
rect 4840 11994 4864 11996
rect 4920 11994 4944 11996
rect 5000 11994 5006 11996
rect 4760 11942 4762 11994
rect 4942 11942 4944 11994
rect 4698 11940 4704 11942
rect 4760 11940 4784 11942
rect 4840 11940 4864 11942
rect 4920 11940 4944 11942
rect 5000 11940 5006 11942
rect 4698 11931 5006 11940
rect 4698 10908 5006 10917
rect 4698 10906 4704 10908
rect 4760 10906 4784 10908
rect 4840 10906 4864 10908
rect 4920 10906 4944 10908
rect 5000 10906 5006 10908
rect 4760 10854 4762 10906
rect 4942 10854 4944 10906
rect 4698 10852 4704 10854
rect 4760 10852 4784 10854
rect 4840 10852 4864 10854
rect 4920 10852 4944 10854
rect 5000 10852 5006 10854
rect 4698 10843 5006 10852
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 4698 9820 5006 9829
rect 4698 9818 4704 9820
rect 4760 9818 4784 9820
rect 4840 9818 4864 9820
rect 4920 9818 4944 9820
rect 5000 9818 5006 9820
rect 4760 9766 4762 9818
rect 4942 9766 4944 9818
rect 4698 9764 4704 9766
rect 4760 9764 4784 9766
rect 4840 9764 4864 9766
rect 4920 9764 4944 9766
rect 5000 9764 5006 9766
rect 4698 9755 5006 9764
rect 4434 9480 4490 9489
rect 4434 9415 4490 9424
rect 4698 8732 5006 8741
rect 4698 8730 4704 8732
rect 4760 8730 4784 8732
rect 4840 8730 4864 8732
rect 4920 8730 4944 8732
rect 5000 8730 5006 8732
rect 4760 8678 4762 8730
rect 4942 8678 4944 8730
rect 4698 8676 4704 8678
rect 4760 8676 4784 8678
rect 4840 8676 4864 8678
rect 4920 8676 4944 8678
rect 5000 8676 5006 8678
rect 4698 8667 5006 8676
rect 4698 7644 5006 7653
rect 4698 7642 4704 7644
rect 4760 7642 4784 7644
rect 4840 7642 4864 7644
rect 4920 7642 4944 7644
rect 5000 7642 5006 7644
rect 4760 7590 4762 7642
rect 4942 7590 4944 7642
rect 4698 7588 4704 7590
rect 4760 7588 4784 7590
rect 4840 7588 4864 7590
rect 4920 7588 4944 7590
rect 5000 7588 5006 7590
rect 4698 7579 5006 7588
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4632 2650 4660 7142
rect 4698 6556 5006 6565
rect 4698 6554 4704 6556
rect 4760 6554 4784 6556
rect 4840 6554 4864 6556
rect 4920 6554 4944 6556
rect 5000 6554 5006 6556
rect 4760 6502 4762 6554
rect 4942 6502 4944 6554
rect 4698 6500 4704 6502
rect 4760 6500 4784 6502
rect 4840 6500 4864 6502
rect 4920 6500 4944 6502
rect 5000 6500 5006 6502
rect 4698 6491 5006 6500
rect 4698 5468 5006 5477
rect 4698 5466 4704 5468
rect 4760 5466 4784 5468
rect 4840 5466 4864 5468
rect 4920 5466 4944 5468
rect 5000 5466 5006 5468
rect 4760 5414 4762 5466
rect 4942 5414 4944 5466
rect 4698 5412 4704 5414
rect 4760 5412 4784 5414
rect 4840 5412 4864 5414
rect 4920 5412 4944 5414
rect 5000 5412 5006 5414
rect 4698 5403 5006 5412
rect 4698 4380 5006 4389
rect 4698 4378 4704 4380
rect 4760 4378 4784 4380
rect 4840 4378 4864 4380
rect 4920 4378 4944 4380
rect 5000 4378 5006 4380
rect 4760 4326 4762 4378
rect 4942 4326 4944 4378
rect 4698 4324 4704 4326
rect 4760 4324 4784 4326
rect 4840 4324 4864 4326
rect 4920 4324 4944 4326
rect 5000 4324 5006 4326
rect 4698 4315 5006 4324
rect 4698 3292 5006 3301
rect 4698 3290 4704 3292
rect 4760 3290 4784 3292
rect 4840 3290 4864 3292
rect 4920 3290 4944 3292
rect 5000 3290 5006 3292
rect 4760 3238 4762 3290
rect 4942 3238 4944 3290
rect 4698 3236 4704 3238
rect 4760 3236 4784 3238
rect 4840 3236 4864 3238
rect 4920 3236 4944 3238
rect 5000 3236 5006 3238
rect 4698 3227 5006 3236
rect 5092 2774 5120 10474
rect 5276 10062 5304 16730
rect 5460 12442 5488 17138
rect 5724 17060 5776 17066
rect 5724 17002 5776 17008
rect 5540 16720 5592 16726
rect 5540 16662 5592 16668
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5552 10810 5580 16662
rect 5736 12986 5764 17002
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5552 10198 5580 10610
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5172 7268 5224 7274
rect 5172 7210 5224 7216
rect 5000 2746 5120 2774
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 5000 2378 5028 2746
rect 5184 2446 5212 7210
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 4344 2304 4396 2310
rect 4344 2246 4396 2252
rect 4620 2304 4672 2310
rect 4620 2246 4672 2252
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 4356 800 4384 2246
rect 4632 1170 4660 2246
rect 4698 2204 5006 2213
rect 4698 2202 4704 2204
rect 4760 2202 4784 2204
rect 4840 2202 4864 2204
rect 4920 2202 4944 2204
rect 5000 2202 5006 2204
rect 4760 2150 4762 2202
rect 4942 2150 4944 2202
rect 4698 2148 4704 2150
rect 4760 2148 4784 2150
rect 4840 2148 4864 2150
rect 4920 2148 4944 2150
rect 5000 2148 5006 2150
rect 4698 2139 5006 2148
rect 4632 1142 4752 1170
rect 4724 800 4752 1142
rect 5092 800 5120 2246
rect 5368 1970 5396 9522
rect 5552 8634 5580 9862
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5644 2774 5672 10542
rect 5736 10130 5764 11630
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5828 10130 5856 10406
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5920 10062 5948 11494
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5828 9722 5856 9930
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 6012 9466 6040 10610
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 5828 9438 6040 9466
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5552 2746 5672 2774
rect 5446 2544 5502 2553
rect 5446 2479 5502 2488
rect 5460 2446 5488 2479
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5356 1964 5408 1970
rect 5356 1906 5408 1912
rect 5460 800 5488 2246
rect 5552 2106 5580 2746
rect 5540 2100 5592 2106
rect 5540 2042 5592 2048
rect 5736 1902 5764 9318
rect 5828 2446 5856 9438
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5724 1896 5776 1902
rect 5724 1838 5776 1844
rect 5828 800 5856 2246
rect 6012 2038 6040 9318
rect 6104 8974 6132 9522
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6196 8838 6224 17138
rect 6288 9761 6316 17138
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 6380 11626 6408 16934
rect 6472 11830 6500 17070
rect 6572 16892 6880 16901
rect 6572 16890 6578 16892
rect 6634 16890 6658 16892
rect 6714 16890 6738 16892
rect 6794 16890 6818 16892
rect 6874 16890 6880 16892
rect 6634 16838 6636 16890
rect 6816 16838 6818 16890
rect 6572 16836 6578 16838
rect 6634 16836 6658 16838
rect 6714 16836 6738 16838
rect 6794 16836 6818 16838
rect 6874 16836 6880 16838
rect 6572 16827 6880 16836
rect 7196 16584 7248 16590
rect 7196 16526 7248 16532
rect 6572 15804 6880 15813
rect 6572 15802 6578 15804
rect 6634 15802 6658 15804
rect 6714 15802 6738 15804
rect 6794 15802 6818 15804
rect 6874 15802 6880 15804
rect 6634 15750 6636 15802
rect 6816 15750 6818 15802
rect 6572 15748 6578 15750
rect 6634 15748 6658 15750
rect 6714 15748 6738 15750
rect 6794 15748 6818 15750
rect 6874 15748 6880 15750
rect 6572 15739 6880 15748
rect 6572 14716 6880 14725
rect 6572 14714 6578 14716
rect 6634 14714 6658 14716
rect 6714 14714 6738 14716
rect 6794 14714 6818 14716
rect 6874 14714 6880 14716
rect 6634 14662 6636 14714
rect 6816 14662 6818 14714
rect 6572 14660 6578 14662
rect 6634 14660 6658 14662
rect 6714 14660 6738 14662
rect 6794 14660 6818 14662
rect 6874 14660 6880 14662
rect 6572 14651 6880 14660
rect 6572 13628 6880 13637
rect 6572 13626 6578 13628
rect 6634 13626 6658 13628
rect 6714 13626 6738 13628
rect 6794 13626 6818 13628
rect 6874 13626 6880 13628
rect 6634 13574 6636 13626
rect 6816 13574 6818 13626
rect 6572 13572 6578 13574
rect 6634 13572 6658 13574
rect 6714 13572 6738 13574
rect 6794 13572 6818 13574
rect 6874 13572 6880 13574
rect 6572 13563 6880 13572
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 6572 12540 6880 12549
rect 6572 12538 6578 12540
rect 6634 12538 6658 12540
rect 6714 12538 6738 12540
rect 6794 12538 6818 12540
rect 6874 12538 6880 12540
rect 6634 12486 6636 12538
rect 6816 12486 6818 12538
rect 6572 12484 6578 12486
rect 6634 12484 6658 12486
rect 6714 12484 6738 12486
rect 6794 12484 6818 12486
rect 6874 12484 6880 12486
rect 6572 12475 6880 12484
rect 6460 11824 6512 11830
rect 6460 11766 6512 11772
rect 6368 11620 6420 11626
rect 6368 11562 6420 11568
rect 7024 11506 7052 12650
rect 7116 11642 7144 12718
rect 7208 11898 7236 16526
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7116 11614 7236 11642
rect 7024 11478 7144 11506
rect 6572 11452 6880 11461
rect 6572 11450 6578 11452
rect 6634 11450 6658 11452
rect 6714 11450 6738 11452
rect 6794 11450 6818 11452
rect 6874 11450 6880 11452
rect 6634 11398 6636 11450
rect 6816 11398 6818 11450
rect 6572 11396 6578 11398
rect 6634 11396 6658 11398
rect 6714 11396 6738 11398
rect 6794 11396 6818 11398
rect 6874 11396 6880 11398
rect 6572 11387 6880 11396
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6826 10704 6882 10713
rect 6826 10639 6828 10648
rect 6880 10639 6882 10648
rect 6828 10610 6880 10616
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6368 10192 6420 10198
rect 6368 10134 6420 10140
rect 6274 9752 6330 9761
rect 6274 9687 6330 9696
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6380 4010 6408 10134
rect 6368 4004 6420 4010
rect 6368 3946 6420 3952
rect 6472 3058 6500 10406
rect 6572 10364 6880 10373
rect 6572 10362 6578 10364
rect 6634 10362 6658 10364
rect 6714 10362 6738 10364
rect 6794 10362 6818 10364
rect 6874 10362 6880 10364
rect 6634 10310 6636 10362
rect 6816 10310 6818 10362
rect 6572 10308 6578 10310
rect 6634 10308 6658 10310
rect 6714 10308 6738 10310
rect 6794 10308 6818 10310
rect 6874 10308 6880 10310
rect 6572 10299 6880 10308
rect 6932 9518 6960 11018
rect 7024 9586 7052 11290
rect 7116 10674 7144 11478
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7116 10130 7144 10610
rect 7208 10606 7236 11614
rect 7300 10674 7328 16390
rect 7484 12434 7512 17138
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7668 12918 7696 13670
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7484 12406 7604 12434
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7116 9586 7144 10066
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6572 9276 6880 9285
rect 6572 9274 6578 9276
rect 6634 9274 6658 9276
rect 6714 9274 6738 9276
rect 6794 9274 6818 9276
rect 6874 9274 6880 9276
rect 6634 9222 6636 9274
rect 6816 9222 6818 9274
rect 6572 9220 6578 9222
rect 6634 9220 6658 9222
rect 6714 9220 6738 9222
rect 6794 9220 6818 9222
rect 6874 9220 6880 9222
rect 6572 9211 6880 9220
rect 6932 9178 6960 9454
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 7116 9178 7144 9386
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 6932 8498 6960 9114
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6572 8188 6880 8197
rect 6572 8186 6578 8188
rect 6634 8186 6658 8188
rect 6714 8186 6738 8188
rect 6794 8186 6818 8188
rect 6874 8186 6880 8188
rect 6634 8134 6636 8186
rect 6816 8134 6818 8186
rect 6572 8132 6578 8134
rect 6634 8132 6658 8134
rect 6714 8132 6738 8134
rect 6794 8132 6818 8134
rect 6874 8132 6880 8134
rect 6572 8123 6880 8132
rect 6572 7100 6880 7109
rect 6572 7098 6578 7100
rect 6634 7098 6658 7100
rect 6714 7098 6738 7100
rect 6794 7098 6818 7100
rect 6874 7098 6880 7100
rect 6634 7046 6636 7098
rect 6816 7046 6818 7098
rect 6572 7044 6578 7046
rect 6634 7044 6658 7046
rect 6714 7044 6738 7046
rect 6794 7044 6818 7046
rect 6874 7044 6880 7046
rect 6572 7035 6880 7044
rect 6572 6012 6880 6021
rect 6572 6010 6578 6012
rect 6634 6010 6658 6012
rect 6714 6010 6738 6012
rect 6794 6010 6818 6012
rect 6874 6010 6880 6012
rect 6634 5958 6636 6010
rect 6816 5958 6818 6010
rect 6572 5956 6578 5958
rect 6634 5956 6658 5958
rect 6714 5956 6738 5958
rect 6794 5956 6818 5958
rect 6874 5956 6880 5958
rect 6572 5947 6880 5956
rect 6572 4924 6880 4933
rect 6572 4922 6578 4924
rect 6634 4922 6658 4924
rect 6714 4922 6738 4924
rect 6794 4922 6818 4924
rect 6874 4922 6880 4924
rect 6634 4870 6636 4922
rect 6816 4870 6818 4922
rect 6572 4868 6578 4870
rect 6634 4868 6658 4870
rect 6714 4868 6738 4870
rect 6794 4868 6818 4870
rect 6874 4868 6880 4870
rect 6572 4859 6880 4868
rect 6572 3836 6880 3845
rect 6572 3834 6578 3836
rect 6634 3834 6658 3836
rect 6714 3834 6738 3836
rect 6794 3834 6818 3836
rect 6874 3834 6880 3836
rect 6634 3782 6636 3834
rect 6816 3782 6818 3834
rect 6572 3780 6578 3782
rect 6634 3780 6658 3782
rect 6714 3780 6738 3782
rect 6794 3780 6818 3782
rect 6874 3780 6880 3782
rect 6572 3771 6880 3780
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6572 2748 6880 2757
rect 6572 2746 6578 2748
rect 6634 2746 6658 2748
rect 6714 2746 6738 2748
rect 6794 2746 6818 2748
rect 6874 2746 6880 2748
rect 6634 2694 6636 2746
rect 6816 2694 6818 2746
rect 6572 2692 6578 2694
rect 6634 2692 6658 2694
rect 6714 2692 6738 2694
rect 6794 2692 6818 2694
rect 6874 2692 6880 2694
rect 6572 2683 6880 2692
rect 7208 2650 7236 10542
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7300 7410 7328 9862
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 6000 2032 6052 2038
rect 6000 1974 6052 1980
rect 6196 800 6224 2246
rect 6472 1834 6500 2382
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 6460 1828 6512 1834
rect 6460 1770 6512 1776
rect 6564 800 6592 2246
rect 6932 800 6960 2246
rect 7300 800 7328 2246
rect 7392 1834 7420 11698
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7484 7546 7512 10610
rect 7576 10554 7604 12406
rect 7668 10810 7696 12854
rect 8220 12434 8248 17138
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 8312 12442 8340 17070
rect 8446 16348 8754 16357
rect 8446 16346 8452 16348
rect 8508 16346 8532 16348
rect 8588 16346 8612 16348
rect 8668 16346 8692 16348
rect 8748 16346 8754 16348
rect 8508 16294 8510 16346
rect 8690 16294 8692 16346
rect 8446 16292 8452 16294
rect 8508 16292 8532 16294
rect 8588 16292 8612 16294
rect 8668 16292 8692 16294
rect 8748 16292 8754 16294
rect 8446 16283 8754 16292
rect 8446 15260 8754 15269
rect 8446 15258 8452 15260
rect 8508 15258 8532 15260
rect 8588 15258 8612 15260
rect 8668 15258 8692 15260
rect 8748 15258 8754 15260
rect 8508 15206 8510 15258
rect 8690 15206 8692 15258
rect 8446 15204 8452 15206
rect 8508 15204 8532 15206
rect 8588 15204 8612 15206
rect 8668 15204 8692 15206
rect 8748 15204 8754 15206
rect 8446 15195 8754 15204
rect 8446 14172 8754 14181
rect 8446 14170 8452 14172
rect 8508 14170 8532 14172
rect 8588 14170 8612 14172
rect 8668 14170 8692 14172
rect 8748 14170 8754 14172
rect 8508 14118 8510 14170
rect 8690 14118 8692 14170
rect 8446 14116 8452 14118
rect 8508 14116 8532 14118
rect 8588 14116 8612 14118
rect 8668 14116 8692 14118
rect 8748 14116 8754 14118
rect 8446 14107 8754 14116
rect 8446 13084 8754 13093
rect 8446 13082 8452 13084
rect 8508 13082 8532 13084
rect 8588 13082 8612 13084
rect 8668 13082 8692 13084
rect 8748 13082 8754 13084
rect 8508 13030 8510 13082
rect 8690 13030 8692 13082
rect 8446 13028 8452 13030
rect 8508 13028 8532 13030
rect 8588 13028 8612 13030
rect 8668 13028 8692 13030
rect 8748 13028 8754 13030
rect 8446 13019 8754 13028
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 7852 12406 8248 12434
rect 8300 12436 8352 12442
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7760 11121 7788 11698
rect 7746 11112 7802 11121
rect 7746 11047 7802 11056
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7852 10690 7880 12406
rect 8300 12378 8352 12384
rect 8116 12164 8168 12170
rect 8404 12152 8432 12786
rect 8864 12434 8892 17138
rect 8956 16658 8984 19200
rect 9220 17740 9272 17746
rect 9220 17682 9272 17688
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9140 17134 9168 17614
rect 9232 17202 9260 17682
rect 9324 17202 9352 19200
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9128 17128 9180 17134
rect 9128 17070 9180 17076
rect 9312 17060 9364 17066
rect 9232 17020 9312 17048
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 8864 12406 8984 12434
rect 8116 12106 8168 12112
rect 8312 12124 8432 12152
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 8036 11121 8064 11698
rect 8022 11112 8078 11121
rect 8128 11098 8156 12106
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8220 11286 8248 11630
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 8128 11070 8248 11098
rect 8022 11047 8078 11056
rect 7852 10662 8156 10690
rect 7576 10526 8064 10554
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7668 10198 7696 10406
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7746 10160 7802 10169
rect 7746 10095 7802 10104
rect 7760 10062 7788 10095
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7564 9988 7616 9994
rect 7564 9930 7616 9936
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7576 7410 7604 9930
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7668 2446 7696 7142
rect 7760 4146 7788 9998
rect 8036 9602 8064 10526
rect 8128 10266 8156 10662
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8220 9874 8248 11070
rect 8312 10130 8340 12124
rect 8446 11996 8754 12005
rect 8446 11994 8452 11996
rect 8508 11994 8532 11996
rect 8588 11994 8612 11996
rect 8668 11994 8692 11996
rect 8748 11994 8754 11996
rect 8508 11942 8510 11994
rect 8690 11942 8692 11994
rect 8446 11940 8452 11942
rect 8508 11940 8532 11942
rect 8588 11940 8612 11942
rect 8668 11940 8692 11942
rect 8748 11940 8754 11942
rect 8446 11931 8754 11940
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8446 10908 8754 10917
rect 8446 10906 8452 10908
rect 8508 10906 8532 10908
rect 8588 10906 8612 10908
rect 8668 10906 8692 10908
rect 8748 10906 8754 10908
rect 8508 10854 8510 10906
rect 8690 10854 8692 10906
rect 8446 10852 8452 10854
rect 8508 10852 8532 10854
rect 8588 10852 8612 10854
rect 8668 10852 8692 10854
rect 8748 10852 8754 10854
rect 8446 10843 8754 10852
rect 8864 10742 8892 11494
rect 8956 10810 8984 12406
rect 9232 11642 9260 17020
rect 9312 17002 9364 17008
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 9416 16794 9444 16934
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9048 11614 9260 11642
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 8852 10736 8904 10742
rect 8852 10678 8904 10684
rect 9048 10305 9076 11614
rect 9128 11076 9180 11082
rect 9128 11018 9180 11024
rect 9140 10606 9168 11018
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 8666 10296 8722 10305
rect 8666 10231 8722 10240
rect 9034 10296 9090 10305
rect 9034 10231 9090 10240
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8312 10033 8340 10066
rect 8298 10024 8354 10033
rect 8298 9959 8354 9968
rect 8404 9926 8432 10066
rect 8680 9926 8708 10231
rect 9048 9976 9076 10231
rect 9232 9994 9260 10950
rect 9220 9988 9272 9994
rect 9048 9948 9168 9976
rect 8392 9920 8444 9926
rect 8220 9846 8340 9874
rect 8392 9862 8444 9868
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 9034 9888 9090 9897
rect 8036 9574 8248 9602
rect 8220 9450 8248 9574
rect 8312 9518 8340 9846
rect 8446 9820 8754 9829
rect 8446 9818 8452 9820
rect 8508 9818 8532 9820
rect 8588 9818 8612 9820
rect 8668 9818 8692 9820
rect 8748 9818 8754 9820
rect 8508 9766 8510 9818
rect 8690 9766 8692 9818
rect 8446 9764 8452 9766
rect 8508 9764 8532 9766
rect 8588 9764 8612 9766
rect 8668 9764 8692 9766
rect 8748 9764 8754 9766
rect 8446 9755 8754 9764
rect 8850 9752 8906 9761
rect 8668 9716 8720 9722
rect 8496 9676 8668 9704
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8390 9480 8446 9489
rect 8208 9444 8260 9450
rect 8390 9415 8446 9424
rect 8208 9386 8260 9392
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8312 8974 8340 9318
rect 8404 9110 8432 9415
rect 8392 9104 8444 9110
rect 8392 9046 8444 9052
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8312 8566 8340 8910
rect 8496 8906 8524 9676
rect 8850 9687 8906 9696
rect 8668 9658 8720 9664
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8588 9110 8616 9454
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8446 8732 8754 8741
rect 8446 8730 8452 8732
rect 8508 8730 8532 8732
rect 8588 8730 8612 8732
rect 8668 8730 8692 8732
rect 8748 8730 8754 8732
rect 8508 8678 8510 8730
rect 8690 8678 8692 8730
rect 8446 8676 8452 8678
rect 8508 8676 8532 8678
rect 8588 8676 8612 8678
rect 8668 8676 8692 8678
rect 8748 8676 8754 8678
rect 8446 8667 8754 8676
rect 8864 8634 8892 9687
rect 8956 9654 8984 9862
rect 9140 9874 9168 9948
rect 9220 9930 9272 9936
rect 9324 9926 9352 12174
rect 9416 11082 9444 16594
rect 9508 12434 9536 17546
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9600 16658 9628 17274
rect 9692 17202 9720 19200
rect 10060 17202 10088 19200
rect 10428 17202 10456 19200
rect 10796 17202 10824 19200
rect 11164 17202 11192 19200
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 10048 17196 10100 17202
rect 10048 17138 10100 17144
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 11152 17196 11204 17202
rect 11152 17138 11204 17144
rect 9692 16794 9720 17138
rect 9956 17060 10008 17066
rect 9956 17002 10008 17008
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9968 16574 9996 17002
rect 10060 16794 10088 17138
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 10152 16574 10180 16934
rect 10320 16892 10628 16901
rect 10320 16890 10326 16892
rect 10382 16890 10406 16892
rect 10462 16890 10486 16892
rect 10542 16890 10566 16892
rect 10622 16890 10628 16892
rect 10382 16838 10384 16890
rect 10564 16838 10566 16890
rect 10320 16836 10326 16838
rect 10382 16836 10406 16838
rect 10462 16836 10486 16838
rect 10542 16836 10566 16838
rect 10622 16836 10628 16838
rect 10320 16827 10628 16836
rect 10704 16574 10732 16934
rect 10796 16794 10824 17138
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 10980 16810 11008 16934
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10888 16782 11008 16810
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 9692 16546 9996 16574
rect 10060 16546 10180 16574
rect 10244 16546 10732 16574
rect 9508 12406 9628 12434
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9312 9920 9364 9926
rect 9140 9846 9260 9874
rect 9312 9862 9364 9868
rect 9034 9823 9090 9832
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8956 9110 8984 9454
rect 9048 9382 9076 9823
rect 9232 9586 9260 9846
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 8956 8945 8984 9046
rect 9036 8968 9088 8974
rect 8942 8936 8998 8945
rect 9036 8910 9088 8916
rect 8942 8871 8998 8880
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8850 8528 8906 8537
rect 8392 8492 8444 8498
rect 8850 8463 8906 8472
rect 8392 8434 8444 8440
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 8312 2582 8340 8298
rect 8404 8294 8432 8434
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8446 7644 8754 7653
rect 8446 7642 8452 7644
rect 8508 7642 8532 7644
rect 8588 7642 8612 7644
rect 8668 7642 8692 7644
rect 8748 7642 8754 7644
rect 8508 7590 8510 7642
rect 8690 7590 8692 7642
rect 8446 7588 8452 7590
rect 8508 7588 8532 7590
rect 8588 7588 8612 7590
rect 8668 7588 8692 7590
rect 8748 7588 8754 7590
rect 8446 7579 8754 7588
rect 8864 7342 8892 8463
rect 8956 8362 8984 8774
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8446 6556 8754 6565
rect 8446 6554 8452 6556
rect 8508 6554 8532 6556
rect 8588 6554 8612 6556
rect 8668 6554 8692 6556
rect 8748 6554 8754 6556
rect 8508 6502 8510 6554
rect 8690 6502 8692 6554
rect 8446 6500 8452 6502
rect 8508 6500 8532 6502
rect 8588 6500 8612 6502
rect 8668 6500 8692 6502
rect 8748 6500 8754 6502
rect 8446 6491 8754 6500
rect 8446 5468 8754 5477
rect 8446 5466 8452 5468
rect 8508 5466 8532 5468
rect 8588 5466 8612 5468
rect 8668 5466 8692 5468
rect 8748 5466 8754 5468
rect 8508 5414 8510 5466
rect 8690 5414 8692 5466
rect 8446 5412 8452 5414
rect 8508 5412 8532 5414
rect 8588 5412 8612 5414
rect 8668 5412 8692 5414
rect 8748 5412 8754 5414
rect 8446 5403 8754 5412
rect 8446 4380 8754 4389
rect 8446 4378 8452 4380
rect 8508 4378 8532 4380
rect 8588 4378 8612 4380
rect 8668 4378 8692 4380
rect 8748 4378 8754 4380
rect 8508 4326 8510 4378
rect 8690 4326 8692 4378
rect 8446 4324 8452 4326
rect 8508 4324 8532 4326
rect 8588 4324 8612 4326
rect 8668 4324 8692 4326
rect 8748 4324 8754 4326
rect 8446 4315 8754 4324
rect 8446 3292 8754 3301
rect 8446 3290 8452 3292
rect 8508 3290 8532 3292
rect 8588 3290 8612 3292
rect 8668 3290 8692 3292
rect 8748 3290 8754 3292
rect 8508 3238 8510 3290
rect 8690 3238 8692 3290
rect 8446 3236 8452 3238
rect 8508 3236 8532 3238
rect 8588 3236 8612 3238
rect 8668 3236 8692 3238
rect 8748 3236 8754 3238
rect 8446 3227 8754 3236
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 7484 2038 7512 2382
rect 8680 2378 8708 2926
rect 8772 2446 8800 3130
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 8864 2378 8892 2790
rect 8668 2372 8720 2378
rect 8668 2314 8720 2320
rect 8852 2372 8904 2378
rect 8852 2314 8904 2320
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 7472 2032 7524 2038
rect 7472 1974 7524 1980
rect 7380 1828 7432 1834
rect 7380 1770 7432 1776
rect 7668 800 7696 2246
rect 8036 800 8064 2246
rect 8312 1170 8340 2246
rect 8446 2204 8754 2213
rect 8446 2202 8452 2204
rect 8508 2202 8532 2204
rect 8588 2202 8612 2204
rect 8668 2202 8692 2204
rect 8748 2202 8754 2204
rect 8508 2150 8510 2202
rect 8690 2150 8692 2202
rect 8446 2148 8452 2150
rect 8508 2148 8532 2150
rect 8588 2148 8612 2150
rect 8668 2148 8692 2150
rect 8748 2148 8754 2150
rect 8446 2139 8754 2148
rect 8864 1986 8892 2314
rect 8772 1958 8892 1986
rect 8312 1142 8432 1170
rect 8404 800 8432 1142
rect 8772 800 8800 1958
rect 9048 1902 9076 8910
rect 9232 4078 9260 9318
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 9140 2428 9168 2790
rect 9220 2440 9272 2446
rect 9140 2400 9220 2428
rect 9036 1896 9088 1902
rect 9036 1838 9088 1844
rect 9140 800 9168 2400
rect 9220 2382 9272 2388
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9232 1970 9260 2246
rect 9324 1970 9352 9862
rect 9416 7410 9444 11018
rect 9508 10130 9536 11154
rect 9600 11014 9628 12406
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9508 9722 9536 10066
rect 9600 9761 9628 10610
rect 9586 9752 9642 9761
rect 9496 9716 9548 9722
rect 9586 9687 9642 9696
rect 9496 9658 9548 9664
rect 9508 8430 9536 9658
rect 9586 9616 9642 9625
rect 9586 9551 9588 9560
rect 9640 9551 9642 9560
rect 9588 9522 9640 9528
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 8906 9628 9318
rect 9692 9178 9720 16546
rect 10060 12434 10088 16546
rect 10060 12406 10180 12434
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9784 8906 9812 12106
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9586 8800 9642 8809
rect 9586 8735 9642 8744
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9508 2394 9536 2790
rect 9600 2650 9628 8735
rect 9784 8362 9812 8842
rect 9876 8498 9904 9862
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 9784 2650 9812 3946
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9876 2446 9904 2790
rect 9968 2553 9996 10406
rect 10048 10192 10100 10198
rect 10048 10134 10100 10140
rect 9954 2544 10010 2553
rect 9954 2479 10010 2488
rect 9680 2440 9732 2446
rect 9508 2388 9680 2394
rect 9508 2382 9732 2388
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9508 2366 9720 2382
rect 9220 1964 9272 1970
rect 9220 1906 9272 1912
rect 9312 1964 9364 1970
rect 9312 1906 9364 1912
rect 9508 800 9536 2366
rect 9876 800 9904 2382
rect 10060 1766 10088 10134
rect 10152 9042 10180 12406
rect 10244 10010 10272 16546
rect 10320 15804 10628 15813
rect 10320 15802 10326 15804
rect 10382 15802 10406 15804
rect 10462 15802 10486 15804
rect 10542 15802 10566 15804
rect 10622 15802 10628 15804
rect 10382 15750 10384 15802
rect 10564 15750 10566 15802
rect 10320 15748 10326 15750
rect 10382 15748 10406 15750
rect 10462 15748 10486 15750
rect 10542 15748 10566 15750
rect 10622 15748 10628 15750
rect 10320 15739 10628 15748
rect 10320 14716 10628 14725
rect 10320 14714 10326 14716
rect 10382 14714 10406 14716
rect 10462 14714 10486 14716
rect 10542 14714 10566 14716
rect 10622 14714 10628 14716
rect 10382 14662 10384 14714
rect 10564 14662 10566 14714
rect 10320 14660 10326 14662
rect 10382 14660 10406 14662
rect 10462 14660 10486 14662
rect 10542 14660 10566 14662
rect 10622 14660 10628 14662
rect 10320 14651 10628 14660
rect 10320 13628 10628 13637
rect 10320 13626 10326 13628
rect 10382 13626 10406 13628
rect 10462 13626 10486 13628
rect 10542 13626 10566 13628
rect 10622 13626 10628 13628
rect 10382 13574 10384 13626
rect 10564 13574 10566 13626
rect 10320 13572 10326 13574
rect 10382 13572 10406 13574
rect 10462 13572 10486 13574
rect 10542 13572 10566 13574
rect 10622 13572 10628 13574
rect 10320 13563 10628 13572
rect 10796 12730 10824 16594
rect 10704 12702 10824 12730
rect 10320 12540 10628 12549
rect 10320 12538 10326 12540
rect 10382 12538 10406 12540
rect 10462 12538 10486 12540
rect 10542 12538 10566 12540
rect 10622 12538 10628 12540
rect 10382 12486 10384 12538
rect 10564 12486 10566 12538
rect 10320 12484 10326 12486
rect 10382 12484 10406 12486
rect 10462 12484 10486 12486
rect 10542 12484 10566 12486
rect 10622 12484 10628 12486
rect 10320 12475 10628 12484
rect 10320 11452 10628 11461
rect 10320 11450 10326 11452
rect 10382 11450 10406 11452
rect 10462 11450 10486 11452
rect 10542 11450 10566 11452
rect 10622 11450 10628 11452
rect 10382 11398 10384 11450
rect 10564 11398 10566 11450
rect 10320 11396 10326 11398
rect 10382 11396 10406 11398
rect 10462 11396 10486 11398
rect 10542 11396 10566 11398
rect 10622 11396 10628 11398
rect 10320 11387 10628 11396
rect 10320 10364 10628 10373
rect 10320 10362 10326 10364
rect 10382 10362 10406 10364
rect 10462 10362 10486 10364
rect 10542 10362 10566 10364
rect 10622 10362 10628 10364
rect 10382 10310 10384 10362
rect 10564 10310 10566 10362
rect 10320 10308 10326 10310
rect 10382 10308 10406 10310
rect 10462 10308 10486 10310
rect 10542 10308 10566 10310
rect 10622 10308 10628 10310
rect 10320 10299 10628 10308
rect 10244 9994 10364 10010
rect 10244 9988 10376 9994
rect 10244 9982 10324 9988
rect 10324 9930 10376 9936
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 10244 9625 10272 9862
rect 10230 9616 10286 9625
rect 10230 9551 10286 9560
rect 10230 9480 10286 9489
rect 10230 9415 10232 9424
rect 10284 9415 10286 9424
rect 10232 9386 10284 9392
rect 10320 9276 10628 9285
rect 10320 9274 10326 9276
rect 10382 9274 10406 9276
rect 10462 9274 10486 9276
rect 10542 9274 10566 9276
rect 10622 9274 10628 9276
rect 10382 9222 10384 9274
rect 10564 9222 10566 9274
rect 10320 9220 10326 9222
rect 10382 9220 10406 9222
rect 10462 9220 10486 9222
rect 10542 9220 10566 9222
rect 10622 9220 10628 9222
rect 10320 9211 10628 9220
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10704 8974 10732 12702
rect 10888 11286 10916 16782
rect 10966 16688 11022 16697
rect 10966 16623 11022 16632
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 10980 10062 11008 16623
rect 11072 10538 11100 17002
rect 11164 16794 11192 17138
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11244 16720 11296 16726
rect 11244 16662 11296 16668
rect 11256 10674 11284 16662
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10320 8188 10628 8197
rect 10320 8186 10326 8188
rect 10382 8186 10406 8188
rect 10462 8186 10486 8188
rect 10542 8186 10566 8188
rect 10622 8186 10628 8188
rect 10382 8134 10384 8186
rect 10564 8134 10566 8186
rect 10320 8132 10326 8134
rect 10382 8132 10406 8134
rect 10462 8132 10486 8134
rect 10542 8132 10566 8134
rect 10622 8132 10628 8134
rect 10320 8123 10628 8132
rect 10320 7100 10628 7109
rect 10320 7098 10326 7100
rect 10382 7098 10406 7100
rect 10462 7098 10486 7100
rect 10542 7098 10566 7100
rect 10622 7098 10628 7100
rect 10382 7046 10384 7098
rect 10564 7046 10566 7098
rect 10320 7044 10326 7046
rect 10382 7044 10406 7046
rect 10462 7044 10486 7046
rect 10542 7044 10566 7046
rect 10622 7044 10628 7046
rect 10320 7035 10628 7044
rect 10320 6012 10628 6021
rect 10320 6010 10326 6012
rect 10382 6010 10406 6012
rect 10462 6010 10486 6012
rect 10542 6010 10566 6012
rect 10622 6010 10628 6012
rect 10382 5958 10384 6010
rect 10564 5958 10566 6010
rect 10320 5956 10326 5958
rect 10382 5956 10406 5958
rect 10462 5956 10486 5958
rect 10542 5956 10566 5958
rect 10622 5956 10628 5958
rect 10320 5947 10628 5956
rect 10320 4924 10628 4933
rect 10320 4922 10326 4924
rect 10382 4922 10406 4924
rect 10462 4922 10486 4924
rect 10542 4922 10566 4924
rect 10622 4922 10628 4924
rect 10382 4870 10384 4922
rect 10564 4870 10566 4922
rect 10320 4868 10326 4870
rect 10382 4868 10406 4870
rect 10462 4868 10486 4870
rect 10542 4868 10566 4870
rect 10622 4868 10628 4870
rect 10320 4859 10628 4868
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10152 2650 10180 4014
rect 10320 3836 10628 3845
rect 10320 3834 10326 3836
rect 10382 3834 10406 3836
rect 10462 3834 10486 3836
rect 10542 3834 10566 3836
rect 10622 3834 10628 3836
rect 10382 3782 10384 3834
rect 10564 3782 10566 3834
rect 10320 3780 10326 3782
rect 10382 3780 10406 3782
rect 10462 3780 10486 3782
rect 10542 3780 10566 3782
rect 10622 3780 10628 3782
rect 10320 3771 10628 3780
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 10244 2446 10272 2790
rect 10320 2748 10628 2757
rect 10320 2746 10326 2748
rect 10382 2746 10406 2748
rect 10462 2746 10486 2748
rect 10542 2746 10566 2748
rect 10622 2746 10628 2748
rect 10382 2694 10384 2746
rect 10564 2694 10566 2746
rect 10320 2692 10326 2694
rect 10382 2692 10406 2694
rect 10462 2692 10486 2694
rect 10542 2692 10566 2694
rect 10622 2692 10628 2694
rect 10320 2683 10628 2692
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 10600 2440 10652 2446
rect 10704 2428 10732 2790
rect 10652 2400 10732 2428
rect 10600 2382 10652 2388
rect 10048 1760 10100 1766
rect 10048 1702 10100 1708
rect 10244 800 10272 2382
rect 10612 800 10640 2382
rect 10796 2378 10824 9454
rect 10888 2990 10916 9862
rect 11164 8566 11192 10542
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 10980 2428 11008 2790
rect 11256 2774 11284 10066
rect 11348 10062 11376 17478
rect 11532 17270 11560 19200
rect 11520 17264 11572 17270
rect 11520 17206 11572 17212
rect 11428 17128 11480 17134
rect 11428 17070 11480 17076
rect 11440 10266 11468 17070
rect 11532 16794 11560 17206
rect 11900 17134 11928 19200
rect 12268 17626 12296 19200
rect 12084 17598 12296 17626
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 11808 10713 11836 16934
rect 11900 16794 11928 17070
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11992 16658 12020 16934
rect 12084 16794 12112 17598
rect 12194 17436 12502 17445
rect 12194 17434 12200 17436
rect 12256 17434 12280 17436
rect 12336 17434 12360 17436
rect 12416 17434 12440 17436
rect 12496 17434 12502 17436
rect 12256 17382 12258 17434
rect 12438 17382 12440 17434
rect 12194 17380 12200 17382
rect 12256 17380 12280 17382
rect 12336 17380 12360 17382
rect 12416 17380 12440 17382
rect 12496 17380 12502 17382
rect 12194 17371 12502 17380
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12256 17060 12308 17066
rect 12256 17002 12308 17008
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 12268 16726 12296 17002
rect 12452 16794 12480 17138
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12256 16720 12308 16726
rect 12256 16662 12308 16668
rect 12348 16720 12400 16726
rect 12348 16662 12400 16668
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 12360 16574 12388 16662
rect 12084 16546 12388 16574
rect 12084 10742 12112 16546
rect 12194 16348 12502 16357
rect 12194 16346 12200 16348
rect 12256 16346 12280 16348
rect 12336 16346 12360 16348
rect 12416 16346 12440 16348
rect 12496 16346 12502 16348
rect 12256 16294 12258 16346
rect 12438 16294 12440 16346
rect 12194 16292 12200 16294
rect 12256 16292 12280 16294
rect 12336 16292 12360 16294
rect 12416 16292 12440 16294
rect 12496 16292 12502 16294
rect 12194 16283 12502 16292
rect 12194 15260 12502 15269
rect 12194 15258 12200 15260
rect 12256 15258 12280 15260
rect 12336 15258 12360 15260
rect 12416 15258 12440 15260
rect 12496 15258 12502 15260
rect 12256 15206 12258 15258
rect 12438 15206 12440 15258
rect 12194 15204 12200 15206
rect 12256 15204 12280 15206
rect 12336 15204 12360 15206
rect 12416 15204 12440 15206
rect 12496 15204 12502 15206
rect 12194 15195 12502 15204
rect 12194 14172 12502 14181
rect 12194 14170 12200 14172
rect 12256 14170 12280 14172
rect 12336 14170 12360 14172
rect 12416 14170 12440 14172
rect 12496 14170 12502 14172
rect 12256 14118 12258 14170
rect 12438 14118 12440 14170
rect 12194 14116 12200 14118
rect 12256 14116 12280 14118
rect 12336 14116 12360 14118
rect 12416 14116 12440 14118
rect 12496 14116 12502 14118
rect 12194 14107 12502 14116
rect 12194 13084 12502 13093
rect 12194 13082 12200 13084
rect 12256 13082 12280 13084
rect 12336 13082 12360 13084
rect 12416 13082 12440 13084
rect 12496 13082 12502 13084
rect 12256 13030 12258 13082
rect 12438 13030 12440 13082
rect 12194 13028 12200 13030
rect 12256 13028 12280 13030
rect 12336 13028 12360 13030
rect 12416 13028 12440 13030
rect 12496 13028 12502 13030
rect 12194 13019 12502 13028
rect 12194 11996 12502 12005
rect 12194 11994 12200 11996
rect 12256 11994 12280 11996
rect 12336 11994 12360 11996
rect 12416 11994 12440 11996
rect 12496 11994 12502 11996
rect 12256 11942 12258 11994
rect 12438 11942 12440 11994
rect 12194 11940 12200 11942
rect 12256 11940 12280 11942
rect 12336 11940 12360 11942
rect 12416 11940 12440 11942
rect 12496 11940 12502 11942
rect 12194 11931 12502 11940
rect 12194 10908 12502 10917
rect 12194 10906 12200 10908
rect 12256 10906 12280 10908
rect 12336 10906 12360 10908
rect 12416 10906 12440 10908
rect 12496 10906 12502 10908
rect 12256 10854 12258 10906
rect 12438 10854 12440 10906
rect 12194 10852 12200 10854
rect 12256 10852 12280 10854
rect 12336 10852 12360 10854
rect 12416 10852 12440 10854
rect 12496 10852 12502 10854
rect 12194 10843 12502 10852
rect 12072 10736 12124 10742
rect 11794 10704 11850 10713
rect 12072 10678 12124 10684
rect 11794 10639 11850 10648
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11612 10192 11664 10198
rect 11612 10134 11664 10140
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11164 2746 11284 2774
rect 11060 2440 11112 2446
rect 10980 2400 11060 2428
rect 10784 2372 10836 2378
rect 10784 2314 10836 2320
rect 10692 2304 10744 2310
rect 10692 2246 10744 2252
rect 10704 2106 10732 2246
rect 10692 2100 10744 2106
rect 10692 2042 10744 2048
rect 10980 800 11008 2400
rect 11060 2382 11112 2388
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11072 1834 11100 2246
rect 11164 2106 11192 2746
rect 11348 2446 11376 2790
rect 11336 2440 11388 2446
rect 11336 2382 11388 2388
rect 11152 2100 11204 2106
rect 11152 2042 11204 2048
rect 11060 1828 11112 1834
rect 11060 1770 11112 1776
rect 11348 800 11376 2382
rect 11440 2038 11468 9862
rect 11532 9722 11560 9998
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 11532 2553 11560 2586
rect 11518 2544 11574 2553
rect 11624 2514 11652 10134
rect 11716 10062 11744 10406
rect 12544 10266 12572 17614
rect 12636 17202 12664 19200
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 12636 16794 12664 17138
rect 12728 16998 12756 17546
rect 13004 17202 13032 19200
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12820 16697 12848 16934
rect 12806 16688 12862 16697
rect 12806 16623 12862 16632
rect 13188 10266 13216 17682
rect 13372 17202 13400 19200
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 13372 16794 13400 17138
rect 13360 16788 13412 16794
rect 13360 16730 13412 16736
rect 13464 16726 13492 17274
rect 13740 17218 13768 19200
rect 14108 17270 14136 19200
rect 14476 17762 14504 19200
rect 14476 17734 14688 17762
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14384 17338 14412 17478
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 14096 17264 14148 17270
rect 13740 17202 13860 17218
rect 14096 17206 14148 17212
rect 14464 17264 14516 17270
rect 14464 17206 14516 17212
rect 13740 17196 13872 17202
rect 13740 17190 13820 17196
rect 13820 17138 13872 17144
rect 13832 16794 13860 17138
rect 14068 16892 14376 16901
rect 14068 16890 14074 16892
rect 14130 16890 14154 16892
rect 14210 16890 14234 16892
rect 14290 16890 14314 16892
rect 14370 16890 14376 16892
rect 14130 16838 14132 16890
rect 14312 16838 14314 16890
rect 14068 16836 14074 16838
rect 14130 16836 14154 16838
rect 14210 16836 14234 16838
rect 14290 16836 14314 16838
rect 14370 16836 14376 16838
rect 14068 16827 14376 16836
rect 14476 16794 14504 17206
rect 14660 17202 14688 17734
rect 14844 17218 14872 19200
rect 14844 17202 14964 17218
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14844 17196 14976 17202
rect 14844 17190 14924 17196
rect 14740 17128 14792 17134
rect 14740 17070 14792 17076
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 14068 15804 14376 15813
rect 14068 15802 14074 15804
rect 14130 15802 14154 15804
rect 14210 15802 14234 15804
rect 14290 15802 14314 15804
rect 14370 15802 14376 15804
rect 14130 15750 14132 15802
rect 14312 15750 14314 15802
rect 14068 15748 14074 15750
rect 14130 15748 14154 15750
rect 14210 15748 14234 15750
rect 14290 15748 14314 15750
rect 14370 15748 14376 15750
rect 14068 15739 14376 15748
rect 14068 14716 14376 14725
rect 14068 14714 14074 14716
rect 14130 14714 14154 14716
rect 14210 14714 14234 14716
rect 14290 14714 14314 14716
rect 14370 14714 14376 14716
rect 14130 14662 14132 14714
rect 14312 14662 14314 14714
rect 14068 14660 14074 14662
rect 14130 14660 14154 14662
rect 14210 14660 14234 14662
rect 14290 14660 14314 14662
rect 14370 14660 14376 14662
rect 14068 14651 14376 14660
rect 14068 13628 14376 13637
rect 14068 13626 14074 13628
rect 14130 13626 14154 13628
rect 14210 13626 14234 13628
rect 14290 13626 14314 13628
rect 14370 13626 14376 13628
rect 14130 13574 14132 13626
rect 14312 13574 14314 13626
rect 14068 13572 14074 13574
rect 14130 13572 14154 13574
rect 14210 13572 14234 13574
rect 14290 13572 14314 13574
rect 14370 13572 14376 13574
rect 14068 13563 14376 13572
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13924 10169 13952 12582
rect 14068 12540 14376 12549
rect 14068 12538 14074 12540
rect 14130 12538 14154 12540
rect 14210 12538 14234 12540
rect 14290 12538 14314 12540
rect 14370 12538 14376 12540
rect 14130 12486 14132 12538
rect 14312 12486 14314 12538
rect 14068 12484 14074 12486
rect 14130 12484 14154 12486
rect 14210 12484 14234 12486
rect 14290 12484 14314 12486
rect 14370 12484 14376 12486
rect 14068 12475 14376 12484
rect 14068 11452 14376 11461
rect 14068 11450 14074 11452
rect 14130 11450 14154 11452
rect 14210 11450 14234 11452
rect 14290 11450 14314 11452
rect 14370 11450 14376 11452
rect 14130 11398 14132 11450
rect 14312 11398 14314 11450
rect 14068 11396 14074 11398
rect 14130 11396 14154 11398
rect 14210 11396 14234 11398
rect 14290 11396 14314 11398
rect 14370 11396 14376 11398
rect 14068 11387 14376 11396
rect 14660 10470 14688 16934
rect 14752 12986 14780 17070
rect 14844 16794 14872 17190
rect 14924 17138 14976 17144
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 15212 16674 15240 19200
rect 15580 17490 15608 19200
rect 15488 17462 15608 17490
rect 15212 16658 15332 16674
rect 15212 16652 15344 16658
rect 15212 16646 15292 16652
rect 15292 16594 15344 16600
rect 15384 16584 15436 16590
rect 15488 16574 15516 17462
rect 15566 17368 15622 17377
rect 15566 17303 15568 17312
rect 15620 17303 15622 17312
rect 15568 17274 15620 17280
rect 15436 16546 15516 16574
rect 15384 16526 15436 16532
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 14648 10464 14700 10470
rect 14648 10406 14700 10412
rect 14068 10364 14376 10373
rect 14068 10362 14074 10364
rect 14130 10362 14154 10364
rect 14210 10362 14234 10364
rect 14290 10362 14314 10364
rect 14370 10362 14376 10364
rect 14130 10310 14132 10362
rect 14312 10310 14314 10362
rect 14068 10308 14074 10310
rect 14130 10308 14154 10310
rect 14210 10308 14234 10310
rect 14290 10308 14314 10310
rect 14370 10308 14376 10310
rect 14068 10299 14376 10308
rect 15028 10198 15056 16390
rect 15016 10192 15068 10198
rect 13910 10160 13966 10169
rect 15016 10134 15068 10140
rect 13910 10095 13966 10104
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11716 2582 11744 9862
rect 12194 9820 12502 9829
rect 12194 9818 12200 9820
rect 12256 9818 12280 9820
rect 12336 9818 12360 9820
rect 12416 9818 12440 9820
rect 12496 9818 12502 9820
rect 12256 9766 12258 9818
rect 12438 9766 12440 9818
rect 12194 9764 12200 9766
rect 12256 9764 12280 9766
rect 12336 9764 12360 9766
rect 12416 9764 12440 9766
rect 12496 9764 12502 9766
rect 12194 9755 12502 9764
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11704 2576 11756 2582
rect 11704 2518 11756 2524
rect 11518 2479 11574 2488
rect 11612 2508 11664 2514
rect 11612 2450 11664 2456
rect 11808 2446 11836 2790
rect 11900 2514 11928 9522
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11992 2582 12020 9454
rect 12624 8900 12676 8906
rect 12624 8842 12676 8848
rect 12194 8732 12502 8741
rect 12194 8730 12200 8732
rect 12256 8730 12280 8732
rect 12336 8730 12360 8732
rect 12416 8730 12440 8732
rect 12496 8730 12502 8732
rect 12256 8678 12258 8730
rect 12438 8678 12440 8730
rect 12194 8676 12200 8678
rect 12256 8676 12280 8678
rect 12336 8676 12360 8678
rect 12416 8676 12440 8678
rect 12496 8676 12502 8678
rect 12194 8667 12502 8676
rect 12194 7644 12502 7653
rect 12194 7642 12200 7644
rect 12256 7642 12280 7644
rect 12336 7642 12360 7644
rect 12416 7642 12440 7644
rect 12496 7642 12502 7644
rect 12256 7590 12258 7642
rect 12438 7590 12440 7642
rect 12194 7588 12200 7590
rect 12256 7588 12280 7590
rect 12336 7588 12360 7590
rect 12416 7588 12440 7590
rect 12496 7588 12502 7590
rect 12194 7579 12502 7588
rect 12194 6556 12502 6565
rect 12194 6554 12200 6556
rect 12256 6554 12280 6556
rect 12336 6554 12360 6556
rect 12416 6554 12440 6556
rect 12496 6554 12502 6556
rect 12256 6502 12258 6554
rect 12438 6502 12440 6554
rect 12194 6500 12200 6502
rect 12256 6500 12280 6502
rect 12336 6500 12360 6502
rect 12416 6500 12440 6502
rect 12496 6500 12502 6502
rect 12194 6491 12502 6500
rect 12194 5468 12502 5477
rect 12194 5466 12200 5468
rect 12256 5466 12280 5468
rect 12336 5466 12360 5468
rect 12416 5466 12440 5468
rect 12496 5466 12502 5468
rect 12256 5414 12258 5466
rect 12438 5414 12440 5466
rect 12194 5412 12200 5414
rect 12256 5412 12280 5414
rect 12336 5412 12360 5414
rect 12416 5412 12440 5414
rect 12496 5412 12502 5414
rect 12194 5403 12502 5412
rect 12194 4380 12502 4389
rect 12194 4378 12200 4380
rect 12256 4378 12280 4380
rect 12336 4378 12360 4380
rect 12416 4378 12440 4380
rect 12496 4378 12502 4380
rect 12256 4326 12258 4378
rect 12438 4326 12440 4378
rect 12194 4324 12200 4326
rect 12256 4324 12280 4326
rect 12336 4324 12360 4326
rect 12416 4324 12440 4326
rect 12496 4324 12502 4326
rect 12194 4315 12502 4324
rect 12194 3292 12502 3301
rect 12194 3290 12200 3292
rect 12256 3290 12280 3292
rect 12336 3290 12360 3292
rect 12416 3290 12440 3292
rect 12496 3290 12502 3292
rect 12256 3238 12258 3290
rect 12438 3238 12440 3290
rect 12194 3236 12200 3238
rect 12256 3236 12280 3238
rect 12336 3236 12360 3238
rect 12416 3236 12440 3238
rect 12496 3236 12502 3238
rect 12194 3227 12502 3236
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 12532 2848 12584 2854
rect 12532 2790 12584 2796
rect 11980 2576 12032 2582
rect 11980 2518 12032 2524
rect 11888 2508 11940 2514
rect 11888 2450 11940 2456
rect 12084 2446 12112 2790
rect 12544 2446 12572 2790
rect 12636 2650 12664 8842
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12728 7585 12756 8298
rect 12714 7576 12770 7585
rect 12714 7511 12770 7520
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 12728 2553 12756 4082
rect 12898 2952 12954 2961
rect 12898 2887 12954 2896
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 12714 2544 12770 2553
rect 12714 2479 12770 2488
rect 12820 2446 12848 2790
rect 12912 2650 12940 2887
rect 13004 2650 13032 9998
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13096 3194 13124 9862
rect 13372 3194 13400 9998
rect 15120 9994 15148 16390
rect 15948 16114 15976 19200
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15488 10130 15516 15846
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15580 12481 15608 12582
rect 15566 12472 15622 12481
rect 15566 12407 15622 12416
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15108 9988 15160 9994
rect 15108 9930 15160 9936
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 13188 2446 13216 2790
rect 11796 2440 11848 2446
rect 11518 2408 11574 2417
rect 11518 2343 11574 2352
rect 11716 2400 11796 2428
rect 11532 2310 11560 2343
rect 11520 2304 11572 2310
rect 11520 2246 11572 2252
rect 11428 2032 11480 2038
rect 11428 1974 11480 1980
rect 11716 800 11744 2400
rect 11796 2382 11848 2388
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11992 1902 12020 2246
rect 11980 1896 12032 1902
rect 11980 1838 12032 1844
rect 12084 800 12112 2382
rect 12194 2204 12502 2213
rect 12194 2202 12200 2204
rect 12256 2202 12280 2204
rect 12336 2202 12360 2204
rect 12416 2202 12440 2204
rect 12496 2202 12502 2204
rect 12256 2150 12258 2202
rect 12438 2150 12440 2202
rect 12194 2148 12200 2150
rect 12256 2148 12280 2150
rect 12336 2148 12360 2150
rect 12416 2148 12440 2150
rect 12496 2148 12502 2150
rect 12194 2139 12502 2148
rect 12544 1986 12572 2382
rect 12452 1958 12572 1986
rect 12452 800 12480 1958
rect 12820 800 12848 2382
rect 13188 800 13216 2382
rect 13740 2310 13768 9658
rect 14068 9276 14376 9285
rect 14068 9274 14074 9276
rect 14130 9274 14154 9276
rect 14210 9274 14234 9276
rect 14290 9274 14314 9276
rect 14370 9274 14376 9276
rect 14130 9222 14132 9274
rect 14312 9222 14314 9274
rect 14068 9220 14074 9222
rect 14130 9220 14154 9222
rect 14210 9220 14234 9222
rect 14290 9220 14314 9222
rect 14370 9220 14376 9222
rect 14068 9211 14376 9220
rect 14068 8188 14376 8197
rect 14068 8186 14074 8188
rect 14130 8186 14154 8188
rect 14210 8186 14234 8188
rect 14290 8186 14314 8188
rect 14370 8186 14376 8188
rect 14130 8134 14132 8186
rect 14312 8134 14314 8186
rect 14068 8132 14074 8134
rect 14130 8132 14154 8134
rect 14210 8132 14234 8134
rect 14290 8132 14314 8134
rect 14370 8132 14376 8134
rect 14068 8123 14376 8132
rect 14068 7100 14376 7109
rect 14068 7098 14074 7100
rect 14130 7098 14154 7100
rect 14210 7098 14234 7100
rect 14290 7098 14314 7100
rect 14370 7098 14376 7100
rect 14130 7046 14132 7098
rect 14312 7046 14314 7098
rect 14068 7044 14074 7046
rect 14130 7044 14154 7046
rect 14210 7044 14234 7046
rect 14290 7044 14314 7046
rect 14370 7044 14376 7046
rect 14068 7035 14376 7044
rect 14068 6012 14376 6021
rect 14068 6010 14074 6012
rect 14130 6010 14154 6012
rect 14210 6010 14234 6012
rect 14290 6010 14314 6012
rect 14370 6010 14376 6012
rect 14130 5958 14132 6010
rect 14312 5958 14314 6010
rect 14068 5956 14074 5958
rect 14130 5956 14154 5958
rect 14210 5956 14234 5958
rect 14290 5956 14314 5958
rect 14370 5956 14376 5958
rect 14068 5947 14376 5956
rect 14068 4924 14376 4933
rect 14068 4922 14074 4924
rect 14130 4922 14154 4924
rect 14210 4922 14234 4924
rect 14290 4922 14314 4924
rect 14370 4922 14376 4924
rect 14130 4870 14132 4922
rect 14312 4870 14314 4922
rect 14068 4868 14074 4870
rect 14130 4868 14154 4870
rect 14210 4868 14234 4870
rect 14290 4868 14314 4870
rect 14370 4868 14376 4870
rect 14068 4859 14376 4868
rect 14068 3836 14376 3845
rect 14068 3834 14074 3836
rect 14130 3834 14154 3836
rect 14210 3834 14234 3836
rect 14290 3834 14314 3836
rect 14370 3834 14376 3836
rect 14130 3782 14132 3834
rect 14312 3782 14314 3834
rect 14068 3780 14074 3782
rect 14130 3780 14154 3782
rect 14210 3780 14234 3782
rect 14290 3780 14314 3782
rect 14370 3780 14376 3782
rect 14068 3771 14376 3780
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 13832 2446 13860 2790
rect 13924 2446 13952 2790
rect 14068 2748 14376 2757
rect 14068 2746 14074 2748
rect 14130 2746 14154 2748
rect 14210 2746 14234 2748
rect 14290 2746 14314 2748
rect 14370 2746 14376 2748
rect 14130 2694 14132 2746
rect 14312 2694 14314 2746
rect 14068 2692 14074 2694
rect 14130 2692 14154 2694
rect 14210 2692 14234 2694
rect 14290 2692 14314 2694
rect 14370 2692 14376 2694
rect 14068 2683 14376 2692
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 13912 2440 13964 2446
rect 14372 2440 14424 2446
rect 13912 2382 13964 2388
rect 14292 2400 14372 2428
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 13832 1816 13860 2382
rect 13556 1788 13860 1816
rect 13556 800 13584 1788
rect 13924 800 13952 2382
rect 14292 800 14320 2400
rect 14476 2428 14504 2790
rect 14660 2446 14688 2790
rect 14424 2400 14504 2428
rect 14648 2440 14700 2446
rect 14372 2382 14424 2388
rect 14648 2382 14700 2388
rect 15028 2394 15056 2790
rect 15396 2446 15424 2790
rect 15200 2440 15252 2446
rect 15028 2388 15200 2394
rect 15028 2382 15252 2388
rect 15384 2440 15436 2446
rect 15384 2382 15436 2388
rect 14660 800 14688 2382
rect 15028 2366 15240 2382
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14752 1970 14780 2246
rect 14740 1964 14792 1970
rect 14740 1906 14792 1912
rect 15028 800 15056 2366
rect 15108 2304 15160 2310
rect 15108 2246 15160 2252
rect 15120 2106 15148 2246
rect 15108 2100 15160 2106
rect 15108 2042 15160 2048
rect 15396 800 15424 2382
rect 15764 800 15792 2994
rect 1398 0 1454 800
rect 1766 0 1822 800
rect 2134 0 2190 800
rect 2502 0 2558 800
rect 2870 0 2926 800
rect 3238 0 3294 800
rect 3606 0 3662 800
rect 3974 0 4030 800
rect 4342 0 4398 800
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11702 0 11758 800
rect 12070 0 12126 800
rect 12438 0 12494 800
rect 12806 0 12862 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 13910 0 13966 800
rect 14278 0 14334 800
rect 14646 0 14702 800
rect 15014 0 15070 800
rect 15382 0 15438 800
rect 15750 0 15806 800
<< via2 >>
rect 1674 18128 1730 18184
rect 1490 14864 1546 14920
rect 1398 11600 1454 11656
rect 2830 16890 2886 16892
rect 2910 16890 2966 16892
rect 2990 16890 3046 16892
rect 3070 16890 3126 16892
rect 2830 16838 2876 16890
rect 2876 16838 2886 16890
rect 2910 16838 2940 16890
rect 2940 16838 2952 16890
rect 2952 16838 2966 16890
rect 2990 16838 3004 16890
rect 3004 16838 3016 16890
rect 3016 16838 3046 16890
rect 3070 16838 3080 16890
rect 3080 16838 3126 16890
rect 2830 16836 2886 16838
rect 2910 16836 2966 16838
rect 2990 16836 3046 16838
rect 3070 16836 3126 16838
rect 2830 15802 2886 15804
rect 2910 15802 2966 15804
rect 2990 15802 3046 15804
rect 3070 15802 3126 15804
rect 2830 15750 2876 15802
rect 2876 15750 2886 15802
rect 2910 15750 2940 15802
rect 2940 15750 2952 15802
rect 2952 15750 2966 15802
rect 2990 15750 3004 15802
rect 3004 15750 3016 15802
rect 3016 15750 3046 15802
rect 3070 15750 3080 15802
rect 3080 15750 3126 15802
rect 2830 15748 2886 15750
rect 2910 15748 2966 15750
rect 2990 15748 3046 15750
rect 3070 15748 3126 15750
rect 2830 14714 2886 14716
rect 2910 14714 2966 14716
rect 2990 14714 3046 14716
rect 3070 14714 3126 14716
rect 2830 14662 2876 14714
rect 2876 14662 2886 14714
rect 2910 14662 2940 14714
rect 2940 14662 2952 14714
rect 2952 14662 2966 14714
rect 2990 14662 3004 14714
rect 3004 14662 3016 14714
rect 3016 14662 3046 14714
rect 3070 14662 3080 14714
rect 3080 14662 3126 14714
rect 2830 14660 2886 14662
rect 2910 14660 2966 14662
rect 2990 14660 3046 14662
rect 3070 14660 3126 14662
rect 2830 13626 2886 13628
rect 2910 13626 2966 13628
rect 2990 13626 3046 13628
rect 3070 13626 3126 13628
rect 2830 13574 2876 13626
rect 2876 13574 2886 13626
rect 2910 13574 2940 13626
rect 2940 13574 2952 13626
rect 2952 13574 2966 13626
rect 2990 13574 3004 13626
rect 3004 13574 3016 13626
rect 3016 13574 3046 13626
rect 3070 13574 3080 13626
rect 3080 13574 3126 13626
rect 2830 13572 2886 13574
rect 2910 13572 2966 13574
rect 2990 13572 3046 13574
rect 3070 13572 3126 13574
rect 2830 12538 2886 12540
rect 2910 12538 2966 12540
rect 2990 12538 3046 12540
rect 3070 12538 3126 12540
rect 2830 12486 2876 12538
rect 2876 12486 2886 12538
rect 2910 12486 2940 12538
rect 2940 12486 2952 12538
rect 2952 12486 2966 12538
rect 2990 12486 3004 12538
rect 3004 12486 3016 12538
rect 3016 12486 3046 12538
rect 3070 12486 3080 12538
rect 3080 12486 3126 12538
rect 2830 12484 2886 12486
rect 2910 12484 2966 12486
rect 2990 12484 3046 12486
rect 3070 12484 3126 12486
rect 2830 11450 2886 11452
rect 2910 11450 2966 11452
rect 2990 11450 3046 11452
rect 3070 11450 3126 11452
rect 2830 11398 2876 11450
rect 2876 11398 2886 11450
rect 2910 11398 2940 11450
rect 2940 11398 2952 11450
rect 2952 11398 2966 11450
rect 2990 11398 3004 11450
rect 3004 11398 3016 11450
rect 3016 11398 3046 11450
rect 3070 11398 3080 11450
rect 3080 11398 3126 11450
rect 2830 11396 2886 11398
rect 2910 11396 2966 11398
rect 2990 11396 3046 11398
rect 3070 11396 3126 11398
rect 4704 17434 4760 17436
rect 4784 17434 4840 17436
rect 4864 17434 4920 17436
rect 4944 17434 5000 17436
rect 4704 17382 4750 17434
rect 4750 17382 4760 17434
rect 4784 17382 4814 17434
rect 4814 17382 4826 17434
rect 4826 17382 4840 17434
rect 4864 17382 4878 17434
rect 4878 17382 4890 17434
rect 4890 17382 4920 17434
rect 4944 17382 4954 17434
rect 4954 17382 5000 17434
rect 4704 17380 4760 17382
rect 4784 17380 4840 17382
rect 4864 17380 4920 17382
rect 4944 17380 5000 17382
rect 8452 17434 8508 17436
rect 8532 17434 8588 17436
rect 8612 17434 8668 17436
rect 8692 17434 8748 17436
rect 8452 17382 8498 17434
rect 8498 17382 8508 17434
rect 8532 17382 8562 17434
rect 8562 17382 8574 17434
rect 8574 17382 8588 17434
rect 8612 17382 8626 17434
rect 8626 17382 8638 17434
rect 8638 17382 8668 17434
rect 8692 17382 8702 17434
rect 8702 17382 8748 17434
rect 8452 17380 8508 17382
rect 8532 17380 8588 17382
rect 8612 17380 8668 17382
rect 8692 17380 8748 17382
rect 2830 10362 2886 10364
rect 2910 10362 2966 10364
rect 2990 10362 3046 10364
rect 3070 10362 3126 10364
rect 2830 10310 2876 10362
rect 2876 10310 2886 10362
rect 2910 10310 2940 10362
rect 2940 10310 2952 10362
rect 2952 10310 2966 10362
rect 2990 10310 3004 10362
rect 3004 10310 3016 10362
rect 3016 10310 3046 10362
rect 3070 10310 3080 10362
rect 3080 10310 3126 10362
rect 2830 10308 2886 10310
rect 2910 10308 2966 10310
rect 2990 10308 3046 10310
rect 3070 10308 3126 10310
rect 2830 9274 2886 9276
rect 2910 9274 2966 9276
rect 2990 9274 3046 9276
rect 3070 9274 3126 9276
rect 2830 9222 2876 9274
rect 2876 9222 2886 9274
rect 2910 9222 2940 9274
rect 2940 9222 2952 9274
rect 2952 9222 2966 9274
rect 2990 9222 3004 9274
rect 3004 9222 3016 9274
rect 3016 9222 3046 9274
rect 3070 9222 3080 9274
rect 3080 9222 3126 9274
rect 2830 9220 2886 9222
rect 2910 9220 2966 9222
rect 2990 9220 3046 9222
rect 3070 9220 3126 9222
rect 1490 8356 1546 8392
rect 1490 8336 1492 8356
rect 1492 8336 1544 8356
rect 1544 8336 1546 8356
rect 2830 8186 2886 8188
rect 2910 8186 2966 8188
rect 2990 8186 3046 8188
rect 3070 8186 3126 8188
rect 2830 8134 2876 8186
rect 2876 8134 2886 8186
rect 2910 8134 2940 8186
rect 2940 8134 2952 8186
rect 2952 8134 2966 8186
rect 2990 8134 3004 8186
rect 3004 8134 3016 8186
rect 3016 8134 3046 8186
rect 3070 8134 3080 8186
rect 3080 8134 3126 8186
rect 2830 8132 2886 8134
rect 2910 8132 2966 8134
rect 2990 8132 3046 8134
rect 3070 8132 3126 8134
rect 2830 7098 2886 7100
rect 2910 7098 2966 7100
rect 2990 7098 3046 7100
rect 3070 7098 3126 7100
rect 2830 7046 2876 7098
rect 2876 7046 2886 7098
rect 2910 7046 2940 7098
rect 2940 7046 2952 7098
rect 2952 7046 2966 7098
rect 2990 7046 3004 7098
rect 3004 7046 3016 7098
rect 3016 7046 3046 7098
rect 3070 7046 3080 7098
rect 3080 7046 3126 7098
rect 2830 7044 2886 7046
rect 2910 7044 2966 7046
rect 2990 7044 3046 7046
rect 3070 7044 3126 7046
rect 2830 6010 2886 6012
rect 2910 6010 2966 6012
rect 2990 6010 3046 6012
rect 3070 6010 3126 6012
rect 2830 5958 2876 6010
rect 2876 5958 2886 6010
rect 2910 5958 2940 6010
rect 2940 5958 2952 6010
rect 2952 5958 2966 6010
rect 2990 5958 3004 6010
rect 3004 5958 3016 6010
rect 3016 5958 3046 6010
rect 3070 5958 3080 6010
rect 3080 5958 3126 6010
rect 2830 5956 2886 5958
rect 2910 5956 2966 5958
rect 2990 5956 3046 5958
rect 3070 5956 3126 5958
rect 1490 5092 1546 5128
rect 1490 5072 1492 5092
rect 1492 5072 1544 5092
rect 1544 5072 1546 5092
rect 2830 4922 2886 4924
rect 2910 4922 2966 4924
rect 2990 4922 3046 4924
rect 3070 4922 3126 4924
rect 2830 4870 2876 4922
rect 2876 4870 2886 4922
rect 2910 4870 2940 4922
rect 2940 4870 2952 4922
rect 2952 4870 2966 4922
rect 2990 4870 3004 4922
rect 3004 4870 3016 4922
rect 3016 4870 3046 4922
rect 3070 4870 3080 4922
rect 3080 4870 3126 4922
rect 2830 4868 2886 4870
rect 2910 4868 2966 4870
rect 2990 4868 3046 4870
rect 3070 4868 3126 4870
rect 2830 3834 2886 3836
rect 2910 3834 2966 3836
rect 2990 3834 3046 3836
rect 3070 3834 3126 3836
rect 2830 3782 2876 3834
rect 2876 3782 2886 3834
rect 2910 3782 2940 3834
rect 2940 3782 2952 3834
rect 2952 3782 2966 3834
rect 2990 3782 3004 3834
rect 3004 3782 3016 3834
rect 3016 3782 3046 3834
rect 3070 3782 3080 3834
rect 3080 3782 3126 3834
rect 2830 3780 2886 3782
rect 2910 3780 2966 3782
rect 2990 3780 3046 3782
rect 3070 3780 3126 3782
rect 2830 2746 2886 2748
rect 2910 2746 2966 2748
rect 2990 2746 3046 2748
rect 3070 2746 3126 2748
rect 2830 2694 2876 2746
rect 2876 2694 2886 2746
rect 2910 2694 2940 2746
rect 2940 2694 2952 2746
rect 2952 2694 2966 2746
rect 2990 2694 3004 2746
rect 3004 2694 3016 2746
rect 3016 2694 3046 2746
rect 3070 2694 3080 2746
rect 3080 2694 3126 2746
rect 2830 2692 2886 2694
rect 2910 2692 2966 2694
rect 2990 2692 3046 2694
rect 3070 2692 3126 2694
rect 1858 1808 1914 1864
rect 4704 16346 4760 16348
rect 4784 16346 4840 16348
rect 4864 16346 4920 16348
rect 4944 16346 5000 16348
rect 4704 16294 4750 16346
rect 4750 16294 4760 16346
rect 4784 16294 4814 16346
rect 4814 16294 4826 16346
rect 4826 16294 4840 16346
rect 4864 16294 4878 16346
rect 4878 16294 4890 16346
rect 4890 16294 4920 16346
rect 4944 16294 4954 16346
rect 4954 16294 5000 16346
rect 4704 16292 4760 16294
rect 4784 16292 4840 16294
rect 4864 16292 4920 16294
rect 4944 16292 5000 16294
rect 4704 15258 4760 15260
rect 4784 15258 4840 15260
rect 4864 15258 4920 15260
rect 4944 15258 5000 15260
rect 4704 15206 4750 15258
rect 4750 15206 4760 15258
rect 4784 15206 4814 15258
rect 4814 15206 4826 15258
rect 4826 15206 4840 15258
rect 4864 15206 4878 15258
rect 4878 15206 4890 15258
rect 4890 15206 4920 15258
rect 4944 15206 4954 15258
rect 4954 15206 5000 15258
rect 4704 15204 4760 15206
rect 4784 15204 4840 15206
rect 4864 15204 4920 15206
rect 4944 15204 5000 15206
rect 4704 14170 4760 14172
rect 4784 14170 4840 14172
rect 4864 14170 4920 14172
rect 4944 14170 5000 14172
rect 4704 14118 4750 14170
rect 4750 14118 4760 14170
rect 4784 14118 4814 14170
rect 4814 14118 4826 14170
rect 4826 14118 4840 14170
rect 4864 14118 4878 14170
rect 4878 14118 4890 14170
rect 4890 14118 4920 14170
rect 4944 14118 4954 14170
rect 4954 14118 5000 14170
rect 4704 14116 4760 14118
rect 4784 14116 4840 14118
rect 4864 14116 4920 14118
rect 4944 14116 5000 14118
rect 4704 13082 4760 13084
rect 4784 13082 4840 13084
rect 4864 13082 4920 13084
rect 4944 13082 5000 13084
rect 4704 13030 4750 13082
rect 4750 13030 4760 13082
rect 4784 13030 4814 13082
rect 4814 13030 4826 13082
rect 4826 13030 4840 13082
rect 4864 13030 4878 13082
rect 4878 13030 4890 13082
rect 4890 13030 4920 13082
rect 4944 13030 4954 13082
rect 4954 13030 5000 13082
rect 4704 13028 4760 13030
rect 4784 13028 4840 13030
rect 4864 13028 4920 13030
rect 4944 13028 5000 13030
rect 4704 11994 4760 11996
rect 4784 11994 4840 11996
rect 4864 11994 4920 11996
rect 4944 11994 5000 11996
rect 4704 11942 4750 11994
rect 4750 11942 4760 11994
rect 4784 11942 4814 11994
rect 4814 11942 4826 11994
rect 4826 11942 4840 11994
rect 4864 11942 4878 11994
rect 4878 11942 4890 11994
rect 4890 11942 4920 11994
rect 4944 11942 4954 11994
rect 4954 11942 5000 11994
rect 4704 11940 4760 11942
rect 4784 11940 4840 11942
rect 4864 11940 4920 11942
rect 4944 11940 5000 11942
rect 4704 10906 4760 10908
rect 4784 10906 4840 10908
rect 4864 10906 4920 10908
rect 4944 10906 5000 10908
rect 4704 10854 4750 10906
rect 4750 10854 4760 10906
rect 4784 10854 4814 10906
rect 4814 10854 4826 10906
rect 4826 10854 4840 10906
rect 4864 10854 4878 10906
rect 4878 10854 4890 10906
rect 4890 10854 4920 10906
rect 4944 10854 4954 10906
rect 4954 10854 5000 10906
rect 4704 10852 4760 10854
rect 4784 10852 4840 10854
rect 4864 10852 4920 10854
rect 4944 10852 5000 10854
rect 4704 9818 4760 9820
rect 4784 9818 4840 9820
rect 4864 9818 4920 9820
rect 4944 9818 5000 9820
rect 4704 9766 4750 9818
rect 4750 9766 4760 9818
rect 4784 9766 4814 9818
rect 4814 9766 4826 9818
rect 4826 9766 4840 9818
rect 4864 9766 4878 9818
rect 4878 9766 4890 9818
rect 4890 9766 4920 9818
rect 4944 9766 4954 9818
rect 4954 9766 5000 9818
rect 4704 9764 4760 9766
rect 4784 9764 4840 9766
rect 4864 9764 4920 9766
rect 4944 9764 5000 9766
rect 4434 9424 4490 9480
rect 4704 8730 4760 8732
rect 4784 8730 4840 8732
rect 4864 8730 4920 8732
rect 4944 8730 5000 8732
rect 4704 8678 4750 8730
rect 4750 8678 4760 8730
rect 4784 8678 4814 8730
rect 4814 8678 4826 8730
rect 4826 8678 4840 8730
rect 4864 8678 4878 8730
rect 4878 8678 4890 8730
rect 4890 8678 4920 8730
rect 4944 8678 4954 8730
rect 4954 8678 5000 8730
rect 4704 8676 4760 8678
rect 4784 8676 4840 8678
rect 4864 8676 4920 8678
rect 4944 8676 5000 8678
rect 4704 7642 4760 7644
rect 4784 7642 4840 7644
rect 4864 7642 4920 7644
rect 4944 7642 5000 7644
rect 4704 7590 4750 7642
rect 4750 7590 4760 7642
rect 4784 7590 4814 7642
rect 4814 7590 4826 7642
rect 4826 7590 4840 7642
rect 4864 7590 4878 7642
rect 4878 7590 4890 7642
rect 4890 7590 4920 7642
rect 4944 7590 4954 7642
rect 4954 7590 5000 7642
rect 4704 7588 4760 7590
rect 4784 7588 4840 7590
rect 4864 7588 4920 7590
rect 4944 7588 5000 7590
rect 4704 6554 4760 6556
rect 4784 6554 4840 6556
rect 4864 6554 4920 6556
rect 4944 6554 5000 6556
rect 4704 6502 4750 6554
rect 4750 6502 4760 6554
rect 4784 6502 4814 6554
rect 4814 6502 4826 6554
rect 4826 6502 4840 6554
rect 4864 6502 4878 6554
rect 4878 6502 4890 6554
rect 4890 6502 4920 6554
rect 4944 6502 4954 6554
rect 4954 6502 5000 6554
rect 4704 6500 4760 6502
rect 4784 6500 4840 6502
rect 4864 6500 4920 6502
rect 4944 6500 5000 6502
rect 4704 5466 4760 5468
rect 4784 5466 4840 5468
rect 4864 5466 4920 5468
rect 4944 5466 5000 5468
rect 4704 5414 4750 5466
rect 4750 5414 4760 5466
rect 4784 5414 4814 5466
rect 4814 5414 4826 5466
rect 4826 5414 4840 5466
rect 4864 5414 4878 5466
rect 4878 5414 4890 5466
rect 4890 5414 4920 5466
rect 4944 5414 4954 5466
rect 4954 5414 5000 5466
rect 4704 5412 4760 5414
rect 4784 5412 4840 5414
rect 4864 5412 4920 5414
rect 4944 5412 5000 5414
rect 4704 4378 4760 4380
rect 4784 4378 4840 4380
rect 4864 4378 4920 4380
rect 4944 4378 5000 4380
rect 4704 4326 4750 4378
rect 4750 4326 4760 4378
rect 4784 4326 4814 4378
rect 4814 4326 4826 4378
rect 4826 4326 4840 4378
rect 4864 4326 4878 4378
rect 4878 4326 4890 4378
rect 4890 4326 4920 4378
rect 4944 4326 4954 4378
rect 4954 4326 5000 4378
rect 4704 4324 4760 4326
rect 4784 4324 4840 4326
rect 4864 4324 4920 4326
rect 4944 4324 5000 4326
rect 4704 3290 4760 3292
rect 4784 3290 4840 3292
rect 4864 3290 4920 3292
rect 4944 3290 5000 3292
rect 4704 3238 4750 3290
rect 4750 3238 4760 3290
rect 4784 3238 4814 3290
rect 4814 3238 4826 3290
rect 4826 3238 4840 3290
rect 4864 3238 4878 3290
rect 4878 3238 4890 3290
rect 4890 3238 4920 3290
rect 4944 3238 4954 3290
rect 4954 3238 5000 3290
rect 4704 3236 4760 3238
rect 4784 3236 4840 3238
rect 4864 3236 4920 3238
rect 4944 3236 5000 3238
rect 4704 2202 4760 2204
rect 4784 2202 4840 2204
rect 4864 2202 4920 2204
rect 4944 2202 5000 2204
rect 4704 2150 4750 2202
rect 4750 2150 4760 2202
rect 4784 2150 4814 2202
rect 4814 2150 4826 2202
rect 4826 2150 4840 2202
rect 4864 2150 4878 2202
rect 4878 2150 4890 2202
rect 4890 2150 4920 2202
rect 4944 2150 4954 2202
rect 4954 2150 5000 2202
rect 4704 2148 4760 2150
rect 4784 2148 4840 2150
rect 4864 2148 4920 2150
rect 4944 2148 5000 2150
rect 5446 2488 5502 2544
rect 6578 16890 6634 16892
rect 6658 16890 6714 16892
rect 6738 16890 6794 16892
rect 6818 16890 6874 16892
rect 6578 16838 6624 16890
rect 6624 16838 6634 16890
rect 6658 16838 6688 16890
rect 6688 16838 6700 16890
rect 6700 16838 6714 16890
rect 6738 16838 6752 16890
rect 6752 16838 6764 16890
rect 6764 16838 6794 16890
rect 6818 16838 6828 16890
rect 6828 16838 6874 16890
rect 6578 16836 6634 16838
rect 6658 16836 6714 16838
rect 6738 16836 6794 16838
rect 6818 16836 6874 16838
rect 6578 15802 6634 15804
rect 6658 15802 6714 15804
rect 6738 15802 6794 15804
rect 6818 15802 6874 15804
rect 6578 15750 6624 15802
rect 6624 15750 6634 15802
rect 6658 15750 6688 15802
rect 6688 15750 6700 15802
rect 6700 15750 6714 15802
rect 6738 15750 6752 15802
rect 6752 15750 6764 15802
rect 6764 15750 6794 15802
rect 6818 15750 6828 15802
rect 6828 15750 6874 15802
rect 6578 15748 6634 15750
rect 6658 15748 6714 15750
rect 6738 15748 6794 15750
rect 6818 15748 6874 15750
rect 6578 14714 6634 14716
rect 6658 14714 6714 14716
rect 6738 14714 6794 14716
rect 6818 14714 6874 14716
rect 6578 14662 6624 14714
rect 6624 14662 6634 14714
rect 6658 14662 6688 14714
rect 6688 14662 6700 14714
rect 6700 14662 6714 14714
rect 6738 14662 6752 14714
rect 6752 14662 6764 14714
rect 6764 14662 6794 14714
rect 6818 14662 6828 14714
rect 6828 14662 6874 14714
rect 6578 14660 6634 14662
rect 6658 14660 6714 14662
rect 6738 14660 6794 14662
rect 6818 14660 6874 14662
rect 6578 13626 6634 13628
rect 6658 13626 6714 13628
rect 6738 13626 6794 13628
rect 6818 13626 6874 13628
rect 6578 13574 6624 13626
rect 6624 13574 6634 13626
rect 6658 13574 6688 13626
rect 6688 13574 6700 13626
rect 6700 13574 6714 13626
rect 6738 13574 6752 13626
rect 6752 13574 6764 13626
rect 6764 13574 6794 13626
rect 6818 13574 6828 13626
rect 6828 13574 6874 13626
rect 6578 13572 6634 13574
rect 6658 13572 6714 13574
rect 6738 13572 6794 13574
rect 6818 13572 6874 13574
rect 6578 12538 6634 12540
rect 6658 12538 6714 12540
rect 6738 12538 6794 12540
rect 6818 12538 6874 12540
rect 6578 12486 6624 12538
rect 6624 12486 6634 12538
rect 6658 12486 6688 12538
rect 6688 12486 6700 12538
rect 6700 12486 6714 12538
rect 6738 12486 6752 12538
rect 6752 12486 6764 12538
rect 6764 12486 6794 12538
rect 6818 12486 6828 12538
rect 6828 12486 6874 12538
rect 6578 12484 6634 12486
rect 6658 12484 6714 12486
rect 6738 12484 6794 12486
rect 6818 12484 6874 12486
rect 6578 11450 6634 11452
rect 6658 11450 6714 11452
rect 6738 11450 6794 11452
rect 6818 11450 6874 11452
rect 6578 11398 6624 11450
rect 6624 11398 6634 11450
rect 6658 11398 6688 11450
rect 6688 11398 6700 11450
rect 6700 11398 6714 11450
rect 6738 11398 6752 11450
rect 6752 11398 6764 11450
rect 6764 11398 6794 11450
rect 6818 11398 6828 11450
rect 6828 11398 6874 11450
rect 6578 11396 6634 11398
rect 6658 11396 6714 11398
rect 6738 11396 6794 11398
rect 6818 11396 6874 11398
rect 6826 10668 6882 10704
rect 6826 10648 6828 10668
rect 6828 10648 6880 10668
rect 6880 10648 6882 10668
rect 6274 9696 6330 9752
rect 6578 10362 6634 10364
rect 6658 10362 6714 10364
rect 6738 10362 6794 10364
rect 6818 10362 6874 10364
rect 6578 10310 6624 10362
rect 6624 10310 6634 10362
rect 6658 10310 6688 10362
rect 6688 10310 6700 10362
rect 6700 10310 6714 10362
rect 6738 10310 6752 10362
rect 6752 10310 6764 10362
rect 6764 10310 6794 10362
rect 6818 10310 6828 10362
rect 6828 10310 6874 10362
rect 6578 10308 6634 10310
rect 6658 10308 6714 10310
rect 6738 10308 6794 10310
rect 6818 10308 6874 10310
rect 6578 9274 6634 9276
rect 6658 9274 6714 9276
rect 6738 9274 6794 9276
rect 6818 9274 6874 9276
rect 6578 9222 6624 9274
rect 6624 9222 6634 9274
rect 6658 9222 6688 9274
rect 6688 9222 6700 9274
rect 6700 9222 6714 9274
rect 6738 9222 6752 9274
rect 6752 9222 6764 9274
rect 6764 9222 6794 9274
rect 6818 9222 6828 9274
rect 6828 9222 6874 9274
rect 6578 9220 6634 9222
rect 6658 9220 6714 9222
rect 6738 9220 6794 9222
rect 6818 9220 6874 9222
rect 6578 8186 6634 8188
rect 6658 8186 6714 8188
rect 6738 8186 6794 8188
rect 6818 8186 6874 8188
rect 6578 8134 6624 8186
rect 6624 8134 6634 8186
rect 6658 8134 6688 8186
rect 6688 8134 6700 8186
rect 6700 8134 6714 8186
rect 6738 8134 6752 8186
rect 6752 8134 6764 8186
rect 6764 8134 6794 8186
rect 6818 8134 6828 8186
rect 6828 8134 6874 8186
rect 6578 8132 6634 8134
rect 6658 8132 6714 8134
rect 6738 8132 6794 8134
rect 6818 8132 6874 8134
rect 6578 7098 6634 7100
rect 6658 7098 6714 7100
rect 6738 7098 6794 7100
rect 6818 7098 6874 7100
rect 6578 7046 6624 7098
rect 6624 7046 6634 7098
rect 6658 7046 6688 7098
rect 6688 7046 6700 7098
rect 6700 7046 6714 7098
rect 6738 7046 6752 7098
rect 6752 7046 6764 7098
rect 6764 7046 6794 7098
rect 6818 7046 6828 7098
rect 6828 7046 6874 7098
rect 6578 7044 6634 7046
rect 6658 7044 6714 7046
rect 6738 7044 6794 7046
rect 6818 7044 6874 7046
rect 6578 6010 6634 6012
rect 6658 6010 6714 6012
rect 6738 6010 6794 6012
rect 6818 6010 6874 6012
rect 6578 5958 6624 6010
rect 6624 5958 6634 6010
rect 6658 5958 6688 6010
rect 6688 5958 6700 6010
rect 6700 5958 6714 6010
rect 6738 5958 6752 6010
rect 6752 5958 6764 6010
rect 6764 5958 6794 6010
rect 6818 5958 6828 6010
rect 6828 5958 6874 6010
rect 6578 5956 6634 5958
rect 6658 5956 6714 5958
rect 6738 5956 6794 5958
rect 6818 5956 6874 5958
rect 6578 4922 6634 4924
rect 6658 4922 6714 4924
rect 6738 4922 6794 4924
rect 6818 4922 6874 4924
rect 6578 4870 6624 4922
rect 6624 4870 6634 4922
rect 6658 4870 6688 4922
rect 6688 4870 6700 4922
rect 6700 4870 6714 4922
rect 6738 4870 6752 4922
rect 6752 4870 6764 4922
rect 6764 4870 6794 4922
rect 6818 4870 6828 4922
rect 6828 4870 6874 4922
rect 6578 4868 6634 4870
rect 6658 4868 6714 4870
rect 6738 4868 6794 4870
rect 6818 4868 6874 4870
rect 6578 3834 6634 3836
rect 6658 3834 6714 3836
rect 6738 3834 6794 3836
rect 6818 3834 6874 3836
rect 6578 3782 6624 3834
rect 6624 3782 6634 3834
rect 6658 3782 6688 3834
rect 6688 3782 6700 3834
rect 6700 3782 6714 3834
rect 6738 3782 6752 3834
rect 6752 3782 6764 3834
rect 6764 3782 6794 3834
rect 6818 3782 6828 3834
rect 6828 3782 6874 3834
rect 6578 3780 6634 3782
rect 6658 3780 6714 3782
rect 6738 3780 6794 3782
rect 6818 3780 6874 3782
rect 6578 2746 6634 2748
rect 6658 2746 6714 2748
rect 6738 2746 6794 2748
rect 6818 2746 6874 2748
rect 6578 2694 6624 2746
rect 6624 2694 6634 2746
rect 6658 2694 6688 2746
rect 6688 2694 6700 2746
rect 6700 2694 6714 2746
rect 6738 2694 6752 2746
rect 6752 2694 6764 2746
rect 6764 2694 6794 2746
rect 6818 2694 6828 2746
rect 6828 2694 6874 2746
rect 6578 2692 6634 2694
rect 6658 2692 6714 2694
rect 6738 2692 6794 2694
rect 6818 2692 6874 2694
rect 8452 16346 8508 16348
rect 8532 16346 8588 16348
rect 8612 16346 8668 16348
rect 8692 16346 8748 16348
rect 8452 16294 8498 16346
rect 8498 16294 8508 16346
rect 8532 16294 8562 16346
rect 8562 16294 8574 16346
rect 8574 16294 8588 16346
rect 8612 16294 8626 16346
rect 8626 16294 8638 16346
rect 8638 16294 8668 16346
rect 8692 16294 8702 16346
rect 8702 16294 8748 16346
rect 8452 16292 8508 16294
rect 8532 16292 8588 16294
rect 8612 16292 8668 16294
rect 8692 16292 8748 16294
rect 8452 15258 8508 15260
rect 8532 15258 8588 15260
rect 8612 15258 8668 15260
rect 8692 15258 8748 15260
rect 8452 15206 8498 15258
rect 8498 15206 8508 15258
rect 8532 15206 8562 15258
rect 8562 15206 8574 15258
rect 8574 15206 8588 15258
rect 8612 15206 8626 15258
rect 8626 15206 8638 15258
rect 8638 15206 8668 15258
rect 8692 15206 8702 15258
rect 8702 15206 8748 15258
rect 8452 15204 8508 15206
rect 8532 15204 8588 15206
rect 8612 15204 8668 15206
rect 8692 15204 8748 15206
rect 8452 14170 8508 14172
rect 8532 14170 8588 14172
rect 8612 14170 8668 14172
rect 8692 14170 8748 14172
rect 8452 14118 8498 14170
rect 8498 14118 8508 14170
rect 8532 14118 8562 14170
rect 8562 14118 8574 14170
rect 8574 14118 8588 14170
rect 8612 14118 8626 14170
rect 8626 14118 8638 14170
rect 8638 14118 8668 14170
rect 8692 14118 8702 14170
rect 8702 14118 8748 14170
rect 8452 14116 8508 14118
rect 8532 14116 8588 14118
rect 8612 14116 8668 14118
rect 8692 14116 8748 14118
rect 8452 13082 8508 13084
rect 8532 13082 8588 13084
rect 8612 13082 8668 13084
rect 8692 13082 8748 13084
rect 8452 13030 8498 13082
rect 8498 13030 8508 13082
rect 8532 13030 8562 13082
rect 8562 13030 8574 13082
rect 8574 13030 8588 13082
rect 8612 13030 8626 13082
rect 8626 13030 8638 13082
rect 8638 13030 8668 13082
rect 8692 13030 8702 13082
rect 8702 13030 8748 13082
rect 8452 13028 8508 13030
rect 8532 13028 8588 13030
rect 8612 13028 8668 13030
rect 8692 13028 8748 13030
rect 7746 11056 7802 11112
rect 8022 11056 8078 11112
rect 7746 10104 7802 10160
rect 8452 11994 8508 11996
rect 8532 11994 8588 11996
rect 8612 11994 8668 11996
rect 8692 11994 8748 11996
rect 8452 11942 8498 11994
rect 8498 11942 8508 11994
rect 8532 11942 8562 11994
rect 8562 11942 8574 11994
rect 8574 11942 8588 11994
rect 8612 11942 8626 11994
rect 8626 11942 8638 11994
rect 8638 11942 8668 11994
rect 8692 11942 8702 11994
rect 8702 11942 8748 11994
rect 8452 11940 8508 11942
rect 8532 11940 8588 11942
rect 8612 11940 8668 11942
rect 8692 11940 8748 11942
rect 8452 10906 8508 10908
rect 8532 10906 8588 10908
rect 8612 10906 8668 10908
rect 8692 10906 8748 10908
rect 8452 10854 8498 10906
rect 8498 10854 8508 10906
rect 8532 10854 8562 10906
rect 8562 10854 8574 10906
rect 8574 10854 8588 10906
rect 8612 10854 8626 10906
rect 8626 10854 8638 10906
rect 8638 10854 8668 10906
rect 8692 10854 8702 10906
rect 8702 10854 8748 10906
rect 8452 10852 8508 10854
rect 8532 10852 8588 10854
rect 8612 10852 8668 10854
rect 8692 10852 8748 10854
rect 8666 10240 8722 10296
rect 9034 10240 9090 10296
rect 8298 9968 8354 10024
rect 8452 9818 8508 9820
rect 8532 9818 8588 9820
rect 8612 9818 8668 9820
rect 8692 9818 8748 9820
rect 8452 9766 8498 9818
rect 8498 9766 8508 9818
rect 8532 9766 8562 9818
rect 8562 9766 8574 9818
rect 8574 9766 8588 9818
rect 8612 9766 8626 9818
rect 8626 9766 8638 9818
rect 8638 9766 8668 9818
rect 8692 9766 8702 9818
rect 8702 9766 8748 9818
rect 8452 9764 8508 9766
rect 8532 9764 8588 9766
rect 8612 9764 8668 9766
rect 8692 9764 8748 9766
rect 8390 9424 8446 9480
rect 8850 9696 8906 9752
rect 8452 8730 8508 8732
rect 8532 8730 8588 8732
rect 8612 8730 8668 8732
rect 8692 8730 8748 8732
rect 8452 8678 8498 8730
rect 8498 8678 8508 8730
rect 8532 8678 8562 8730
rect 8562 8678 8574 8730
rect 8574 8678 8588 8730
rect 8612 8678 8626 8730
rect 8626 8678 8638 8730
rect 8638 8678 8668 8730
rect 8692 8678 8702 8730
rect 8702 8678 8748 8730
rect 8452 8676 8508 8678
rect 8532 8676 8588 8678
rect 8612 8676 8668 8678
rect 8692 8676 8748 8678
rect 9034 9832 9090 9888
rect 10326 16890 10382 16892
rect 10406 16890 10462 16892
rect 10486 16890 10542 16892
rect 10566 16890 10622 16892
rect 10326 16838 10372 16890
rect 10372 16838 10382 16890
rect 10406 16838 10436 16890
rect 10436 16838 10448 16890
rect 10448 16838 10462 16890
rect 10486 16838 10500 16890
rect 10500 16838 10512 16890
rect 10512 16838 10542 16890
rect 10566 16838 10576 16890
rect 10576 16838 10622 16890
rect 10326 16836 10382 16838
rect 10406 16836 10462 16838
rect 10486 16836 10542 16838
rect 10566 16836 10622 16838
rect 8942 8880 8998 8936
rect 8850 8472 8906 8528
rect 8452 7642 8508 7644
rect 8532 7642 8588 7644
rect 8612 7642 8668 7644
rect 8692 7642 8748 7644
rect 8452 7590 8498 7642
rect 8498 7590 8508 7642
rect 8532 7590 8562 7642
rect 8562 7590 8574 7642
rect 8574 7590 8588 7642
rect 8612 7590 8626 7642
rect 8626 7590 8638 7642
rect 8638 7590 8668 7642
rect 8692 7590 8702 7642
rect 8702 7590 8748 7642
rect 8452 7588 8508 7590
rect 8532 7588 8588 7590
rect 8612 7588 8668 7590
rect 8692 7588 8748 7590
rect 8452 6554 8508 6556
rect 8532 6554 8588 6556
rect 8612 6554 8668 6556
rect 8692 6554 8748 6556
rect 8452 6502 8498 6554
rect 8498 6502 8508 6554
rect 8532 6502 8562 6554
rect 8562 6502 8574 6554
rect 8574 6502 8588 6554
rect 8612 6502 8626 6554
rect 8626 6502 8638 6554
rect 8638 6502 8668 6554
rect 8692 6502 8702 6554
rect 8702 6502 8748 6554
rect 8452 6500 8508 6502
rect 8532 6500 8588 6502
rect 8612 6500 8668 6502
rect 8692 6500 8748 6502
rect 8452 5466 8508 5468
rect 8532 5466 8588 5468
rect 8612 5466 8668 5468
rect 8692 5466 8748 5468
rect 8452 5414 8498 5466
rect 8498 5414 8508 5466
rect 8532 5414 8562 5466
rect 8562 5414 8574 5466
rect 8574 5414 8588 5466
rect 8612 5414 8626 5466
rect 8626 5414 8638 5466
rect 8638 5414 8668 5466
rect 8692 5414 8702 5466
rect 8702 5414 8748 5466
rect 8452 5412 8508 5414
rect 8532 5412 8588 5414
rect 8612 5412 8668 5414
rect 8692 5412 8748 5414
rect 8452 4378 8508 4380
rect 8532 4378 8588 4380
rect 8612 4378 8668 4380
rect 8692 4378 8748 4380
rect 8452 4326 8498 4378
rect 8498 4326 8508 4378
rect 8532 4326 8562 4378
rect 8562 4326 8574 4378
rect 8574 4326 8588 4378
rect 8612 4326 8626 4378
rect 8626 4326 8638 4378
rect 8638 4326 8668 4378
rect 8692 4326 8702 4378
rect 8702 4326 8748 4378
rect 8452 4324 8508 4326
rect 8532 4324 8588 4326
rect 8612 4324 8668 4326
rect 8692 4324 8748 4326
rect 8452 3290 8508 3292
rect 8532 3290 8588 3292
rect 8612 3290 8668 3292
rect 8692 3290 8748 3292
rect 8452 3238 8498 3290
rect 8498 3238 8508 3290
rect 8532 3238 8562 3290
rect 8562 3238 8574 3290
rect 8574 3238 8588 3290
rect 8612 3238 8626 3290
rect 8626 3238 8638 3290
rect 8638 3238 8668 3290
rect 8692 3238 8702 3290
rect 8702 3238 8748 3290
rect 8452 3236 8508 3238
rect 8532 3236 8588 3238
rect 8612 3236 8668 3238
rect 8692 3236 8748 3238
rect 8452 2202 8508 2204
rect 8532 2202 8588 2204
rect 8612 2202 8668 2204
rect 8692 2202 8748 2204
rect 8452 2150 8498 2202
rect 8498 2150 8508 2202
rect 8532 2150 8562 2202
rect 8562 2150 8574 2202
rect 8574 2150 8588 2202
rect 8612 2150 8626 2202
rect 8626 2150 8638 2202
rect 8638 2150 8668 2202
rect 8692 2150 8702 2202
rect 8702 2150 8748 2202
rect 8452 2148 8508 2150
rect 8532 2148 8588 2150
rect 8612 2148 8668 2150
rect 8692 2148 8748 2150
rect 9586 9696 9642 9752
rect 9586 9580 9642 9616
rect 9586 9560 9588 9580
rect 9588 9560 9640 9580
rect 9640 9560 9642 9580
rect 9586 8744 9642 8800
rect 9954 2488 10010 2544
rect 10326 15802 10382 15804
rect 10406 15802 10462 15804
rect 10486 15802 10542 15804
rect 10566 15802 10622 15804
rect 10326 15750 10372 15802
rect 10372 15750 10382 15802
rect 10406 15750 10436 15802
rect 10436 15750 10448 15802
rect 10448 15750 10462 15802
rect 10486 15750 10500 15802
rect 10500 15750 10512 15802
rect 10512 15750 10542 15802
rect 10566 15750 10576 15802
rect 10576 15750 10622 15802
rect 10326 15748 10382 15750
rect 10406 15748 10462 15750
rect 10486 15748 10542 15750
rect 10566 15748 10622 15750
rect 10326 14714 10382 14716
rect 10406 14714 10462 14716
rect 10486 14714 10542 14716
rect 10566 14714 10622 14716
rect 10326 14662 10372 14714
rect 10372 14662 10382 14714
rect 10406 14662 10436 14714
rect 10436 14662 10448 14714
rect 10448 14662 10462 14714
rect 10486 14662 10500 14714
rect 10500 14662 10512 14714
rect 10512 14662 10542 14714
rect 10566 14662 10576 14714
rect 10576 14662 10622 14714
rect 10326 14660 10382 14662
rect 10406 14660 10462 14662
rect 10486 14660 10542 14662
rect 10566 14660 10622 14662
rect 10326 13626 10382 13628
rect 10406 13626 10462 13628
rect 10486 13626 10542 13628
rect 10566 13626 10622 13628
rect 10326 13574 10372 13626
rect 10372 13574 10382 13626
rect 10406 13574 10436 13626
rect 10436 13574 10448 13626
rect 10448 13574 10462 13626
rect 10486 13574 10500 13626
rect 10500 13574 10512 13626
rect 10512 13574 10542 13626
rect 10566 13574 10576 13626
rect 10576 13574 10622 13626
rect 10326 13572 10382 13574
rect 10406 13572 10462 13574
rect 10486 13572 10542 13574
rect 10566 13572 10622 13574
rect 10326 12538 10382 12540
rect 10406 12538 10462 12540
rect 10486 12538 10542 12540
rect 10566 12538 10622 12540
rect 10326 12486 10372 12538
rect 10372 12486 10382 12538
rect 10406 12486 10436 12538
rect 10436 12486 10448 12538
rect 10448 12486 10462 12538
rect 10486 12486 10500 12538
rect 10500 12486 10512 12538
rect 10512 12486 10542 12538
rect 10566 12486 10576 12538
rect 10576 12486 10622 12538
rect 10326 12484 10382 12486
rect 10406 12484 10462 12486
rect 10486 12484 10542 12486
rect 10566 12484 10622 12486
rect 10326 11450 10382 11452
rect 10406 11450 10462 11452
rect 10486 11450 10542 11452
rect 10566 11450 10622 11452
rect 10326 11398 10372 11450
rect 10372 11398 10382 11450
rect 10406 11398 10436 11450
rect 10436 11398 10448 11450
rect 10448 11398 10462 11450
rect 10486 11398 10500 11450
rect 10500 11398 10512 11450
rect 10512 11398 10542 11450
rect 10566 11398 10576 11450
rect 10576 11398 10622 11450
rect 10326 11396 10382 11398
rect 10406 11396 10462 11398
rect 10486 11396 10542 11398
rect 10566 11396 10622 11398
rect 10326 10362 10382 10364
rect 10406 10362 10462 10364
rect 10486 10362 10542 10364
rect 10566 10362 10622 10364
rect 10326 10310 10372 10362
rect 10372 10310 10382 10362
rect 10406 10310 10436 10362
rect 10436 10310 10448 10362
rect 10448 10310 10462 10362
rect 10486 10310 10500 10362
rect 10500 10310 10512 10362
rect 10512 10310 10542 10362
rect 10566 10310 10576 10362
rect 10576 10310 10622 10362
rect 10326 10308 10382 10310
rect 10406 10308 10462 10310
rect 10486 10308 10542 10310
rect 10566 10308 10622 10310
rect 10230 9560 10286 9616
rect 10230 9444 10286 9480
rect 10230 9424 10232 9444
rect 10232 9424 10284 9444
rect 10284 9424 10286 9444
rect 10326 9274 10382 9276
rect 10406 9274 10462 9276
rect 10486 9274 10542 9276
rect 10566 9274 10622 9276
rect 10326 9222 10372 9274
rect 10372 9222 10382 9274
rect 10406 9222 10436 9274
rect 10436 9222 10448 9274
rect 10448 9222 10462 9274
rect 10486 9222 10500 9274
rect 10500 9222 10512 9274
rect 10512 9222 10542 9274
rect 10566 9222 10576 9274
rect 10576 9222 10622 9274
rect 10326 9220 10382 9222
rect 10406 9220 10462 9222
rect 10486 9220 10542 9222
rect 10566 9220 10622 9222
rect 10966 16632 11022 16688
rect 10326 8186 10382 8188
rect 10406 8186 10462 8188
rect 10486 8186 10542 8188
rect 10566 8186 10622 8188
rect 10326 8134 10372 8186
rect 10372 8134 10382 8186
rect 10406 8134 10436 8186
rect 10436 8134 10448 8186
rect 10448 8134 10462 8186
rect 10486 8134 10500 8186
rect 10500 8134 10512 8186
rect 10512 8134 10542 8186
rect 10566 8134 10576 8186
rect 10576 8134 10622 8186
rect 10326 8132 10382 8134
rect 10406 8132 10462 8134
rect 10486 8132 10542 8134
rect 10566 8132 10622 8134
rect 10326 7098 10382 7100
rect 10406 7098 10462 7100
rect 10486 7098 10542 7100
rect 10566 7098 10622 7100
rect 10326 7046 10372 7098
rect 10372 7046 10382 7098
rect 10406 7046 10436 7098
rect 10436 7046 10448 7098
rect 10448 7046 10462 7098
rect 10486 7046 10500 7098
rect 10500 7046 10512 7098
rect 10512 7046 10542 7098
rect 10566 7046 10576 7098
rect 10576 7046 10622 7098
rect 10326 7044 10382 7046
rect 10406 7044 10462 7046
rect 10486 7044 10542 7046
rect 10566 7044 10622 7046
rect 10326 6010 10382 6012
rect 10406 6010 10462 6012
rect 10486 6010 10542 6012
rect 10566 6010 10622 6012
rect 10326 5958 10372 6010
rect 10372 5958 10382 6010
rect 10406 5958 10436 6010
rect 10436 5958 10448 6010
rect 10448 5958 10462 6010
rect 10486 5958 10500 6010
rect 10500 5958 10512 6010
rect 10512 5958 10542 6010
rect 10566 5958 10576 6010
rect 10576 5958 10622 6010
rect 10326 5956 10382 5958
rect 10406 5956 10462 5958
rect 10486 5956 10542 5958
rect 10566 5956 10622 5958
rect 10326 4922 10382 4924
rect 10406 4922 10462 4924
rect 10486 4922 10542 4924
rect 10566 4922 10622 4924
rect 10326 4870 10372 4922
rect 10372 4870 10382 4922
rect 10406 4870 10436 4922
rect 10436 4870 10448 4922
rect 10448 4870 10462 4922
rect 10486 4870 10500 4922
rect 10500 4870 10512 4922
rect 10512 4870 10542 4922
rect 10566 4870 10576 4922
rect 10576 4870 10622 4922
rect 10326 4868 10382 4870
rect 10406 4868 10462 4870
rect 10486 4868 10542 4870
rect 10566 4868 10622 4870
rect 10326 3834 10382 3836
rect 10406 3834 10462 3836
rect 10486 3834 10542 3836
rect 10566 3834 10622 3836
rect 10326 3782 10372 3834
rect 10372 3782 10382 3834
rect 10406 3782 10436 3834
rect 10436 3782 10448 3834
rect 10448 3782 10462 3834
rect 10486 3782 10500 3834
rect 10500 3782 10512 3834
rect 10512 3782 10542 3834
rect 10566 3782 10576 3834
rect 10576 3782 10622 3834
rect 10326 3780 10382 3782
rect 10406 3780 10462 3782
rect 10486 3780 10542 3782
rect 10566 3780 10622 3782
rect 10326 2746 10382 2748
rect 10406 2746 10462 2748
rect 10486 2746 10542 2748
rect 10566 2746 10622 2748
rect 10326 2694 10372 2746
rect 10372 2694 10382 2746
rect 10406 2694 10436 2746
rect 10436 2694 10448 2746
rect 10448 2694 10462 2746
rect 10486 2694 10500 2746
rect 10500 2694 10512 2746
rect 10512 2694 10542 2746
rect 10566 2694 10576 2746
rect 10576 2694 10622 2746
rect 10326 2692 10382 2694
rect 10406 2692 10462 2694
rect 10486 2692 10542 2694
rect 10566 2692 10622 2694
rect 12200 17434 12256 17436
rect 12280 17434 12336 17436
rect 12360 17434 12416 17436
rect 12440 17434 12496 17436
rect 12200 17382 12246 17434
rect 12246 17382 12256 17434
rect 12280 17382 12310 17434
rect 12310 17382 12322 17434
rect 12322 17382 12336 17434
rect 12360 17382 12374 17434
rect 12374 17382 12386 17434
rect 12386 17382 12416 17434
rect 12440 17382 12450 17434
rect 12450 17382 12496 17434
rect 12200 17380 12256 17382
rect 12280 17380 12336 17382
rect 12360 17380 12416 17382
rect 12440 17380 12496 17382
rect 12200 16346 12256 16348
rect 12280 16346 12336 16348
rect 12360 16346 12416 16348
rect 12440 16346 12496 16348
rect 12200 16294 12246 16346
rect 12246 16294 12256 16346
rect 12280 16294 12310 16346
rect 12310 16294 12322 16346
rect 12322 16294 12336 16346
rect 12360 16294 12374 16346
rect 12374 16294 12386 16346
rect 12386 16294 12416 16346
rect 12440 16294 12450 16346
rect 12450 16294 12496 16346
rect 12200 16292 12256 16294
rect 12280 16292 12336 16294
rect 12360 16292 12416 16294
rect 12440 16292 12496 16294
rect 12200 15258 12256 15260
rect 12280 15258 12336 15260
rect 12360 15258 12416 15260
rect 12440 15258 12496 15260
rect 12200 15206 12246 15258
rect 12246 15206 12256 15258
rect 12280 15206 12310 15258
rect 12310 15206 12322 15258
rect 12322 15206 12336 15258
rect 12360 15206 12374 15258
rect 12374 15206 12386 15258
rect 12386 15206 12416 15258
rect 12440 15206 12450 15258
rect 12450 15206 12496 15258
rect 12200 15204 12256 15206
rect 12280 15204 12336 15206
rect 12360 15204 12416 15206
rect 12440 15204 12496 15206
rect 12200 14170 12256 14172
rect 12280 14170 12336 14172
rect 12360 14170 12416 14172
rect 12440 14170 12496 14172
rect 12200 14118 12246 14170
rect 12246 14118 12256 14170
rect 12280 14118 12310 14170
rect 12310 14118 12322 14170
rect 12322 14118 12336 14170
rect 12360 14118 12374 14170
rect 12374 14118 12386 14170
rect 12386 14118 12416 14170
rect 12440 14118 12450 14170
rect 12450 14118 12496 14170
rect 12200 14116 12256 14118
rect 12280 14116 12336 14118
rect 12360 14116 12416 14118
rect 12440 14116 12496 14118
rect 12200 13082 12256 13084
rect 12280 13082 12336 13084
rect 12360 13082 12416 13084
rect 12440 13082 12496 13084
rect 12200 13030 12246 13082
rect 12246 13030 12256 13082
rect 12280 13030 12310 13082
rect 12310 13030 12322 13082
rect 12322 13030 12336 13082
rect 12360 13030 12374 13082
rect 12374 13030 12386 13082
rect 12386 13030 12416 13082
rect 12440 13030 12450 13082
rect 12450 13030 12496 13082
rect 12200 13028 12256 13030
rect 12280 13028 12336 13030
rect 12360 13028 12416 13030
rect 12440 13028 12496 13030
rect 12200 11994 12256 11996
rect 12280 11994 12336 11996
rect 12360 11994 12416 11996
rect 12440 11994 12496 11996
rect 12200 11942 12246 11994
rect 12246 11942 12256 11994
rect 12280 11942 12310 11994
rect 12310 11942 12322 11994
rect 12322 11942 12336 11994
rect 12360 11942 12374 11994
rect 12374 11942 12386 11994
rect 12386 11942 12416 11994
rect 12440 11942 12450 11994
rect 12450 11942 12496 11994
rect 12200 11940 12256 11942
rect 12280 11940 12336 11942
rect 12360 11940 12416 11942
rect 12440 11940 12496 11942
rect 12200 10906 12256 10908
rect 12280 10906 12336 10908
rect 12360 10906 12416 10908
rect 12440 10906 12496 10908
rect 12200 10854 12246 10906
rect 12246 10854 12256 10906
rect 12280 10854 12310 10906
rect 12310 10854 12322 10906
rect 12322 10854 12336 10906
rect 12360 10854 12374 10906
rect 12374 10854 12386 10906
rect 12386 10854 12416 10906
rect 12440 10854 12450 10906
rect 12450 10854 12496 10906
rect 12200 10852 12256 10854
rect 12280 10852 12336 10854
rect 12360 10852 12416 10854
rect 12440 10852 12496 10854
rect 11794 10648 11850 10704
rect 11518 2488 11574 2544
rect 12806 16632 12862 16688
rect 14074 16890 14130 16892
rect 14154 16890 14210 16892
rect 14234 16890 14290 16892
rect 14314 16890 14370 16892
rect 14074 16838 14120 16890
rect 14120 16838 14130 16890
rect 14154 16838 14184 16890
rect 14184 16838 14196 16890
rect 14196 16838 14210 16890
rect 14234 16838 14248 16890
rect 14248 16838 14260 16890
rect 14260 16838 14290 16890
rect 14314 16838 14324 16890
rect 14324 16838 14370 16890
rect 14074 16836 14130 16838
rect 14154 16836 14210 16838
rect 14234 16836 14290 16838
rect 14314 16836 14370 16838
rect 14074 15802 14130 15804
rect 14154 15802 14210 15804
rect 14234 15802 14290 15804
rect 14314 15802 14370 15804
rect 14074 15750 14120 15802
rect 14120 15750 14130 15802
rect 14154 15750 14184 15802
rect 14184 15750 14196 15802
rect 14196 15750 14210 15802
rect 14234 15750 14248 15802
rect 14248 15750 14260 15802
rect 14260 15750 14290 15802
rect 14314 15750 14324 15802
rect 14324 15750 14370 15802
rect 14074 15748 14130 15750
rect 14154 15748 14210 15750
rect 14234 15748 14290 15750
rect 14314 15748 14370 15750
rect 14074 14714 14130 14716
rect 14154 14714 14210 14716
rect 14234 14714 14290 14716
rect 14314 14714 14370 14716
rect 14074 14662 14120 14714
rect 14120 14662 14130 14714
rect 14154 14662 14184 14714
rect 14184 14662 14196 14714
rect 14196 14662 14210 14714
rect 14234 14662 14248 14714
rect 14248 14662 14260 14714
rect 14260 14662 14290 14714
rect 14314 14662 14324 14714
rect 14324 14662 14370 14714
rect 14074 14660 14130 14662
rect 14154 14660 14210 14662
rect 14234 14660 14290 14662
rect 14314 14660 14370 14662
rect 14074 13626 14130 13628
rect 14154 13626 14210 13628
rect 14234 13626 14290 13628
rect 14314 13626 14370 13628
rect 14074 13574 14120 13626
rect 14120 13574 14130 13626
rect 14154 13574 14184 13626
rect 14184 13574 14196 13626
rect 14196 13574 14210 13626
rect 14234 13574 14248 13626
rect 14248 13574 14260 13626
rect 14260 13574 14290 13626
rect 14314 13574 14324 13626
rect 14324 13574 14370 13626
rect 14074 13572 14130 13574
rect 14154 13572 14210 13574
rect 14234 13572 14290 13574
rect 14314 13572 14370 13574
rect 14074 12538 14130 12540
rect 14154 12538 14210 12540
rect 14234 12538 14290 12540
rect 14314 12538 14370 12540
rect 14074 12486 14120 12538
rect 14120 12486 14130 12538
rect 14154 12486 14184 12538
rect 14184 12486 14196 12538
rect 14196 12486 14210 12538
rect 14234 12486 14248 12538
rect 14248 12486 14260 12538
rect 14260 12486 14290 12538
rect 14314 12486 14324 12538
rect 14324 12486 14370 12538
rect 14074 12484 14130 12486
rect 14154 12484 14210 12486
rect 14234 12484 14290 12486
rect 14314 12484 14370 12486
rect 14074 11450 14130 11452
rect 14154 11450 14210 11452
rect 14234 11450 14290 11452
rect 14314 11450 14370 11452
rect 14074 11398 14120 11450
rect 14120 11398 14130 11450
rect 14154 11398 14184 11450
rect 14184 11398 14196 11450
rect 14196 11398 14210 11450
rect 14234 11398 14248 11450
rect 14248 11398 14260 11450
rect 14260 11398 14290 11450
rect 14314 11398 14324 11450
rect 14324 11398 14370 11450
rect 14074 11396 14130 11398
rect 14154 11396 14210 11398
rect 14234 11396 14290 11398
rect 14314 11396 14370 11398
rect 15566 17332 15622 17368
rect 15566 17312 15568 17332
rect 15568 17312 15620 17332
rect 15620 17312 15622 17332
rect 14074 10362 14130 10364
rect 14154 10362 14210 10364
rect 14234 10362 14290 10364
rect 14314 10362 14370 10364
rect 14074 10310 14120 10362
rect 14120 10310 14130 10362
rect 14154 10310 14184 10362
rect 14184 10310 14196 10362
rect 14196 10310 14210 10362
rect 14234 10310 14248 10362
rect 14248 10310 14260 10362
rect 14260 10310 14290 10362
rect 14314 10310 14324 10362
rect 14324 10310 14370 10362
rect 14074 10308 14130 10310
rect 14154 10308 14210 10310
rect 14234 10308 14290 10310
rect 14314 10308 14370 10310
rect 13910 10104 13966 10160
rect 12200 9818 12256 9820
rect 12280 9818 12336 9820
rect 12360 9818 12416 9820
rect 12440 9818 12496 9820
rect 12200 9766 12246 9818
rect 12246 9766 12256 9818
rect 12280 9766 12310 9818
rect 12310 9766 12322 9818
rect 12322 9766 12336 9818
rect 12360 9766 12374 9818
rect 12374 9766 12386 9818
rect 12386 9766 12416 9818
rect 12440 9766 12450 9818
rect 12450 9766 12496 9818
rect 12200 9764 12256 9766
rect 12280 9764 12336 9766
rect 12360 9764 12416 9766
rect 12440 9764 12496 9766
rect 12200 8730 12256 8732
rect 12280 8730 12336 8732
rect 12360 8730 12416 8732
rect 12440 8730 12496 8732
rect 12200 8678 12246 8730
rect 12246 8678 12256 8730
rect 12280 8678 12310 8730
rect 12310 8678 12322 8730
rect 12322 8678 12336 8730
rect 12360 8678 12374 8730
rect 12374 8678 12386 8730
rect 12386 8678 12416 8730
rect 12440 8678 12450 8730
rect 12450 8678 12496 8730
rect 12200 8676 12256 8678
rect 12280 8676 12336 8678
rect 12360 8676 12416 8678
rect 12440 8676 12496 8678
rect 12200 7642 12256 7644
rect 12280 7642 12336 7644
rect 12360 7642 12416 7644
rect 12440 7642 12496 7644
rect 12200 7590 12246 7642
rect 12246 7590 12256 7642
rect 12280 7590 12310 7642
rect 12310 7590 12322 7642
rect 12322 7590 12336 7642
rect 12360 7590 12374 7642
rect 12374 7590 12386 7642
rect 12386 7590 12416 7642
rect 12440 7590 12450 7642
rect 12450 7590 12496 7642
rect 12200 7588 12256 7590
rect 12280 7588 12336 7590
rect 12360 7588 12416 7590
rect 12440 7588 12496 7590
rect 12200 6554 12256 6556
rect 12280 6554 12336 6556
rect 12360 6554 12416 6556
rect 12440 6554 12496 6556
rect 12200 6502 12246 6554
rect 12246 6502 12256 6554
rect 12280 6502 12310 6554
rect 12310 6502 12322 6554
rect 12322 6502 12336 6554
rect 12360 6502 12374 6554
rect 12374 6502 12386 6554
rect 12386 6502 12416 6554
rect 12440 6502 12450 6554
rect 12450 6502 12496 6554
rect 12200 6500 12256 6502
rect 12280 6500 12336 6502
rect 12360 6500 12416 6502
rect 12440 6500 12496 6502
rect 12200 5466 12256 5468
rect 12280 5466 12336 5468
rect 12360 5466 12416 5468
rect 12440 5466 12496 5468
rect 12200 5414 12246 5466
rect 12246 5414 12256 5466
rect 12280 5414 12310 5466
rect 12310 5414 12322 5466
rect 12322 5414 12336 5466
rect 12360 5414 12374 5466
rect 12374 5414 12386 5466
rect 12386 5414 12416 5466
rect 12440 5414 12450 5466
rect 12450 5414 12496 5466
rect 12200 5412 12256 5414
rect 12280 5412 12336 5414
rect 12360 5412 12416 5414
rect 12440 5412 12496 5414
rect 12200 4378 12256 4380
rect 12280 4378 12336 4380
rect 12360 4378 12416 4380
rect 12440 4378 12496 4380
rect 12200 4326 12246 4378
rect 12246 4326 12256 4378
rect 12280 4326 12310 4378
rect 12310 4326 12322 4378
rect 12322 4326 12336 4378
rect 12360 4326 12374 4378
rect 12374 4326 12386 4378
rect 12386 4326 12416 4378
rect 12440 4326 12450 4378
rect 12450 4326 12496 4378
rect 12200 4324 12256 4326
rect 12280 4324 12336 4326
rect 12360 4324 12416 4326
rect 12440 4324 12496 4326
rect 12200 3290 12256 3292
rect 12280 3290 12336 3292
rect 12360 3290 12416 3292
rect 12440 3290 12496 3292
rect 12200 3238 12246 3290
rect 12246 3238 12256 3290
rect 12280 3238 12310 3290
rect 12310 3238 12322 3290
rect 12322 3238 12336 3290
rect 12360 3238 12374 3290
rect 12374 3238 12386 3290
rect 12386 3238 12416 3290
rect 12440 3238 12450 3290
rect 12450 3238 12496 3290
rect 12200 3236 12256 3238
rect 12280 3236 12336 3238
rect 12360 3236 12416 3238
rect 12440 3236 12496 3238
rect 12714 7520 12770 7576
rect 12898 2896 12954 2952
rect 12714 2488 12770 2544
rect 15566 12416 15622 12472
rect 11518 2352 11574 2408
rect 12200 2202 12256 2204
rect 12280 2202 12336 2204
rect 12360 2202 12416 2204
rect 12440 2202 12496 2204
rect 12200 2150 12246 2202
rect 12246 2150 12256 2202
rect 12280 2150 12310 2202
rect 12310 2150 12322 2202
rect 12322 2150 12336 2202
rect 12360 2150 12374 2202
rect 12374 2150 12386 2202
rect 12386 2150 12416 2202
rect 12440 2150 12450 2202
rect 12450 2150 12496 2202
rect 12200 2148 12256 2150
rect 12280 2148 12336 2150
rect 12360 2148 12416 2150
rect 12440 2148 12496 2150
rect 14074 9274 14130 9276
rect 14154 9274 14210 9276
rect 14234 9274 14290 9276
rect 14314 9274 14370 9276
rect 14074 9222 14120 9274
rect 14120 9222 14130 9274
rect 14154 9222 14184 9274
rect 14184 9222 14196 9274
rect 14196 9222 14210 9274
rect 14234 9222 14248 9274
rect 14248 9222 14260 9274
rect 14260 9222 14290 9274
rect 14314 9222 14324 9274
rect 14324 9222 14370 9274
rect 14074 9220 14130 9222
rect 14154 9220 14210 9222
rect 14234 9220 14290 9222
rect 14314 9220 14370 9222
rect 14074 8186 14130 8188
rect 14154 8186 14210 8188
rect 14234 8186 14290 8188
rect 14314 8186 14370 8188
rect 14074 8134 14120 8186
rect 14120 8134 14130 8186
rect 14154 8134 14184 8186
rect 14184 8134 14196 8186
rect 14196 8134 14210 8186
rect 14234 8134 14248 8186
rect 14248 8134 14260 8186
rect 14260 8134 14290 8186
rect 14314 8134 14324 8186
rect 14324 8134 14370 8186
rect 14074 8132 14130 8134
rect 14154 8132 14210 8134
rect 14234 8132 14290 8134
rect 14314 8132 14370 8134
rect 14074 7098 14130 7100
rect 14154 7098 14210 7100
rect 14234 7098 14290 7100
rect 14314 7098 14370 7100
rect 14074 7046 14120 7098
rect 14120 7046 14130 7098
rect 14154 7046 14184 7098
rect 14184 7046 14196 7098
rect 14196 7046 14210 7098
rect 14234 7046 14248 7098
rect 14248 7046 14260 7098
rect 14260 7046 14290 7098
rect 14314 7046 14324 7098
rect 14324 7046 14370 7098
rect 14074 7044 14130 7046
rect 14154 7044 14210 7046
rect 14234 7044 14290 7046
rect 14314 7044 14370 7046
rect 14074 6010 14130 6012
rect 14154 6010 14210 6012
rect 14234 6010 14290 6012
rect 14314 6010 14370 6012
rect 14074 5958 14120 6010
rect 14120 5958 14130 6010
rect 14154 5958 14184 6010
rect 14184 5958 14196 6010
rect 14196 5958 14210 6010
rect 14234 5958 14248 6010
rect 14248 5958 14260 6010
rect 14260 5958 14290 6010
rect 14314 5958 14324 6010
rect 14324 5958 14370 6010
rect 14074 5956 14130 5958
rect 14154 5956 14210 5958
rect 14234 5956 14290 5958
rect 14314 5956 14370 5958
rect 14074 4922 14130 4924
rect 14154 4922 14210 4924
rect 14234 4922 14290 4924
rect 14314 4922 14370 4924
rect 14074 4870 14120 4922
rect 14120 4870 14130 4922
rect 14154 4870 14184 4922
rect 14184 4870 14196 4922
rect 14196 4870 14210 4922
rect 14234 4870 14248 4922
rect 14248 4870 14260 4922
rect 14260 4870 14290 4922
rect 14314 4870 14324 4922
rect 14324 4870 14370 4922
rect 14074 4868 14130 4870
rect 14154 4868 14210 4870
rect 14234 4868 14290 4870
rect 14314 4868 14370 4870
rect 14074 3834 14130 3836
rect 14154 3834 14210 3836
rect 14234 3834 14290 3836
rect 14314 3834 14370 3836
rect 14074 3782 14120 3834
rect 14120 3782 14130 3834
rect 14154 3782 14184 3834
rect 14184 3782 14196 3834
rect 14196 3782 14210 3834
rect 14234 3782 14248 3834
rect 14248 3782 14260 3834
rect 14260 3782 14290 3834
rect 14314 3782 14324 3834
rect 14324 3782 14370 3834
rect 14074 3780 14130 3782
rect 14154 3780 14210 3782
rect 14234 3780 14290 3782
rect 14314 3780 14370 3782
rect 14074 2746 14130 2748
rect 14154 2746 14210 2748
rect 14234 2746 14290 2748
rect 14314 2746 14370 2748
rect 14074 2694 14120 2746
rect 14120 2694 14130 2746
rect 14154 2694 14184 2746
rect 14184 2694 14196 2746
rect 14196 2694 14210 2746
rect 14234 2694 14248 2746
rect 14248 2694 14260 2746
rect 14260 2694 14290 2746
rect 14314 2694 14324 2746
rect 14324 2694 14370 2746
rect 14074 2692 14130 2694
rect 14154 2692 14210 2694
rect 14234 2692 14290 2694
rect 14314 2692 14370 2694
<< metal3 >>
rect 0 18186 800 18216
rect 1669 18186 1735 18189
rect 0 18184 1735 18186
rect 0 18128 1674 18184
rect 1730 18128 1735 18184
rect 0 18126 1735 18128
rect 0 18096 800 18126
rect 1669 18123 1735 18126
rect 4694 17440 5010 17441
rect 4694 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5010 17440
rect 4694 17375 5010 17376
rect 8442 17440 8758 17441
rect 8442 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8758 17440
rect 8442 17375 8758 17376
rect 12190 17440 12506 17441
rect 12190 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12506 17440
rect 12190 17375 12506 17376
rect 15561 17370 15627 17373
rect 16400 17370 17200 17400
rect 15561 17368 17200 17370
rect 15561 17312 15566 17368
rect 15622 17312 17200 17368
rect 15561 17310 17200 17312
rect 15561 17307 15627 17310
rect 16400 17280 17200 17310
rect 2820 16896 3136 16897
rect 2820 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3136 16896
rect 2820 16831 3136 16832
rect 6568 16896 6884 16897
rect 6568 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6884 16896
rect 6568 16831 6884 16832
rect 10316 16896 10632 16897
rect 10316 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10632 16896
rect 10316 16831 10632 16832
rect 14064 16896 14380 16897
rect 14064 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14380 16896
rect 14064 16831 14380 16832
rect 10961 16690 11027 16693
rect 12801 16690 12867 16693
rect 10961 16688 12867 16690
rect 10961 16632 10966 16688
rect 11022 16632 12806 16688
rect 12862 16632 12867 16688
rect 10961 16630 12867 16632
rect 10961 16627 11027 16630
rect 12801 16627 12867 16630
rect 4694 16352 5010 16353
rect 4694 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5010 16352
rect 4694 16287 5010 16288
rect 8442 16352 8758 16353
rect 8442 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8758 16352
rect 8442 16287 8758 16288
rect 12190 16352 12506 16353
rect 12190 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12506 16352
rect 12190 16287 12506 16288
rect 2820 15808 3136 15809
rect 2820 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3136 15808
rect 2820 15743 3136 15744
rect 6568 15808 6884 15809
rect 6568 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6884 15808
rect 6568 15743 6884 15744
rect 10316 15808 10632 15809
rect 10316 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10632 15808
rect 10316 15743 10632 15744
rect 14064 15808 14380 15809
rect 14064 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14380 15808
rect 14064 15743 14380 15744
rect 4694 15264 5010 15265
rect 4694 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5010 15264
rect 4694 15199 5010 15200
rect 8442 15264 8758 15265
rect 8442 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8758 15264
rect 8442 15199 8758 15200
rect 12190 15264 12506 15265
rect 12190 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12506 15264
rect 12190 15199 12506 15200
rect 0 14922 800 14952
rect 1485 14922 1551 14925
rect 0 14920 1551 14922
rect 0 14864 1490 14920
rect 1546 14864 1551 14920
rect 0 14862 1551 14864
rect 0 14832 800 14862
rect 1485 14859 1551 14862
rect 2820 14720 3136 14721
rect 2820 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3136 14720
rect 2820 14655 3136 14656
rect 6568 14720 6884 14721
rect 6568 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6884 14720
rect 6568 14655 6884 14656
rect 10316 14720 10632 14721
rect 10316 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10632 14720
rect 10316 14655 10632 14656
rect 14064 14720 14380 14721
rect 14064 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14380 14720
rect 14064 14655 14380 14656
rect 4694 14176 5010 14177
rect 4694 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5010 14176
rect 4694 14111 5010 14112
rect 8442 14176 8758 14177
rect 8442 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8758 14176
rect 8442 14111 8758 14112
rect 12190 14176 12506 14177
rect 12190 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12506 14176
rect 12190 14111 12506 14112
rect 2820 13632 3136 13633
rect 2820 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3136 13632
rect 2820 13567 3136 13568
rect 6568 13632 6884 13633
rect 6568 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6884 13632
rect 6568 13567 6884 13568
rect 10316 13632 10632 13633
rect 10316 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10632 13632
rect 10316 13567 10632 13568
rect 14064 13632 14380 13633
rect 14064 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14380 13632
rect 14064 13567 14380 13568
rect 4694 13088 5010 13089
rect 4694 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5010 13088
rect 4694 13023 5010 13024
rect 8442 13088 8758 13089
rect 8442 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8758 13088
rect 8442 13023 8758 13024
rect 12190 13088 12506 13089
rect 12190 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12506 13088
rect 12190 13023 12506 13024
rect 2820 12544 3136 12545
rect 2820 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3136 12544
rect 2820 12479 3136 12480
rect 6568 12544 6884 12545
rect 6568 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6884 12544
rect 6568 12479 6884 12480
rect 10316 12544 10632 12545
rect 10316 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10632 12544
rect 10316 12479 10632 12480
rect 14064 12544 14380 12545
rect 14064 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14380 12544
rect 14064 12479 14380 12480
rect 15561 12474 15627 12477
rect 16400 12474 17200 12504
rect 15561 12472 17200 12474
rect 15561 12416 15566 12472
rect 15622 12416 17200 12472
rect 15561 12414 17200 12416
rect 15561 12411 15627 12414
rect 16400 12384 17200 12414
rect 4694 12000 5010 12001
rect 4694 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5010 12000
rect 4694 11935 5010 11936
rect 8442 12000 8758 12001
rect 8442 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8758 12000
rect 8442 11935 8758 11936
rect 12190 12000 12506 12001
rect 12190 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12506 12000
rect 12190 11935 12506 11936
rect 0 11658 800 11688
rect 1393 11658 1459 11661
rect 0 11656 1459 11658
rect 0 11600 1398 11656
rect 1454 11600 1459 11656
rect 0 11598 1459 11600
rect 0 11568 800 11598
rect 1393 11595 1459 11598
rect 2820 11456 3136 11457
rect 2820 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3136 11456
rect 2820 11391 3136 11392
rect 6568 11456 6884 11457
rect 6568 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6884 11456
rect 6568 11391 6884 11392
rect 10316 11456 10632 11457
rect 10316 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10632 11456
rect 10316 11391 10632 11392
rect 14064 11456 14380 11457
rect 14064 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14380 11456
rect 14064 11391 14380 11392
rect 7741 11116 7807 11117
rect 7741 11112 7788 11116
rect 7852 11114 7858 11116
rect 8017 11114 8083 11117
rect 8150 11114 8156 11116
rect 7741 11056 7746 11112
rect 7741 11052 7788 11056
rect 7852 11054 7898 11114
rect 8017 11112 8156 11114
rect 8017 11056 8022 11112
rect 8078 11056 8156 11112
rect 8017 11054 8156 11056
rect 7852 11052 7858 11054
rect 7741 11051 7807 11052
rect 8017 11051 8083 11054
rect 8150 11052 8156 11054
rect 8220 11052 8226 11116
rect 4694 10912 5010 10913
rect 4694 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5010 10912
rect 4694 10847 5010 10848
rect 8442 10912 8758 10913
rect 8442 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8758 10912
rect 8442 10847 8758 10848
rect 12190 10912 12506 10913
rect 12190 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12506 10912
rect 12190 10847 12506 10848
rect 6821 10706 6887 10709
rect 11789 10706 11855 10709
rect 6821 10704 11855 10706
rect 6821 10648 6826 10704
rect 6882 10648 11794 10704
rect 11850 10648 11855 10704
rect 6821 10646 11855 10648
rect 6821 10643 6887 10646
rect 11789 10643 11855 10646
rect 2820 10368 3136 10369
rect 2820 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3136 10368
rect 2820 10303 3136 10304
rect 6568 10368 6884 10369
rect 6568 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6884 10368
rect 6568 10303 6884 10304
rect 10316 10368 10632 10369
rect 10316 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10632 10368
rect 10316 10303 10632 10304
rect 14064 10368 14380 10369
rect 14064 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14380 10368
rect 14064 10303 14380 10304
rect 8661 10298 8727 10301
rect 9029 10300 9095 10301
rect 8886 10298 8892 10300
rect 8661 10296 8892 10298
rect 8661 10240 8666 10296
rect 8722 10240 8892 10296
rect 8661 10238 8892 10240
rect 8661 10235 8727 10238
rect 8886 10236 8892 10238
rect 8956 10236 8962 10300
rect 9029 10296 9076 10300
rect 9140 10298 9146 10300
rect 9029 10240 9034 10296
rect 9029 10236 9076 10240
rect 9140 10238 9186 10298
rect 9140 10236 9146 10238
rect 9029 10235 9095 10236
rect 7741 10162 7807 10165
rect 13905 10162 13971 10165
rect 7741 10160 13971 10162
rect 7741 10104 7746 10160
rect 7802 10104 13910 10160
rect 13966 10104 13971 10160
rect 7741 10102 13971 10104
rect 7741 10099 7807 10102
rect 13905 10099 13971 10102
rect 8293 10026 8359 10029
rect 8293 10024 8954 10026
rect 8293 9968 8298 10024
rect 8354 9968 8954 10024
rect 8293 9966 8954 9968
rect 8293 9963 8359 9966
rect 8894 9890 8954 9966
rect 9029 9890 9095 9893
rect 8894 9888 9095 9890
rect 8894 9832 9034 9888
rect 9090 9832 9095 9888
rect 8894 9830 9095 9832
rect 9029 9827 9095 9830
rect 4694 9824 5010 9825
rect 4694 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5010 9824
rect 4694 9759 5010 9760
rect 8442 9824 8758 9825
rect 8442 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8758 9824
rect 8442 9759 8758 9760
rect 12190 9824 12506 9825
rect 12190 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12506 9824
rect 12190 9759 12506 9760
rect 6269 9754 6335 9757
rect 8845 9756 8911 9757
rect 9581 9756 9647 9757
rect 6269 9752 8218 9754
rect 6269 9696 6274 9752
rect 6330 9696 8218 9752
rect 6269 9694 8218 9696
rect 6269 9691 6335 9694
rect 8158 9618 8218 9694
rect 8845 9752 8892 9756
rect 8956 9754 8962 9756
rect 8845 9696 8850 9752
rect 8845 9692 8892 9696
rect 8956 9694 9002 9754
rect 9581 9752 9628 9756
rect 9692 9754 9698 9756
rect 9581 9696 9586 9752
rect 8956 9692 8962 9694
rect 9581 9692 9628 9696
rect 9692 9694 9738 9754
rect 9692 9692 9698 9694
rect 8845 9691 8911 9692
rect 9581 9691 9647 9692
rect 9581 9618 9647 9621
rect 10225 9618 10291 9621
rect 8158 9558 9184 9618
rect 4429 9482 4495 9485
rect 8385 9482 8451 9485
rect 4429 9480 8451 9482
rect 4429 9424 4434 9480
rect 4490 9424 8390 9480
rect 8446 9424 8451 9480
rect 4429 9422 8451 9424
rect 9124 9482 9184 9558
rect 9581 9616 10291 9618
rect 9581 9560 9586 9616
rect 9642 9560 10230 9616
rect 10286 9560 10291 9616
rect 9581 9558 10291 9560
rect 9581 9555 9647 9558
rect 10225 9555 10291 9558
rect 10225 9482 10291 9485
rect 9124 9480 10291 9482
rect 9124 9424 10230 9480
rect 10286 9424 10291 9480
rect 9124 9422 10291 9424
rect 4429 9419 4495 9422
rect 8385 9419 8451 9422
rect 10225 9419 10291 9422
rect 2820 9280 3136 9281
rect 2820 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3136 9280
rect 2820 9215 3136 9216
rect 6568 9280 6884 9281
rect 6568 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6884 9280
rect 6568 9215 6884 9216
rect 10316 9280 10632 9281
rect 10316 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10632 9280
rect 10316 9215 10632 9216
rect 14064 9280 14380 9281
rect 14064 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14380 9280
rect 14064 9215 14380 9216
rect 8937 8938 9003 8941
rect 8937 8936 9138 8938
rect 8937 8880 8942 8936
rect 8998 8880 9138 8936
rect 8937 8878 9138 8880
rect 8937 8875 9003 8878
rect 9078 8802 9138 8878
rect 9581 8802 9647 8805
rect 9078 8800 9647 8802
rect 9078 8744 9586 8800
rect 9642 8744 9647 8800
rect 9078 8742 9647 8744
rect 9581 8739 9647 8742
rect 4694 8736 5010 8737
rect 4694 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5010 8736
rect 4694 8671 5010 8672
rect 8442 8736 8758 8737
rect 8442 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8758 8736
rect 8442 8671 8758 8672
rect 12190 8736 12506 8737
rect 12190 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12506 8736
rect 12190 8671 12506 8672
rect 8845 8530 8911 8533
rect 9070 8530 9076 8532
rect 8845 8528 9076 8530
rect 8845 8472 8850 8528
rect 8906 8472 9076 8528
rect 8845 8470 9076 8472
rect 8845 8467 8911 8470
rect 9070 8468 9076 8470
rect 9140 8468 9146 8532
rect 0 8394 800 8424
rect 1485 8394 1551 8397
rect 0 8392 1551 8394
rect 0 8336 1490 8392
rect 1546 8336 1551 8392
rect 0 8334 1551 8336
rect 0 8304 800 8334
rect 1485 8331 1551 8334
rect 2820 8192 3136 8193
rect 2820 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3136 8192
rect 2820 8127 3136 8128
rect 6568 8192 6884 8193
rect 6568 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6884 8192
rect 6568 8127 6884 8128
rect 10316 8192 10632 8193
rect 10316 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10632 8192
rect 10316 8127 10632 8128
rect 14064 8192 14380 8193
rect 14064 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14380 8192
rect 14064 8127 14380 8128
rect 4694 7648 5010 7649
rect 4694 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5010 7648
rect 4694 7583 5010 7584
rect 8442 7648 8758 7649
rect 8442 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8758 7648
rect 8442 7583 8758 7584
rect 12190 7648 12506 7649
rect 12190 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12506 7648
rect 12190 7583 12506 7584
rect 12709 7578 12775 7581
rect 16400 7578 17200 7608
rect 12709 7576 17200 7578
rect 12709 7520 12714 7576
rect 12770 7520 17200 7576
rect 12709 7518 17200 7520
rect 12709 7515 12775 7518
rect 16400 7488 17200 7518
rect 2820 7104 3136 7105
rect 2820 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3136 7104
rect 2820 7039 3136 7040
rect 6568 7104 6884 7105
rect 6568 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6884 7104
rect 6568 7039 6884 7040
rect 10316 7104 10632 7105
rect 10316 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10632 7104
rect 10316 7039 10632 7040
rect 14064 7104 14380 7105
rect 14064 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14380 7104
rect 14064 7039 14380 7040
rect 4694 6560 5010 6561
rect 4694 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5010 6560
rect 4694 6495 5010 6496
rect 8442 6560 8758 6561
rect 8442 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8758 6560
rect 8442 6495 8758 6496
rect 12190 6560 12506 6561
rect 12190 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12506 6560
rect 12190 6495 12506 6496
rect 2820 6016 3136 6017
rect 2820 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3136 6016
rect 2820 5951 3136 5952
rect 6568 6016 6884 6017
rect 6568 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6884 6016
rect 6568 5951 6884 5952
rect 10316 6016 10632 6017
rect 10316 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10632 6016
rect 10316 5951 10632 5952
rect 14064 6016 14380 6017
rect 14064 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14380 6016
rect 14064 5951 14380 5952
rect 4694 5472 5010 5473
rect 4694 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5010 5472
rect 4694 5407 5010 5408
rect 8442 5472 8758 5473
rect 8442 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8758 5472
rect 8442 5407 8758 5408
rect 12190 5472 12506 5473
rect 12190 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12506 5472
rect 12190 5407 12506 5408
rect 0 5130 800 5160
rect 1485 5130 1551 5133
rect 0 5128 1551 5130
rect 0 5072 1490 5128
rect 1546 5072 1551 5128
rect 0 5070 1551 5072
rect 0 5040 800 5070
rect 1485 5067 1551 5070
rect 2820 4928 3136 4929
rect 2820 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3136 4928
rect 2820 4863 3136 4864
rect 6568 4928 6884 4929
rect 6568 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6884 4928
rect 6568 4863 6884 4864
rect 10316 4928 10632 4929
rect 10316 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10632 4928
rect 10316 4863 10632 4864
rect 14064 4928 14380 4929
rect 14064 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14380 4928
rect 14064 4863 14380 4864
rect 4694 4384 5010 4385
rect 4694 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5010 4384
rect 4694 4319 5010 4320
rect 8442 4384 8758 4385
rect 8442 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8758 4384
rect 8442 4319 8758 4320
rect 12190 4384 12506 4385
rect 12190 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12506 4384
rect 12190 4319 12506 4320
rect 2820 3840 3136 3841
rect 2820 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3136 3840
rect 2820 3775 3136 3776
rect 6568 3840 6884 3841
rect 6568 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6884 3840
rect 6568 3775 6884 3776
rect 10316 3840 10632 3841
rect 10316 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10632 3840
rect 10316 3775 10632 3776
rect 14064 3840 14380 3841
rect 14064 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14380 3840
rect 14064 3775 14380 3776
rect 4694 3296 5010 3297
rect 4694 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5010 3296
rect 4694 3231 5010 3232
rect 8442 3296 8758 3297
rect 8442 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8758 3296
rect 8442 3231 8758 3232
rect 12190 3296 12506 3297
rect 12190 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12506 3296
rect 12190 3231 12506 3232
rect 9622 2892 9628 2956
rect 9692 2954 9698 2956
rect 12893 2954 12959 2957
rect 9692 2952 12959 2954
rect 9692 2896 12898 2952
rect 12954 2896 12959 2952
rect 9692 2894 12959 2896
rect 9692 2892 9698 2894
rect 12893 2891 12959 2894
rect 2820 2752 3136 2753
rect 2820 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3136 2752
rect 2820 2687 3136 2688
rect 6568 2752 6884 2753
rect 6568 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6884 2752
rect 6568 2687 6884 2688
rect 10316 2752 10632 2753
rect 10316 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10632 2752
rect 10316 2687 10632 2688
rect 14064 2752 14380 2753
rect 14064 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14380 2752
rect 14064 2687 14380 2688
rect 8150 2620 8156 2684
rect 8220 2682 8226 2684
rect 16400 2682 17200 2712
rect 8220 2622 10242 2682
rect 8220 2620 8226 2622
rect 5441 2546 5507 2549
rect 9949 2546 10015 2549
rect 5441 2544 10015 2546
rect 5441 2488 5446 2544
rect 5502 2488 9954 2544
rect 10010 2488 10015 2544
rect 5441 2486 10015 2488
rect 10182 2546 10242 2622
rect 14598 2622 17200 2682
rect 11513 2546 11579 2549
rect 10182 2544 11579 2546
rect 10182 2488 11518 2544
rect 11574 2488 11579 2544
rect 10182 2486 11579 2488
rect 5441 2483 5507 2486
rect 9949 2483 10015 2486
rect 11513 2483 11579 2486
rect 12709 2546 12775 2549
rect 14598 2546 14658 2622
rect 16400 2592 17200 2622
rect 12709 2544 14658 2546
rect 12709 2488 12714 2544
rect 12770 2488 14658 2544
rect 12709 2486 14658 2488
rect 12709 2483 12775 2486
rect 7782 2348 7788 2412
rect 7852 2410 7858 2412
rect 11513 2410 11579 2413
rect 7852 2408 11579 2410
rect 7852 2352 11518 2408
rect 11574 2352 11579 2408
rect 7852 2350 11579 2352
rect 7852 2348 7858 2350
rect 11513 2347 11579 2350
rect 4694 2208 5010 2209
rect 4694 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5010 2208
rect 4694 2143 5010 2144
rect 8442 2208 8758 2209
rect 8442 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8758 2208
rect 8442 2143 8758 2144
rect 12190 2208 12506 2209
rect 12190 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12506 2208
rect 12190 2143 12506 2144
rect 0 1866 800 1896
rect 1853 1866 1919 1869
rect 0 1864 1919 1866
rect 0 1808 1858 1864
rect 1914 1808 1919 1864
rect 0 1806 1919 1808
rect 0 1776 800 1806
rect 1853 1803 1919 1806
<< via3 >>
rect 4700 17436 4764 17440
rect 4700 17380 4704 17436
rect 4704 17380 4760 17436
rect 4760 17380 4764 17436
rect 4700 17376 4764 17380
rect 4780 17436 4844 17440
rect 4780 17380 4784 17436
rect 4784 17380 4840 17436
rect 4840 17380 4844 17436
rect 4780 17376 4844 17380
rect 4860 17436 4924 17440
rect 4860 17380 4864 17436
rect 4864 17380 4920 17436
rect 4920 17380 4924 17436
rect 4860 17376 4924 17380
rect 4940 17436 5004 17440
rect 4940 17380 4944 17436
rect 4944 17380 5000 17436
rect 5000 17380 5004 17436
rect 4940 17376 5004 17380
rect 8448 17436 8512 17440
rect 8448 17380 8452 17436
rect 8452 17380 8508 17436
rect 8508 17380 8512 17436
rect 8448 17376 8512 17380
rect 8528 17436 8592 17440
rect 8528 17380 8532 17436
rect 8532 17380 8588 17436
rect 8588 17380 8592 17436
rect 8528 17376 8592 17380
rect 8608 17436 8672 17440
rect 8608 17380 8612 17436
rect 8612 17380 8668 17436
rect 8668 17380 8672 17436
rect 8608 17376 8672 17380
rect 8688 17436 8752 17440
rect 8688 17380 8692 17436
rect 8692 17380 8748 17436
rect 8748 17380 8752 17436
rect 8688 17376 8752 17380
rect 12196 17436 12260 17440
rect 12196 17380 12200 17436
rect 12200 17380 12256 17436
rect 12256 17380 12260 17436
rect 12196 17376 12260 17380
rect 12276 17436 12340 17440
rect 12276 17380 12280 17436
rect 12280 17380 12336 17436
rect 12336 17380 12340 17436
rect 12276 17376 12340 17380
rect 12356 17436 12420 17440
rect 12356 17380 12360 17436
rect 12360 17380 12416 17436
rect 12416 17380 12420 17436
rect 12356 17376 12420 17380
rect 12436 17436 12500 17440
rect 12436 17380 12440 17436
rect 12440 17380 12496 17436
rect 12496 17380 12500 17436
rect 12436 17376 12500 17380
rect 2826 16892 2890 16896
rect 2826 16836 2830 16892
rect 2830 16836 2886 16892
rect 2886 16836 2890 16892
rect 2826 16832 2890 16836
rect 2906 16892 2970 16896
rect 2906 16836 2910 16892
rect 2910 16836 2966 16892
rect 2966 16836 2970 16892
rect 2906 16832 2970 16836
rect 2986 16892 3050 16896
rect 2986 16836 2990 16892
rect 2990 16836 3046 16892
rect 3046 16836 3050 16892
rect 2986 16832 3050 16836
rect 3066 16892 3130 16896
rect 3066 16836 3070 16892
rect 3070 16836 3126 16892
rect 3126 16836 3130 16892
rect 3066 16832 3130 16836
rect 6574 16892 6638 16896
rect 6574 16836 6578 16892
rect 6578 16836 6634 16892
rect 6634 16836 6638 16892
rect 6574 16832 6638 16836
rect 6654 16892 6718 16896
rect 6654 16836 6658 16892
rect 6658 16836 6714 16892
rect 6714 16836 6718 16892
rect 6654 16832 6718 16836
rect 6734 16892 6798 16896
rect 6734 16836 6738 16892
rect 6738 16836 6794 16892
rect 6794 16836 6798 16892
rect 6734 16832 6798 16836
rect 6814 16892 6878 16896
rect 6814 16836 6818 16892
rect 6818 16836 6874 16892
rect 6874 16836 6878 16892
rect 6814 16832 6878 16836
rect 10322 16892 10386 16896
rect 10322 16836 10326 16892
rect 10326 16836 10382 16892
rect 10382 16836 10386 16892
rect 10322 16832 10386 16836
rect 10402 16892 10466 16896
rect 10402 16836 10406 16892
rect 10406 16836 10462 16892
rect 10462 16836 10466 16892
rect 10402 16832 10466 16836
rect 10482 16892 10546 16896
rect 10482 16836 10486 16892
rect 10486 16836 10542 16892
rect 10542 16836 10546 16892
rect 10482 16832 10546 16836
rect 10562 16892 10626 16896
rect 10562 16836 10566 16892
rect 10566 16836 10622 16892
rect 10622 16836 10626 16892
rect 10562 16832 10626 16836
rect 14070 16892 14134 16896
rect 14070 16836 14074 16892
rect 14074 16836 14130 16892
rect 14130 16836 14134 16892
rect 14070 16832 14134 16836
rect 14150 16892 14214 16896
rect 14150 16836 14154 16892
rect 14154 16836 14210 16892
rect 14210 16836 14214 16892
rect 14150 16832 14214 16836
rect 14230 16892 14294 16896
rect 14230 16836 14234 16892
rect 14234 16836 14290 16892
rect 14290 16836 14294 16892
rect 14230 16832 14294 16836
rect 14310 16892 14374 16896
rect 14310 16836 14314 16892
rect 14314 16836 14370 16892
rect 14370 16836 14374 16892
rect 14310 16832 14374 16836
rect 4700 16348 4764 16352
rect 4700 16292 4704 16348
rect 4704 16292 4760 16348
rect 4760 16292 4764 16348
rect 4700 16288 4764 16292
rect 4780 16348 4844 16352
rect 4780 16292 4784 16348
rect 4784 16292 4840 16348
rect 4840 16292 4844 16348
rect 4780 16288 4844 16292
rect 4860 16348 4924 16352
rect 4860 16292 4864 16348
rect 4864 16292 4920 16348
rect 4920 16292 4924 16348
rect 4860 16288 4924 16292
rect 4940 16348 5004 16352
rect 4940 16292 4944 16348
rect 4944 16292 5000 16348
rect 5000 16292 5004 16348
rect 4940 16288 5004 16292
rect 8448 16348 8512 16352
rect 8448 16292 8452 16348
rect 8452 16292 8508 16348
rect 8508 16292 8512 16348
rect 8448 16288 8512 16292
rect 8528 16348 8592 16352
rect 8528 16292 8532 16348
rect 8532 16292 8588 16348
rect 8588 16292 8592 16348
rect 8528 16288 8592 16292
rect 8608 16348 8672 16352
rect 8608 16292 8612 16348
rect 8612 16292 8668 16348
rect 8668 16292 8672 16348
rect 8608 16288 8672 16292
rect 8688 16348 8752 16352
rect 8688 16292 8692 16348
rect 8692 16292 8748 16348
rect 8748 16292 8752 16348
rect 8688 16288 8752 16292
rect 12196 16348 12260 16352
rect 12196 16292 12200 16348
rect 12200 16292 12256 16348
rect 12256 16292 12260 16348
rect 12196 16288 12260 16292
rect 12276 16348 12340 16352
rect 12276 16292 12280 16348
rect 12280 16292 12336 16348
rect 12336 16292 12340 16348
rect 12276 16288 12340 16292
rect 12356 16348 12420 16352
rect 12356 16292 12360 16348
rect 12360 16292 12416 16348
rect 12416 16292 12420 16348
rect 12356 16288 12420 16292
rect 12436 16348 12500 16352
rect 12436 16292 12440 16348
rect 12440 16292 12496 16348
rect 12496 16292 12500 16348
rect 12436 16288 12500 16292
rect 2826 15804 2890 15808
rect 2826 15748 2830 15804
rect 2830 15748 2886 15804
rect 2886 15748 2890 15804
rect 2826 15744 2890 15748
rect 2906 15804 2970 15808
rect 2906 15748 2910 15804
rect 2910 15748 2966 15804
rect 2966 15748 2970 15804
rect 2906 15744 2970 15748
rect 2986 15804 3050 15808
rect 2986 15748 2990 15804
rect 2990 15748 3046 15804
rect 3046 15748 3050 15804
rect 2986 15744 3050 15748
rect 3066 15804 3130 15808
rect 3066 15748 3070 15804
rect 3070 15748 3126 15804
rect 3126 15748 3130 15804
rect 3066 15744 3130 15748
rect 6574 15804 6638 15808
rect 6574 15748 6578 15804
rect 6578 15748 6634 15804
rect 6634 15748 6638 15804
rect 6574 15744 6638 15748
rect 6654 15804 6718 15808
rect 6654 15748 6658 15804
rect 6658 15748 6714 15804
rect 6714 15748 6718 15804
rect 6654 15744 6718 15748
rect 6734 15804 6798 15808
rect 6734 15748 6738 15804
rect 6738 15748 6794 15804
rect 6794 15748 6798 15804
rect 6734 15744 6798 15748
rect 6814 15804 6878 15808
rect 6814 15748 6818 15804
rect 6818 15748 6874 15804
rect 6874 15748 6878 15804
rect 6814 15744 6878 15748
rect 10322 15804 10386 15808
rect 10322 15748 10326 15804
rect 10326 15748 10382 15804
rect 10382 15748 10386 15804
rect 10322 15744 10386 15748
rect 10402 15804 10466 15808
rect 10402 15748 10406 15804
rect 10406 15748 10462 15804
rect 10462 15748 10466 15804
rect 10402 15744 10466 15748
rect 10482 15804 10546 15808
rect 10482 15748 10486 15804
rect 10486 15748 10542 15804
rect 10542 15748 10546 15804
rect 10482 15744 10546 15748
rect 10562 15804 10626 15808
rect 10562 15748 10566 15804
rect 10566 15748 10622 15804
rect 10622 15748 10626 15804
rect 10562 15744 10626 15748
rect 14070 15804 14134 15808
rect 14070 15748 14074 15804
rect 14074 15748 14130 15804
rect 14130 15748 14134 15804
rect 14070 15744 14134 15748
rect 14150 15804 14214 15808
rect 14150 15748 14154 15804
rect 14154 15748 14210 15804
rect 14210 15748 14214 15804
rect 14150 15744 14214 15748
rect 14230 15804 14294 15808
rect 14230 15748 14234 15804
rect 14234 15748 14290 15804
rect 14290 15748 14294 15804
rect 14230 15744 14294 15748
rect 14310 15804 14374 15808
rect 14310 15748 14314 15804
rect 14314 15748 14370 15804
rect 14370 15748 14374 15804
rect 14310 15744 14374 15748
rect 4700 15260 4764 15264
rect 4700 15204 4704 15260
rect 4704 15204 4760 15260
rect 4760 15204 4764 15260
rect 4700 15200 4764 15204
rect 4780 15260 4844 15264
rect 4780 15204 4784 15260
rect 4784 15204 4840 15260
rect 4840 15204 4844 15260
rect 4780 15200 4844 15204
rect 4860 15260 4924 15264
rect 4860 15204 4864 15260
rect 4864 15204 4920 15260
rect 4920 15204 4924 15260
rect 4860 15200 4924 15204
rect 4940 15260 5004 15264
rect 4940 15204 4944 15260
rect 4944 15204 5000 15260
rect 5000 15204 5004 15260
rect 4940 15200 5004 15204
rect 8448 15260 8512 15264
rect 8448 15204 8452 15260
rect 8452 15204 8508 15260
rect 8508 15204 8512 15260
rect 8448 15200 8512 15204
rect 8528 15260 8592 15264
rect 8528 15204 8532 15260
rect 8532 15204 8588 15260
rect 8588 15204 8592 15260
rect 8528 15200 8592 15204
rect 8608 15260 8672 15264
rect 8608 15204 8612 15260
rect 8612 15204 8668 15260
rect 8668 15204 8672 15260
rect 8608 15200 8672 15204
rect 8688 15260 8752 15264
rect 8688 15204 8692 15260
rect 8692 15204 8748 15260
rect 8748 15204 8752 15260
rect 8688 15200 8752 15204
rect 12196 15260 12260 15264
rect 12196 15204 12200 15260
rect 12200 15204 12256 15260
rect 12256 15204 12260 15260
rect 12196 15200 12260 15204
rect 12276 15260 12340 15264
rect 12276 15204 12280 15260
rect 12280 15204 12336 15260
rect 12336 15204 12340 15260
rect 12276 15200 12340 15204
rect 12356 15260 12420 15264
rect 12356 15204 12360 15260
rect 12360 15204 12416 15260
rect 12416 15204 12420 15260
rect 12356 15200 12420 15204
rect 12436 15260 12500 15264
rect 12436 15204 12440 15260
rect 12440 15204 12496 15260
rect 12496 15204 12500 15260
rect 12436 15200 12500 15204
rect 2826 14716 2890 14720
rect 2826 14660 2830 14716
rect 2830 14660 2886 14716
rect 2886 14660 2890 14716
rect 2826 14656 2890 14660
rect 2906 14716 2970 14720
rect 2906 14660 2910 14716
rect 2910 14660 2966 14716
rect 2966 14660 2970 14716
rect 2906 14656 2970 14660
rect 2986 14716 3050 14720
rect 2986 14660 2990 14716
rect 2990 14660 3046 14716
rect 3046 14660 3050 14716
rect 2986 14656 3050 14660
rect 3066 14716 3130 14720
rect 3066 14660 3070 14716
rect 3070 14660 3126 14716
rect 3126 14660 3130 14716
rect 3066 14656 3130 14660
rect 6574 14716 6638 14720
rect 6574 14660 6578 14716
rect 6578 14660 6634 14716
rect 6634 14660 6638 14716
rect 6574 14656 6638 14660
rect 6654 14716 6718 14720
rect 6654 14660 6658 14716
rect 6658 14660 6714 14716
rect 6714 14660 6718 14716
rect 6654 14656 6718 14660
rect 6734 14716 6798 14720
rect 6734 14660 6738 14716
rect 6738 14660 6794 14716
rect 6794 14660 6798 14716
rect 6734 14656 6798 14660
rect 6814 14716 6878 14720
rect 6814 14660 6818 14716
rect 6818 14660 6874 14716
rect 6874 14660 6878 14716
rect 6814 14656 6878 14660
rect 10322 14716 10386 14720
rect 10322 14660 10326 14716
rect 10326 14660 10382 14716
rect 10382 14660 10386 14716
rect 10322 14656 10386 14660
rect 10402 14716 10466 14720
rect 10402 14660 10406 14716
rect 10406 14660 10462 14716
rect 10462 14660 10466 14716
rect 10402 14656 10466 14660
rect 10482 14716 10546 14720
rect 10482 14660 10486 14716
rect 10486 14660 10542 14716
rect 10542 14660 10546 14716
rect 10482 14656 10546 14660
rect 10562 14716 10626 14720
rect 10562 14660 10566 14716
rect 10566 14660 10622 14716
rect 10622 14660 10626 14716
rect 10562 14656 10626 14660
rect 14070 14716 14134 14720
rect 14070 14660 14074 14716
rect 14074 14660 14130 14716
rect 14130 14660 14134 14716
rect 14070 14656 14134 14660
rect 14150 14716 14214 14720
rect 14150 14660 14154 14716
rect 14154 14660 14210 14716
rect 14210 14660 14214 14716
rect 14150 14656 14214 14660
rect 14230 14716 14294 14720
rect 14230 14660 14234 14716
rect 14234 14660 14290 14716
rect 14290 14660 14294 14716
rect 14230 14656 14294 14660
rect 14310 14716 14374 14720
rect 14310 14660 14314 14716
rect 14314 14660 14370 14716
rect 14370 14660 14374 14716
rect 14310 14656 14374 14660
rect 4700 14172 4764 14176
rect 4700 14116 4704 14172
rect 4704 14116 4760 14172
rect 4760 14116 4764 14172
rect 4700 14112 4764 14116
rect 4780 14172 4844 14176
rect 4780 14116 4784 14172
rect 4784 14116 4840 14172
rect 4840 14116 4844 14172
rect 4780 14112 4844 14116
rect 4860 14172 4924 14176
rect 4860 14116 4864 14172
rect 4864 14116 4920 14172
rect 4920 14116 4924 14172
rect 4860 14112 4924 14116
rect 4940 14172 5004 14176
rect 4940 14116 4944 14172
rect 4944 14116 5000 14172
rect 5000 14116 5004 14172
rect 4940 14112 5004 14116
rect 8448 14172 8512 14176
rect 8448 14116 8452 14172
rect 8452 14116 8508 14172
rect 8508 14116 8512 14172
rect 8448 14112 8512 14116
rect 8528 14172 8592 14176
rect 8528 14116 8532 14172
rect 8532 14116 8588 14172
rect 8588 14116 8592 14172
rect 8528 14112 8592 14116
rect 8608 14172 8672 14176
rect 8608 14116 8612 14172
rect 8612 14116 8668 14172
rect 8668 14116 8672 14172
rect 8608 14112 8672 14116
rect 8688 14172 8752 14176
rect 8688 14116 8692 14172
rect 8692 14116 8748 14172
rect 8748 14116 8752 14172
rect 8688 14112 8752 14116
rect 12196 14172 12260 14176
rect 12196 14116 12200 14172
rect 12200 14116 12256 14172
rect 12256 14116 12260 14172
rect 12196 14112 12260 14116
rect 12276 14172 12340 14176
rect 12276 14116 12280 14172
rect 12280 14116 12336 14172
rect 12336 14116 12340 14172
rect 12276 14112 12340 14116
rect 12356 14172 12420 14176
rect 12356 14116 12360 14172
rect 12360 14116 12416 14172
rect 12416 14116 12420 14172
rect 12356 14112 12420 14116
rect 12436 14172 12500 14176
rect 12436 14116 12440 14172
rect 12440 14116 12496 14172
rect 12496 14116 12500 14172
rect 12436 14112 12500 14116
rect 2826 13628 2890 13632
rect 2826 13572 2830 13628
rect 2830 13572 2886 13628
rect 2886 13572 2890 13628
rect 2826 13568 2890 13572
rect 2906 13628 2970 13632
rect 2906 13572 2910 13628
rect 2910 13572 2966 13628
rect 2966 13572 2970 13628
rect 2906 13568 2970 13572
rect 2986 13628 3050 13632
rect 2986 13572 2990 13628
rect 2990 13572 3046 13628
rect 3046 13572 3050 13628
rect 2986 13568 3050 13572
rect 3066 13628 3130 13632
rect 3066 13572 3070 13628
rect 3070 13572 3126 13628
rect 3126 13572 3130 13628
rect 3066 13568 3130 13572
rect 6574 13628 6638 13632
rect 6574 13572 6578 13628
rect 6578 13572 6634 13628
rect 6634 13572 6638 13628
rect 6574 13568 6638 13572
rect 6654 13628 6718 13632
rect 6654 13572 6658 13628
rect 6658 13572 6714 13628
rect 6714 13572 6718 13628
rect 6654 13568 6718 13572
rect 6734 13628 6798 13632
rect 6734 13572 6738 13628
rect 6738 13572 6794 13628
rect 6794 13572 6798 13628
rect 6734 13568 6798 13572
rect 6814 13628 6878 13632
rect 6814 13572 6818 13628
rect 6818 13572 6874 13628
rect 6874 13572 6878 13628
rect 6814 13568 6878 13572
rect 10322 13628 10386 13632
rect 10322 13572 10326 13628
rect 10326 13572 10382 13628
rect 10382 13572 10386 13628
rect 10322 13568 10386 13572
rect 10402 13628 10466 13632
rect 10402 13572 10406 13628
rect 10406 13572 10462 13628
rect 10462 13572 10466 13628
rect 10402 13568 10466 13572
rect 10482 13628 10546 13632
rect 10482 13572 10486 13628
rect 10486 13572 10542 13628
rect 10542 13572 10546 13628
rect 10482 13568 10546 13572
rect 10562 13628 10626 13632
rect 10562 13572 10566 13628
rect 10566 13572 10622 13628
rect 10622 13572 10626 13628
rect 10562 13568 10626 13572
rect 14070 13628 14134 13632
rect 14070 13572 14074 13628
rect 14074 13572 14130 13628
rect 14130 13572 14134 13628
rect 14070 13568 14134 13572
rect 14150 13628 14214 13632
rect 14150 13572 14154 13628
rect 14154 13572 14210 13628
rect 14210 13572 14214 13628
rect 14150 13568 14214 13572
rect 14230 13628 14294 13632
rect 14230 13572 14234 13628
rect 14234 13572 14290 13628
rect 14290 13572 14294 13628
rect 14230 13568 14294 13572
rect 14310 13628 14374 13632
rect 14310 13572 14314 13628
rect 14314 13572 14370 13628
rect 14370 13572 14374 13628
rect 14310 13568 14374 13572
rect 4700 13084 4764 13088
rect 4700 13028 4704 13084
rect 4704 13028 4760 13084
rect 4760 13028 4764 13084
rect 4700 13024 4764 13028
rect 4780 13084 4844 13088
rect 4780 13028 4784 13084
rect 4784 13028 4840 13084
rect 4840 13028 4844 13084
rect 4780 13024 4844 13028
rect 4860 13084 4924 13088
rect 4860 13028 4864 13084
rect 4864 13028 4920 13084
rect 4920 13028 4924 13084
rect 4860 13024 4924 13028
rect 4940 13084 5004 13088
rect 4940 13028 4944 13084
rect 4944 13028 5000 13084
rect 5000 13028 5004 13084
rect 4940 13024 5004 13028
rect 8448 13084 8512 13088
rect 8448 13028 8452 13084
rect 8452 13028 8508 13084
rect 8508 13028 8512 13084
rect 8448 13024 8512 13028
rect 8528 13084 8592 13088
rect 8528 13028 8532 13084
rect 8532 13028 8588 13084
rect 8588 13028 8592 13084
rect 8528 13024 8592 13028
rect 8608 13084 8672 13088
rect 8608 13028 8612 13084
rect 8612 13028 8668 13084
rect 8668 13028 8672 13084
rect 8608 13024 8672 13028
rect 8688 13084 8752 13088
rect 8688 13028 8692 13084
rect 8692 13028 8748 13084
rect 8748 13028 8752 13084
rect 8688 13024 8752 13028
rect 12196 13084 12260 13088
rect 12196 13028 12200 13084
rect 12200 13028 12256 13084
rect 12256 13028 12260 13084
rect 12196 13024 12260 13028
rect 12276 13084 12340 13088
rect 12276 13028 12280 13084
rect 12280 13028 12336 13084
rect 12336 13028 12340 13084
rect 12276 13024 12340 13028
rect 12356 13084 12420 13088
rect 12356 13028 12360 13084
rect 12360 13028 12416 13084
rect 12416 13028 12420 13084
rect 12356 13024 12420 13028
rect 12436 13084 12500 13088
rect 12436 13028 12440 13084
rect 12440 13028 12496 13084
rect 12496 13028 12500 13084
rect 12436 13024 12500 13028
rect 2826 12540 2890 12544
rect 2826 12484 2830 12540
rect 2830 12484 2886 12540
rect 2886 12484 2890 12540
rect 2826 12480 2890 12484
rect 2906 12540 2970 12544
rect 2906 12484 2910 12540
rect 2910 12484 2966 12540
rect 2966 12484 2970 12540
rect 2906 12480 2970 12484
rect 2986 12540 3050 12544
rect 2986 12484 2990 12540
rect 2990 12484 3046 12540
rect 3046 12484 3050 12540
rect 2986 12480 3050 12484
rect 3066 12540 3130 12544
rect 3066 12484 3070 12540
rect 3070 12484 3126 12540
rect 3126 12484 3130 12540
rect 3066 12480 3130 12484
rect 6574 12540 6638 12544
rect 6574 12484 6578 12540
rect 6578 12484 6634 12540
rect 6634 12484 6638 12540
rect 6574 12480 6638 12484
rect 6654 12540 6718 12544
rect 6654 12484 6658 12540
rect 6658 12484 6714 12540
rect 6714 12484 6718 12540
rect 6654 12480 6718 12484
rect 6734 12540 6798 12544
rect 6734 12484 6738 12540
rect 6738 12484 6794 12540
rect 6794 12484 6798 12540
rect 6734 12480 6798 12484
rect 6814 12540 6878 12544
rect 6814 12484 6818 12540
rect 6818 12484 6874 12540
rect 6874 12484 6878 12540
rect 6814 12480 6878 12484
rect 10322 12540 10386 12544
rect 10322 12484 10326 12540
rect 10326 12484 10382 12540
rect 10382 12484 10386 12540
rect 10322 12480 10386 12484
rect 10402 12540 10466 12544
rect 10402 12484 10406 12540
rect 10406 12484 10462 12540
rect 10462 12484 10466 12540
rect 10402 12480 10466 12484
rect 10482 12540 10546 12544
rect 10482 12484 10486 12540
rect 10486 12484 10542 12540
rect 10542 12484 10546 12540
rect 10482 12480 10546 12484
rect 10562 12540 10626 12544
rect 10562 12484 10566 12540
rect 10566 12484 10622 12540
rect 10622 12484 10626 12540
rect 10562 12480 10626 12484
rect 14070 12540 14134 12544
rect 14070 12484 14074 12540
rect 14074 12484 14130 12540
rect 14130 12484 14134 12540
rect 14070 12480 14134 12484
rect 14150 12540 14214 12544
rect 14150 12484 14154 12540
rect 14154 12484 14210 12540
rect 14210 12484 14214 12540
rect 14150 12480 14214 12484
rect 14230 12540 14294 12544
rect 14230 12484 14234 12540
rect 14234 12484 14290 12540
rect 14290 12484 14294 12540
rect 14230 12480 14294 12484
rect 14310 12540 14374 12544
rect 14310 12484 14314 12540
rect 14314 12484 14370 12540
rect 14370 12484 14374 12540
rect 14310 12480 14374 12484
rect 4700 11996 4764 12000
rect 4700 11940 4704 11996
rect 4704 11940 4760 11996
rect 4760 11940 4764 11996
rect 4700 11936 4764 11940
rect 4780 11996 4844 12000
rect 4780 11940 4784 11996
rect 4784 11940 4840 11996
rect 4840 11940 4844 11996
rect 4780 11936 4844 11940
rect 4860 11996 4924 12000
rect 4860 11940 4864 11996
rect 4864 11940 4920 11996
rect 4920 11940 4924 11996
rect 4860 11936 4924 11940
rect 4940 11996 5004 12000
rect 4940 11940 4944 11996
rect 4944 11940 5000 11996
rect 5000 11940 5004 11996
rect 4940 11936 5004 11940
rect 8448 11996 8512 12000
rect 8448 11940 8452 11996
rect 8452 11940 8508 11996
rect 8508 11940 8512 11996
rect 8448 11936 8512 11940
rect 8528 11996 8592 12000
rect 8528 11940 8532 11996
rect 8532 11940 8588 11996
rect 8588 11940 8592 11996
rect 8528 11936 8592 11940
rect 8608 11996 8672 12000
rect 8608 11940 8612 11996
rect 8612 11940 8668 11996
rect 8668 11940 8672 11996
rect 8608 11936 8672 11940
rect 8688 11996 8752 12000
rect 8688 11940 8692 11996
rect 8692 11940 8748 11996
rect 8748 11940 8752 11996
rect 8688 11936 8752 11940
rect 12196 11996 12260 12000
rect 12196 11940 12200 11996
rect 12200 11940 12256 11996
rect 12256 11940 12260 11996
rect 12196 11936 12260 11940
rect 12276 11996 12340 12000
rect 12276 11940 12280 11996
rect 12280 11940 12336 11996
rect 12336 11940 12340 11996
rect 12276 11936 12340 11940
rect 12356 11996 12420 12000
rect 12356 11940 12360 11996
rect 12360 11940 12416 11996
rect 12416 11940 12420 11996
rect 12356 11936 12420 11940
rect 12436 11996 12500 12000
rect 12436 11940 12440 11996
rect 12440 11940 12496 11996
rect 12496 11940 12500 11996
rect 12436 11936 12500 11940
rect 2826 11452 2890 11456
rect 2826 11396 2830 11452
rect 2830 11396 2886 11452
rect 2886 11396 2890 11452
rect 2826 11392 2890 11396
rect 2906 11452 2970 11456
rect 2906 11396 2910 11452
rect 2910 11396 2966 11452
rect 2966 11396 2970 11452
rect 2906 11392 2970 11396
rect 2986 11452 3050 11456
rect 2986 11396 2990 11452
rect 2990 11396 3046 11452
rect 3046 11396 3050 11452
rect 2986 11392 3050 11396
rect 3066 11452 3130 11456
rect 3066 11396 3070 11452
rect 3070 11396 3126 11452
rect 3126 11396 3130 11452
rect 3066 11392 3130 11396
rect 6574 11452 6638 11456
rect 6574 11396 6578 11452
rect 6578 11396 6634 11452
rect 6634 11396 6638 11452
rect 6574 11392 6638 11396
rect 6654 11452 6718 11456
rect 6654 11396 6658 11452
rect 6658 11396 6714 11452
rect 6714 11396 6718 11452
rect 6654 11392 6718 11396
rect 6734 11452 6798 11456
rect 6734 11396 6738 11452
rect 6738 11396 6794 11452
rect 6794 11396 6798 11452
rect 6734 11392 6798 11396
rect 6814 11452 6878 11456
rect 6814 11396 6818 11452
rect 6818 11396 6874 11452
rect 6874 11396 6878 11452
rect 6814 11392 6878 11396
rect 10322 11452 10386 11456
rect 10322 11396 10326 11452
rect 10326 11396 10382 11452
rect 10382 11396 10386 11452
rect 10322 11392 10386 11396
rect 10402 11452 10466 11456
rect 10402 11396 10406 11452
rect 10406 11396 10462 11452
rect 10462 11396 10466 11452
rect 10402 11392 10466 11396
rect 10482 11452 10546 11456
rect 10482 11396 10486 11452
rect 10486 11396 10542 11452
rect 10542 11396 10546 11452
rect 10482 11392 10546 11396
rect 10562 11452 10626 11456
rect 10562 11396 10566 11452
rect 10566 11396 10622 11452
rect 10622 11396 10626 11452
rect 10562 11392 10626 11396
rect 14070 11452 14134 11456
rect 14070 11396 14074 11452
rect 14074 11396 14130 11452
rect 14130 11396 14134 11452
rect 14070 11392 14134 11396
rect 14150 11452 14214 11456
rect 14150 11396 14154 11452
rect 14154 11396 14210 11452
rect 14210 11396 14214 11452
rect 14150 11392 14214 11396
rect 14230 11452 14294 11456
rect 14230 11396 14234 11452
rect 14234 11396 14290 11452
rect 14290 11396 14294 11452
rect 14230 11392 14294 11396
rect 14310 11452 14374 11456
rect 14310 11396 14314 11452
rect 14314 11396 14370 11452
rect 14370 11396 14374 11452
rect 14310 11392 14374 11396
rect 7788 11112 7852 11116
rect 7788 11056 7802 11112
rect 7802 11056 7852 11112
rect 7788 11052 7852 11056
rect 8156 11052 8220 11116
rect 4700 10908 4764 10912
rect 4700 10852 4704 10908
rect 4704 10852 4760 10908
rect 4760 10852 4764 10908
rect 4700 10848 4764 10852
rect 4780 10908 4844 10912
rect 4780 10852 4784 10908
rect 4784 10852 4840 10908
rect 4840 10852 4844 10908
rect 4780 10848 4844 10852
rect 4860 10908 4924 10912
rect 4860 10852 4864 10908
rect 4864 10852 4920 10908
rect 4920 10852 4924 10908
rect 4860 10848 4924 10852
rect 4940 10908 5004 10912
rect 4940 10852 4944 10908
rect 4944 10852 5000 10908
rect 5000 10852 5004 10908
rect 4940 10848 5004 10852
rect 8448 10908 8512 10912
rect 8448 10852 8452 10908
rect 8452 10852 8508 10908
rect 8508 10852 8512 10908
rect 8448 10848 8512 10852
rect 8528 10908 8592 10912
rect 8528 10852 8532 10908
rect 8532 10852 8588 10908
rect 8588 10852 8592 10908
rect 8528 10848 8592 10852
rect 8608 10908 8672 10912
rect 8608 10852 8612 10908
rect 8612 10852 8668 10908
rect 8668 10852 8672 10908
rect 8608 10848 8672 10852
rect 8688 10908 8752 10912
rect 8688 10852 8692 10908
rect 8692 10852 8748 10908
rect 8748 10852 8752 10908
rect 8688 10848 8752 10852
rect 12196 10908 12260 10912
rect 12196 10852 12200 10908
rect 12200 10852 12256 10908
rect 12256 10852 12260 10908
rect 12196 10848 12260 10852
rect 12276 10908 12340 10912
rect 12276 10852 12280 10908
rect 12280 10852 12336 10908
rect 12336 10852 12340 10908
rect 12276 10848 12340 10852
rect 12356 10908 12420 10912
rect 12356 10852 12360 10908
rect 12360 10852 12416 10908
rect 12416 10852 12420 10908
rect 12356 10848 12420 10852
rect 12436 10908 12500 10912
rect 12436 10852 12440 10908
rect 12440 10852 12496 10908
rect 12496 10852 12500 10908
rect 12436 10848 12500 10852
rect 2826 10364 2890 10368
rect 2826 10308 2830 10364
rect 2830 10308 2886 10364
rect 2886 10308 2890 10364
rect 2826 10304 2890 10308
rect 2906 10364 2970 10368
rect 2906 10308 2910 10364
rect 2910 10308 2966 10364
rect 2966 10308 2970 10364
rect 2906 10304 2970 10308
rect 2986 10364 3050 10368
rect 2986 10308 2990 10364
rect 2990 10308 3046 10364
rect 3046 10308 3050 10364
rect 2986 10304 3050 10308
rect 3066 10364 3130 10368
rect 3066 10308 3070 10364
rect 3070 10308 3126 10364
rect 3126 10308 3130 10364
rect 3066 10304 3130 10308
rect 6574 10364 6638 10368
rect 6574 10308 6578 10364
rect 6578 10308 6634 10364
rect 6634 10308 6638 10364
rect 6574 10304 6638 10308
rect 6654 10364 6718 10368
rect 6654 10308 6658 10364
rect 6658 10308 6714 10364
rect 6714 10308 6718 10364
rect 6654 10304 6718 10308
rect 6734 10364 6798 10368
rect 6734 10308 6738 10364
rect 6738 10308 6794 10364
rect 6794 10308 6798 10364
rect 6734 10304 6798 10308
rect 6814 10364 6878 10368
rect 6814 10308 6818 10364
rect 6818 10308 6874 10364
rect 6874 10308 6878 10364
rect 6814 10304 6878 10308
rect 10322 10364 10386 10368
rect 10322 10308 10326 10364
rect 10326 10308 10382 10364
rect 10382 10308 10386 10364
rect 10322 10304 10386 10308
rect 10402 10364 10466 10368
rect 10402 10308 10406 10364
rect 10406 10308 10462 10364
rect 10462 10308 10466 10364
rect 10402 10304 10466 10308
rect 10482 10364 10546 10368
rect 10482 10308 10486 10364
rect 10486 10308 10542 10364
rect 10542 10308 10546 10364
rect 10482 10304 10546 10308
rect 10562 10364 10626 10368
rect 10562 10308 10566 10364
rect 10566 10308 10622 10364
rect 10622 10308 10626 10364
rect 10562 10304 10626 10308
rect 14070 10364 14134 10368
rect 14070 10308 14074 10364
rect 14074 10308 14130 10364
rect 14130 10308 14134 10364
rect 14070 10304 14134 10308
rect 14150 10364 14214 10368
rect 14150 10308 14154 10364
rect 14154 10308 14210 10364
rect 14210 10308 14214 10364
rect 14150 10304 14214 10308
rect 14230 10364 14294 10368
rect 14230 10308 14234 10364
rect 14234 10308 14290 10364
rect 14290 10308 14294 10364
rect 14230 10304 14294 10308
rect 14310 10364 14374 10368
rect 14310 10308 14314 10364
rect 14314 10308 14370 10364
rect 14370 10308 14374 10364
rect 14310 10304 14374 10308
rect 8892 10236 8956 10300
rect 9076 10296 9140 10300
rect 9076 10240 9090 10296
rect 9090 10240 9140 10296
rect 9076 10236 9140 10240
rect 4700 9820 4764 9824
rect 4700 9764 4704 9820
rect 4704 9764 4760 9820
rect 4760 9764 4764 9820
rect 4700 9760 4764 9764
rect 4780 9820 4844 9824
rect 4780 9764 4784 9820
rect 4784 9764 4840 9820
rect 4840 9764 4844 9820
rect 4780 9760 4844 9764
rect 4860 9820 4924 9824
rect 4860 9764 4864 9820
rect 4864 9764 4920 9820
rect 4920 9764 4924 9820
rect 4860 9760 4924 9764
rect 4940 9820 5004 9824
rect 4940 9764 4944 9820
rect 4944 9764 5000 9820
rect 5000 9764 5004 9820
rect 4940 9760 5004 9764
rect 8448 9820 8512 9824
rect 8448 9764 8452 9820
rect 8452 9764 8508 9820
rect 8508 9764 8512 9820
rect 8448 9760 8512 9764
rect 8528 9820 8592 9824
rect 8528 9764 8532 9820
rect 8532 9764 8588 9820
rect 8588 9764 8592 9820
rect 8528 9760 8592 9764
rect 8608 9820 8672 9824
rect 8608 9764 8612 9820
rect 8612 9764 8668 9820
rect 8668 9764 8672 9820
rect 8608 9760 8672 9764
rect 8688 9820 8752 9824
rect 8688 9764 8692 9820
rect 8692 9764 8748 9820
rect 8748 9764 8752 9820
rect 8688 9760 8752 9764
rect 12196 9820 12260 9824
rect 12196 9764 12200 9820
rect 12200 9764 12256 9820
rect 12256 9764 12260 9820
rect 12196 9760 12260 9764
rect 12276 9820 12340 9824
rect 12276 9764 12280 9820
rect 12280 9764 12336 9820
rect 12336 9764 12340 9820
rect 12276 9760 12340 9764
rect 12356 9820 12420 9824
rect 12356 9764 12360 9820
rect 12360 9764 12416 9820
rect 12416 9764 12420 9820
rect 12356 9760 12420 9764
rect 12436 9820 12500 9824
rect 12436 9764 12440 9820
rect 12440 9764 12496 9820
rect 12496 9764 12500 9820
rect 12436 9760 12500 9764
rect 8892 9752 8956 9756
rect 8892 9696 8906 9752
rect 8906 9696 8956 9752
rect 8892 9692 8956 9696
rect 9628 9752 9692 9756
rect 9628 9696 9642 9752
rect 9642 9696 9692 9752
rect 9628 9692 9692 9696
rect 2826 9276 2890 9280
rect 2826 9220 2830 9276
rect 2830 9220 2886 9276
rect 2886 9220 2890 9276
rect 2826 9216 2890 9220
rect 2906 9276 2970 9280
rect 2906 9220 2910 9276
rect 2910 9220 2966 9276
rect 2966 9220 2970 9276
rect 2906 9216 2970 9220
rect 2986 9276 3050 9280
rect 2986 9220 2990 9276
rect 2990 9220 3046 9276
rect 3046 9220 3050 9276
rect 2986 9216 3050 9220
rect 3066 9276 3130 9280
rect 3066 9220 3070 9276
rect 3070 9220 3126 9276
rect 3126 9220 3130 9276
rect 3066 9216 3130 9220
rect 6574 9276 6638 9280
rect 6574 9220 6578 9276
rect 6578 9220 6634 9276
rect 6634 9220 6638 9276
rect 6574 9216 6638 9220
rect 6654 9276 6718 9280
rect 6654 9220 6658 9276
rect 6658 9220 6714 9276
rect 6714 9220 6718 9276
rect 6654 9216 6718 9220
rect 6734 9276 6798 9280
rect 6734 9220 6738 9276
rect 6738 9220 6794 9276
rect 6794 9220 6798 9276
rect 6734 9216 6798 9220
rect 6814 9276 6878 9280
rect 6814 9220 6818 9276
rect 6818 9220 6874 9276
rect 6874 9220 6878 9276
rect 6814 9216 6878 9220
rect 10322 9276 10386 9280
rect 10322 9220 10326 9276
rect 10326 9220 10382 9276
rect 10382 9220 10386 9276
rect 10322 9216 10386 9220
rect 10402 9276 10466 9280
rect 10402 9220 10406 9276
rect 10406 9220 10462 9276
rect 10462 9220 10466 9276
rect 10402 9216 10466 9220
rect 10482 9276 10546 9280
rect 10482 9220 10486 9276
rect 10486 9220 10542 9276
rect 10542 9220 10546 9276
rect 10482 9216 10546 9220
rect 10562 9276 10626 9280
rect 10562 9220 10566 9276
rect 10566 9220 10622 9276
rect 10622 9220 10626 9276
rect 10562 9216 10626 9220
rect 14070 9276 14134 9280
rect 14070 9220 14074 9276
rect 14074 9220 14130 9276
rect 14130 9220 14134 9276
rect 14070 9216 14134 9220
rect 14150 9276 14214 9280
rect 14150 9220 14154 9276
rect 14154 9220 14210 9276
rect 14210 9220 14214 9276
rect 14150 9216 14214 9220
rect 14230 9276 14294 9280
rect 14230 9220 14234 9276
rect 14234 9220 14290 9276
rect 14290 9220 14294 9276
rect 14230 9216 14294 9220
rect 14310 9276 14374 9280
rect 14310 9220 14314 9276
rect 14314 9220 14370 9276
rect 14370 9220 14374 9276
rect 14310 9216 14374 9220
rect 4700 8732 4764 8736
rect 4700 8676 4704 8732
rect 4704 8676 4760 8732
rect 4760 8676 4764 8732
rect 4700 8672 4764 8676
rect 4780 8732 4844 8736
rect 4780 8676 4784 8732
rect 4784 8676 4840 8732
rect 4840 8676 4844 8732
rect 4780 8672 4844 8676
rect 4860 8732 4924 8736
rect 4860 8676 4864 8732
rect 4864 8676 4920 8732
rect 4920 8676 4924 8732
rect 4860 8672 4924 8676
rect 4940 8732 5004 8736
rect 4940 8676 4944 8732
rect 4944 8676 5000 8732
rect 5000 8676 5004 8732
rect 4940 8672 5004 8676
rect 8448 8732 8512 8736
rect 8448 8676 8452 8732
rect 8452 8676 8508 8732
rect 8508 8676 8512 8732
rect 8448 8672 8512 8676
rect 8528 8732 8592 8736
rect 8528 8676 8532 8732
rect 8532 8676 8588 8732
rect 8588 8676 8592 8732
rect 8528 8672 8592 8676
rect 8608 8732 8672 8736
rect 8608 8676 8612 8732
rect 8612 8676 8668 8732
rect 8668 8676 8672 8732
rect 8608 8672 8672 8676
rect 8688 8732 8752 8736
rect 8688 8676 8692 8732
rect 8692 8676 8748 8732
rect 8748 8676 8752 8732
rect 8688 8672 8752 8676
rect 12196 8732 12260 8736
rect 12196 8676 12200 8732
rect 12200 8676 12256 8732
rect 12256 8676 12260 8732
rect 12196 8672 12260 8676
rect 12276 8732 12340 8736
rect 12276 8676 12280 8732
rect 12280 8676 12336 8732
rect 12336 8676 12340 8732
rect 12276 8672 12340 8676
rect 12356 8732 12420 8736
rect 12356 8676 12360 8732
rect 12360 8676 12416 8732
rect 12416 8676 12420 8732
rect 12356 8672 12420 8676
rect 12436 8732 12500 8736
rect 12436 8676 12440 8732
rect 12440 8676 12496 8732
rect 12496 8676 12500 8732
rect 12436 8672 12500 8676
rect 9076 8468 9140 8532
rect 2826 8188 2890 8192
rect 2826 8132 2830 8188
rect 2830 8132 2886 8188
rect 2886 8132 2890 8188
rect 2826 8128 2890 8132
rect 2906 8188 2970 8192
rect 2906 8132 2910 8188
rect 2910 8132 2966 8188
rect 2966 8132 2970 8188
rect 2906 8128 2970 8132
rect 2986 8188 3050 8192
rect 2986 8132 2990 8188
rect 2990 8132 3046 8188
rect 3046 8132 3050 8188
rect 2986 8128 3050 8132
rect 3066 8188 3130 8192
rect 3066 8132 3070 8188
rect 3070 8132 3126 8188
rect 3126 8132 3130 8188
rect 3066 8128 3130 8132
rect 6574 8188 6638 8192
rect 6574 8132 6578 8188
rect 6578 8132 6634 8188
rect 6634 8132 6638 8188
rect 6574 8128 6638 8132
rect 6654 8188 6718 8192
rect 6654 8132 6658 8188
rect 6658 8132 6714 8188
rect 6714 8132 6718 8188
rect 6654 8128 6718 8132
rect 6734 8188 6798 8192
rect 6734 8132 6738 8188
rect 6738 8132 6794 8188
rect 6794 8132 6798 8188
rect 6734 8128 6798 8132
rect 6814 8188 6878 8192
rect 6814 8132 6818 8188
rect 6818 8132 6874 8188
rect 6874 8132 6878 8188
rect 6814 8128 6878 8132
rect 10322 8188 10386 8192
rect 10322 8132 10326 8188
rect 10326 8132 10382 8188
rect 10382 8132 10386 8188
rect 10322 8128 10386 8132
rect 10402 8188 10466 8192
rect 10402 8132 10406 8188
rect 10406 8132 10462 8188
rect 10462 8132 10466 8188
rect 10402 8128 10466 8132
rect 10482 8188 10546 8192
rect 10482 8132 10486 8188
rect 10486 8132 10542 8188
rect 10542 8132 10546 8188
rect 10482 8128 10546 8132
rect 10562 8188 10626 8192
rect 10562 8132 10566 8188
rect 10566 8132 10622 8188
rect 10622 8132 10626 8188
rect 10562 8128 10626 8132
rect 14070 8188 14134 8192
rect 14070 8132 14074 8188
rect 14074 8132 14130 8188
rect 14130 8132 14134 8188
rect 14070 8128 14134 8132
rect 14150 8188 14214 8192
rect 14150 8132 14154 8188
rect 14154 8132 14210 8188
rect 14210 8132 14214 8188
rect 14150 8128 14214 8132
rect 14230 8188 14294 8192
rect 14230 8132 14234 8188
rect 14234 8132 14290 8188
rect 14290 8132 14294 8188
rect 14230 8128 14294 8132
rect 14310 8188 14374 8192
rect 14310 8132 14314 8188
rect 14314 8132 14370 8188
rect 14370 8132 14374 8188
rect 14310 8128 14374 8132
rect 4700 7644 4764 7648
rect 4700 7588 4704 7644
rect 4704 7588 4760 7644
rect 4760 7588 4764 7644
rect 4700 7584 4764 7588
rect 4780 7644 4844 7648
rect 4780 7588 4784 7644
rect 4784 7588 4840 7644
rect 4840 7588 4844 7644
rect 4780 7584 4844 7588
rect 4860 7644 4924 7648
rect 4860 7588 4864 7644
rect 4864 7588 4920 7644
rect 4920 7588 4924 7644
rect 4860 7584 4924 7588
rect 4940 7644 5004 7648
rect 4940 7588 4944 7644
rect 4944 7588 5000 7644
rect 5000 7588 5004 7644
rect 4940 7584 5004 7588
rect 8448 7644 8512 7648
rect 8448 7588 8452 7644
rect 8452 7588 8508 7644
rect 8508 7588 8512 7644
rect 8448 7584 8512 7588
rect 8528 7644 8592 7648
rect 8528 7588 8532 7644
rect 8532 7588 8588 7644
rect 8588 7588 8592 7644
rect 8528 7584 8592 7588
rect 8608 7644 8672 7648
rect 8608 7588 8612 7644
rect 8612 7588 8668 7644
rect 8668 7588 8672 7644
rect 8608 7584 8672 7588
rect 8688 7644 8752 7648
rect 8688 7588 8692 7644
rect 8692 7588 8748 7644
rect 8748 7588 8752 7644
rect 8688 7584 8752 7588
rect 12196 7644 12260 7648
rect 12196 7588 12200 7644
rect 12200 7588 12256 7644
rect 12256 7588 12260 7644
rect 12196 7584 12260 7588
rect 12276 7644 12340 7648
rect 12276 7588 12280 7644
rect 12280 7588 12336 7644
rect 12336 7588 12340 7644
rect 12276 7584 12340 7588
rect 12356 7644 12420 7648
rect 12356 7588 12360 7644
rect 12360 7588 12416 7644
rect 12416 7588 12420 7644
rect 12356 7584 12420 7588
rect 12436 7644 12500 7648
rect 12436 7588 12440 7644
rect 12440 7588 12496 7644
rect 12496 7588 12500 7644
rect 12436 7584 12500 7588
rect 2826 7100 2890 7104
rect 2826 7044 2830 7100
rect 2830 7044 2886 7100
rect 2886 7044 2890 7100
rect 2826 7040 2890 7044
rect 2906 7100 2970 7104
rect 2906 7044 2910 7100
rect 2910 7044 2966 7100
rect 2966 7044 2970 7100
rect 2906 7040 2970 7044
rect 2986 7100 3050 7104
rect 2986 7044 2990 7100
rect 2990 7044 3046 7100
rect 3046 7044 3050 7100
rect 2986 7040 3050 7044
rect 3066 7100 3130 7104
rect 3066 7044 3070 7100
rect 3070 7044 3126 7100
rect 3126 7044 3130 7100
rect 3066 7040 3130 7044
rect 6574 7100 6638 7104
rect 6574 7044 6578 7100
rect 6578 7044 6634 7100
rect 6634 7044 6638 7100
rect 6574 7040 6638 7044
rect 6654 7100 6718 7104
rect 6654 7044 6658 7100
rect 6658 7044 6714 7100
rect 6714 7044 6718 7100
rect 6654 7040 6718 7044
rect 6734 7100 6798 7104
rect 6734 7044 6738 7100
rect 6738 7044 6794 7100
rect 6794 7044 6798 7100
rect 6734 7040 6798 7044
rect 6814 7100 6878 7104
rect 6814 7044 6818 7100
rect 6818 7044 6874 7100
rect 6874 7044 6878 7100
rect 6814 7040 6878 7044
rect 10322 7100 10386 7104
rect 10322 7044 10326 7100
rect 10326 7044 10382 7100
rect 10382 7044 10386 7100
rect 10322 7040 10386 7044
rect 10402 7100 10466 7104
rect 10402 7044 10406 7100
rect 10406 7044 10462 7100
rect 10462 7044 10466 7100
rect 10402 7040 10466 7044
rect 10482 7100 10546 7104
rect 10482 7044 10486 7100
rect 10486 7044 10542 7100
rect 10542 7044 10546 7100
rect 10482 7040 10546 7044
rect 10562 7100 10626 7104
rect 10562 7044 10566 7100
rect 10566 7044 10622 7100
rect 10622 7044 10626 7100
rect 10562 7040 10626 7044
rect 14070 7100 14134 7104
rect 14070 7044 14074 7100
rect 14074 7044 14130 7100
rect 14130 7044 14134 7100
rect 14070 7040 14134 7044
rect 14150 7100 14214 7104
rect 14150 7044 14154 7100
rect 14154 7044 14210 7100
rect 14210 7044 14214 7100
rect 14150 7040 14214 7044
rect 14230 7100 14294 7104
rect 14230 7044 14234 7100
rect 14234 7044 14290 7100
rect 14290 7044 14294 7100
rect 14230 7040 14294 7044
rect 14310 7100 14374 7104
rect 14310 7044 14314 7100
rect 14314 7044 14370 7100
rect 14370 7044 14374 7100
rect 14310 7040 14374 7044
rect 4700 6556 4764 6560
rect 4700 6500 4704 6556
rect 4704 6500 4760 6556
rect 4760 6500 4764 6556
rect 4700 6496 4764 6500
rect 4780 6556 4844 6560
rect 4780 6500 4784 6556
rect 4784 6500 4840 6556
rect 4840 6500 4844 6556
rect 4780 6496 4844 6500
rect 4860 6556 4924 6560
rect 4860 6500 4864 6556
rect 4864 6500 4920 6556
rect 4920 6500 4924 6556
rect 4860 6496 4924 6500
rect 4940 6556 5004 6560
rect 4940 6500 4944 6556
rect 4944 6500 5000 6556
rect 5000 6500 5004 6556
rect 4940 6496 5004 6500
rect 8448 6556 8512 6560
rect 8448 6500 8452 6556
rect 8452 6500 8508 6556
rect 8508 6500 8512 6556
rect 8448 6496 8512 6500
rect 8528 6556 8592 6560
rect 8528 6500 8532 6556
rect 8532 6500 8588 6556
rect 8588 6500 8592 6556
rect 8528 6496 8592 6500
rect 8608 6556 8672 6560
rect 8608 6500 8612 6556
rect 8612 6500 8668 6556
rect 8668 6500 8672 6556
rect 8608 6496 8672 6500
rect 8688 6556 8752 6560
rect 8688 6500 8692 6556
rect 8692 6500 8748 6556
rect 8748 6500 8752 6556
rect 8688 6496 8752 6500
rect 12196 6556 12260 6560
rect 12196 6500 12200 6556
rect 12200 6500 12256 6556
rect 12256 6500 12260 6556
rect 12196 6496 12260 6500
rect 12276 6556 12340 6560
rect 12276 6500 12280 6556
rect 12280 6500 12336 6556
rect 12336 6500 12340 6556
rect 12276 6496 12340 6500
rect 12356 6556 12420 6560
rect 12356 6500 12360 6556
rect 12360 6500 12416 6556
rect 12416 6500 12420 6556
rect 12356 6496 12420 6500
rect 12436 6556 12500 6560
rect 12436 6500 12440 6556
rect 12440 6500 12496 6556
rect 12496 6500 12500 6556
rect 12436 6496 12500 6500
rect 2826 6012 2890 6016
rect 2826 5956 2830 6012
rect 2830 5956 2886 6012
rect 2886 5956 2890 6012
rect 2826 5952 2890 5956
rect 2906 6012 2970 6016
rect 2906 5956 2910 6012
rect 2910 5956 2966 6012
rect 2966 5956 2970 6012
rect 2906 5952 2970 5956
rect 2986 6012 3050 6016
rect 2986 5956 2990 6012
rect 2990 5956 3046 6012
rect 3046 5956 3050 6012
rect 2986 5952 3050 5956
rect 3066 6012 3130 6016
rect 3066 5956 3070 6012
rect 3070 5956 3126 6012
rect 3126 5956 3130 6012
rect 3066 5952 3130 5956
rect 6574 6012 6638 6016
rect 6574 5956 6578 6012
rect 6578 5956 6634 6012
rect 6634 5956 6638 6012
rect 6574 5952 6638 5956
rect 6654 6012 6718 6016
rect 6654 5956 6658 6012
rect 6658 5956 6714 6012
rect 6714 5956 6718 6012
rect 6654 5952 6718 5956
rect 6734 6012 6798 6016
rect 6734 5956 6738 6012
rect 6738 5956 6794 6012
rect 6794 5956 6798 6012
rect 6734 5952 6798 5956
rect 6814 6012 6878 6016
rect 6814 5956 6818 6012
rect 6818 5956 6874 6012
rect 6874 5956 6878 6012
rect 6814 5952 6878 5956
rect 10322 6012 10386 6016
rect 10322 5956 10326 6012
rect 10326 5956 10382 6012
rect 10382 5956 10386 6012
rect 10322 5952 10386 5956
rect 10402 6012 10466 6016
rect 10402 5956 10406 6012
rect 10406 5956 10462 6012
rect 10462 5956 10466 6012
rect 10402 5952 10466 5956
rect 10482 6012 10546 6016
rect 10482 5956 10486 6012
rect 10486 5956 10542 6012
rect 10542 5956 10546 6012
rect 10482 5952 10546 5956
rect 10562 6012 10626 6016
rect 10562 5956 10566 6012
rect 10566 5956 10622 6012
rect 10622 5956 10626 6012
rect 10562 5952 10626 5956
rect 14070 6012 14134 6016
rect 14070 5956 14074 6012
rect 14074 5956 14130 6012
rect 14130 5956 14134 6012
rect 14070 5952 14134 5956
rect 14150 6012 14214 6016
rect 14150 5956 14154 6012
rect 14154 5956 14210 6012
rect 14210 5956 14214 6012
rect 14150 5952 14214 5956
rect 14230 6012 14294 6016
rect 14230 5956 14234 6012
rect 14234 5956 14290 6012
rect 14290 5956 14294 6012
rect 14230 5952 14294 5956
rect 14310 6012 14374 6016
rect 14310 5956 14314 6012
rect 14314 5956 14370 6012
rect 14370 5956 14374 6012
rect 14310 5952 14374 5956
rect 4700 5468 4764 5472
rect 4700 5412 4704 5468
rect 4704 5412 4760 5468
rect 4760 5412 4764 5468
rect 4700 5408 4764 5412
rect 4780 5468 4844 5472
rect 4780 5412 4784 5468
rect 4784 5412 4840 5468
rect 4840 5412 4844 5468
rect 4780 5408 4844 5412
rect 4860 5468 4924 5472
rect 4860 5412 4864 5468
rect 4864 5412 4920 5468
rect 4920 5412 4924 5468
rect 4860 5408 4924 5412
rect 4940 5468 5004 5472
rect 4940 5412 4944 5468
rect 4944 5412 5000 5468
rect 5000 5412 5004 5468
rect 4940 5408 5004 5412
rect 8448 5468 8512 5472
rect 8448 5412 8452 5468
rect 8452 5412 8508 5468
rect 8508 5412 8512 5468
rect 8448 5408 8512 5412
rect 8528 5468 8592 5472
rect 8528 5412 8532 5468
rect 8532 5412 8588 5468
rect 8588 5412 8592 5468
rect 8528 5408 8592 5412
rect 8608 5468 8672 5472
rect 8608 5412 8612 5468
rect 8612 5412 8668 5468
rect 8668 5412 8672 5468
rect 8608 5408 8672 5412
rect 8688 5468 8752 5472
rect 8688 5412 8692 5468
rect 8692 5412 8748 5468
rect 8748 5412 8752 5468
rect 8688 5408 8752 5412
rect 12196 5468 12260 5472
rect 12196 5412 12200 5468
rect 12200 5412 12256 5468
rect 12256 5412 12260 5468
rect 12196 5408 12260 5412
rect 12276 5468 12340 5472
rect 12276 5412 12280 5468
rect 12280 5412 12336 5468
rect 12336 5412 12340 5468
rect 12276 5408 12340 5412
rect 12356 5468 12420 5472
rect 12356 5412 12360 5468
rect 12360 5412 12416 5468
rect 12416 5412 12420 5468
rect 12356 5408 12420 5412
rect 12436 5468 12500 5472
rect 12436 5412 12440 5468
rect 12440 5412 12496 5468
rect 12496 5412 12500 5468
rect 12436 5408 12500 5412
rect 2826 4924 2890 4928
rect 2826 4868 2830 4924
rect 2830 4868 2886 4924
rect 2886 4868 2890 4924
rect 2826 4864 2890 4868
rect 2906 4924 2970 4928
rect 2906 4868 2910 4924
rect 2910 4868 2966 4924
rect 2966 4868 2970 4924
rect 2906 4864 2970 4868
rect 2986 4924 3050 4928
rect 2986 4868 2990 4924
rect 2990 4868 3046 4924
rect 3046 4868 3050 4924
rect 2986 4864 3050 4868
rect 3066 4924 3130 4928
rect 3066 4868 3070 4924
rect 3070 4868 3126 4924
rect 3126 4868 3130 4924
rect 3066 4864 3130 4868
rect 6574 4924 6638 4928
rect 6574 4868 6578 4924
rect 6578 4868 6634 4924
rect 6634 4868 6638 4924
rect 6574 4864 6638 4868
rect 6654 4924 6718 4928
rect 6654 4868 6658 4924
rect 6658 4868 6714 4924
rect 6714 4868 6718 4924
rect 6654 4864 6718 4868
rect 6734 4924 6798 4928
rect 6734 4868 6738 4924
rect 6738 4868 6794 4924
rect 6794 4868 6798 4924
rect 6734 4864 6798 4868
rect 6814 4924 6878 4928
rect 6814 4868 6818 4924
rect 6818 4868 6874 4924
rect 6874 4868 6878 4924
rect 6814 4864 6878 4868
rect 10322 4924 10386 4928
rect 10322 4868 10326 4924
rect 10326 4868 10382 4924
rect 10382 4868 10386 4924
rect 10322 4864 10386 4868
rect 10402 4924 10466 4928
rect 10402 4868 10406 4924
rect 10406 4868 10462 4924
rect 10462 4868 10466 4924
rect 10402 4864 10466 4868
rect 10482 4924 10546 4928
rect 10482 4868 10486 4924
rect 10486 4868 10542 4924
rect 10542 4868 10546 4924
rect 10482 4864 10546 4868
rect 10562 4924 10626 4928
rect 10562 4868 10566 4924
rect 10566 4868 10622 4924
rect 10622 4868 10626 4924
rect 10562 4864 10626 4868
rect 14070 4924 14134 4928
rect 14070 4868 14074 4924
rect 14074 4868 14130 4924
rect 14130 4868 14134 4924
rect 14070 4864 14134 4868
rect 14150 4924 14214 4928
rect 14150 4868 14154 4924
rect 14154 4868 14210 4924
rect 14210 4868 14214 4924
rect 14150 4864 14214 4868
rect 14230 4924 14294 4928
rect 14230 4868 14234 4924
rect 14234 4868 14290 4924
rect 14290 4868 14294 4924
rect 14230 4864 14294 4868
rect 14310 4924 14374 4928
rect 14310 4868 14314 4924
rect 14314 4868 14370 4924
rect 14370 4868 14374 4924
rect 14310 4864 14374 4868
rect 4700 4380 4764 4384
rect 4700 4324 4704 4380
rect 4704 4324 4760 4380
rect 4760 4324 4764 4380
rect 4700 4320 4764 4324
rect 4780 4380 4844 4384
rect 4780 4324 4784 4380
rect 4784 4324 4840 4380
rect 4840 4324 4844 4380
rect 4780 4320 4844 4324
rect 4860 4380 4924 4384
rect 4860 4324 4864 4380
rect 4864 4324 4920 4380
rect 4920 4324 4924 4380
rect 4860 4320 4924 4324
rect 4940 4380 5004 4384
rect 4940 4324 4944 4380
rect 4944 4324 5000 4380
rect 5000 4324 5004 4380
rect 4940 4320 5004 4324
rect 8448 4380 8512 4384
rect 8448 4324 8452 4380
rect 8452 4324 8508 4380
rect 8508 4324 8512 4380
rect 8448 4320 8512 4324
rect 8528 4380 8592 4384
rect 8528 4324 8532 4380
rect 8532 4324 8588 4380
rect 8588 4324 8592 4380
rect 8528 4320 8592 4324
rect 8608 4380 8672 4384
rect 8608 4324 8612 4380
rect 8612 4324 8668 4380
rect 8668 4324 8672 4380
rect 8608 4320 8672 4324
rect 8688 4380 8752 4384
rect 8688 4324 8692 4380
rect 8692 4324 8748 4380
rect 8748 4324 8752 4380
rect 8688 4320 8752 4324
rect 12196 4380 12260 4384
rect 12196 4324 12200 4380
rect 12200 4324 12256 4380
rect 12256 4324 12260 4380
rect 12196 4320 12260 4324
rect 12276 4380 12340 4384
rect 12276 4324 12280 4380
rect 12280 4324 12336 4380
rect 12336 4324 12340 4380
rect 12276 4320 12340 4324
rect 12356 4380 12420 4384
rect 12356 4324 12360 4380
rect 12360 4324 12416 4380
rect 12416 4324 12420 4380
rect 12356 4320 12420 4324
rect 12436 4380 12500 4384
rect 12436 4324 12440 4380
rect 12440 4324 12496 4380
rect 12496 4324 12500 4380
rect 12436 4320 12500 4324
rect 2826 3836 2890 3840
rect 2826 3780 2830 3836
rect 2830 3780 2886 3836
rect 2886 3780 2890 3836
rect 2826 3776 2890 3780
rect 2906 3836 2970 3840
rect 2906 3780 2910 3836
rect 2910 3780 2966 3836
rect 2966 3780 2970 3836
rect 2906 3776 2970 3780
rect 2986 3836 3050 3840
rect 2986 3780 2990 3836
rect 2990 3780 3046 3836
rect 3046 3780 3050 3836
rect 2986 3776 3050 3780
rect 3066 3836 3130 3840
rect 3066 3780 3070 3836
rect 3070 3780 3126 3836
rect 3126 3780 3130 3836
rect 3066 3776 3130 3780
rect 6574 3836 6638 3840
rect 6574 3780 6578 3836
rect 6578 3780 6634 3836
rect 6634 3780 6638 3836
rect 6574 3776 6638 3780
rect 6654 3836 6718 3840
rect 6654 3780 6658 3836
rect 6658 3780 6714 3836
rect 6714 3780 6718 3836
rect 6654 3776 6718 3780
rect 6734 3836 6798 3840
rect 6734 3780 6738 3836
rect 6738 3780 6794 3836
rect 6794 3780 6798 3836
rect 6734 3776 6798 3780
rect 6814 3836 6878 3840
rect 6814 3780 6818 3836
rect 6818 3780 6874 3836
rect 6874 3780 6878 3836
rect 6814 3776 6878 3780
rect 10322 3836 10386 3840
rect 10322 3780 10326 3836
rect 10326 3780 10382 3836
rect 10382 3780 10386 3836
rect 10322 3776 10386 3780
rect 10402 3836 10466 3840
rect 10402 3780 10406 3836
rect 10406 3780 10462 3836
rect 10462 3780 10466 3836
rect 10402 3776 10466 3780
rect 10482 3836 10546 3840
rect 10482 3780 10486 3836
rect 10486 3780 10542 3836
rect 10542 3780 10546 3836
rect 10482 3776 10546 3780
rect 10562 3836 10626 3840
rect 10562 3780 10566 3836
rect 10566 3780 10622 3836
rect 10622 3780 10626 3836
rect 10562 3776 10626 3780
rect 14070 3836 14134 3840
rect 14070 3780 14074 3836
rect 14074 3780 14130 3836
rect 14130 3780 14134 3836
rect 14070 3776 14134 3780
rect 14150 3836 14214 3840
rect 14150 3780 14154 3836
rect 14154 3780 14210 3836
rect 14210 3780 14214 3836
rect 14150 3776 14214 3780
rect 14230 3836 14294 3840
rect 14230 3780 14234 3836
rect 14234 3780 14290 3836
rect 14290 3780 14294 3836
rect 14230 3776 14294 3780
rect 14310 3836 14374 3840
rect 14310 3780 14314 3836
rect 14314 3780 14370 3836
rect 14370 3780 14374 3836
rect 14310 3776 14374 3780
rect 4700 3292 4764 3296
rect 4700 3236 4704 3292
rect 4704 3236 4760 3292
rect 4760 3236 4764 3292
rect 4700 3232 4764 3236
rect 4780 3292 4844 3296
rect 4780 3236 4784 3292
rect 4784 3236 4840 3292
rect 4840 3236 4844 3292
rect 4780 3232 4844 3236
rect 4860 3292 4924 3296
rect 4860 3236 4864 3292
rect 4864 3236 4920 3292
rect 4920 3236 4924 3292
rect 4860 3232 4924 3236
rect 4940 3292 5004 3296
rect 4940 3236 4944 3292
rect 4944 3236 5000 3292
rect 5000 3236 5004 3292
rect 4940 3232 5004 3236
rect 8448 3292 8512 3296
rect 8448 3236 8452 3292
rect 8452 3236 8508 3292
rect 8508 3236 8512 3292
rect 8448 3232 8512 3236
rect 8528 3292 8592 3296
rect 8528 3236 8532 3292
rect 8532 3236 8588 3292
rect 8588 3236 8592 3292
rect 8528 3232 8592 3236
rect 8608 3292 8672 3296
rect 8608 3236 8612 3292
rect 8612 3236 8668 3292
rect 8668 3236 8672 3292
rect 8608 3232 8672 3236
rect 8688 3292 8752 3296
rect 8688 3236 8692 3292
rect 8692 3236 8748 3292
rect 8748 3236 8752 3292
rect 8688 3232 8752 3236
rect 12196 3292 12260 3296
rect 12196 3236 12200 3292
rect 12200 3236 12256 3292
rect 12256 3236 12260 3292
rect 12196 3232 12260 3236
rect 12276 3292 12340 3296
rect 12276 3236 12280 3292
rect 12280 3236 12336 3292
rect 12336 3236 12340 3292
rect 12276 3232 12340 3236
rect 12356 3292 12420 3296
rect 12356 3236 12360 3292
rect 12360 3236 12416 3292
rect 12416 3236 12420 3292
rect 12356 3232 12420 3236
rect 12436 3292 12500 3296
rect 12436 3236 12440 3292
rect 12440 3236 12496 3292
rect 12496 3236 12500 3292
rect 12436 3232 12500 3236
rect 9628 2892 9692 2956
rect 2826 2748 2890 2752
rect 2826 2692 2830 2748
rect 2830 2692 2886 2748
rect 2886 2692 2890 2748
rect 2826 2688 2890 2692
rect 2906 2748 2970 2752
rect 2906 2692 2910 2748
rect 2910 2692 2966 2748
rect 2966 2692 2970 2748
rect 2906 2688 2970 2692
rect 2986 2748 3050 2752
rect 2986 2692 2990 2748
rect 2990 2692 3046 2748
rect 3046 2692 3050 2748
rect 2986 2688 3050 2692
rect 3066 2748 3130 2752
rect 3066 2692 3070 2748
rect 3070 2692 3126 2748
rect 3126 2692 3130 2748
rect 3066 2688 3130 2692
rect 6574 2748 6638 2752
rect 6574 2692 6578 2748
rect 6578 2692 6634 2748
rect 6634 2692 6638 2748
rect 6574 2688 6638 2692
rect 6654 2748 6718 2752
rect 6654 2692 6658 2748
rect 6658 2692 6714 2748
rect 6714 2692 6718 2748
rect 6654 2688 6718 2692
rect 6734 2748 6798 2752
rect 6734 2692 6738 2748
rect 6738 2692 6794 2748
rect 6794 2692 6798 2748
rect 6734 2688 6798 2692
rect 6814 2748 6878 2752
rect 6814 2692 6818 2748
rect 6818 2692 6874 2748
rect 6874 2692 6878 2748
rect 6814 2688 6878 2692
rect 10322 2748 10386 2752
rect 10322 2692 10326 2748
rect 10326 2692 10382 2748
rect 10382 2692 10386 2748
rect 10322 2688 10386 2692
rect 10402 2748 10466 2752
rect 10402 2692 10406 2748
rect 10406 2692 10462 2748
rect 10462 2692 10466 2748
rect 10402 2688 10466 2692
rect 10482 2748 10546 2752
rect 10482 2692 10486 2748
rect 10486 2692 10542 2748
rect 10542 2692 10546 2748
rect 10482 2688 10546 2692
rect 10562 2748 10626 2752
rect 10562 2692 10566 2748
rect 10566 2692 10622 2748
rect 10622 2692 10626 2748
rect 10562 2688 10626 2692
rect 14070 2748 14134 2752
rect 14070 2692 14074 2748
rect 14074 2692 14130 2748
rect 14130 2692 14134 2748
rect 14070 2688 14134 2692
rect 14150 2748 14214 2752
rect 14150 2692 14154 2748
rect 14154 2692 14210 2748
rect 14210 2692 14214 2748
rect 14150 2688 14214 2692
rect 14230 2748 14294 2752
rect 14230 2692 14234 2748
rect 14234 2692 14290 2748
rect 14290 2692 14294 2748
rect 14230 2688 14294 2692
rect 14310 2748 14374 2752
rect 14310 2692 14314 2748
rect 14314 2692 14370 2748
rect 14370 2692 14374 2748
rect 14310 2688 14374 2692
rect 8156 2620 8220 2684
rect 7788 2348 7852 2412
rect 4700 2204 4764 2208
rect 4700 2148 4704 2204
rect 4704 2148 4760 2204
rect 4760 2148 4764 2204
rect 4700 2144 4764 2148
rect 4780 2204 4844 2208
rect 4780 2148 4784 2204
rect 4784 2148 4840 2204
rect 4840 2148 4844 2204
rect 4780 2144 4844 2148
rect 4860 2204 4924 2208
rect 4860 2148 4864 2204
rect 4864 2148 4920 2204
rect 4920 2148 4924 2204
rect 4860 2144 4924 2148
rect 4940 2204 5004 2208
rect 4940 2148 4944 2204
rect 4944 2148 5000 2204
rect 5000 2148 5004 2204
rect 4940 2144 5004 2148
rect 8448 2204 8512 2208
rect 8448 2148 8452 2204
rect 8452 2148 8508 2204
rect 8508 2148 8512 2204
rect 8448 2144 8512 2148
rect 8528 2204 8592 2208
rect 8528 2148 8532 2204
rect 8532 2148 8588 2204
rect 8588 2148 8592 2204
rect 8528 2144 8592 2148
rect 8608 2204 8672 2208
rect 8608 2148 8612 2204
rect 8612 2148 8668 2204
rect 8668 2148 8672 2204
rect 8608 2144 8672 2148
rect 8688 2204 8752 2208
rect 8688 2148 8692 2204
rect 8692 2148 8748 2204
rect 8748 2148 8752 2204
rect 8688 2144 8752 2148
rect 12196 2204 12260 2208
rect 12196 2148 12200 2204
rect 12200 2148 12256 2204
rect 12256 2148 12260 2204
rect 12196 2144 12260 2148
rect 12276 2204 12340 2208
rect 12276 2148 12280 2204
rect 12280 2148 12336 2204
rect 12336 2148 12340 2204
rect 12276 2144 12340 2148
rect 12356 2204 12420 2208
rect 12356 2148 12360 2204
rect 12360 2148 12416 2204
rect 12416 2148 12420 2204
rect 12356 2144 12420 2148
rect 12436 2204 12500 2208
rect 12436 2148 12440 2204
rect 12440 2148 12496 2204
rect 12496 2148 12500 2204
rect 12436 2144 12500 2148
<< metal4 >>
rect 2818 16896 3138 17456
rect 2818 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3138 16896
rect 2818 15808 3138 16832
rect 2818 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3138 15808
rect 2818 14720 3138 15744
rect 2818 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3138 14720
rect 2818 13632 3138 14656
rect 2818 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3138 13632
rect 2818 12544 3138 13568
rect 2818 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3138 12544
rect 2818 11456 3138 12480
rect 2818 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3138 11456
rect 2818 10368 3138 11392
rect 2818 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3138 10368
rect 2818 9280 3138 10304
rect 2818 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3138 9280
rect 2818 8192 3138 9216
rect 2818 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3138 8192
rect 2818 7104 3138 8128
rect 2818 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3138 7104
rect 2818 6016 3138 7040
rect 2818 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3138 6016
rect 2818 4928 3138 5952
rect 2818 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3138 4928
rect 2818 3840 3138 4864
rect 2818 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3138 3840
rect 2818 2752 3138 3776
rect 2818 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3138 2752
rect 2818 2128 3138 2688
rect 4692 17440 5012 17456
rect 4692 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5012 17440
rect 4692 16352 5012 17376
rect 4692 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5012 16352
rect 4692 15264 5012 16288
rect 4692 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5012 15264
rect 4692 14176 5012 15200
rect 4692 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5012 14176
rect 4692 13088 5012 14112
rect 4692 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5012 13088
rect 4692 12000 5012 13024
rect 4692 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5012 12000
rect 4692 10912 5012 11936
rect 4692 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5012 10912
rect 4692 9824 5012 10848
rect 4692 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5012 9824
rect 4692 8736 5012 9760
rect 4692 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5012 8736
rect 4692 7648 5012 8672
rect 4692 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5012 7648
rect 4692 6560 5012 7584
rect 4692 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5012 6560
rect 4692 5472 5012 6496
rect 4692 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5012 5472
rect 4692 4384 5012 5408
rect 4692 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5012 4384
rect 4692 3296 5012 4320
rect 4692 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5012 3296
rect 4692 2208 5012 3232
rect 4692 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5012 2208
rect 4692 2128 5012 2144
rect 6566 16896 6886 17456
rect 6566 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6886 16896
rect 6566 15808 6886 16832
rect 6566 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6886 15808
rect 6566 14720 6886 15744
rect 6566 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6886 14720
rect 6566 13632 6886 14656
rect 6566 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6886 13632
rect 6566 12544 6886 13568
rect 6566 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6886 12544
rect 6566 11456 6886 12480
rect 6566 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6886 11456
rect 6566 10368 6886 11392
rect 8440 17440 8760 17456
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 16352 8760 17376
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 15264 8760 16288
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 14176 8760 15200
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 13088 8760 14112
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 12000 8760 13024
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 7787 11116 7853 11117
rect 7787 11052 7788 11116
rect 7852 11052 7853 11116
rect 7787 11051 7853 11052
rect 8155 11116 8221 11117
rect 8155 11052 8156 11116
rect 8220 11052 8221 11116
rect 8155 11051 8221 11052
rect 6566 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6886 10368
rect 6566 9280 6886 10304
rect 6566 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6886 9280
rect 6566 8192 6886 9216
rect 6566 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6886 8192
rect 6566 7104 6886 8128
rect 6566 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6886 7104
rect 6566 6016 6886 7040
rect 6566 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6886 6016
rect 6566 4928 6886 5952
rect 6566 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6886 4928
rect 6566 3840 6886 4864
rect 6566 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6886 3840
rect 6566 2752 6886 3776
rect 6566 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6886 2752
rect 6566 2128 6886 2688
rect 7790 2413 7850 11051
rect 8158 2685 8218 11051
rect 8440 10912 8760 11936
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 9824 8760 10848
rect 10314 16896 10634 17456
rect 10314 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10634 16896
rect 10314 15808 10634 16832
rect 10314 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10634 15808
rect 10314 14720 10634 15744
rect 10314 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10634 14720
rect 10314 13632 10634 14656
rect 10314 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10634 13632
rect 10314 12544 10634 13568
rect 10314 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10634 12544
rect 10314 11456 10634 12480
rect 10314 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10634 11456
rect 10314 10368 10634 11392
rect 10314 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10634 10368
rect 8891 10300 8957 10301
rect 8891 10236 8892 10300
rect 8956 10236 8957 10300
rect 8891 10235 8957 10236
rect 9075 10300 9141 10301
rect 9075 10236 9076 10300
rect 9140 10236 9141 10300
rect 9075 10235 9141 10236
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 8736 8760 9760
rect 8894 9757 8954 10235
rect 8891 9756 8957 9757
rect 8891 9692 8892 9756
rect 8956 9692 8957 9756
rect 8891 9691 8957 9692
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 7648 8760 8672
rect 9078 8533 9138 10235
rect 9627 9756 9693 9757
rect 9627 9692 9628 9756
rect 9692 9692 9693 9756
rect 9627 9691 9693 9692
rect 9075 8532 9141 8533
rect 9075 8468 9076 8532
rect 9140 8468 9141 8532
rect 9075 8467 9141 8468
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 6560 8760 7584
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 5472 8760 6496
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 4384 8760 5408
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 3296 8760 4320
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8155 2684 8221 2685
rect 8155 2620 8156 2684
rect 8220 2620 8221 2684
rect 8155 2619 8221 2620
rect 7787 2412 7853 2413
rect 7787 2348 7788 2412
rect 7852 2348 7853 2412
rect 7787 2347 7853 2348
rect 8440 2208 8760 3232
rect 9630 2957 9690 9691
rect 10314 9280 10634 10304
rect 10314 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10634 9280
rect 10314 8192 10634 9216
rect 10314 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10634 8192
rect 10314 7104 10634 8128
rect 10314 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10634 7104
rect 10314 6016 10634 7040
rect 10314 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10634 6016
rect 10314 4928 10634 5952
rect 10314 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10634 4928
rect 10314 3840 10634 4864
rect 10314 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10634 3840
rect 9627 2956 9693 2957
rect 9627 2892 9628 2956
rect 9692 2892 9693 2956
rect 9627 2891 9693 2892
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2128 8760 2144
rect 10314 2752 10634 3776
rect 10314 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10634 2752
rect 10314 2128 10634 2688
rect 12188 17440 12508 17456
rect 12188 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12508 17440
rect 12188 16352 12508 17376
rect 12188 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12508 16352
rect 12188 15264 12508 16288
rect 12188 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12508 15264
rect 12188 14176 12508 15200
rect 12188 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12508 14176
rect 12188 13088 12508 14112
rect 12188 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12508 13088
rect 12188 12000 12508 13024
rect 12188 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12508 12000
rect 12188 10912 12508 11936
rect 12188 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12508 10912
rect 12188 9824 12508 10848
rect 12188 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12508 9824
rect 12188 8736 12508 9760
rect 12188 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12508 8736
rect 12188 7648 12508 8672
rect 12188 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12508 7648
rect 12188 6560 12508 7584
rect 12188 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12508 6560
rect 12188 5472 12508 6496
rect 12188 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12508 5472
rect 12188 4384 12508 5408
rect 12188 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12508 4384
rect 12188 3296 12508 4320
rect 12188 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12508 3296
rect 12188 2208 12508 3232
rect 12188 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12508 2208
rect 12188 2128 12508 2144
rect 14062 16896 14382 17456
rect 14062 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14382 16896
rect 14062 15808 14382 16832
rect 14062 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14382 15808
rect 14062 14720 14382 15744
rect 14062 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14382 14720
rect 14062 13632 14382 14656
rect 14062 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14382 13632
rect 14062 12544 14382 13568
rect 14062 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14382 12544
rect 14062 11456 14382 12480
rect 14062 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14382 11456
rect 14062 10368 14382 11392
rect 14062 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14382 10368
rect 14062 9280 14382 10304
rect 14062 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14382 9280
rect 14062 8192 14382 9216
rect 14062 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14382 8192
rect 14062 7104 14382 8128
rect 14062 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14382 7104
rect 14062 6016 14382 7040
rect 14062 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14382 6016
rect 14062 4928 14382 5952
rect 14062 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14382 4928
rect 14062 3840 14382 4864
rect 14062 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14382 3840
rect 14062 2752 14382 3776
rect 14062 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14382 2752
rect 14062 2128 14382 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 1564 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 2116 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 8924 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 12512 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 12880 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 13248 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 13616 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 14076 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 14352 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 14720 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 15088 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 15272 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 15456 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 9200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 9568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 9936 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 10304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 10672 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 11040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 11684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 11868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 12144 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 9476 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 12696 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 13892 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 13432 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 14260 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 14444 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 15364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 14904 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 15732 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 14720 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 15456 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 8832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 9752 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 11316 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 10856 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 11500 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 11776 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 12052 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 12328 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 1840 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91
timestamp 1649977179
transform 1 0 9476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95
timestamp 1649977179
transform 1 0 9844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99
timestamp 1649977179
transform 1 0 10212 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103
timestamp 1649977179
transform 1 0 10580 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107
timestamp 1649977179
transform 1 0 10948 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119
timestamp 1649977179
transform 1 0 12052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123
timestamp 1649977179
transform 1 0 12420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_127
timestamp 1649977179
transform 1 0 12788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131
timestamp 1649977179
transform 1 0 13156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_135
timestamp 1649977179
transform 1 0 13524 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1649977179
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_147
timestamp 1649977179
transform 1 0 14628 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_151
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_155
timestamp 1649977179
transform 1 0 15364 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_13 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_25 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3404 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_31
timestamp 1649977179
transform 1 0 3956 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_36
timestamp 1649977179
transform 1 0 4416 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_48 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_85
timestamp 1649977179
transform 1 0 8924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_88
timestamp 1649977179
transform 1 0 9200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_92
timestamp 1649977179
transform 1 0 9568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_96
timestamp 1649977179
transform 1 0 9936 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_100
timestamp 1649977179
transform 1 0 10304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_104
timestamp 1649977179
transform 1 0 10672 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1649977179
transform 1 0 12144 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_124
timestamp 1649977179
transform 1 0 12512 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_128
timestamp 1649977179
transform 1 0 12880 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1649977179
transform 1 0 13248 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_136
timestamp 1649977179
transform 1 0 13616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_141
timestamp 1649977179
transform 1 0 14076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_144
timestamp 1649977179
transform 1 0 14352 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_148
timestamp 1649977179
transform 1 0 14720 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_157
timestamp 1649977179
transform 1 0 15548 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_19
timestamp 1649977179
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_31
timestamp 1649977179
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_43
timestamp 1649977179
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_157
timestamp 1649977179
transform 1 0 15548 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_157
timestamp 1649977179
transform 1 0 15548 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_24
timestamp 1649977179
transform 1 0 3312 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_36
timestamp 1649977179
transform 1 0 4416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_40
timestamp 1649977179
transform 1 0 4784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_46
timestamp 1649977179
transform 1 0 5336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_65
timestamp 1649977179
transform 1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_71
timestamp 1649977179
transform 1 0 7636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_83
timestamp 1649977179
transform 1 0 8740 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_87
timestamp 1649977179
transform 1 0 9108 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_91
timestamp 1649977179
transform 1 0 9476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1649977179
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_157
timestamp 1649977179
transform 1 0 15548 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_7
timestamp 1649977179
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_19
timestamp 1649977179
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_31
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_43
timestamp 1649977179
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_74
timestamp 1649977179
transform 1 0 7912 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_84
timestamp 1649977179
transform 1 0 8832 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_96
timestamp 1649977179
transform 1 0 9936 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1649977179
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_127
timestamp 1649977179
transform 1 0 12788 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_139
timestamp 1649977179
transform 1 0 13892 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_151
timestamp 1649977179
transform 1 0 14996 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_61
timestamp 1649977179
transform 1 0 6716 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_88
timestamp 1649977179
transform 1 0 9200 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_100
timestamp 1649977179
transform 1 0 10304 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_112
timestamp 1649977179
transform 1 0 11408 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_124
timestamp 1649977179
transform 1 0 12512 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_24
timestamp 1649977179
transform 1 0 3312 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_36
timestamp 1649977179
transform 1 0 4416 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_47
timestamp 1649977179
transform 1 0 5428 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_91
timestamp 1649977179
transform 1 0 9476 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_95
timestamp 1649977179
transform 1 0 9844 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_100
timestamp 1649977179
transform 1 0 10304 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_104
timestamp 1649977179
transform 1 0 10672 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_157
timestamp 1649977179
transform 1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_37
timestamp 1649977179
transform 1 0 4508 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_73
timestamp 1649977179
transform 1 0 7820 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_134
timestamp 1649977179
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_23
timestamp 1649977179
transform 1 0 3220 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_28
timestamp 1649977179
transform 1 0 3680 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_40
timestamp 1649977179
transform 1 0 4784 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1649977179
transform 1 0 5520 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_91
timestamp 1649977179
transform 1 0 9476 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_98
timestamp 1649977179
transform 1 0 10120 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1649977179
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_157
timestamp 1649977179
transform 1 0 15548 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_61
timestamp 1649977179
transform 1 0 6716 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_94
timestamp 1649977179
transform 1 0 9752 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_106
timestamp 1649977179
transform 1 0 10856 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_118
timestamp 1649977179
transform 1 0 11960 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_130
timestamp 1649977179
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_8
timestamp 1649977179
transform 1 0 1840 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_20
timestamp 1649977179
transform 1 0 2944 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_32
timestamp 1649977179
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_44
timestamp 1649977179
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_65
timestamp 1649977179
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_84
timestamp 1649977179
transform 1 0 8832 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_96
timestamp 1649977179
transform 1 0 9936 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1649977179
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_157
timestamp 1649977179
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_46
timestamp 1649977179
transform 1 0 5336 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_58
timestamp 1649977179
transform 1 0 6440 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_66
timestamp 1649977179
transform 1 0 7176 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_71
timestamp 1649977179
transform 1 0 7636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_92
timestamp 1649977179
transform 1 0 9568 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_104
timestamp 1649977179
transform 1 0 10672 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_116
timestamp 1649977179
transform 1 0 11776 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_128
timestamp 1649977179
transform 1 0 12880 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_31
timestamp 1649977179
transform 1 0 3956 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1649977179
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_146
timestamp 1649977179
transform 1 0 14536 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_154
timestamp 1649977179
transform 1 0 15272 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_35
timestamp 1649977179
transform 1 0 4324 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_44
timestamp 1649977179
transform 1 0 5152 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_157
timestamp 1649977179
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_157
timestamp 1649977179
transform 1 0 15548 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_5
timestamp 1649977179
transform 1 0 1564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_17
timestamp 1649977179
transform 1 0 2668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_29
timestamp 1649977179
transform 1 0 3772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_41
timestamp 1649977179
transform 1 0 4876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1649977179
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_153
timestamp 1649977179
transform 1 0 15180 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_11
timestamp 1649977179
transform 1 0 2116 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1649977179
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_34
timestamp 1649977179
transform 1 0 4232 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_46
timestamp 1649977179
transform 1 0 5336 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_58
timestamp 1649977179
transform 1 0 6440 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_70
timestamp 1649977179
transform 1 0 7544 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1649977179
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1649977179
transform 1 0 9476 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_94
timestamp 1649977179
transform 1 0 9752 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_98
timestamp 1649977179
transform 1 0 10120 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_106
timestamp 1649977179
transform 1 0 10856 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_110
timestamp 1649977179
transform 1 0 11224 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_113
timestamp 1649977179
transform 1 0 11500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_116
timestamp 1649977179
transform 1 0 11776 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_119
timestamp 1649977179
transform 1 0 12052 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_122
timestamp 1649977179
transform 1 0 12328 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_126
timestamp 1649977179
transform 1 0 12696 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_134
timestamp 1649977179
transform 1 0 13432 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_145
timestamp 1649977179
transform 1 0 14444 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_150
timestamp 1649977179
transform 1 0 14904 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_29
timestamp 1649977179
transform 1 0 3772 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_89
timestamp 1649977179
transform 1 0 9292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_97
timestamp 1649977179
transform 1 0 10028 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_101
timestamp 1649977179
transform 1 0 10396 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_129
timestamp 1649977179
transform 1 0 12972 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_133
timestamp 1649977179
transform 1 0 13340 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_139
timestamp 1649977179
transform 1 0 13892 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 16008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 16008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 16008 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 16008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 16008 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 16008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 16008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 16008 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 16008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 16008 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 16008 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 16008 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 16008 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 16008 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 16008 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _02_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _03_
timestamp 1649977179
transform 1 0 5060 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _04_
timestamp 1649977179
transform 1 0 5704 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _05_
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _06_
timestamp 1649977179
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _07_
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _08_
timestamp 1649977179
transform 1 0 7544 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _09_
timestamp 1649977179
transform 1 0 7820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _10_
timestamp 1649977179
transform 1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _11_
timestamp 1649977179
transform 1 0 7360 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp 1649977179
transform 1 0 9200 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _13_
timestamp 1649977179
transform 1 0 9568 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _14_
timestamp 1649977179
transform 1 0 10028 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1649977179
transform 1 0 11224 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _16_
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 1649977179
transform 1 0 9292 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _18_
timestamp 1649977179
transform 1 0 12052 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1649977179
transform 1 0 12604 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1649977179
transform 1 0 13156 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _21_
timestamp 1649977179
transform -1 0 14536 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1649977179
transform 1 0 4508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1649977179
transform 1 0 4784 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp 1649977179
transform 1 0 5060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1649977179
transform 1 0 5704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _26_
timestamp 1649977179
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 1649977179
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _28_
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _29_
timestamp 1649977179
transform 1 0 6624 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp 1649977179
transform 1 0 8280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _31_
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1649977179
transform 1 0 7360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1649977179
transform 1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1649977179
transform 1 0 9568 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1649977179
transform 1 0 10672 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1649977179
transform 1 0 10948 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1649977179
transform 1 0 11500 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1649977179
transform 1 0 9200 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1649977179
transform 1 0 11776 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1649977179
transform 1 0 12328 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1649977179
transform 1 0 12880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1649977179
transform 1 0 4048 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8096 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 1932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 12512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform 1 0 13248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform 1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 14720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform 1 0 15088 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform 1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform 1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform 1 0 9568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform 1 0 9936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform 1 0 10672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform 1 0 12144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform 1 0 9016 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform 1 0 12696 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform 1 0 13064 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform 1 0 13432 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform 1 0 14352 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform 1 0 14628 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform 1 0 14904 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 15272 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform 1 0 14996 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform 1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform 1 0 9384 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform 1 0 9752 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform 1 0 10120 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 10488 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform 1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform 1 0 11776 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform 1 0 12052 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform 1 0 12328 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform -1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform -1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5888 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_2  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5152 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform -1 0 3312 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9200 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8372 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6808 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7728 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform -1 0 9476 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform -1 0 8832 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9844 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8004 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9016 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_0.mux_l2_in_3__89 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8832 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7084 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5060 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output45 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15364 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1649977179
transform -1 0 1840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1649977179
transform -1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1649977179
transform -1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1649977179
transform -1 0 6256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1649977179
transform -1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1649977179
transform -1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform -1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform -1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform -1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform -1 0 8832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform -1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform -1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform -1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform -1 0 2944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform -1 0 3680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform -1 0 4416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform -1 0 4416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform -1 0 1840 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform -1 0 5520 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform -1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform -1 0 6256 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform -1 0 6808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 7176 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform -1 0 7544 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 7912 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 8280 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 8648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform -1 0 9292 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 2208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform -1 0 2576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform -1 0 2944 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform -1 0 3312 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform -1 0 3680 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform -1 0 4232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform -1 0 4416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform -1 0 4784 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 5152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 15364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12604 0 -1 8704
box -38 -48 1142 592
<< labels >>
flabel metal2 s 1214 19200 1270 20000 0 FreeSans 224 90 0 0 IO_ISOL_N
port 0 nsew signal input
flabel metal4 s 4692 2128 5012 17456 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 8440 2128 8760 17456 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 12188 2128 12508 17456 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 2818 2128 3138 17456 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 6566 2128 6886 17456 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 10314 2128 10634 17456 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 14062 2128 14382 17456 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal3 s 0 18096 800 18216 0 FreeSans 480 0 0 0 ccff_head
port 3 nsew signal input
flabel metal3 s 16400 12384 17200 12504 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 5 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 6 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 7 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 8 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 9 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 10 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 11 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 12 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 13 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 14 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 15 nsew signal input
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 16 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 17 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 18 nsew signal input
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 19 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 20 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 21 nsew signal input
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 22 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 23 nsew signal input
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 24 nsew signal input
flabel metal2 s 1398 0 1454 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 25 nsew signal tristate
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 26 nsew signal tristate
flabel metal2 s 5446 0 5502 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 27 nsew signal tristate
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 28 nsew signal tristate
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 29 nsew signal tristate
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 30 nsew signal tristate
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 31 nsew signal tristate
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 32 nsew signal tristate
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 33 nsew signal tristate
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 34 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 35 nsew signal tristate
flabel metal2 s 1766 0 1822 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 36 nsew signal tristate
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 37 nsew signal tristate
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 38 nsew signal tristate
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 39 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 40 nsew signal tristate
flabel metal2 s 3606 0 3662 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 41 nsew signal tristate
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 42 nsew signal tristate
flabel metal2 s 4342 0 4398 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 43 nsew signal tristate
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 44 nsew signal tristate
flabel metal2 s 8942 19200 8998 20000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 45 nsew signal input
flabel metal2 s 12622 19200 12678 20000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 46 nsew signal input
flabel metal2 s 12990 19200 13046 20000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 47 nsew signal input
flabel metal2 s 13358 19200 13414 20000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 48 nsew signal input
flabel metal2 s 13726 19200 13782 20000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 49 nsew signal input
flabel metal2 s 14094 19200 14150 20000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 50 nsew signal input
flabel metal2 s 14462 19200 14518 20000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 51 nsew signal input
flabel metal2 s 14830 19200 14886 20000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 52 nsew signal input
flabel metal2 s 15198 19200 15254 20000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 53 nsew signal input
flabel metal2 s 15566 19200 15622 20000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 54 nsew signal input
flabel metal2 s 15934 19200 15990 20000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 55 nsew signal input
flabel metal2 s 9310 19200 9366 20000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 56 nsew signal input
flabel metal2 s 9678 19200 9734 20000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 57 nsew signal input
flabel metal2 s 10046 19200 10102 20000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 58 nsew signal input
flabel metal2 s 10414 19200 10470 20000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 59 nsew signal input
flabel metal2 s 10782 19200 10838 20000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 60 nsew signal input
flabel metal2 s 11150 19200 11206 20000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 61 nsew signal input
flabel metal2 s 11518 19200 11574 20000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 62 nsew signal input
flabel metal2 s 11886 19200 11942 20000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 63 nsew signal input
flabel metal2 s 12254 19200 12310 20000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 64 nsew signal input
flabel metal2 s 1582 19200 1638 20000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 65 nsew signal tristate
flabel metal2 s 5262 19200 5318 20000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 66 nsew signal tristate
flabel metal2 s 5630 19200 5686 20000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 67 nsew signal tristate
flabel metal2 s 5998 19200 6054 20000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 68 nsew signal tristate
flabel metal2 s 6366 19200 6422 20000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 69 nsew signal tristate
flabel metal2 s 6734 19200 6790 20000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 70 nsew signal tristate
flabel metal2 s 7102 19200 7158 20000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 71 nsew signal tristate
flabel metal2 s 7470 19200 7526 20000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 72 nsew signal tristate
flabel metal2 s 7838 19200 7894 20000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 73 nsew signal tristate
flabel metal2 s 8206 19200 8262 20000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 74 nsew signal tristate
flabel metal2 s 8574 19200 8630 20000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 75 nsew signal tristate
flabel metal2 s 1950 19200 2006 20000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 76 nsew signal tristate
flabel metal2 s 2318 19200 2374 20000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 77 nsew signal tristate
flabel metal2 s 2686 19200 2742 20000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 78 nsew signal tristate
flabel metal2 s 3054 19200 3110 20000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 79 nsew signal tristate
flabel metal2 s 3422 19200 3478 20000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 80 nsew signal tristate
flabel metal2 s 3790 19200 3846 20000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 81 nsew signal tristate
flabel metal2 s 4158 19200 4214 20000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 82 nsew signal tristate
flabel metal2 s 4526 19200 4582 20000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 83 nsew signal tristate
flabel metal2 s 4894 19200 4950 20000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 84 nsew signal tristate
flabel metal3 s 0 8304 800 8424 0 FreeSans 480 0 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 85 nsew signal tristate
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 86 nsew signal input
flabel metal3 s 0 14832 800 14952 0 FreeSans 480 0 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 87 nsew signal tristate
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 left_grid_pin_0_
port 88 nsew signal tristate
flabel metal3 s 16400 7488 17200 7608 0 FreeSans 480 0 0 0 prog_clk_0_E_in
port 89 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_0_
port 90 nsew signal input
flabel metal3 s 16400 2592 17200 2712 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_1_lower
port 91 nsew signal tristate
flabel metal3 s 16400 17280 17200 17400 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_1_upper
port 92 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 17200 20000
<< end >>
